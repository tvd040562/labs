* NGSPICE file created from cust_rom.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

.subckt cust_rom VGND VPWR addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6]
+ addr0[7] clk0 cs0 dout0[0] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15]
+ dout0[16] dout0[17] dout0[18] dout0[19] dout0[1] dout0[20] dout0[21] dout0[22] dout0[23]
+ dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[2] dout0[30] dout0[31]
+ dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[32]
XFILLER_0_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1270_ _0539_ _0541_ _0546_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_14_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0985_ net112 net78 net76 net116 VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout127 addr0_reg\[3\] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
Xfanout105 _0697_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_4
Xfanout116 _0667_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dlymetal6s2s_1
X_1399_ net42 _0658_ _0666_ net151 net137 VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__o32a_1
Xfanout138 net139 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_37_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0770_ net124 net119 net122 net126 VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__nor4b_1
X_1322_ _0096_ _0193_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__or2_1
X_1253_ _0191_ _0193_ _0234_ _0405_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__or4_1
X_1184_ _0060_ _0228_ _0446_ _0466_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__or4_1
X_0968_ _0065_ _0259_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0899_ _0115_ _0185_ _0186_ _0187_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__or4_2
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0822_ net106 net90 net85 net98 VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_31_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0753_ _0040_ _0043_ _0044_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__or3_1
X_1236_ _0119_ _0199_ _0209_ _0514_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__or4_1
X_1305_ _0158_ _0576_ _0577_ _0578_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__or4_1
X_1167_ _0141_ _0205_ _0230_ _0248_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__or4_1
X_1098_ _0099_ _0102_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_22_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire100 _0699_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
X_1021_ _0136_ _0142_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0805_ net78 net49 net47 net76 VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__a22o_2
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0736_ net91 net89 net84 net94 VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__a22o_2
XFILLER_0_24_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1219_ _0166_ _0489_ _0497_ _0499_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold30 net23 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_5 _0060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1004_ _0069_ _0295_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0719_ net117 net115 net113 net111 VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__a22o_2
Xoutput20 net20 VGND VGND VPWR VPWR dout0[19] sky130_fd_sc_hd__clkbuf_4
Xoutput31 net31 VGND VGND VPWR VPWR dout0[29] sky130_fd_sc_hd__buf_2
XFILLER_0_27_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0984_ net116 net113 net112 net117 VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout128 addr0_reg\[3\] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_1
Xfanout106 _0697_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_2
Xfanout139 net9 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__buf_2
X_1467_ clknet_2_0__leaf_clk0 net8 VGND VGND VPWR VPWR addr0_reg\[7\] sky130_fd_sc_hd__dfxtp_1
X_1398_ _0163_ _0659_ _0662_ _0665_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__or4_1
Xfanout117 _0657_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_37_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1321_ _0201_ _0231_ _0366_ _0548_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__or4_1
X_1252_ _0487_ _0489_ _0527_ _0529_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__or4_1
X_1183_ _0049_ _0389_ _0414_ _0459_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0967_ net58 net55 _0046_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__o21ba_1
X_0898_ _0185_ _0186_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0821_ _0110_ _0112_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__or2_1
X_0752_ net79 net74 net72 net77 VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__a22o_2
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1235_ _0090_ _0161_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__or2_2
X_1166_ _0069_ _0272_ _0297_ _0411_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1304_ _0165_ _0171_ _0219_ _0250_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__or4_1
X_1097_ net44 _0381_ _0384_ net163 net139 VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__o32a_1
XFILLER_0_35_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1020_ _0086_ _0310_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__or2_1
X_0735_ net132 net130 net128 net134 VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__nor4b_1
X_0804_ _0093_ _0094_ _0095_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1149_ net135 _0082_ _0431_ _0432_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1218_ _0068_ _0268_ _0307_ _0498_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold31 net27 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 net32 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_6 _0060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1003_ net66 net59 net56 net68 VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__a22o_2
XFILLER_0_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0718_ net126 net124 net119 net122 VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__nor4_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput32 net32 VGND VGND VPWR VPWR dout0[2] sky130_fd_sc_hd__clkbuf_4
Xoutput10 net10 VGND VGND VPWR VPWR dout0[0] sky130_fd_sc_hd__buf_2
Xoutput21 net21 VGND VGND VPWR VPWR dout0[1] sky130_fd_sc_hd__buf_2
XFILLER_0_26_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0983_ _0109_ _0274_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_14_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout129 addr0_reg\[2\] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
Xfanout118 _0657_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
Xfanout107 _0695_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_2
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1466_ clknet_2_0__leaf_clk0 net7 VGND VGND VPWR VPWR addr0_reg\[6\] sky130_fd_sc_hd__dfxtp_1
X_1397_ _0430_ _0573_ _0663_ _0664_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_37_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1320_ _0074_ _0076_ _0221_ _0244_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__or4_1
X_1182_ _0252_ _0300_ _0406_ _0460_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_19_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1251_ _0069_ _0149_ _0297_ _0491_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0966_ net109 net58 net55 net107 VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__a22o_1
X_0897_ _0115_ _0186_ _0187_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__or3_1
X_1449_ clknet_2_3__leaf_clk0 _0021_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_2_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0751_ net75 net69 net67 net73 VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__a22o_2
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0820_ _0702_ _0111_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__nor2_1
X_1303_ _0180_ _0288_ _0305_ _0308_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__or4_1
X_1165_ _0149_ _0446_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__or2_1
X_1234_ _0107_ _0225_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__or2_1
X_1096_ _0370_ _0375_ _0382_ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__or4_1
X_0949_ _0239_ _0240_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__or2_2
XFILLER_0_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0734_ net134 net131 net129 net128 VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__and4_1
X_0803_ net95 net58 net56 net101 VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1079_ _0058_ _0171_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__or2_1
X_1148_ _0100_ _0194_ _0238_ _0314_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__or4_1
X_1217_ _0705_ _0711_ _0301_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold32 net34 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 net29 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 net16 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_7 _0082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1002_ _0696_ _0105_ _0290_ _0292_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__or4_1
X_0717_ net133 net129 net127 net131 VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput22 net22 VGND VGND VPWR VPWR dout0[20] sky130_fd_sc_hd__buf_2
Xoutput33 net33 VGND VGND VPWR VPWR dout0[30] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput11 net11 VGND VGND VPWR VPWR dout0[10] sky130_fd_sc_hd__buf_2
XFILLER_0_41_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0982_ net111 net68 net66 net116 VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_14_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout108 _0695_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout119 net120 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
X_1465_ clknet_2_0__leaf_clk0 net6 VGND VGND VPWR VPWR addr0_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1396_ _0710_ _0131_ _0282_ _0285_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_37_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1250_ _0693_ _0221_ _0274_ _0285_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__or4_1
X_1181_ _0355_ _0457_ _0461_ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0896_ _0186_ _0187_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__or2_1
X_0965_ _0144_ _0216_ _0255_ _0256_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__or4_2
X_1448_ clknet_2_3__leaf_clk0 _0020_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1379_ net43 _0643_ _0646_ net149 net139 VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_25_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout90 _0708_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
X_0750_ net134 net132 net130 net128 VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1233_ _0094_ _0095_ _0261_ _0511_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__or4_2
XFILLER_0_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1302_ _0101_ _0262_ _0574_ _0575_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_47_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1164_ _0057_ _0171_ _0246_ _0447_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__or4_1
X_1095_ _0240_ _0365_ _0368_ _0373_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0948_ net74 net54 net52 net72 VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__a22o_2
X_0879_ _0059_ _0170_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__or2_2
XFILLER_0_33_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0802_ net89 net58 net55 net84 VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__a22o_2
XFILLER_0_21_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0733_ net102 net94 net92 net96 VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__a22o_2
X_1216_ _0189_ _0371_ _0428_ _0490_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1147_ _0140_ _0229_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__or2_1
X_1078_ _0189_ _0296_ _0297_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__or3_2
XFILLER_0_30_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_45_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold22 net35 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 net28 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_8 _0130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1001_ _0696_ _0292_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0716_ net119 net122 net126 net124 VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__and4b_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput23 net23 VGND VGND VPWR VPWR dout0[21] sky130_fd_sc_hd__buf_2
Xoutput34 net34 VGND VGND VPWR VPWR dout0[31] sky130_fd_sc_hd__buf_2
Xoutput12 net12 VGND VGND VPWR VPWR dout0[11] sky130_fd_sc_hd__buf_2
XFILLER_0_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_32_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0981_ _0093_ _0094_ _0095_ _0270_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__or4_2
XFILLER_0_38_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1464_ clknet_2_0__leaf_clk0 net5 VGND VGND VPWR VPWR addr0_reg\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1395_ _0705_ _0203_ _0275_ _0277_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__or4_1
Xfanout109 _0694_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_11_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1180_ _0053_ _0275_ _0462_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0964_ _0218_ _0224_ _0228_ _0231_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0895_ net114 net106 net98 net118 VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__a22o_2
XFILLER_0_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1447_ clknet_2_1__leaf_clk0 _0019_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfxtp_1
X_1378_ _0425_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout91 _0706_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
Xfanout80 net81 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_2
X_1232_ _0693_ _0696_ _0130_ _0192_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1301_ _0076_ _0090_ _0181_ _0264_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_47_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1094_ _0169_ _0206_ _0371_ _0374_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__or4_1
X_1163_ net135 _0693_ net46 _0329_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0947_ net102 net74 net72 net96 VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0878_ net66 net62 net60 net68 VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__a22o_2
Xwire104 _0698_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
Xclkload0 clknet_2_0__leaf_clk0 VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_44_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0801_ net115 net55 _0702_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_24_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0732_ net125 net123 net120 net121 VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__and4b_1
XFILLER_0_21_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1146_ _0707_ _0118_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__or2_1
X_1215_ _0235_ _0492_ _0494_ _0495_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__or4_2
X_1077_ _0236_ _0239_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__or2_1
Xhold23 net36 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 net12 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_9 _0132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1000_ net115 net112 _0046_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0715_ net133 net127 net129 net131 VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_12_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1129_ _0105_ _0259_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput35 net35 VGND VGND VPWR VPWR dout0[3] sky130_fd_sc_hd__clkbuf_4
Xoutput24 net24 VGND VGND VPWR VPWR dout0[22] sky130_fd_sc_hd__buf_2
Xoutput13 net13 VGND VGND VPWR VPWR dout0[12] sky130_fd_sc_hd__buf_2
XFILLER_0_11_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0980_ _0093_ _0270_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1463_ clknet_2_1__leaf_clk0 net4 VGND VGND VPWR VPWR addr0_reg\[3\] sky130_fd_sc_hd__dfxtp_1
X_1394_ _0149_ _0326_ _0660_ _0661_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0894_ net98 net79 net77 net106 VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0963_ _0235_ _0243_ _0247_ _0254_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1377_ _0200_ _0228_ _0231_ _0644_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__or4_1
X_1446_ clknet_2_3__leaf_clk0 _0018_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout81 _0713_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_2
Xfanout92 _0706_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_1
XFILLER_0_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1162_ _0185_ _0186_ _0187_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__or3_1
X_1231_ net43 _0509_ _0510_ net141 net138 VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__o32a_1
X_1300_ _0088_ _0125_ _0134_ _0225_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1093_ _0377_ _0378_ _0379_ _0380_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__or4_1
X_0946_ _0236_ _0237_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_30_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0877_ _0122_ _0164_ _0166_ _0167_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1429_ clknet_2_2__leaf_clk0 _0001_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfxtp_1
Xclkload1 clknet_2_1__leaf_clk0 VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__bufinv_16
Xcust_rom_140 VGND VGND VPWR VPWR cust_rom_140/HI dout0[32] sky130_fd_sc_hd__conb_1
XFILLER_0_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0731_ _0701_ _0704_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__or2_2
XFILLER_0_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0800_ _0088_ _0089_ _0090_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1145_ _0064_ _0258_ _0259_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__or3_2
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1214_ _0049_ _0102_ _0270_ _0282_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1076_ net44 _0359_ _0364_ net162 net139 VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__o32a_1
XFILLER_0_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0929_ net117 net93 net91 net113 VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a22o_2
Xhold13 net33 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 net17 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0714_ net138 VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1059_ _0043_ _0220_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__or2_1
X_1128_ _0064_ _0068_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput36 net36 VGND VGND VPWR VPWR dout0[4] sky130_fd_sc_hd__clkbuf_4
Xoutput14 net14 VGND VGND VPWR VPWR dout0[13] sky130_fd_sc_hd__clkbuf_4
Xoutput25 net25 VGND VGND VPWR VPWR dout0[23] sky130_fd_sc_hd__buf_2
XFILLER_0_26_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1462_ clknet_2_1__leaf_clk0 net3 VGND VGND VPWR VPWR addr0_reg\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1393_ _0102_ _0103_ _0241_ _0308_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_19_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0893_ net106 net98 _0046_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__o21ba_2
X_0962_ _0117_ _0248_ _0249_ _0250_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__or4_1
X_1445_ clknet_2_2__leaf_clk0 _0017_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfxtp_1
X_1376_ _0094_ _0137_ _0142_ _0270_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout82 net83 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_2
Xfanout60 _0048_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
Xfanout93 net94 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_2
XFILLER_0_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1092_ _0710_ _0121_ _0142_ _0250_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__or4_1
X_1230_ _0306_ _0407_ _0445_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__or3_1
X_1161_ _0056_ _0065_ _0263_ _0444_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__or4_2
XFILLER_0_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0876_ _0166_ _0167_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__or2_1
X_0945_ net80 net75 _0702_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_30_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1428_ clknet_2_0__leaf_clk0 _0000_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfxtp_1
X_1359_ _0079_ _0159_ _0279_ _0617_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload2 clknet_2_3__leaf_clk0 VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0730_ net105 net94 _0702_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__o21ba_1
X_1213_ _0288_ _0291_ _0493_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1075_ _0360_ _0361_ _0362_ _0363_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__or4_1
X_1144_ _0064_ _0258_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0928_ _0040_ _0219_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0859_ _0108_ _0115_ _0117_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__or3_1
Xhold14 net41 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 net38 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_7_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1127_ _0137_ _0412_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__or2_1
X_1058_ _0711_ _0244_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput26 net26 VGND VGND VPWR VPWR dout0[24] sky130_fd_sc_hd__buf_2
Xoutput37 net37 VGND VGND VPWR VPWR dout0[5] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR dout0[14] sky130_fd_sc_hd__buf_2
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1461_ clknet_2_1__leaf_clk0 net2 VGND VGND VPWR VPWR addr0_reg\[1\] sky130_fd_sc_hd__dfxtp_1
X_1392_ _0209_ _0230_ _0281_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0961_ _0117_ _0248_ _0249_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_20_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0892_ _0079_ _0159_ _0173_ _0183_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1375_ _0526_ _0639_ _0641_ _0642_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__or4_1
X_1444_ clknet_2_0__leaf_clk0 _0016_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout50 _0070_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout94 _0703_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout83 _0712_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
Xfanout72 _0039_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_2
Xfanout61 _0048_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_0_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1091_ _0076_ _0110_ _0178_ _0210_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__or4_1
X_1160_ _0040_ _0208_ _0210_ _0213_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__or4_1
X_0944_ net85 net75 net73 net90 VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_30_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0875_ net60 net53 net51 net62 VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__a22o_2
XFILLER_0_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1427_ net135 _0207_ _0257_ _0692_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__o31a_1
X_1358_ _0234_ _0242_ _0458_ _0626_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__or4_1
X_1289_ _0096_ _0243_ _0514_ _0563_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_44_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1212_ _0040_ _0123_ _0212_ _0236_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__or4_1
X_1143_ _0181_ _0404_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1074_ _0068_ _0093_ _0104_ _0211_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_23_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0927_ net118 net74 net72 net114 VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__a22o_1
X_0789_ net90 net74 net73 net85 VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__a22o_1
X_0858_ _0705_ _0065_ _0113_ _0149_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__or4_1
Xhold26 net39 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 net31 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_41_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1126_ _0136_ _0140_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__or2_1
X_1057_ net139 net160 net44 _0346_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput38 net38 VGND VGND VPWR VPWR dout0[6] sky130_fd_sc_hd__clkbuf_4
Xoutput27 net27 VGND VGND VPWR VPWR dout0[25] sky130_fd_sc_hd__buf_2
Xoutput16 net16 VGND VGND VPWR VPWR dout0[15] sky130_fd_sc_hd__buf_2
Xclkbuf_2_3__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_3__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_17_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ _0055_ _0253_ _0262_ _0332_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1460_ clknet_2_1__leaf_clk0 net1 VGND VGND VPWR VPWR addr0_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1391_ _0226_ _0473_ _0603_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0960_ _0117_ _0249_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0891_ _0177_ _0180_ _0182_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__or3_1
X_1374_ _0560_ _0605_ _0636_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__or3_1
X_1443_ clknet_2_2__leaf_clk0 _0015_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout73 _0039_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_1
Xfanout62 net65 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
Xfanout51 _0067_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_2
XFILLER_0_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout84 net86 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_2
Xfanout95 _0700_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1090_ _0051_ _0065_ _0135_ _0271_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__or4_1
X_0874_ net60 net50 _0702_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__o21ba_4
X_0943_ _0032_ _0033_ _0036_ _0232_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1426_ net136 net172 VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__or2_1
X_1288_ _0058_ _0129_ _0167_ _0202_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__or4_1
X_1357_ _0114_ _0122_ _0167_ _0197_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1142_ _0052_ _0054_ _0162_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__or3_1
X_1211_ _0469_ _0470_ _0487_ _0491_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__or4_1
X_1073_ _0055_ _0079_ _0328_ _0356_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0857_ _0114_ _0121_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__or2_2
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0926_ _0043_ _0044_ _0107_ _0217_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__or4_1
Xhold16 net14 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dlygate4sd3_1
X_0788_ net96 net75 net73 net102 VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__a22o_2
Xhold27 net18 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ _0201_ _0231_ _0273_ _0296_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_41_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1125_ _0232_ _0240_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__or2_1
X_1056_ _0331_ _0343_ _0345_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__or3_1
Xoutput39 net39 VGND VGND VPWR VPWR dout0[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0909_ _0114_ _0121_ _0196_ _0197_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__or4_4
Xoutput28 net28 VGND VGND VPWR VPWR dout0[26] sky130_fd_sc_hd__buf_2
Xoutput17 net17 VGND VGND VPWR VPWR dout0[16] sky130_fd_sc_hd__buf_2
XFILLER_0_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1108_ _0241_ _0386_ _0388_ _0391_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__or4_1
X_1039_ _0102_ _0103_ _0156_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1390_ _0166_ _0489_ _0592_ _0656_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_13_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0890_ _0120_ _0181_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_10_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1442_ clknet_2_2__leaf_clk0 _0014_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfxtp_1
X_1373_ _0162_ _0203_ _0305_ _0640_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout96 _0700_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_2
Xfanout85 net87 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout74 _0038_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout63 net64 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_1
Xfanout52 _0067_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_0_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0942_ _0032_ _0036_ _0232_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__or3_2
X_0873_ _0122_ _0164_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1425_ net136 net153 net42 _0691_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1356_ net139 net169 net44 _0625_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__o22a_1
X_1287_ _0275_ _0277_ _0559_ _0560_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1072_ _0347_ _0348_ _0355_ _0357_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__or4_1
X_1141_ _0221_ _0222_ _0244_ _0245_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1210_ net135 _0118_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__or2_1
X_0787_ _0075_ _0078_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__or2_2
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0856_ _0693_ _0696_ _0144_ _0147_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0925_ net93 net91 _0046_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold28 net22 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 net37 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ net136 net161 net42 _0675_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__o22a_1
X_1339_ _0200_ _0385_ _0404_ _0412_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_41_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1055_ _0325_ _0334_ _0338_ _0344_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__or4_1
X_1124_ _0406_ _0407_ _0408_ _0409_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0908_ _0196_ _0197_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__or2_1
X_0839_ net109 net105 net97 net107 VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__a22o_2
Xoutput18 net18 VGND VGND VPWR VPWR dout0[17] sky130_fd_sc_hd__buf_2
Xoutput29 net29 VGND VGND VPWR VPWR dout0[27] sky130_fd_sc_hd__buf_2
XFILLER_0_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap71 _0041_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1038_ _0089_ _0133_ _0141_ _0160_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__or4_1
X_1107_ _0208_ _0222_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1441_ clknet_2_1__leaf_clk0 _0013_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1372_ _0693_ _0052_ _0063_ _0104_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout75 _0038_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout42 net45 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
Xfanout97 net100 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_24_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout53 _0066_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_47_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0941_ _0032_ _0232_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0872_ net89 net62 net60 net84 VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__a22o_2
X_1355_ _0331_ _0619_ _0621_ _0624_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__or4_1
X_1424_ _0184_ _0207_ _0690_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__or3_1
X_1286_ _0647_ _0044_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1140_ _0252_ _0267_ _0424_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__or3_1
X_1071_ _0126_ _0286_ _0291_ _0358_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0924_ _0211_ _0213_ _0215_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__or3_2
XFILLER_0_11_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0855_ _0068_ _0069_ _0118_ _0119_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__or4_1
X_0786_ _0072_ _0076_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__or2_2
Xhold29 net24 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 net20 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1338_ _0097_ _0156_ _0416_ _0603_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__or4_1
X_1407_ _0668_ _0671_ _0672_ _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_41_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1269_ _0337_ _0542_ _0543_ _0545_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__or4_1
XFILLER_0_21_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_27_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1123_ _0696_ _0052_ _0054_ _0281_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__or4_1
X_1054_ _0326_ _0335_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_11_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0907_ _0197_ _0198_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput19 net19 VGND VGND VPWR VPWR dout0[18] sky130_fd_sc_hd__buf_2
X_0838_ net105 net68 net66 net97 VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__a22o_2
X_0769_ net126 net119 net122 net124 VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1106_ _0198_ _0233_ _0296_ _0298_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__or4_1
X_1037_ _0133_ _0141_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1440_ clknet_2_3__leaf_clk0 _0012_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1371_ _0215_ _0308_ _0637_ _0638_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout98 net99 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout76 _0035_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_2
Xfanout43 net44 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
Xfanout54 _0066_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_47_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0940_ net83 net69 net67 net81 VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0871_ _0056_ _0162_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__or2_1
X_1354_ _0175_ _0367_ _0622_ _0623_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__or4_1
X_1285_ _0098_ _0174_ _0473_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__or3_1
X_1423_ _0108_ _0247_ _0269_ _0299_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_41_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1070_ _0311_ _0351_ _0354_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0854_ _0037_ _0084_ _0101_ _0145_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__or4_1
X_0923_ _0112_ _0214_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__or2_2
X_0785_ _0075_ _0076_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1337_ _0514_ _0607_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__or2_1
X_1268_ _0431_ _0474_ _0475_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__or4_1
Xhold19 net25 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dlygate4sd3_1
X_1406_ _0226_ _0296_ _0308_ _0673_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__or4_1
X_1199_ _0476_ _0477_ _0480_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1122_ _0116_ _0251_ _0295_ _0299_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__or4_1
X_1053_ _0337_ _0340_ _0341_ _0342_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__or4_1
X_0906_ _0121_ _0196_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__or2_2
X_0837_ net117 net105 net97 net113 VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0768_ _0057_ _0058_ _0059_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_44_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1105_ _0284_ _0290_ _0292_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__or3_2
X_1036_ _0105_ _0179_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_16_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1019_ _0109_ _0274_ _0276_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1370_ _0033_ _0036_ _0044_ _0222_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout44 net45 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
Xfanout55 net57 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout66 _0042_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_2
Xfanout77 _0035_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0870_ _0088_ _0089_ _0090_ _0160_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__or4_2
XFILLER_0_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1422_ _0173_ net42 _0689_ net155 net136 VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__o32a_1
X_1284_ _0075_ _0081_ _0082_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__or3_1
X_1353_ _0081_ _0160_ _0196_ _0292_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0999_ _0105_ _0290_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0922_ net94 net89 net84 net91 VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__a22o_2
X_0853_ _0045_ _0060_ _0092_ _0106_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__or4_1
X_0784_ net89 net50 net48 net84 VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__a22o_2
X_1405_ _0127_ _0188_ _0213_ _0275_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__or4_1
Xinput1 addr0[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_1267_ _0114_ _0130_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__or2_1
X_1336_ _0573_ _0602_ _0604_ _0605_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__or4_1
X_1198_ _0299_ _0478_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1052_ _0078_ _0176_ _0190_ _0227_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__or4_1
X_1121_ _0274_ _0278_ _0286_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0905_ net102 net97 net96 net105 VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__a22o_2
X_0836_ _0124_ _0127_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__or2_1
X_0767_ net107 net62 net60 net109 VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1319_ net139 net158 net44 _0591_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1104_ _0236_ _0390_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__or2_1
X_1035_ _0068_ _0253_ _0268_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_16_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0819_ net125 net123 net120 VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_39_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1018_ _0217_ _0244_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout67 _0042_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
Xfanout56 net57 VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout45 _0304_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
Xfanout89 _0708_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout78 _0034_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_2
XFILLER_0_44_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1421_ _0072_ _0201_ _0216_ _0688_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__or4_1
X_1352_ _0107_ _0141_ _0142_ _0217_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__or4_1
X_1283_ net138 net164 net43 _0558_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_21_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0998_ net115 net53 net51 net111 VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0921_ _0110_ _0212_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__or2_2
X_0852_ _0138_ _0143_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__or2_1
X_0783_ net46 _0074_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__or2_2
XFILLER_0_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1335_ _0710_ _0080_ _0123_ _0187_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__or4_1
X_1404_ _0177_ _0386_ _0604_ _0626_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput2 addr0[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_1266_ _0113_ _0205_ _0290_ _0297_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__or4_1
X_1197_ _0051_ _0170_ _0194_ _0210_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1051_ _0261_ _0278_ _0288_ _0293_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__or4_1
X_1120_ _0209_ _0210_ _0405_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0904_ net97 net69 net67 net106 VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0835_ _0123_ _0125_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__or2_2
X_0766_ net76 net62 net60 net78 VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__a22o_2
XFILLER_0_11_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1318_ _0586_ _0587_ _0590_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1249_ _0040_ _0094_ _0272_ _0389_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap64 net65 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1103_ _0043_ _0044_ _0219_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_74 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1034_ net136 net148 net42 _0324_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_16_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0749_ net134 net132 net128 net130 VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__nor4b_1
X_0818_ net91 net53 net51 net94 VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1017_ net135 _0043_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout79 _0034_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_2
Xfanout68 net70 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_2
XFILLER_0_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1351_ _0408_ _0617_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__or3_1
X_1420_ _0183_ _0684_ _0685_ _0686_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1282_ _0549_ _0551_ _0552_ _0557_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0997_ _0085_ _0284_ _0288_ _0287_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__or4b_1
XFILLER_0_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0920_ net95 net93 net92 net101 VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__a22o_1
X_0851_ _0139_ _0140_ _0141_ _0142_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__or4_1
X_0782_ net95 net49 net47 net101 VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__a22o_2
X_1265_ _0295_ _0327_ _0411_ _0412_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__or4_1
X_1334_ _0087_ _0109_ _0277_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__or3_1
X_1403_ _0172_ _0243_ _0670_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 addr0[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_1196_ _0696_ _0074_ _0181_ _0201_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1050_ _0194_ _0205_ _0328_ _0339_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__or4_1
X_0834_ _0124_ _0125_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__or2_1
X_0903_ _0129_ _0191_ _0193_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__or3_1
X_0765_ net113 net62 net60 net117 VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__a22o_2
XFILLER_0_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1317_ _0083_ _0351_ _0588_ _0589_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1248_ _0240_ _0245_ _0501_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1179_ _0033_ _0098_ _0157_ _0167_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__or4_1
Xmax_cap87 net88 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_6_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1102_ _0044_ _0219_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1033_ _0306_ _0315_ _0316_ _0323_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__or4_1
X_0817_ net111 net109 net107 net116 VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0748_ net110 net74 net72 net108 VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_39_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1016_ _0097_ _0099_ _0198_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_4_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout69 net71 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout47 net48 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
Xfanout58 _0061_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_35_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1350_ _0072_ _0074_ _0365_ _0561_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__or4_1
X_1281_ _0370_ _0553_ _0554_ _0556_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__or4_1
X_0996_ _0086_ _0285_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_21_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0850_ net114 net82 net80 net118 VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__a22o_1
X_0781_ net126 net119 _0702_ net124 VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1402_ _0711_ _0208_ _0248_ _0669_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__or4_1
Xinput4 addr0[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1333_ _0065_ _0258_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__or2_1
X_1264_ _0373_ _0405_ _0430_ _0540_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1195_ _0045_ _0128_ _0260_ _0373_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0979_ _0095_ _0270_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_40_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0833_ net108 net75 net72 net110 VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__a22o_1
X_0902_ _0129_ _0192_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__or2_2
XFILLER_0_44_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0764_ _0049_ _0050_ _0052_ _0053_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__or4_2
X_1316_ _0043_ _0044_ _0209_ _0327_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1247_ _0701_ _0202_ _0203_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_22_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1178_ _0705_ _0203_ _0458_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__or3_1
XANTENNA_20 _0283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap99 net100 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1101_ _0109_ _0276_ _0288_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__or3_2
XFILLER_0_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1032_ _0317_ _0319_ _0321_ _0322_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0816_ _0647_ _0107_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__or2_1
X_0747_ net125 net121 net120 net123 VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_39_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1015_ _0193_ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout48 _0071_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_2
Xfanout59 _0061_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_1
XFILLER_0_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1280_ _0069_ _0074_ _0093_ _0555_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_46_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0995_ net125 net123 net121 _0702_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_21_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0780_ net51 net50 net48 net53 VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1401_ _0085_ _0157_ _0263_ _0270_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput5 addr0[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_1332_ _0095_ _0264_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__or2_1
X_1194_ _0246_ _0457_ _0471_ _0472_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__or4_1
X_1263_ _0158_ _0286_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0978_ net55 net53 net51 net58 VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_40_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0832_ net74 net72 _0046_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__o21ba_1
X_0901_ _0130_ _0131_ _0192_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__or3_2
X_0763_ _0049_ _0050_ _0053_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1315_ _0299_ _0387_ _0424_ _0513_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1246_ net44 _0519_ _0524_ net156 net139 VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__o32a_1
X_1177_ net135 _0133_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_21 _0288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_10 _0156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1100_ _0068_ _0072_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1031_ _0135_ _0232_ _0284_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__or3_1
XFILLER_0_33_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0746_ net123 net120 net121 net125 VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__and4b_1
X_0815_ net110 net94 net92 net108 VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__a22o_2
X_1229_ _0504_ _0506_ _0508_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__or3_1
Xclkbuf_2_2__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_2__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1014_ _0704_ _0202_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__or2_2
XFILLER_0_8_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0729_ net123 net121 net119 net125 VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_4_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout49 net50 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_2
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0994_ _0085_ _0285_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__or2_2
XFILLER_0_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1331_ _0647_ _0251_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__or2_1
X_1400_ _0077_ _0163_ _0370_ _0392_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput6 addr0[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_1193_ _0058_ _0122_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__or2_1
X_1262_ _0527_ _0535_ _0538_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0977_ _0262_ _0265_ _0268_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ net105 net78 net76 net97 VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0831_ net114 net75 net72 net118 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0762_ _0050_ _0053_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__or2_2
XFILLER_0_47_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1314_ _0175_ _0354_ _0430_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__or3_1
X_1245_ _0515_ _0520_ _0523_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1176_ _0086_ _0094_ _0280_ _0282_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__or4_1
XANTENNA_11 _0205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _0292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1030_ _0052_ _0103_ _0170_ _0320_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0814_ _0102_ _0103_ _0104_ _0105_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__or4_1
X_0745_ _0032_ _0033_ _0036_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__or3_2
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1228_ _0336_ _0470_ _0501_ _0507_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1159_ _0117_ _0137_ _0217_ _0221_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_13_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1013_ _0154_ _0155_ net45 net137 net144 VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__o32a_1
X_0728_ net133 net131 net129 net127 VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__or4_4
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0993_ net112 net101 net95 net116 VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__a22o_2
XFILLER_0_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1330_ net138 net168 net43 _0601_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__o22a_1
X_1261_ _0189_ _0228_ _0536_ _0537_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__or4_1
X_1192_ _0107_ _0250_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__or2_1
Xinput7 addr0[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0976_ _0263_ _0266_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__or2_2
X_1459_ clknet_2_2__leaf_clk0 _0031_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dfxtp_1
X_0830_ net95 net62 net60 net101 VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0761_ net78 net63 net61 net76 VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__a22o_1
X_1244_ _0188_ _0231_ _0521_ _0522_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__or4_1
X_1313_ _0056_ _0243_ _0583_ _0585_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_19_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1175_ _0107_ _0217_ _0222_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_12 _0205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0959_ _0117_ _0250_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__or2_1
XANTENNA_23 _0292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0813_ net115 net68 net66 net111 VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__a22o_2
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0744_ net83 net79 net77 net81 VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__a22o_1
X_1158_ net138 net166 net43 _0442_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__o22a_1
X_1227_ _0116_ _0161_ _0300_ _0349_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__or4_1
X_1089_ _0126_ _0288_ _0366_ _0376_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_38_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1012_ _0184_ _0207_ _0257_ _0303_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__nor4_1
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0727_ net105 net101 net97 net95 VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0992_ _0693_ _0104_ _0280_ _0282_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 addr0[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
X_1260_ _0248_ _0249_ _0274_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__or3_1
X_1191_ _0185_ _0187_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__or2_1
X_0975_ _0068_ _0264_ _0266_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_40_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1458_ clknet_2_2__leaf_clk0 _0030_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dfxtp_1
X_1389_ _0098_ _0176_ _0296_ _0297_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0760_ net109 net62 net60 net107 VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__a22o_2
X_1243_ _0086_ _0109_ _0292_ _0295_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__or4_1
X_1312_ _0085_ _0089_ _0229_ _0584_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__or4_1
X_1174_ _0089_ _0161_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__or2_1
XANTENNA_13 _0205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_24 _0421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0889_ net53 net50 net48 net51 VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__a22o_2
X_0958_ net81 net53 net51 net83 VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__a22o_2
XFILLER_0_10_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0743_ net131 net129 net127 net133 VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0812_ net115 net101 net95 net111 VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__a22o_2
X_1157_ _0435_ _0436_ _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__or3_1
XFILLER_0_35_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1226_ _0138_ _0241_ _0254_ _0505_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__or4_1
X_1088_ _0043_ _0245_ _0369_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_43_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1011_ _0269_ _0279_ _0289_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__or4_1
X_0726_ net134 net132 net130 net128 VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__and4b_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1209_ _0072_ _0075_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0991_ _0104_ _0282_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__or2_2
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 cs0 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
X_1190_ _0113_ _0164_ _0166_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__or3_1
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0974_ net68 net59 net56 net66 VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__a22o_1
X_1457_ clknet_2_2__leaf_clk0 _0029_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dfxtp_1
X_1388_ net43 _0650_ _0655_ net171 net139 VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__o32a_1
XFILLER_0_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1311_ _0114_ _0197_ _0232_ _0245_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__or4_1
X_1242_ _0214_ _0223_ _0244_ _0513_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1173_ net42 _0448_ _0456_ net147 net136 VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__o32a_1
XANTENNA_25 _0466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_14 _0215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0957_ net80 net69 net67 net82 VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__a22o_1
X_0888_ _0178_ _0179_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0742_ net127 net129 net131 net133 VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__and4b_1
X_0811_ net113 net49 net47 net117 VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__a22o_2
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1156_ _0199_ _0437_ _0438_ _0440_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__or4_2
X_1225_ _0099_ _0127_ _0157_ _0179_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__or4_1
X_1087_ _0098_ _0176_ _0234_ _0367_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1010_ _0294_ _0301_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__or2_1
X_0725_ net126 net124 net122 net120 VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1208_ _0136_ _0250_ _0252_ _0488_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__or4_2
XFILLER_0_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1139_ _0164_ _0167_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1 net13 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_1_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0990_ net111 net89 net84 net115 VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0973_ _0068_ _0264_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__or2_2
X_1387_ _0649_ _0651_ _0653_ _0654_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__or4_1
X_1456_ clknet_2_2__leaf_clk0 _0028_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1241_ _0079_ _0253_ _0348_ _0413_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__or4_1
X_1310_ _0106_ _0273_ _0310_ _0332_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1172_ _0445_ _0450_ _0453_ _0455_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0956_ net90 net83 net81 net85 VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__a22o_2
XANTENNA_15 _0216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_26 _0496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0887_ net84 net49 net47 net89 VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1439_ clknet_2_0__leaf_clk0 _0011_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfxtp_1
X_0810_ net107 net49 net47 net109 VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__a22o_2
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0741_ net118 net83 net81 net114 VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1224_ _0390_ _0458_ _0490_ _0503_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__or4_1
X_1155_ _0127_ _0389_ _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__or3_1
X_1086_ net135 net46 _0105_ _0274_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__or4_1
X_0939_ _0123_ _0124_ _0125_ _0229_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__or4_4
XFILLER_0_15_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire70 _0041_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0724_ net133 net130 net128 net132 VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_12_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1207_ _0057_ _0058_ _0164_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1138_ net44 _0410_ _0423_ net165 net138 VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__o32a_1
XFILLER_0_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1069_ _0097_ _0236_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2 net11 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0972_ net101 net58 net56 net95 VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__a22o_2
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1386_ _0164_ _0166_ _0356_ _0550_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__or4_1
X_1455_ clknet_2_2__leaf_clk0 _0027_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1240_ _0512_ _0516_ _0517_ _0518_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__or4_1
X_1171_ _0084_ _0193_ _0290_ _0454_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_27 _0654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_16 _0261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0886_ net101 net50 net48 net95 VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__a22o_2
X_0955_ _0707_ _0710_ _0244_ _0245_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__or4_2
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1369_ _0131_ _0192_ _0335_ _0415_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1438_ clknet_2_2__leaf_clk0 _0010_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0740_ net110 net83 net81 net108 VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1223_ _0094_ _0270_ _0502_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__or3_1
X_1154_ _0130_ _0156_ _0157_ _0214_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__or4_1
X_1085_ _0264_ _0268_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__or2_1
X_0938_ _0124_ _0229_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__or2_1
X_0869_ _0088_ _0160_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0723_ net126 net124 net120 net122 VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_12_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1137_ _0417_ _0420_ _0421_ _0422_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__or4_1
X_1206_ _0135_ _0141_ _0430_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1068_ _0107_ _0217_ _0221_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_35_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_31_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3 net15 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0971_ net84 net59 net56 net89 VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__a22o_1
X_1454_ clknet_2_2__leaf_clk0 _0026_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1385_ _0704_ _0171_ _0203_ _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1170_ _0275_ _0285_ _0405_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_28 _0441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 _0267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0885_ _0097_ _0098_ _0099_ _0174_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__or4_1
X_0954_ _0711_ _0245_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__or2_1
X_1437_ clknet_2_1__leaf_clk0 _0009_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1299_ _0113_ _0214_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__or2_1
X_1368_ _0119_ _0180_ _0210_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__or3_1
XFILLER_0_33_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1153_ _0696_ _0086_ _0104_ _0191_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__or4_1
X_1222_ _0104_ _0290_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__or2_1
X_1084_ _0263_ _0264_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__or2_1
X_0799_ _0089_ _0090_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0868_ net68 net63 net61 net66 VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__a22o_1
X_0937_ net76 net74 net72 net78 VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_7_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0722_ net115 net109 net107 net111 VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_12_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1136_ _0108_ _0220_ _0283_ _0372_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__or4_1
X_1067_ _0103_ _0156_ _0212_ _0214_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1205_ net45 _0481_ _0486_ net142 net136 VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_35_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold4 net10 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1119_ _0120_ _0178_ _0179_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0970_ _0063_ _0064_ _0258_ _0259_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__or4_4
X_1453_ clknet_2_3__leaf_clk0 _0025_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1384_ _0068_ _0069_ _0283_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_18 _0274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0884_ _0097_ _0174_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0953_ net93 net69 net67 net91 VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__a22o_2
X_1367_ net42 _0628_ _0635_ net159 net136 VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__o32a_1
XFILLER_0_10_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1436_ clknet_2_2__leaf_clk0 _0008_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dfxtp_1
X_1298_ _0137_ _0140_ _0142_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_18_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1221_ _0707_ _0237_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__or2_1
X_1083_ _0131_ _0192_ _0349_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__or3_1
X_1152_ _0060_ _0203_ _0305_ _0430_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__or4_1
X_0936_ _0080_ _0081_ _0082_ _0225_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__or4_2
X_0867_ _0102_ _0103_ _0156_ _0157_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0798_ net85 net62 net61 net90 VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__a22o_1
X_1419_ net135 _0696_ _0159_ _0370_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0721_ net129 net127 net133 net131 VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_12_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1204_ _0469_ _0482_ _0484_ _0485_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1135_ _0411_ _0414_ _0415_ _0416_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__or4_1
X_1066_ _0032_ _0164_ _0166_ _0240_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0919_ _0118_ _0119_ _0208_ _0210_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_26_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 net19 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1049_ _0115_ _0124_ _0137_ _0274_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__or4_1
X_1118_ _0120_ _0178_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1383_ _0190_ _0198_ _0388_ _0648_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__or4_1
X_1452_ clknet_2_3__leaf_clk0 _0024_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_19 _0283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0952_ net93 net54 net52 net91 VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__a22o_2
XFILLER_0_27_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0883_ _0100_ _0174_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__or2_1
X_1435_ clknet_2_3__leaf_clk0 _0007_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfxtp_1
X_1366_ _0627_ _0631_ _0634_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__or3_1
X_1297_ net136 net167 net42 _0571_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_18_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1151_ _0077_ _0426_ _0428_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__or3_1
X_1220_ net43 _0496_ _0500_ net152 net138 VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__o32a_1
X_1082_ _0217_ _0221_ _0222_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__or3_2
X_0935_ _0080_ _0225_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__or2_1
X_0866_ _0103_ _0157_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0797_ net101 net63 net61 net95 VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1349_ _0278_ _0286_ _0472_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1418_ _0083_ _0194_ _0283_ _0291_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0720_ net131 net127 net129 net133 VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_12_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1134_ _0128_ _0347_ _0418_ _0419_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__or4_1
X_1203_ _0272_ _0365_ _0460_ _0473_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_35_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1065_ _0204_ _0352_ _0353_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__or3_1
X_0849_ net82 net54 net52 net80 VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__a22o_2
X_0918_ net107 net93 net91 net109 VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__a22o_2
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_1__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
Xhold6 net30 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap103 net104 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1117_ net138 net157 net43 _0403_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_0_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1048_ _0220_ _0242_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1382_ _0391_ _0427_ _0512_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__or3_1
X_1451_ clknet_2_2__leaf_clk0 _0023_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0882_ net117 net49 net47 net113 VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__a22o_2
X_0951_ _0236_ _0237_ _0239_ _0240_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__or4_2
X_1434_ clknet_2_3__leaf_clk0 _0006_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dfxtp_1
X_1296_ _0562_ _0564_ _0567_ _0570_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__or4_1
X_1365_ _0092_ _0313_ _0633_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_18_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1150_ _0425_ _0427_ _0433_ _0434_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__or4_1
X_1081_ _0088_ _0103_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__or2_1
X_0934_ _0082_ _0225_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__or2_1
X_0865_ net76 net49 net47 net78 VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__a22o_2
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1417_ _0191_ _0273_ _0296_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__or3_1
X_0796_ net63 net54 net52 net61 VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__a22o_1
X_1348_ _0091_ _0333_ _0372_ _0432_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__or4_1
X_1279_ _0130_ _0140_ _0166_ _0203_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__or4_1
Xwire86 net88 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1133_ _0057_ _0076_ _0097_ _0164_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__or4_1
X_1064_ _0117_ _0131_ _0137_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__or3_1
X_1202_ _0204_ _0312_ _0483_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_25_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0848_ net82 net80 _0046_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__o21ba_1
X_0917_ _0118_ _0208_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__or2_2
X_0779_ net125 net119 net121 net123 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_11_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold7 net40 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1047_ _0166_ _0221_ _0336_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__or3_1
X_1116_ _0395_ _0400_ _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_0_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk0 clk0 VGND VGND VPWR VPWR clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1450_ clknet_2_3__leaf_clk0 _0022_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1381_ _0549_ _0559_ _0572_ _0602_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0881_ _0056_ _0162_ _0169_ _0172_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__or4_1
X_0950_ _0236_ _0237_ _0240_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__or3_1
X_1433_ clknet_2_3__leaf_clk0 _0005_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dfxtp_1
X_1364_ _0063_ _0258_ _0292_ _0632_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__or4_1
X_1295_ _0301_ _0540_ _0568_ _0569_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_18_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1080_ _0080_ _0226_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__or2_1
X_0933_ net73 net69 net67 net74 VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0864_ net66 net49 net47 net68 VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__a22o_2
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0795_ _0085_ _0086_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1347_ _0129_ _0193_ _0525_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__or3_1
X_1416_ _0173_ net42 _0683_ net146 net136 VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__o32a_1
Xwire65 _0047_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
X_1278_ _0369_ _0429_ _0491_ _0550_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__or4_1
Xfanout130 addr0_reg\[2\] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1201_ _0032_ _0036_ _0104_ _0105_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1063_ net135 _0186_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__or2_1
X_1132_ _0112_ _0185_ _0203_ _0237_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0916_ net91 net68 net66 net93 VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__a22o_2
X_0847_ _0702_ net82 VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__and2b_1
X_0778_ net123 net119 net121 net125 VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold8 net21 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1046_ net135 _0057_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__or2_1
X_1115_ _0392_ _0393_ _0401_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_0_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1029_ _0125_ _0137_ _0187_ _0212_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1380_ _0119_ _0209_ _0426_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0880_ _0057_ _0058_ _0059_ _0170_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1432_ clknet_2_3__leaf_clk0 _0004_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dfxtp_1
X_1363_ _0058_ _0174_ _0214_ _0298_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1294_ _0696_ _0156_ _0280_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_18_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0932_ _0040_ _0219_ _0221_ _0222_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__or4_1
X_0794_ net116 net89 net84 net112 VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__a22o_1
X_0863_ _0132_ _0146_ _0148_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__or3_1
X_1346_ net43 _0608_ _0616_ net170 net138 VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__o32a_1
X_1415_ _0636_ _0678_ _0680_ _0682_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__or4_1
Xwire88 _0709_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_1
X_1277_ _0135_ _0172_ _0232_ _0247_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__or4_1
Xfanout131 addr0_reg\[1\] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout120 addr0_reg\[7\] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_29_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1200_ _0109_ _0277_ _0474_ _0475_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__or4_1
X_1131_ _0135_ _0141_ _0368_ _0413_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1062_ _0057_ _0171_ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0915_ _0195_ _0201_ _0206_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__or3_1
X_0846_ _0133_ _0134_ _0136_ _0137_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__or4_1
X_0777_ net107 net58 net55 net109 VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__a22o_2
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1329_ _0593_ _0595_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_34_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold9 net26 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1114_ _0100_ _0168_ _0387_ _0394_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1045_ _0049_ _0059_ _0069_ _0298_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_23_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0829_ net98 net54 net52 net106 VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1028_ _0051_ _0161_ _0318_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1431_ clknet_2_1__leaf_clk0 _0003_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1293_ _0049_ _0118_ _0120_ _0212_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__or4_1
X_1362_ _0051_ _0265_ _0629_ _0630_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0931_ _0221_ _0222_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__or2_1
X_0862_ _0079_ _0096_ _0152_ _0153_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_15_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0793_ net111 net53 net51 net115 VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__a22o_1
X_1345_ _0611_ _0612_ _0615_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__or3_1
X_1276_ _0391_ _0409_ _0449_ _0548_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1414_ _0265_ _0268_ _0679_ _0681_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__or4_1
Xfanout110 _0694_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
Xfanout132 addr0_reg\[1\] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout121 addr0_reg\[6\] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_29_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1130_ _0093_ _0170_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1061_ _0693_ _0280_ _0292_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__or3_1
X_0845_ net80 net79 net77 net82 VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__a22o_2
X_0914_ _0705_ _0204_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__or2_1
X_0776_ net59 net53 net51 net55 VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__a22o_2
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1328_ _0594_ _0596_ _0598_ _0599_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__or4_1
X_1259_ _0033_ _0052_ _0053_ _0089_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_34_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_29_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1044_ _0121_ _0197_ _0332_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__or4_1
X_1113_ _0352_ _0396_ _0397_ _0399_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0828_ net68 net50 net48 net66 VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__a22o_1
X_0759_ _0049_ _0050_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__or2_2
XFILLER_0_19_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1027_ _0036_ _0040_ _0080_ _0112_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1430_ clknet_2_1__leaf_clk0 _0002_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1292_ _0325_ _0516_ _0565_ _0566_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__or4_1
X_1361_ _0040_ _0121_ _0124_ _0245_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0861_ _0056_ _0109_ _0120_ _0122_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_15_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0792_ _0082_ _0083_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__or2_1
X_0930_ net93 net79 net77 net91 VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__a22o_2
XFILLER_0_2_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1413_ _0182_ _0226_ _0278_ _0491_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1344_ _0078_ _0606_ _0613_ _0614_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__or4_1
X_1275_ _0267_ _0275_ _0285_ _0471_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__or4_1
Xwire46 _0073_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_1
Xwire57 _0062_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout133 addr0_reg\[0\] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout122 addr0_reg\[6\] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_1
Xfanout111 _0687_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1060_ _0693_ _0292_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0844_ net108 net82 net80 net110 VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__a22o_1
X_0913_ _0701_ _0202_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__or2_2
X_0775_ net131 net129 net127 net133 VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_3_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1258_ _0281_ _0293_ _0385_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__or3_1
X_1327_ _0141_ _0203_ _0238_ _0262_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__or4_1
X_1189_ _0082_ _0470_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1043_ _0707_ _0244_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__or2_1
X_1112_ _0711_ _0057_ _0058_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0827_ net114 net93 net92 net118 VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__a22o_2
X_0758_ net117 net63 net61 net113 VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_46_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1026_ _0078_ _0165_ _0265_ _0271_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1009_ _0069_ _0295_ _0297_ _0298_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1360_ _0119_ _0208_ _0404_ _0561_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1291_ _0502_ _0544_ _0561_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0791_ _0080_ _0081_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__or2_1
X_0860_ _0711_ _0087_ _0150_ _0151_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_15_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1412_ _0040_ _0350_ _0389_ _0525_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__or4_1
X_1343_ _0157_ _0266_ _0297_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__or3_1
X_1274_ _0125_ _0229_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0989_ _0693_ _0280_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__or2_1
Xfanout134 addr0_reg\[0\] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_1
Xfanout112 _0687_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_1
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout123 addr0_reg\[5\] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
Xfanout101 net103 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_29_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0912_ _0202_ _0203_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__or2_1
X_0843_ _0133_ _0134_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__or2_2
X_0774_ net129 net127 net133 net131 VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1326_ _0054_ _0178_ _0181_ _0597_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_3_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1188_ _0081_ _0225_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__or2_1
X_1257_ net45 _0530_ _0534_ net143 net137 VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__o32a_1
XFILLER_0_46_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1111_ _0088_ _0123_ _0136_ _0270_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__or4_1
X_1042_ _0112_ _0212_ _0214_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__or3_2
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0757_ net62 net60 _0046_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_10_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0826_ net92 net79 net77 net93 VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1309_ net43 _0580_ _0582_ net145 net138 VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_22_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1025_ _0260_ _0307_ _0313_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__or3_1
X_0809_ _0097_ _0098_ _0099_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1 _0051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1008_ _0295_ _0298_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1290_ _0126_ _0309_ _0312_ _0429_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0790_ net72 net54 net52 net74 VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__a22o_2
X_1342_ _0194_ _0205_ _0357_ _0488_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__or4_1
X_1273_ _0100_ _0178_ _0181_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__or3_1
X_1411_ _0115_ _0130_ _0131_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0988_ net115 net78 net76 net111 VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout102 net104 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout113 _0677_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_2
Xfanout135 _0647_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_2
Xfanout124 addr0_reg\[5\] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0842_ net102 net82 net80 net96 VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__a22o_1
X_0911_ net105 net53 net51 net97 VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__a22o_4
X_0773_ _0063_ _0064_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__or2_2
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1325_ _0647_ _0082_ _0098_ _0156_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_3_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1256_ _0471_ _0525_ _0526_ _0533_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_34_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1187_ _0157_ _0174_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1110_ _0083_ _0102_ _0135_ _0156_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1041_ _0037_ _0182_ _0330_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0825_ net96 net82 net80 net102 VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_31_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0756_ net119 net121 net126 net124 VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1239_ _0178_ _0181_ _0336_ _0502_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1308_ _0195_ _0393_ _0501_ _0581_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1024_ _0308_ _0309_ _0311_ _0314_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__or4_1
X_0808_ _0098_ _0099_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__or2_1
X_0739_ net121 net120 net123 net125 VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__and4b_1
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_2 _0057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1007_ _0297_ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1410_ _0077_ _0370_ _0676_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__or3_1
X_1272_ _0215_ _0248_ _0251_ _0283_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__or4_1
X_1341_ _0244_ _0245_ _0294_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0987_ _0273_ _0275_ _0278_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout114 _0677_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
Xfanout125 addr0_reg\[4\] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
Xfanout136 net137 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__buf_2
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0841_ net85 net82 net80 net90 VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__a22o_1
X_0910_ net97 net89 net84 net105 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__a22o_1
X_0772_ net117 net58 net55 net113 VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1186_ net44 _0464_ _0468_ net154 net139 VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__o32a_1
X_1324_ _0091_ _0171_ _0233_ _0349_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1255_ _0231_ _0528_ _0531_ _0532_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1040_ _0093_ _0094_ _0211_ _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0824_ _0114_ _0115_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0755_ net126 net124 net119 net122 VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__nor4b_1
X_1169_ _0091_ _0449_ _0451_ _0452_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__or4_1
X_1238_ _0168_ _0265_ _0305_ _0358_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__or4_1
X_1307_ _0054_ _0072_ _0074_ _0394_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1023_ _0069_ _0094_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0738_ net125 net123 net120 net121 VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__and4bb_1
X_0807_ net49 net47 _0046_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__o21ba_2
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_3 _0057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1006_ net113 net58 net55 net117 VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__a22o_2
XFILLER_0_32_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput40 net40 VGND VGND VPWR VPWR dout0[8] sky130_fd_sc_hd__buf_2
XFILLER_0_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1340_ _0338_ _0516_ _0609_ _0610_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1271_ net137 net150 net42 _0547_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_14_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0986_ _0276_ _0277_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__or2_2
Xfanout126 addr0_reg\[4\] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
Xfanout137 net9 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
Xfanout115 _0667_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_2
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0771_ net78 net58 net55 net76 VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__a22o_1
X_0840_ _0128_ _0129_ _0130_ _0131_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__or4_1
X_1323_ _0267_ _0390_ _0572_ _0592_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1185_ _0132_ _0334_ _0465_ _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__or4_1
X_1254_ _0051_ _0075_ _0213_ _0268_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0969_ _0258_ _0259_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0754_ net134 net132 net130 net127 VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__or4b_4
X_0823_ net108 net105 net97 net110 VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__a22o_2
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1306_ _0503_ _0572_ _0573_ _0579_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__or4_1
X_1168_ _0168_ _0176_ _0443_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__or3_1
X_1237_ _0037_ _0134_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__or2_1
X_1099_ _0704_ _0130_ _0131_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_45_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1022_ _0248_ _0249_ _0312_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__or3_1
X_0737_ _0707_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__or2_2
X_0806_ net109 net49 net47 net107 VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__a22o_2
XFILLER_0_24_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 _0057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1005_ net76 net59 net56 net78 VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__a22o_2
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput41 net41 VGND VGND VPWR VPWR dout0[9] sky130_fd_sc_hd__clkbuf_4
Xoutput30 net30 VGND VGND VPWR VPWR dout0[28] sky130_fd_sc_hd__buf_2
XFILLER_0_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
.ends

