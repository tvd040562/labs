logic [0:(ROM_DEPTH/8)-1] [DATA_WIDTH-1:0] table1 = {
32'h00000000,
32'h003243f1,
32'h006487c4,
32'h0096cb58,
32'h00c90e90,
32'h00fb514b,
32'h012d936c,
32'h015fd4d2,
32'h0192155f,
32'h01c454f5,
32'h01f69373,
32'h0228d0bb,
32'h025b0caf,
32'h028d472e,
32'h02bf801a,
32'h02f1b755,
32'h0323ecbe,
32'h03562038,
32'h038851a2,
32'h03ba80df,
32'h03ecadcf,
32'h041ed854,
32'h0451004d,
32'h0483259d,
32'h04b54825,
32'h04e767c5,
32'h0519845e,
32'h054b9dd3,
32'h057db403,
32'h05afc6d0,
32'h05e1d61b,
32'h0613e1c5,
32'h0645e9af,
32'h0677edbb,
32'h06a9edc9,
32'h06dbe9bb,
32'h070de172,
32'h073fd4cf,
32'h0771c3b3,
32'h07a3adff,
32'h07d59396,
32'h08077457,
32'h08395024,
32'h086b26de,
32'h089cf867,
32'h08cec4a0,
32'h09008b6a,
32'h09324ca7,
32'h09640837,
32'h0995bdfd,
32'h09c76dd8,
32'h09f917ac,
32'h0a2abb59,
32'h0a5c58c0,
32'h0a8defc3,
32'h0abf8043,
32'h0af10a22,
32'h0b228d42,
32'h0b540982,
32'h0b857ec7,
32'h0bb6ecef,
32'h0be853de,
32'h0c19b374,
32'h0c4b0b94,
32'h0c7c5c1e,
32'h0cada4f5,
32'h0cdee5f9,
32'h0d101f0e,
32'h0d415013,
32'h0d7278eb,
32'h0da39978,
32'h0dd4b19a,
32'h0e05c135,
32'h0e36c82a,
32'h0e67c65a,
32'h0e98bba7,
32'h0ec9a7f3,
32'h0efa8b20,
32'h0f2b650f,
32'h0f5c35a3,
32'h0f8cfcbe,
32'h0fbdba40,
32'h0fee6e0d,
32'h101f1807,
32'h104fb80e,
32'h10804e06,
32'h10b0d9d0,
32'h10e15b4e,
32'h1111d263,
32'h11423ef0,
32'h1172a0d7,
32'h11a2f7fc,
32'h11d3443f,
32'h12038584,
32'h1233bbac,
32'h1263e699,
32'h1294062f,
32'h12c41a4f,
32'h12f422db,
32'h13241fb6,
32'h135410c3,
32'h1383f5e3,
32'h13b3cefa,
32'h13e39be9,
32'h14135c94,
32'h144310dd,
32'h1472b8a5,
32'h14a253d1,
32'h14d1e242,
32'h150163dc,
32'h1530d881,
32'h15604013,
32'h158f9a76,
32'h15bee78c,
32'h15ee2738,
32'h161d595d,
32'h164c7ddd,
32'h167b949d,
32'h16aa9d7e,
32'h16d99864,
32'h17088531,
32'h173763c9,
32'h1766340f,
32'h1794f5e6,
32'h17c3a931,
32'h17f24dd3,
32'h1820e3b0,
32'h184f6aab,
32'h187de2a7,
32'h18ac4b87,
32'h18daa52f,
32'h1908ef82,
32'h19372a64,
32'h196555b8,
32'h19937161,
32'h19c17d44,
32'h19ef7944,
32'h1a1d6544,
32'h1a4b4128,
32'h1a790cd4,
32'h1aa6c82b,
32'h1ad47312,
32'h1b020d6c,
32'h1b2f971e,
32'h1b5d100a,
32'h1b8a7815,
32'h1bb7cf23,
32'h1be51518,
32'h1c1249d8,
32'h1c3f6d47,
32'h1c6c7f4a,
32'h1c997fc4,
32'h1cc66e99,
32'h1cf34baf,
32'h1d2016e9,
32'h1d4cd02c,
32'h1d79775c,
32'h1da60c5d,
32'h1dd28f15,
32'h1dfeff67,
32'h1e2b5d38,
32'h1e57a86d,
32'h1e83e0eb,
32'h1eb00696,
32'h1edc1953,
32'h1f081907,
32'h1f340596,
32'h1f5fdee6,
32'h1f8ba4dc,
32'h1fb7575c,
32'h1fe2f64c,
32'h200e8190,
32'h2039f90f,
32'h20655cac,
32'h2090ac4d,
32'h20bbe7d8,
32'h20e70f32,
32'h21122240,
32'h213d20e8,
32'h21680b0f,
32'h2192e09b,
32'h21bda171,
32'h21e84d76,
32'h2212e492,
32'h223d66a8,
32'h2267d3a0,
32'h22922b5e,
32'h22bc6dca,
32'h22e69ac8,
32'h2310b23e,
32'h233ab414,
32'h2364a02e,
32'h238e7673,
32'h23b836ca,
32'h23e1e117,
32'h240b7543,
32'h2434f332,
32'h245e5acc,
32'h2487abf7,
32'h24b0e699,
32'h24da0a9a,
32'h250317df,
32'h252c0e4f,
32'h2554edd1,
32'h257db64c,
32'h25a667a7,
32'h25cf01c8,
32'h25f78497,
32'h261feffa,
32'h264843d9,
32'h2670801a,
32'h2698a4a6,
32'h26c0b162,
32'h26e8a637,
32'h2710830c,
32'h273847c8,
32'h275ff452,
32'h27878893,
32'h27af0472,
32'h27d667d5,
32'h27fdb2a7,
32'h2824e4cc,
32'h284bfe2f,
32'h2872feb6,
32'h2899e64a,
32'h28c0b4d2,
32'h28e76a37,
32'h290e0661,
32'h29348937,
32'h295af2a3,
32'h2981428c,
32'h29a778db,
32'h29cd9578,
32'h29f3984c,
32'h2a19813f,
32'h2a3f503a,
32'h2a650525,
32'h2a8a9fea,
32'h2ab02071,
32'h2ad586a3,
32'h2afad269,
32'h2b2003ac,
32'h2b451a55,
32'h2b6a164d,
32'h2b8ef77d,
32'h2bb3bdce,
32'h2bd8692b,
32'h2bfcf97c,
32'h2c216eaa,
32'h2c45c8a0,
32'h2c6a0746,
32'h2c8e2a87,
32'h2cb2324c,
32'h2cd61e7f,
32'h2cf9ef09,
32'h2d1da3d5
};
