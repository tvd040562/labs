module cust_rom (clk0,
    cs0,
    addr0,
    dout0);
 input clk0;
 input cs0;
 input [7:0] addr0;
 output [32:0] dout0;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire \addr0_reg[0] ;
 wire \addr0_reg[1] ;
 wire \addr0_reg[2] ;
 wire \addr0_reg[3] ;
 wire \addr0_reg[4] ;
 wire \addr0_reg[5] ;
 wire \addr0_reg[6] ;
 wire \addr0_reg[7] ;
 wire clknet_0_clk0;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire clknet_2_0__leaf_clk0;
 wire clknet_2_1__leaf_clk0;
 wire clknet_2_2__leaf_clk0;
 wire clknet_2_3__leaf_clk0;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;

 sky130_fd_sc_hd__inv_2 _0714_ (.A(net138),
    .Y(_0647_));
 sky130_fd_sc_hd__and4bb_1 _0715_ (.A_N(net133),
    .B_N(net127),
    .C(net129),
    .D(net131),
    .X(_0657_));
 sky130_fd_sc_hd__and4b_1 _0716_ (.A_N(net119),
    .B(net122),
    .C(net126),
    .D(net124),
    .X(_0667_));
 sky130_fd_sc_hd__and4bb_1 _0717_ (.A_N(net133),
    .B_N(net129),
    .C(net127),
    .D(net131),
    .X(_0677_));
 sky130_fd_sc_hd__nor4_1 _0718_ (.A(net126),
    .B(net124),
    .C(net119),
    .D(net122),
    .Y(_0687_));
 sky130_fd_sc_hd__a22o_2 _0719_ (.A1(net117),
    .A2(net115),
    .B1(net113),
    .B2(net111),
    .X(_0693_));
 sky130_fd_sc_hd__and4bb_1 _0720_ (.A_N(net131),
    .B_N(net127),
    .C(net129),
    .D(net133),
    .X(_0694_));
 sky130_fd_sc_hd__and4b_1 _0721_ (.A_N(net129),
    .B(net127),
    .C(net133),
    .D(net131),
    .X(_0695_));
 sky130_fd_sc_hd__a22o_2 _0722_ (.A1(net115),
    .A2(net109),
    .B1(net107),
    .B2(net111),
    .X(_0696_));
 sky130_fd_sc_hd__and4_1 _0723_ (.A(net126),
    .B(net124),
    .C(net120),
    .D(net122),
    .X(_0697_));
 sky130_fd_sc_hd__nor4b_1 _0724_ (.A(net133),
    .B(net130),
    .C(net128),
    .D_N(net132),
    .Y(_0698_));
 sky130_fd_sc_hd__nor4b_1 _0725_ (.A(net126),
    .B(net124),
    .C(net122),
    .D_N(net120),
    .Y(_0699_));
 sky130_fd_sc_hd__and4b_1 _0726_ (.A_N(net134),
    .B(net132),
    .C(net130),
    .D(net128),
    .X(_0700_));
 sky130_fd_sc_hd__a22o_1 _0727_ (.A1(net105),
    .A2(net101),
    .B1(net97),
    .B2(net95),
    .X(_0701_));
 sky130_fd_sc_hd__or4_4 _0728_ (.A(net133),
    .B(net131),
    .C(net129),
    .D(net127),
    .X(_0702_));
 sky130_fd_sc_hd__and4bb_1 _0729_ (.A_N(net123),
    .B_N(net121),
    .C(net119),
    .D(net125),
    .X(_0703_));
 sky130_fd_sc_hd__o21ba_1 _0730_ (.A1(net105),
    .A2(net94),
    .B1_N(_0702_),
    .X(_0704_));
 sky130_fd_sc_hd__or2_2 _0731_ (.A(_0701_),
    .B(_0704_),
    .X(_0705_));
 sky130_fd_sc_hd__and4b_1 _0732_ (.A_N(net125),
    .B(net123),
    .C(net120),
    .D(net121),
    .X(_0706_));
 sky130_fd_sc_hd__a22o_2 _0733_ (.A1(net102),
    .A2(net94),
    .B1(net92),
    .B2(net96),
    .X(_0707_));
 sky130_fd_sc_hd__and4_1 _0734_ (.A(net134),
    .B(net131),
    .C(net129),
    .D(net128),
    .X(_0708_));
 sky130_fd_sc_hd__nor4b_1 _0735_ (.A(net132),
    .B(net130),
    .C(net128),
    .D_N(net134),
    .Y(_0709_));
 sky130_fd_sc_hd__a22o_2 _0736_ (.A1(net91),
    .A2(net89),
    .B1(net84),
    .B2(net94),
    .X(_0710_));
 sky130_fd_sc_hd__or2_2 _0737_ (.A(_0707_),
    .B(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__and4bb_1 _0738_ (.A_N(net125),
    .B_N(net123),
    .C(net120),
    .D(net121),
    .X(_0712_));
 sky130_fd_sc_hd__and4b_1 _0739_ (.A_N(net121),
    .B(net120),
    .C(net123),
    .D(net125),
    .X(_0713_));
 sky130_fd_sc_hd__a22o_1 _0740_ (.A1(net110),
    .A2(net83),
    .B1(net81),
    .B2(net108),
    .X(_0032_));
 sky130_fd_sc_hd__a22o_1 _0741_ (.A1(net118),
    .A2(net83),
    .B1(net81),
    .B2(net114),
    .X(_0033_));
 sky130_fd_sc_hd__and4b_1 _0742_ (.A_N(net127),
    .B(net129),
    .C(net131),
    .D(net133),
    .X(_0034_));
 sky130_fd_sc_hd__and4bb_1 _0743_ (.A_N(net131),
    .B_N(net129),
    .C(net127),
    .D(net133),
    .X(_0035_));
 sky130_fd_sc_hd__a22o_1 _0744_ (.A1(net83),
    .A2(net79),
    .B1(net77),
    .B2(net81),
    .X(_0036_));
 sky130_fd_sc_hd__or3_2 _0745_ (.A(_0032_),
    .B(_0033_),
    .C(_0036_),
    .X(_0037_));
 sky130_fd_sc_hd__and4b_1 _0746_ (.A_N(net123),
    .B(net120),
    .C(net121),
    .D(net125),
    .X(_0038_));
 sky130_fd_sc_hd__and4bb_1 _0747_ (.A_N(net125),
    .B_N(net121),
    .C(net120),
    .D(net123),
    .X(_0039_));
 sky130_fd_sc_hd__a22o_2 _0748_ (.A1(net110),
    .A2(net74),
    .B1(net72),
    .B2(net108),
    .X(_0040_));
 sky130_fd_sc_hd__nor4b_1 _0749_ (.A(net134),
    .B(net132),
    .C(net128),
    .D_N(net130),
    .Y(_0041_));
 sky130_fd_sc_hd__and4bb_1 _0750_ (.A_N(net134),
    .B_N(net132),
    .C(net130),
    .D(net128),
    .X(_0042_));
 sky130_fd_sc_hd__a22o_2 _0751_ (.A1(net75),
    .A2(net69),
    .B1(net67),
    .B2(net73),
    .X(_0043_));
 sky130_fd_sc_hd__a22o_2 _0752_ (.A1(net79),
    .A2(net74),
    .B1(net72),
    .B2(net77),
    .X(_0044_));
 sky130_fd_sc_hd__or3_1 _0753_ (.A(_0040_),
    .B(_0043_),
    .C(_0044_),
    .X(_0045_));
 sky130_fd_sc_hd__or4b_4 _0754_ (.A(net134),
    .B(net132),
    .C(net130),
    .D_N(net127),
    .X(_0046_));
 sky130_fd_sc_hd__nor4b_1 _0755_ (.A(net126),
    .B(net124),
    .C(net119),
    .D_N(net122),
    .Y(_0047_));
 sky130_fd_sc_hd__and4bb_1 _0756_ (.A_N(net119),
    .B_N(net121),
    .C(net126),
    .D(net124),
    .X(_0048_));
 sky130_fd_sc_hd__o21ba_1 _0757_ (.A1(net62),
    .A2(net60),
    .B1_N(_0046_),
    .X(_0049_));
 sky130_fd_sc_hd__a22o_1 _0758_ (.A1(net117),
    .A2(net63),
    .B1(net61),
    .B2(net113),
    .X(_0050_));
 sky130_fd_sc_hd__or2_2 _0759_ (.A(_0049_),
    .B(_0050_),
    .X(_0051_));
 sky130_fd_sc_hd__a22o_2 _0760_ (.A1(net109),
    .A2(net62),
    .B1(net60),
    .B2(net107),
    .X(_0052_));
 sky130_fd_sc_hd__a22o_1 _0761_ (.A1(net78),
    .A2(net63),
    .B1(net61),
    .B2(net76),
    .X(_0053_));
 sky130_fd_sc_hd__or2_2 _0762_ (.A(_0050_),
    .B(_0053_),
    .X(_0054_));
 sky130_fd_sc_hd__or3_1 _0763_ (.A(_0049_),
    .B(_0050_),
    .C(_0053_),
    .X(_0055_));
 sky130_fd_sc_hd__or4_2 _0764_ (.A(_0049_),
    .B(_0050_),
    .C(_0052_),
    .D(_0053_),
    .X(_0056_));
 sky130_fd_sc_hd__a22o_2 _0765_ (.A1(net113),
    .A2(net62),
    .B1(net60),
    .B2(net117),
    .X(_0057_));
 sky130_fd_sc_hd__a22o_2 _0766_ (.A1(net76),
    .A2(net62),
    .B1(net60),
    .B2(net78),
    .X(_0058_));
 sky130_fd_sc_hd__a22o_1 _0767_ (.A1(net107),
    .A2(net62),
    .B1(net60),
    .B2(net109),
    .X(_0059_));
 sky130_fd_sc_hd__or3_2 _0768_ (.A(_0057_),
    .B(_0058_),
    .C(_0059_),
    .X(_0060_));
 sky130_fd_sc_hd__and4bb_1 _0769_ (.A_N(net126),
    .B_N(net119),
    .C(net122),
    .D(net124),
    .X(_0061_));
 sky130_fd_sc_hd__nor4b_1 _0770_ (.A(net124),
    .B(net119),
    .C(net122),
    .D_N(net126),
    .Y(_0062_));
 sky130_fd_sc_hd__a22o_1 _0771_ (.A1(net78),
    .A2(net58),
    .B1(net55),
    .B2(net76),
    .X(_0063_));
 sky130_fd_sc_hd__a22o_1 _0772_ (.A1(net117),
    .A2(net58),
    .B1(net55),
    .B2(net113),
    .X(_0064_));
 sky130_fd_sc_hd__or2_2 _0773_ (.A(_0063_),
    .B(_0064_),
    .X(_0065_));
 sky130_fd_sc_hd__and4bb_1 _0774_ (.A_N(net129),
    .B_N(net127),
    .C(net133),
    .D(net131),
    .X(_0066_));
 sky130_fd_sc_hd__and4b_1 _0775_ (.A_N(net131),
    .B(net129),
    .C(net127),
    .D(net133),
    .X(_0067_));
 sky130_fd_sc_hd__a22o_2 _0776_ (.A1(net59),
    .A2(net53),
    .B1(net51),
    .B2(net55),
    .X(_0068_));
 sky130_fd_sc_hd__a22o_2 _0777_ (.A1(net107),
    .A2(net58),
    .B1(net55),
    .B2(net109),
    .X(_0069_));
 sky130_fd_sc_hd__and4bb_1 _0778_ (.A_N(net123),
    .B_N(net119),
    .C(net121),
    .D(net125),
    .X(_0070_));
 sky130_fd_sc_hd__nor4b_1 _0779_ (.A(net125),
    .B(net119),
    .C(net121),
    .D_N(net123),
    .Y(_0071_));
 sky130_fd_sc_hd__a22o_2 _0780_ (.A1(net51),
    .A2(net50),
    .B1(net48),
    .B2(net53),
    .X(_0072_));
 sky130_fd_sc_hd__nor4b_1 _0781_ (.A(net126),
    .B(net119),
    .C(_0702_),
    .D_N(net124),
    .Y(_0073_));
 sky130_fd_sc_hd__a22o_2 _0782_ (.A1(net95),
    .A2(net49),
    .B1(net47),
    .B2(net101),
    .X(_0074_));
 sky130_fd_sc_hd__or2_2 _0783_ (.A(net46),
    .B(_0074_),
    .X(_0075_));
 sky130_fd_sc_hd__a22o_2 _0784_ (.A1(net89),
    .A2(net50),
    .B1(net48),
    .B2(net84),
    .X(_0076_));
 sky130_fd_sc_hd__or2_1 _0785_ (.A(_0075_),
    .B(_0076_),
    .X(_0077_));
 sky130_fd_sc_hd__or2_2 _0786_ (.A(_0072_),
    .B(_0076_),
    .X(_0078_));
 sky130_fd_sc_hd__or2_2 _0787_ (.A(_0075_),
    .B(_0078_),
    .X(_0079_));
 sky130_fd_sc_hd__a22o_2 _0788_ (.A1(net96),
    .A2(net75),
    .B1(net73),
    .B2(net102),
    .X(_0080_));
 sky130_fd_sc_hd__a22o_1 _0789_ (.A1(net90),
    .A2(net74),
    .B1(net73),
    .B2(net85),
    .X(_0081_));
 sky130_fd_sc_hd__a22o_2 _0790_ (.A1(net72),
    .A2(net54),
    .B1(net52),
    .B2(net74),
    .X(_0082_));
 sky130_fd_sc_hd__or2_1 _0791_ (.A(_0080_),
    .B(_0081_),
    .X(_0083_));
 sky130_fd_sc_hd__or2_1 _0792_ (.A(_0082_),
    .B(_0083_),
    .X(_0084_));
 sky130_fd_sc_hd__a22o_1 _0793_ (.A1(net111),
    .A2(net53),
    .B1(net51),
    .B2(net115),
    .X(_0085_));
 sky130_fd_sc_hd__a22o_1 _0794_ (.A1(net116),
    .A2(net89),
    .B1(net84),
    .B2(net112),
    .X(_0086_));
 sky130_fd_sc_hd__or2_1 _0795_ (.A(_0085_),
    .B(_0086_),
    .X(_0087_));
 sky130_fd_sc_hd__a22o_1 _0796_ (.A1(net63),
    .A2(net54),
    .B1(net52),
    .B2(net61),
    .X(_0088_));
 sky130_fd_sc_hd__a22o_1 _0797_ (.A1(net101),
    .A2(net63),
    .B1(net61),
    .B2(net95),
    .X(_0089_));
 sky130_fd_sc_hd__a22o_1 _0798_ (.A1(net85),
    .A2(net62),
    .B1(net61),
    .B2(net90),
    .X(_0090_));
 sky130_fd_sc_hd__or2_1 _0799_ (.A(_0089_),
    .B(_0090_),
    .X(_0091_));
 sky130_fd_sc_hd__or3_1 _0800_ (.A(_0088_),
    .B(_0089_),
    .C(_0090_),
    .X(_0092_));
 sky130_fd_sc_hd__o21ba_2 _0801_ (.A1(net115),
    .A2(net55),
    .B1_N(_0702_),
    .X(_0093_));
 sky130_fd_sc_hd__a22o_2 _0802_ (.A1(net89),
    .A2(net58),
    .B1(net55),
    .B2(net84),
    .X(_0094_));
 sky130_fd_sc_hd__a22o_1 _0803_ (.A1(net95),
    .A2(net58),
    .B1(net56),
    .B2(net101),
    .X(_0095_));
 sky130_fd_sc_hd__or3_1 _0804_ (.A(_0093_),
    .B(_0094_),
    .C(_0095_),
    .X(_0096_));
 sky130_fd_sc_hd__a22o_2 _0805_ (.A1(net78),
    .A2(net49),
    .B1(net47),
    .B2(net76),
    .X(_0097_));
 sky130_fd_sc_hd__a22o_2 _0806_ (.A1(net109),
    .A2(net49),
    .B1(net47),
    .B2(net107),
    .X(_0098_));
 sky130_fd_sc_hd__o21ba_2 _0807_ (.A1(net49),
    .A2(net47),
    .B1_N(_0046_),
    .X(_0099_));
 sky130_fd_sc_hd__or2_1 _0808_ (.A(_0098_),
    .B(_0099_),
    .X(_0100_));
 sky130_fd_sc_hd__or3_1 _0809_ (.A(_0097_),
    .B(_0098_),
    .C(_0099_),
    .X(_0101_));
 sky130_fd_sc_hd__a22o_2 _0810_ (.A1(net107),
    .A2(net49),
    .B1(net47),
    .B2(net109),
    .X(_0102_));
 sky130_fd_sc_hd__a22o_2 _0811_ (.A1(net113),
    .A2(net49),
    .B1(net47),
    .B2(net117),
    .X(_0103_));
 sky130_fd_sc_hd__a22o_2 _0812_ (.A1(net115),
    .A2(net101),
    .B1(net95),
    .B2(net111),
    .X(_0104_));
 sky130_fd_sc_hd__a22o_2 _0813_ (.A1(net115),
    .A2(net68),
    .B1(net66),
    .B2(net111),
    .X(_0105_));
 sky130_fd_sc_hd__or4_1 _0814_ (.A(_0102_),
    .B(_0103_),
    .C(_0104_),
    .D(_0105_),
    .X(_0106_));
 sky130_fd_sc_hd__a22o_2 _0815_ (.A1(net110),
    .A2(net94),
    .B1(net92),
    .B2(net108),
    .X(_0107_));
 sky130_fd_sc_hd__or2_1 _0816_ (.A(_0647_),
    .B(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__a22o_1 _0817_ (.A1(net111),
    .A2(net109),
    .B1(net107),
    .B2(net116),
    .X(_0109_));
 sky130_fd_sc_hd__a22o_1 _0818_ (.A1(net91),
    .A2(net53),
    .B1(net51),
    .B2(net94),
    .X(_0110_));
 sky130_fd_sc_hd__nand3b_1 _0819_ (.A_N(net125),
    .B(net123),
    .C(net120),
    .Y(_0111_));
 sky130_fd_sc_hd__nor2_1 _0820_ (.A(_0702_),
    .B(_0111_),
    .Y(_0112_));
 sky130_fd_sc_hd__or2_1 _0821_ (.A(_0110_),
    .B(_0112_),
    .X(_0113_));
 sky130_fd_sc_hd__a22o_2 _0822_ (.A1(net106),
    .A2(net90),
    .B1(net85),
    .B2(net98),
    .X(_0114_));
 sky130_fd_sc_hd__a22o_2 _0823_ (.A1(net108),
    .A2(net105),
    .B1(net97),
    .B2(net110),
    .X(_0115_));
 sky130_fd_sc_hd__or2_1 _0824_ (.A(_0114_),
    .B(_0115_),
    .X(_0116_));
 sky130_fd_sc_hd__a22o_2 _0825_ (.A1(net96),
    .A2(net82),
    .B1(net80),
    .B2(net102),
    .X(_0117_));
 sky130_fd_sc_hd__a22o_1 _0826_ (.A1(net92),
    .A2(net79),
    .B1(net77),
    .B2(net93),
    .X(_0118_));
 sky130_fd_sc_hd__a22o_2 _0827_ (.A1(net114),
    .A2(net93),
    .B1(net92),
    .B2(net118),
    .X(_0119_));
 sky130_fd_sc_hd__a22o_1 _0828_ (.A1(net68),
    .A2(net50),
    .B1(net48),
    .B2(net66),
    .X(_0120_));
 sky130_fd_sc_hd__a22o_1 _0829_ (.A1(net98),
    .A2(net54),
    .B1(net52),
    .B2(net106),
    .X(_0121_));
 sky130_fd_sc_hd__a22o_1 _0830_ (.A1(net95),
    .A2(net62),
    .B1(net60),
    .B2(net101),
    .X(_0122_));
 sky130_fd_sc_hd__a22o_1 _0831_ (.A1(net114),
    .A2(net75),
    .B1(net72),
    .B2(net118),
    .X(_0123_));
 sky130_fd_sc_hd__o21ba_1 _0832_ (.A1(net74),
    .A2(net72),
    .B1_N(_0046_),
    .X(_0124_));
 sky130_fd_sc_hd__a22o_1 _0833_ (.A1(net108),
    .A2(net75),
    .B1(net72),
    .B2(net110),
    .X(_0125_));
 sky130_fd_sc_hd__or2_1 _0834_ (.A(_0124_),
    .B(_0125_),
    .X(_0126_));
 sky130_fd_sc_hd__or2_2 _0835_ (.A(_0123_),
    .B(_0125_),
    .X(_0127_));
 sky130_fd_sc_hd__or2_1 _0836_ (.A(_0124_),
    .B(_0127_),
    .X(_0128_));
 sky130_fd_sc_hd__a22o_1 _0837_ (.A1(net117),
    .A2(net105),
    .B1(net97),
    .B2(net113),
    .X(_0129_));
 sky130_fd_sc_hd__a22o_2 _0838_ (.A1(net105),
    .A2(net68),
    .B1(net66),
    .B2(net97),
    .X(_0130_));
 sky130_fd_sc_hd__a22o_2 _0839_ (.A1(net109),
    .A2(net105),
    .B1(net97),
    .B2(net107),
    .X(_0131_));
 sky130_fd_sc_hd__or4_1 _0840_ (.A(_0128_),
    .B(_0129_),
    .C(_0130_),
    .D(_0131_),
    .X(_0132_));
 sky130_fd_sc_hd__a22o_1 _0841_ (.A1(net85),
    .A2(net82),
    .B1(net80),
    .B2(net90),
    .X(_0133_));
 sky130_fd_sc_hd__a22o_1 _0842_ (.A1(net102),
    .A2(net82),
    .B1(net80),
    .B2(net96),
    .X(_0134_));
 sky130_fd_sc_hd__or2_2 _0843_ (.A(_0133_),
    .B(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__a22o_1 _0844_ (.A1(net108),
    .A2(net82),
    .B1(net80),
    .B2(net110),
    .X(_0136_));
 sky130_fd_sc_hd__a22o_2 _0845_ (.A1(net80),
    .A2(net79),
    .B1(net77),
    .B2(net82),
    .X(_0137_));
 sky130_fd_sc_hd__or4_1 _0846_ (.A(_0133_),
    .B(_0134_),
    .C(_0136_),
    .D(_0137_),
    .X(_0138_));
 sky130_fd_sc_hd__and2b_1 _0847_ (.A_N(_0702_),
    .B(net82),
    .X(_0139_));
 sky130_fd_sc_hd__o21ba_1 _0848_ (.A1(net82),
    .A2(net80),
    .B1_N(_0046_),
    .X(_0140_));
 sky130_fd_sc_hd__a22o_2 _0849_ (.A1(net82),
    .A2(net54),
    .B1(net52),
    .B2(net80),
    .X(_0141_));
 sky130_fd_sc_hd__a22o_1 _0850_ (.A1(net114),
    .A2(net82),
    .B1(net80),
    .B2(net118),
    .X(_0142_));
 sky130_fd_sc_hd__or4_1 _0851_ (.A(_0139_),
    .B(_0140_),
    .C(_0141_),
    .D(_0142_),
    .X(_0143_));
 sky130_fd_sc_hd__or2_1 _0852_ (.A(_0138_),
    .B(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__or4_1 _0853_ (.A(_0045_),
    .B(_0060_),
    .C(_0092_),
    .D(_0106_),
    .X(_0145_));
 sky130_fd_sc_hd__or4_1 _0854_ (.A(_0037_),
    .B(_0084_),
    .C(_0101_),
    .D(_0145_),
    .X(_0146_));
 sky130_fd_sc_hd__or4_1 _0855_ (.A(_0068_),
    .B(_0069_),
    .C(_0118_),
    .D(_0119_),
    .X(_0147_));
 sky130_fd_sc_hd__or4_1 _0856_ (.A(_0693_),
    .B(_0696_),
    .C(_0144_),
    .D(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__or2_2 _0857_ (.A(_0114_),
    .B(_0121_),
    .X(_0149_));
 sky130_fd_sc_hd__or4_1 _0858_ (.A(_0705_),
    .B(_0065_),
    .C(_0113_),
    .D(_0149_),
    .X(_0150_));
 sky130_fd_sc_hd__or3_1 _0859_ (.A(_0108_),
    .B(_0115_),
    .C(_0117_),
    .X(_0151_));
 sky130_fd_sc_hd__or4_1 _0860_ (.A(_0711_),
    .B(_0087_),
    .C(_0150_),
    .D(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__or4_1 _0861_ (.A(_0056_),
    .B(_0109_),
    .C(_0120_),
    .D(_0122_),
    .X(_0153_));
 sky130_fd_sc_hd__or4_1 _0862_ (.A(_0079_),
    .B(_0096_),
    .C(_0152_),
    .D(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__or3_1 _0863_ (.A(_0132_),
    .B(_0146_),
    .C(_0148_),
    .X(_0155_));
 sky130_fd_sc_hd__a22o_2 _0864_ (.A1(net66),
    .A2(net49),
    .B1(net47),
    .B2(net68),
    .X(_0156_));
 sky130_fd_sc_hd__a22o_2 _0865_ (.A1(net76),
    .A2(net49),
    .B1(net47),
    .B2(net78),
    .X(_0157_));
 sky130_fd_sc_hd__or2_1 _0866_ (.A(_0103_),
    .B(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__or4_1 _0867_ (.A(_0102_),
    .B(_0103_),
    .C(_0156_),
    .D(_0157_),
    .X(_0159_));
 sky130_fd_sc_hd__a22o_1 _0868_ (.A1(net68),
    .A2(net63),
    .B1(net61),
    .B2(net66),
    .X(_0160_));
 sky130_fd_sc_hd__or2_1 _0869_ (.A(_0088_),
    .B(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__or4_2 _0870_ (.A(_0088_),
    .B(_0089_),
    .C(_0090_),
    .D(_0160_),
    .X(_0162_));
 sky130_fd_sc_hd__or2_1 _0871_ (.A(_0056_),
    .B(_0162_),
    .X(_0163_));
 sky130_fd_sc_hd__a22o_2 _0872_ (.A1(net89),
    .A2(net62),
    .B1(net60),
    .B2(net84),
    .X(_0164_));
 sky130_fd_sc_hd__or2_1 _0873_ (.A(_0122_),
    .B(_0164_),
    .X(_0165_));
 sky130_fd_sc_hd__o21ba_4 _0874_ (.A1(net60),
    .A2(net50),
    .B1_N(_0702_),
    .X(_0166_));
 sky130_fd_sc_hd__a22o_2 _0875_ (.A1(net60),
    .A2(net53),
    .B1(net51),
    .B2(net62),
    .X(_0167_));
 sky130_fd_sc_hd__or2_1 _0876_ (.A(_0166_),
    .B(_0167_),
    .X(_0168_));
 sky130_fd_sc_hd__or4_1 _0877_ (.A(_0122_),
    .B(_0164_),
    .C(_0166_),
    .D(_0167_),
    .X(_0169_));
 sky130_fd_sc_hd__a22o_2 _0878_ (.A1(net66),
    .A2(net62),
    .B1(net60),
    .B2(net68),
    .X(_0170_));
 sky130_fd_sc_hd__or2_2 _0879_ (.A(_0059_),
    .B(_0170_),
    .X(_0171_));
 sky130_fd_sc_hd__or4_1 _0880_ (.A(_0057_),
    .B(_0058_),
    .C(_0059_),
    .D(_0170_),
    .X(_0172_));
 sky130_fd_sc_hd__or4_1 _0881_ (.A(_0056_),
    .B(_0162_),
    .C(_0169_),
    .D(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__a22o_2 _0882_ (.A1(net117),
    .A2(net49),
    .B1(net47),
    .B2(net113),
    .X(_0174_));
 sky130_fd_sc_hd__or2_1 _0883_ (.A(_0100_),
    .B(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__or2_1 _0884_ (.A(_0097_),
    .B(_0174_),
    .X(_0176_));
 sky130_fd_sc_hd__or4_1 _0885_ (.A(_0097_),
    .B(_0098_),
    .C(_0099_),
    .D(_0174_),
    .X(_0177_));
 sky130_fd_sc_hd__a22o_2 _0886_ (.A1(net101),
    .A2(net50),
    .B1(net48),
    .B2(net95),
    .X(_0178_));
 sky130_fd_sc_hd__a22o_1 _0887_ (.A1(net84),
    .A2(net49),
    .B1(net47),
    .B2(net89),
    .X(_0179_));
 sky130_fd_sc_hd__or2_1 _0888_ (.A(_0178_),
    .B(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__a22o_2 _0889_ (.A1(net53),
    .A2(net50),
    .B1(net48),
    .B2(net51),
    .X(_0181_));
 sky130_fd_sc_hd__or2_1 _0890_ (.A(_0120_),
    .B(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__or3_1 _0891_ (.A(_0177_),
    .B(_0180_),
    .C(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__or4_1 _0892_ (.A(_0079_),
    .B(_0159_),
    .C(_0173_),
    .D(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__o21ba_2 _0893_ (.A1(net106),
    .A2(net98),
    .B1_N(_0046_),
    .X(_0185_));
 sky130_fd_sc_hd__a22o_1 _0894_ (.A1(net98),
    .A2(net79),
    .B1(net77),
    .B2(net106),
    .X(_0186_));
 sky130_fd_sc_hd__a22o_2 _0895_ (.A1(net114),
    .A2(net106),
    .B1(net98),
    .B2(net118),
    .X(_0187_));
 sky130_fd_sc_hd__or2_1 _0896_ (.A(_0186_),
    .B(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__or3_1 _0897_ (.A(_0115_),
    .B(_0186_),
    .C(_0187_),
    .X(_0189_));
 sky130_fd_sc_hd__or2_1 _0898_ (.A(_0185_),
    .B(_0186_),
    .X(_0190_));
 sky130_fd_sc_hd__or4_2 _0899_ (.A(_0115_),
    .B(_0185_),
    .C(_0186_),
    .D(_0187_),
    .X(_0191_));
 sky130_fd_sc_hd__a22o_1 _0900_ (.A1(net105),
    .A2(net78),
    .B1(net76),
    .B2(net97),
    .X(_0192_));
 sky130_fd_sc_hd__or3_2 _0901_ (.A(_0130_),
    .B(_0131_),
    .C(_0192_),
    .X(_0193_));
 sky130_fd_sc_hd__or2_2 _0902_ (.A(_0129_),
    .B(_0192_),
    .X(_0194_));
 sky130_fd_sc_hd__or3_1 _0903_ (.A(_0129_),
    .B(_0191_),
    .C(_0193_),
    .X(_0195_));
 sky130_fd_sc_hd__a22o_1 _0904_ (.A1(net97),
    .A2(net69),
    .B1(net67),
    .B2(net106),
    .X(_0196_));
 sky130_fd_sc_hd__a22o_2 _0905_ (.A1(net102),
    .A2(net97),
    .B1(net96),
    .B2(net105),
    .X(_0197_));
 sky130_fd_sc_hd__or2_2 _0906_ (.A(_0121_),
    .B(_0196_),
    .X(_0198_));
 sky130_fd_sc_hd__or2_1 _0907_ (.A(_0197_),
    .B(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__or2_1 _0908_ (.A(_0196_),
    .B(_0197_),
    .X(_0200_));
 sky130_fd_sc_hd__or4_4 _0909_ (.A(_0114_),
    .B(_0121_),
    .C(_0196_),
    .D(_0197_),
    .X(_0201_));
 sky130_fd_sc_hd__a22o_1 _0910_ (.A1(net97),
    .A2(net89),
    .B1(net84),
    .B2(net105),
    .X(_0202_));
 sky130_fd_sc_hd__a22o_4 _0911_ (.A1(net105),
    .A2(net53),
    .B1(net51),
    .B2(net97),
    .X(_0203_));
 sky130_fd_sc_hd__or2_1 _0912_ (.A(_0202_),
    .B(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__or2_2 _0913_ (.A(_0701_),
    .B(_0202_),
    .X(_0205_));
 sky130_fd_sc_hd__or2_1 _0914_ (.A(_0705_),
    .B(_0204_),
    .X(_0206_));
 sky130_fd_sc_hd__or3_1 _0915_ (.A(_0195_),
    .B(_0201_),
    .C(_0206_),
    .X(_0207_));
 sky130_fd_sc_hd__a22o_2 _0916_ (.A1(net91),
    .A2(net68),
    .B1(net66),
    .B2(net93),
    .X(_0208_));
 sky130_fd_sc_hd__or2_2 _0917_ (.A(_0118_),
    .B(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__a22o_2 _0918_ (.A1(net107),
    .A2(net93),
    .B1(net91),
    .B2(net109),
    .X(_0210_));
 sky130_fd_sc_hd__or4_1 _0919_ (.A(_0118_),
    .B(_0119_),
    .C(_0208_),
    .D(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__a22o_1 _0920_ (.A1(net95),
    .A2(net93),
    .B1(net92),
    .B2(net101),
    .X(_0212_));
 sky130_fd_sc_hd__or2_2 _0921_ (.A(_0110_),
    .B(_0212_),
    .X(_0213_));
 sky130_fd_sc_hd__a22o_2 _0922_ (.A1(net94),
    .A2(net89),
    .B1(net84),
    .B2(net91),
    .X(_0214_));
 sky130_fd_sc_hd__or2_2 _0923_ (.A(_0112_),
    .B(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__or3_2 _0924_ (.A(_0211_),
    .B(_0213_),
    .C(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__o21ba_2 _0925_ (.A1(net93),
    .A2(net91),
    .B1_N(_0046_),
    .X(_0217_));
 sky130_fd_sc_hd__or4_1 _0926_ (.A(_0043_),
    .B(_0044_),
    .C(_0107_),
    .D(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__a22o_1 _0927_ (.A1(net118),
    .A2(net74),
    .B1(net72),
    .B2(net114),
    .X(_0219_));
 sky130_fd_sc_hd__or2_1 _0928_ (.A(_0040_),
    .B(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__a22o_2 _0929_ (.A1(net117),
    .A2(net93),
    .B1(net91),
    .B2(net113),
    .X(_0221_));
 sky130_fd_sc_hd__a22o_2 _0930_ (.A1(net93),
    .A2(net79),
    .B1(net77),
    .B2(net91),
    .X(_0222_));
 sky130_fd_sc_hd__or2_1 _0931_ (.A(_0221_),
    .B(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__or4_1 _0932_ (.A(_0040_),
    .B(_0219_),
    .C(_0221_),
    .D(_0222_),
    .X(_0224_));
 sky130_fd_sc_hd__a22o_1 _0933_ (.A1(net73),
    .A2(net69),
    .B1(net67),
    .B2(net74),
    .X(_0225_));
 sky130_fd_sc_hd__or2_1 _0934_ (.A(_0082_),
    .B(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__or2_1 _0935_ (.A(_0080_),
    .B(_0225_),
    .X(_0227_));
 sky130_fd_sc_hd__or4_2 _0936_ (.A(_0080_),
    .B(_0081_),
    .C(_0082_),
    .D(_0225_),
    .X(_0228_));
 sky130_fd_sc_hd__a22o_1 _0937_ (.A1(net76),
    .A2(net74),
    .B1(net72),
    .B2(net78),
    .X(_0229_));
 sky130_fd_sc_hd__or2_1 _0938_ (.A(_0124_),
    .B(_0229_),
    .X(_0230_));
 sky130_fd_sc_hd__or4_4 _0939_ (.A(_0123_),
    .B(_0124_),
    .C(_0125_),
    .D(_0229_),
    .X(_0231_));
 sky130_fd_sc_hd__a22o_1 _0940_ (.A1(net83),
    .A2(net69),
    .B1(net67),
    .B2(net81),
    .X(_0232_));
 sky130_fd_sc_hd__or2_1 _0941_ (.A(_0032_),
    .B(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__or3_2 _0942_ (.A(_0032_),
    .B(_0036_),
    .C(_0232_),
    .X(_0234_));
 sky130_fd_sc_hd__or4_1 _0943_ (.A(_0032_),
    .B(_0033_),
    .C(_0036_),
    .D(_0232_),
    .X(_0235_));
 sky130_fd_sc_hd__a22o_2 _0944_ (.A1(net85),
    .A2(net75),
    .B1(net73),
    .B2(net90),
    .X(_0236_));
 sky130_fd_sc_hd__o21ba_1 _0945_ (.A1(net80),
    .A2(net75),
    .B1_N(_0702_),
    .X(_0237_));
 sky130_fd_sc_hd__or2_1 _0946_ (.A(_0236_),
    .B(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__a22o_1 _0947_ (.A1(net102),
    .A2(net74),
    .B1(net72),
    .B2(net96),
    .X(_0239_));
 sky130_fd_sc_hd__a22o_2 _0948_ (.A1(net74),
    .A2(net54),
    .B1(net52),
    .B2(net72),
    .X(_0240_));
 sky130_fd_sc_hd__or2_2 _0949_ (.A(_0239_),
    .B(_0240_),
    .X(_0241_));
 sky130_fd_sc_hd__or3_1 _0950_ (.A(_0236_),
    .B(_0237_),
    .C(_0240_),
    .X(_0242_));
 sky130_fd_sc_hd__or4_2 _0951_ (.A(_0236_),
    .B(_0237_),
    .C(_0239_),
    .D(_0240_),
    .X(_0243_));
 sky130_fd_sc_hd__a22o_2 _0952_ (.A1(net93),
    .A2(net54),
    .B1(net52),
    .B2(net91),
    .X(_0244_));
 sky130_fd_sc_hd__a22o_2 _0953_ (.A1(net93),
    .A2(net69),
    .B1(net67),
    .B2(net91),
    .X(_0245_));
 sky130_fd_sc_hd__or2_1 _0954_ (.A(_0711_),
    .B(_0245_),
    .X(_0246_));
 sky130_fd_sc_hd__or4_2 _0955_ (.A(_0707_),
    .B(_0710_),
    .C(_0244_),
    .D(_0245_),
    .X(_0247_));
 sky130_fd_sc_hd__a22o_2 _0956_ (.A1(net90),
    .A2(net83),
    .B1(net81),
    .B2(net85),
    .X(_0248_));
 sky130_fd_sc_hd__a22o_1 _0957_ (.A1(net80),
    .A2(net69),
    .B1(net67),
    .B2(net82),
    .X(_0249_));
 sky130_fd_sc_hd__a22o_2 _0958_ (.A1(net81),
    .A2(net53),
    .B1(net51),
    .B2(net83),
    .X(_0250_));
 sky130_fd_sc_hd__or2_1 _0959_ (.A(_0117_),
    .B(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__or2_1 _0960_ (.A(_0117_),
    .B(_0249_),
    .X(_0252_));
 sky130_fd_sc_hd__or3_1 _0961_ (.A(_0117_),
    .B(_0248_),
    .C(_0249_),
    .X(_0253_));
 sky130_fd_sc_hd__or4_1 _0962_ (.A(_0117_),
    .B(_0248_),
    .C(_0249_),
    .D(_0250_),
    .X(_0254_));
 sky130_fd_sc_hd__or4_1 _0963_ (.A(_0235_),
    .B(_0243_),
    .C(_0247_),
    .D(_0254_),
    .X(_0255_));
 sky130_fd_sc_hd__or4_1 _0964_ (.A(_0218_),
    .B(_0224_),
    .C(_0228_),
    .D(_0231_),
    .X(_0256_));
 sky130_fd_sc_hd__or4_2 _0965_ (.A(_0144_),
    .B(_0216_),
    .C(_0255_),
    .D(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__a22o_1 _0966_ (.A1(net109),
    .A2(net58),
    .B1(net55),
    .B2(net107),
    .X(_0258_));
 sky130_fd_sc_hd__o21ba_1 _0967_ (.A1(net58),
    .A2(net55),
    .B1_N(_0046_),
    .X(_0259_));
 sky130_fd_sc_hd__or2_1 _0968_ (.A(_0065_),
    .B(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__or2_1 _0969_ (.A(_0258_),
    .B(_0259_),
    .X(_0261_));
 sky130_fd_sc_hd__or4_4 _0970_ (.A(_0063_),
    .B(_0064_),
    .C(_0258_),
    .D(_0259_),
    .X(_0262_));
 sky130_fd_sc_hd__a22o_1 _0971_ (.A1(net84),
    .A2(net59),
    .B1(net56),
    .B2(net89),
    .X(_0263_));
 sky130_fd_sc_hd__a22o_2 _0972_ (.A1(net101),
    .A2(net58),
    .B1(net56),
    .B2(net95),
    .X(_0264_));
 sky130_fd_sc_hd__or2_2 _0973_ (.A(_0068_),
    .B(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__a22o_1 _0974_ (.A1(net68),
    .A2(net59),
    .B1(net56),
    .B2(net66),
    .X(_0266_));
 sky130_fd_sc_hd__or3_2 _0975_ (.A(_0068_),
    .B(_0264_),
    .C(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__or2_2 _0976_ (.A(_0263_),
    .B(_0266_),
    .X(_0268_));
 sky130_fd_sc_hd__or3_1 _0977_ (.A(_0262_),
    .B(_0265_),
    .C(_0268_),
    .X(_0269_));
 sky130_fd_sc_hd__a22o_2 _0978_ (.A1(net55),
    .A2(net53),
    .B1(net51),
    .B2(net58),
    .X(_0270_));
 sky130_fd_sc_hd__or2_1 _0979_ (.A(_0095_),
    .B(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__or2_1 _0980_ (.A(_0093_),
    .B(_0270_),
    .X(_0272_));
 sky130_fd_sc_hd__or4_2 _0981_ (.A(_0093_),
    .B(_0094_),
    .C(_0095_),
    .D(_0270_),
    .X(_0273_));
 sky130_fd_sc_hd__a22o_2 _0982_ (.A1(net111),
    .A2(net68),
    .B1(net66),
    .B2(net116),
    .X(_0274_));
 sky130_fd_sc_hd__or2_2 _0983_ (.A(_0109_),
    .B(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__a22o_1 _0984_ (.A1(net116),
    .A2(net113),
    .B1(net112),
    .B2(net117),
    .X(_0276_));
 sky130_fd_sc_hd__a22o_1 _0985_ (.A1(net112),
    .A2(net78),
    .B1(net76),
    .B2(net116),
    .X(_0277_));
 sky130_fd_sc_hd__or2_2 _0986_ (.A(_0276_),
    .B(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__or3_1 _0987_ (.A(_0273_),
    .B(_0275_),
    .C(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__a22o_1 _0988_ (.A1(net115),
    .A2(net78),
    .B1(net76),
    .B2(net111),
    .X(_0280_));
 sky130_fd_sc_hd__or2_1 _0989_ (.A(_0693_),
    .B(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__a22o_1 _0990_ (.A1(net111),
    .A2(net89),
    .B1(net84),
    .B2(net115),
    .X(_0282_));
 sky130_fd_sc_hd__or2_2 _0991_ (.A(_0104_),
    .B(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__or4_1 _0992_ (.A(_0693_),
    .B(_0104_),
    .C(_0280_),
    .D(_0282_),
    .X(_0284_));
 sky130_fd_sc_hd__a22o_2 _0993_ (.A1(net112),
    .A2(net101),
    .B1(net95),
    .B2(net116),
    .X(_0285_));
 sky130_fd_sc_hd__or2_2 _0994_ (.A(_0085_),
    .B(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__or4_1 _0995_ (.A(net125),
    .B(net123),
    .C(net121),
    .D(_0702_),
    .X(_0287_));
 sky130_fd_sc_hd__or2_2 _0996_ (.A(_0086_),
    .B(_0285_),
    .X(_0288_));
 sky130_fd_sc_hd__or4b_1 _0997_ (.A(_0085_),
    .B(_0284_),
    .C(_0288_),
    .D_N(_0287_),
    .X(_0289_));
 sky130_fd_sc_hd__a22o_1 _0998_ (.A1(net115),
    .A2(net53),
    .B1(net51),
    .B2(net111),
    .X(_0290_));
 sky130_fd_sc_hd__or2_1 _0999_ (.A(_0105_),
    .B(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__o21ba_2 _1000_ (.A1(net115),
    .A2(net112),
    .B1_N(_0046_),
    .X(_0292_));
 sky130_fd_sc_hd__or2_1 _1001_ (.A(_0696_),
    .B(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__or4_1 _1002_ (.A(_0696_),
    .B(_0105_),
    .C(_0290_),
    .D(_0292_),
    .X(_0294_));
 sky130_fd_sc_hd__a22o_2 _1003_ (.A1(net66),
    .A2(net59),
    .B1(net56),
    .B2(net68),
    .X(_0295_));
 sky130_fd_sc_hd__or2_1 _1004_ (.A(_0069_),
    .B(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__a22o_2 _1005_ (.A1(net76),
    .A2(net59),
    .B1(net56),
    .B2(net78),
    .X(_0297_));
 sky130_fd_sc_hd__a22o_2 _1006_ (.A1(net113),
    .A2(net58),
    .B1(net55),
    .B2(net117),
    .X(_0298_));
 sky130_fd_sc_hd__or2_1 _1007_ (.A(_0297_),
    .B(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__or2_1 _1008_ (.A(_0295_),
    .B(_0298_),
    .X(_0300_));
 sky130_fd_sc_hd__or4_1 _1009_ (.A(_0069_),
    .B(_0295_),
    .C(_0297_),
    .D(_0298_),
    .X(_0301_));
 sky130_fd_sc_hd__or2_1 _1010_ (.A(_0294_),
    .B(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__or4_1 _1011_ (.A(_0269_),
    .B(_0279_),
    .C(_0289_),
    .D(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__nor4_1 _1012_ (.A(_0184_),
    .B(_0207_),
    .C(_0257_),
    .D(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__o32a_1 _1013_ (.A1(_0154_),
    .A2(_0155_),
    .A3(net45),
    .B1(net137),
    .B2(net144),
    .X(_0000_));
 sky130_fd_sc_hd__or2_2 _1014_ (.A(_0704_),
    .B(_0202_),
    .X(_0305_));
 sky130_fd_sc_hd__or2_1 _1015_ (.A(_0193_),
    .B(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__or3_1 _1016_ (.A(_0097_),
    .B(_0099_),
    .C(_0198_),
    .X(_0307_));
 sky130_fd_sc_hd__or2_1 _1017_ (.A(net135),
    .B(_0043_),
    .X(_0308_));
 sky130_fd_sc_hd__or2_1 _1018_ (.A(_0217_),
    .B(_0244_),
    .X(_0309_));
 sky130_fd_sc_hd__or3_1 _1019_ (.A(_0109_),
    .B(_0274_),
    .C(_0276_),
    .X(_0310_));
 sky130_fd_sc_hd__or2_1 _1020_ (.A(_0086_),
    .B(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__or2_1 _1021_ (.A(_0136_),
    .B(_0142_),
    .X(_0312_));
 sky130_fd_sc_hd__or3_1 _1022_ (.A(_0248_),
    .B(_0249_),
    .C(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__or2_1 _1023_ (.A(_0069_),
    .B(_0094_),
    .X(_0314_));
 sky130_fd_sc_hd__or4_1 _1024_ (.A(_0308_),
    .B(_0309_),
    .C(_0311_),
    .D(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__or3_1 _1025_ (.A(_0260_),
    .B(_0307_),
    .C(_0313_),
    .X(_0316_));
 sky130_fd_sc_hd__or4_1 _1026_ (.A(_0078_),
    .B(_0165_),
    .C(_0265_),
    .D(_0271_),
    .X(_0317_));
 sky130_fd_sc_hd__or4_1 _1027_ (.A(_0036_),
    .B(_0040_),
    .C(_0080_),
    .D(_0112_),
    .X(_0318_));
 sky130_fd_sc_hd__or3_1 _1028_ (.A(_0051_),
    .B(_0161_),
    .C(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__or4_1 _1029_ (.A(_0125_),
    .B(_0137_),
    .C(_0187_),
    .D(_0212_),
    .X(_0320_));
 sky130_fd_sc_hd__or4_1 _1030_ (.A(_0052_),
    .B(_0103_),
    .C(_0170_),
    .D(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__or3_1 _1031_ (.A(_0135_),
    .B(_0232_),
    .C(_0284_),
    .X(_0322_));
 sky130_fd_sc_hd__or4_1 _1032_ (.A(_0317_),
    .B(_0319_),
    .C(_0321_),
    .D(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__or4_1 _1033_ (.A(_0306_),
    .B(_0315_),
    .C(_0316_),
    .D(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__o22a_1 _1034_ (.A1(net136),
    .A2(net148),
    .B1(net42),
    .B2(_0324_),
    .X(_0001_));
 sky130_fd_sc_hd__or3_1 _1035_ (.A(_0068_),
    .B(_0253_),
    .C(_0268_),
    .X(_0325_));
 sky130_fd_sc_hd__or2_1 _1036_ (.A(_0105_),
    .B(_0179_),
    .X(_0326_));
 sky130_fd_sc_hd__or2_1 _1037_ (.A(_0133_),
    .B(_0141_),
    .X(_0327_));
 sky130_fd_sc_hd__or4_1 _1038_ (.A(_0089_),
    .B(_0133_),
    .C(_0141_),
    .D(_0160_),
    .X(_0328_));
 sky130_fd_sc_hd__or3_1 _1039_ (.A(_0102_),
    .B(_0103_),
    .C(_0156_),
    .X(_0329_));
 sky130_fd_sc_hd__or4_1 _1040_ (.A(_0093_),
    .B(_0094_),
    .C(_0211_),
    .D(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__or3_1 _1041_ (.A(_0037_),
    .B(_0182_),
    .C(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__or3_2 _1042_ (.A(_0112_),
    .B(_0212_),
    .C(_0214_),
    .X(_0332_));
 sky130_fd_sc_hd__or2_1 _1043_ (.A(_0707_),
    .B(_0244_),
    .X(_0333_));
 sky130_fd_sc_hd__or4_1 _1044_ (.A(_0121_),
    .B(_0197_),
    .C(_0332_),
    .D(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__or4_1 _1045_ (.A(_0049_),
    .B(_0059_),
    .C(_0069_),
    .D(_0298_),
    .X(_0335_));
 sky130_fd_sc_hd__or2_1 _1046_ (.A(net135),
    .B(_0057_),
    .X(_0336_));
 sky130_fd_sc_hd__or3_1 _1047_ (.A(_0166_),
    .B(_0221_),
    .C(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__or2_1 _1048_ (.A(_0220_),
    .B(_0242_),
    .X(_0338_));
 sky130_fd_sc_hd__or4_1 _1049_ (.A(_0115_),
    .B(_0124_),
    .C(_0137_),
    .D(_0274_),
    .X(_0339_));
 sky130_fd_sc_hd__or4_1 _1050_ (.A(_0194_),
    .B(_0205_),
    .C(_0328_),
    .D(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__or4_1 _1051_ (.A(_0261_),
    .B(_0278_),
    .C(_0288_),
    .D(_0293_),
    .X(_0341_));
 sky130_fd_sc_hd__or4_1 _1052_ (.A(_0078_),
    .B(_0176_),
    .C(_0190_),
    .D(_0227_),
    .X(_0342_));
 sky130_fd_sc_hd__or4_1 _1053_ (.A(_0337_),
    .B(_0340_),
    .C(_0341_),
    .D(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__or2_1 _1054_ (.A(_0326_),
    .B(_0335_),
    .X(_0344_));
 sky130_fd_sc_hd__or4_1 _1055_ (.A(_0325_),
    .B(_0334_),
    .C(_0338_),
    .D(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__or3_1 _1056_ (.A(_0331_),
    .B(_0343_),
    .C(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__o22a_1 _1057_ (.A1(net139),
    .A2(net160),
    .B1(net44),
    .B2(_0346_),
    .X(_0002_));
 sky130_fd_sc_hd__or2_1 _1058_ (.A(_0711_),
    .B(_0244_),
    .X(_0347_));
 sky130_fd_sc_hd__or2_1 _1059_ (.A(_0043_),
    .B(_0220_),
    .X(_0348_));
 sky130_fd_sc_hd__or2_1 _1060_ (.A(_0693_),
    .B(_0292_),
    .X(_0349_));
 sky130_fd_sc_hd__or3_1 _1061_ (.A(_0693_),
    .B(_0280_),
    .C(_0292_),
    .X(_0350_));
 sky130_fd_sc_hd__or3_1 _1062_ (.A(_0057_),
    .B(_0171_),
    .C(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__or2_1 _1063_ (.A(net135),
    .B(_0186_),
    .X(_0352_));
 sky130_fd_sc_hd__or3_1 _1064_ (.A(_0117_),
    .B(_0131_),
    .C(_0137_),
    .X(_0353_));
 sky130_fd_sc_hd__or3_1 _1065_ (.A(_0204_),
    .B(_0352_),
    .C(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__or4_1 _1066_ (.A(_0032_),
    .B(_0164_),
    .C(_0166_),
    .D(_0240_),
    .X(_0355_));
 sky130_fd_sc_hd__or4_1 _1067_ (.A(_0103_),
    .B(_0156_),
    .C(_0212_),
    .D(_0214_),
    .X(_0356_));
 sky130_fd_sc_hd__or3_1 _1068_ (.A(_0107_),
    .B(_0217_),
    .C(_0221_),
    .X(_0357_));
 sky130_fd_sc_hd__or2_1 _1069_ (.A(_0097_),
    .B(_0236_),
    .X(_0358_));
 sky130_fd_sc_hd__or3_1 _1070_ (.A(_0311_),
    .B(_0351_),
    .C(_0354_),
    .X(_0359_));
 sky130_fd_sc_hd__or4_1 _1071_ (.A(_0126_),
    .B(_0286_),
    .C(_0291_),
    .D(_0358_),
    .X(_0360_));
 sky130_fd_sc_hd__or4_1 _1072_ (.A(_0347_),
    .B(_0348_),
    .C(_0355_),
    .D(_0357_),
    .X(_0361_));
 sky130_fd_sc_hd__or4_1 _1073_ (.A(_0055_),
    .B(_0079_),
    .C(_0328_),
    .D(_0356_),
    .X(_0362_));
 sky130_fd_sc_hd__or4_1 _1074_ (.A(_0068_),
    .B(_0093_),
    .C(_0104_),
    .D(_0211_),
    .X(_0363_));
 sky130_fd_sc_hd__or4_1 _1075_ (.A(_0360_),
    .B(_0361_),
    .C(_0362_),
    .D(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__o32a_1 _1076_ (.A1(net44),
    .A2(_0359_),
    .A3(_0364_),
    .B1(net162),
    .B2(net139),
    .X(_0003_));
 sky130_fd_sc_hd__or2_1 _1077_ (.A(_0236_),
    .B(_0239_),
    .X(_0365_));
 sky130_fd_sc_hd__or3_2 _1078_ (.A(_0189_),
    .B(_0296_),
    .C(_0297_),
    .X(_0366_));
 sky130_fd_sc_hd__or2_1 _1079_ (.A(_0058_),
    .B(_0171_),
    .X(_0367_));
 sky130_fd_sc_hd__or2_1 _1080_ (.A(_0080_),
    .B(_0226_),
    .X(_0368_));
 sky130_fd_sc_hd__or2_1 _1081_ (.A(_0088_),
    .B(_0103_),
    .X(_0369_));
 sky130_fd_sc_hd__or3_2 _1082_ (.A(_0217_),
    .B(_0221_),
    .C(_0222_),
    .X(_0370_));
 sky130_fd_sc_hd__or3_1 _1083_ (.A(_0131_),
    .B(_0192_),
    .C(_0349_),
    .X(_0371_));
 sky130_fd_sc_hd__or2_1 _1084_ (.A(_0263_),
    .B(_0264_),
    .X(_0372_));
 sky130_fd_sc_hd__or2_1 _1085_ (.A(_0264_),
    .B(_0268_),
    .X(_0373_));
 sky130_fd_sc_hd__or4_1 _1086_ (.A(net135),
    .B(net46),
    .C(_0105_),
    .D(_0274_),
    .X(_0374_));
 sky130_fd_sc_hd__or4_1 _1087_ (.A(_0098_),
    .B(_0176_),
    .C(_0234_),
    .D(_0367_),
    .X(_0375_));
 sky130_fd_sc_hd__or3_1 _1088_ (.A(_0043_),
    .B(_0245_),
    .C(_0369_),
    .X(_0376_));
 sky130_fd_sc_hd__or4_1 _1089_ (.A(_0126_),
    .B(_0288_),
    .C(_0366_),
    .D(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__or4_1 _1090_ (.A(_0051_),
    .B(_0065_),
    .C(_0135_),
    .D(_0271_),
    .X(_0378_));
 sky130_fd_sc_hd__or4_1 _1091_ (.A(_0076_),
    .B(_0110_),
    .C(_0178_),
    .D(_0210_),
    .X(_0379_));
 sky130_fd_sc_hd__or4_1 _1092_ (.A(_0710_),
    .B(_0121_),
    .C(_0142_),
    .D(_0250_),
    .X(_0380_));
 sky130_fd_sc_hd__or4_1 _1093_ (.A(_0377_),
    .B(_0378_),
    .C(_0379_),
    .D(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__or4_1 _1094_ (.A(_0169_),
    .B(_0206_),
    .C(_0371_),
    .D(_0374_),
    .X(_0382_));
 sky130_fd_sc_hd__or4_1 _1095_ (.A(_0240_),
    .B(_0365_),
    .C(_0368_),
    .D(_0373_),
    .X(_0383_));
 sky130_fd_sc_hd__or4_1 _1096_ (.A(_0370_),
    .B(_0375_),
    .C(_0382_),
    .D(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__o32a_1 _1097_ (.A1(net44),
    .A2(_0381_),
    .A3(_0384_),
    .B1(net163),
    .B2(net139),
    .X(_0004_));
 sky130_fd_sc_hd__or2_1 _1098_ (.A(_0099_),
    .B(_0102_),
    .X(_0385_));
 sky130_fd_sc_hd__or3_1 _1099_ (.A(_0704_),
    .B(_0130_),
    .C(_0131_),
    .X(_0386_));
 sky130_fd_sc_hd__or2_1 _1100_ (.A(_0068_),
    .B(_0072_),
    .X(_0387_));
 sky130_fd_sc_hd__or3_2 _1101_ (.A(_0109_),
    .B(_0276_),
    .C(_0288_),
    .X(_0388_));
 sky130_fd_sc_hd__or2_1 _1102_ (.A(_0044_),
    .B(_0219_),
    .X(_0389_));
 sky130_fd_sc_hd__or3_1 _1103_ (.A(_0043_),
    .B(_0044_),
    .C(_0219_),
    .X(_0390_));
 sky130_fd_sc_hd__or2_1 _1104_ (.A(_0236_),
    .B(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__or3_2 _1105_ (.A(_0284_),
    .B(_0290_),
    .C(_0292_),
    .X(_0392_));
 sky130_fd_sc_hd__or4_1 _1106_ (.A(_0198_),
    .B(_0233_),
    .C(_0296_),
    .D(_0298_),
    .X(_0393_));
 sky130_fd_sc_hd__or2_1 _1107_ (.A(_0208_),
    .B(_0222_),
    .X(_0394_));
 sky130_fd_sc_hd__or4_1 _1108_ (.A(_0241_),
    .B(_0386_),
    .C(_0388_),
    .D(_0391_),
    .X(_0395_));
 sky130_fd_sc_hd__or4_1 _1109_ (.A(_0055_),
    .B(_0253_),
    .C(_0262_),
    .D(_0332_),
    .X(_0396_));
 sky130_fd_sc_hd__or4_1 _1110_ (.A(_0083_),
    .B(_0102_),
    .C(_0135_),
    .D(_0156_),
    .X(_0397_));
 sky130_fd_sc_hd__or4_1 _1111_ (.A(_0088_),
    .B(_0123_),
    .C(_0136_),
    .D(_0270_),
    .X(_0398_));
 sky130_fd_sc_hd__or4_1 _1112_ (.A(_0711_),
    .B(_0057_),
    .C(_0058_),
    .D(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__or4_1 _1113_ (.A(_0352_),
    .B(_0396_),
    .C(_0397_),
    .D(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__or4_1 _1114_ (.A(_0100_),
    .B(_0168_),
    .C(_0387_),
    .D(_0394_),
    .X(_0401_));
 sky130_fd_sc_hd__or3_1 _1115_ (.A(_0392_),
    .B(_0393_),
    .C(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__or3_1 _1116_ (.A(_0395_),
    .B(_0400_),
    .C(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__o22a_1 _1117_ (.A1(net138),
    .A2(net157),
    .B1(net43),
    .B2(_0403_),
    .X(_0005_));
 sky130_fd_sc_hd__or2_1 _1118_ (.A(_0120_),
    .B(_0178_),
    .X(_0404_));
 sky130_fd_sc_hd__or3_1 _1119_ (.A(_0120_),
    .B(_0178_),
    .C(_0179_),
    .X(_0405_));
 sky130_fd_sc_hd__or3_1 _1120_ (.A(_0209_),
    .B(_0210_),
    .C(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__or3_1 _1121_ (.A(_0274_),
    .B(_0278_),
    .C(_0286_),
    .X(_0407_));
 sky130_fd_sc_hd__or4_1 _1122_ (.A(_0116_),
    .B(_0251_),
    .C(_0295_),
    .D(_0299_),
    .X(_0408_));
 sky130_fd_sc_hd__or4_1 _1123_ (.A(_0696_),
    .B(_0052_),
    .C(_0054_),
    .D(_0281_),
    .X(_0409_));
 sky130_fd_sc_hd__or4_1 _1124_ (.A(_0406_),
    .B(_0407_),
    .C(_0408_),
    .D(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__or2_1 _1125_ (.A(_0232_),
    .B(_0240_),
    .X(_0411_));
 sky130_fd_sc_hd__or2_1 _1126_ (.A(_0136_),
    .B(_0140_),
    .X(_0412_));
 sky130_fd_sc_hd__or2_1 _1127_ (.A(_0137_),
    .B(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__or2_1 _1128_ (.A(_0064_),
    .B(_0068_),
    .X(_0414_));
 sky130_fd_sc_hd__or2_1 _1129_ (.A(_0105_),
    .B(_0259_),
    .X(_0415_));
 sky130_fd_sc_hd__or2_1 _1130_ (.A(_0093_),
    .B(_0170_),
    .X(_0416_));
 sky130_fd_sc_hd__or4_1 _1131_ (.A(_0135_),
    .B(_0141_),
    .C(_0368_),
    .D(_0413_),
    .X(_0417_));
 sky130_fd_sc_hd__or4_1 _1132_ (.A(_0112_),
    .B(_0185_),
    .C(_0203_),
    .D(_0237_),
    .X(_0418_));
 sky130_fd_sc_hd__or4_1 _1133_ (.A(_0057_),
    .B(_0076_),
    .C(_0097_),
    .D(_0164_),
    .X(_0419_));
 sky130_fd_sc_hd__or4_1 _1134_ (.A(_0128_),
    .B(_0347_),
    .C(_0418_),
    .D(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__or4_1 _1135_ (.A(_0411_),
    .B(_0414_),
    .C(_0415_),
    .D(_0416_),
    .X(_0421_));
 sky130_fd_sc_hd__or4_1 _1136_ (.A(_0108_),
    .B(_0220_),
    .C(_0283_),
    .D(_0372_),
    .X(_0422_));
 sky130_fd_sc_hd__or4_1 _1137_ (.A(_0417_),
    .B(_0420_),
    .C(_0421_),
    .D(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__o32a_1 _1138_ (.A1(net44),
    .A2(_0410_),
    .A3(_0423_),
    .B1(net165),
    .B2(net138),
    .X(_0006_));
 sky130_fd_sc_hd__or2_1 _1139_ (.A(_0164_),
    .B(_0167_),
    .X(_0424_));
 sky130_fd_sc_hd__or3_1 _1140_ (.A(_0252_),
    .B(_0267_),
    .C(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__or4_1 _1141_ (.A(_0221_),
    .B(_0222_),
    .C(_0244_),
    .D(_0245_),
    .X(_0426_));
 sky130_fd_sc_hd__or3_1 _1142_ (.A(_0052_),
    .B(_0054_),
    .C(_0162_),
    .X(_0427_));
 sky130_fd_sc_hd__or2_1 _1143_ (.A(_0181_),
    .B(_0404_),
    .X(_0428_));
 sky130_fd_sc_hd__or2_1 _1144_ (.A(_0064_),
    .B(_0258_),
    .X(_0429_));
 sky130_fd_sc_hd__or3_2 _1145_ (.A(_0064_),
    .B(_0258_),
    .C(_0259_),
    .X(_0430_));
 sky130_fd_sc_hd__or2_1 _1146_ (.A(_0707_),
    .B(_0118_),
    .X(_0431_));
 sky130_fd_sc_hd__or2_1 _1147_ (.A(_0140_),
    .B(_0229_),
    .X(_0432_));
 sky130_fd_sc_hd__or4_1 _1148_ (.A(_0100_),
    .B(_0194_),
    .C(_0238_),
    .D(_0314_),
    .X(_0433_));
 sky130_fd_sc_hd__or4_1 _1149_ (.A(net135),
    .B(_0082_),
    .C(_0431_),
    .D(_0432_),
    .X(_0434_));
 sky130_fd_sc_hd__or4_1 _1150_ (.A(_0425_),
    .B(_0427_),
    .C(_0433_),
    .D(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__or3_1 _1151_ (.A(_0077_),
    .B(_0426_),
    .C(_0428_),
    .X(_0436_));
 sky130_fd_sc_hd__or4_1 _1152_ (.A(_0060_),
    .B(_0203_),
    .C(_0305_),
    .D(_0430_),
    .X(_0437_));
 sky130_fd_sc_hd__or4_1 _1153_ (.A(_0696_),
    .B(_0086_),
    .C(_0104_),
    .D(_0191_),
    .X(_0438_));
 sky130_fd_sc_hd__or4_1 _1154_ (.A(_0130_),
    .B(_0156_),
    .C(_0157_),
    .D(_0214_),
    .X(_0439_));
 sky130_fd_sc_hd__or3_1 _1155_ (.A(_0127_),
    .B(_0389_),
    .C(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__or4_2 _1156_ (.A(_0199_),
    .B(_0437_),
    .C(_0438_),
    .D(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__or3_1 _1157_ (.A(_0435_),
    .B(_0436_),
    .C(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__o22a_1 _1158_ (.A1(net138),
    .A2(net166),
    .B1(net43),
    .B2(_0442_),
    .X(_0007_));
 sky130_fd_sc_hd__or4_1 _1159_ (.A(_0117_),
    .B(_0137_),
    .C(_0217_),
    .D(_0221_),
    .X(_0443_));
 sky130_fd_sc_hd__or4_1 _1160_ (.A(_0040_),
    .B(_0208_),
    .C(_0210_),
    .D(_0213_),
    .X(_0444_));
 sky130_fd_sc_hd__or4_2 _1161_ (.A(_0056_),
    .B(_0065_),
    .C(_0263_),
    .D(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__or3_1 _1162_ (.A(_0185_),
    .B(_0186_),
    .C(_0187_),
    .X(_0446_));
 sky130_fd_sc_hd__or4_1 _1163_ (.A(net135),
    .B(_0693_),
    .C(net46),
    .D(_0329_),
    .X(_0447_));
 sky130_fd_sc_hd__or4_1 _1164_ (.A(_0057_),
    .B(_0171_),
    .C(_0246_),
    .D(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__or2_1 _1165_ (.A(_0149_),
    .B(_0446_),
    .X(_0449_));
 sky130_fd_sc_hd__or4_1 _1166_ (.A(_0069_),
    .B(_0272_),
    .C(_0297_),
    .D(_0411_),
    .X(_0450_));
 sky130_fd_sc_hd__or4_1 _1167_ (.A(_0141_),
    .B(_0205_),
    .C(_0230_),
    .D(_0248_),
    .X(_0451_));
 sky130_fd_sc_hd__or3_1 _1168_ (.A(_0168_),
    .B(_0176_),
    .C(_0443_),
    .X(_0452_));
 sky130_fd_sc_hd__or4_1 _1169_ (.A(_0091_),
    .B(_0449_),
    .C(_0451_),
    .D(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__or3_1 _1170_ (.A(_0275_),
    .B(_0285_),
    .C(_0405_),
    .X(_0454_));
 sky130_fd_sc_hd__or4_1 _1171_ (.A(_0084_),
    .B(_0193_),
    .C(_0290_),
    .D(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__or4_1 _1172_ (.A(_0445_),
    .B(_0450_),
    .C(_0453_),
    .D(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__o32a_1 _1173_ (.A1(net42),
    .A2(_0448_),
    .A3(_0456_),
    .B1(net147),
    .B2(net136),
    .X(_0008_));
 sky130_fd_sc_hd__or2_1 _1174_ (.A(_0089_),
    .B(_0161_),
    .X(_0457_));
 sky130_fd_sc_hd__or3_1 _1175_ (.A(_0107_),
    .B(_0217_),
    .C(_0222_),
    .X(_0458_));
 sky130_fd_sc_hd__or4_1 _1176_ (.A(_0086_),
    .B(_0094_),
    .C(_0280_),
    .D(_0282_),
    .X(_0459_));
 sky130_fd_sc_hd__or2_1 _1177_ (.A(net135),
    .B(_0133_),
    .X(_0460_));
 sky130_fd_sc_hd__or3_1 _1178_ (.A(_0705_),
    .B(_0203_),
    .C(_0458_),
    .X(_0461_));
 sky130_fd_sc_hd__or4_1 _1179_ (.A(_0033_),
    .B(_0098_),
    .C(_0157_),
    .D(_0167_),
    .X(_0462_));
 sky130_fd_sc_hd__or3_1 _1180_ (.A(_0053_),
    .B(_0275_),
    .C(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__or4_1 _1181_ (.A(_0355_),
    .B(_0457_),
    .C(_0461_),
    .D(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__or4_1 _1182_ (.A(_0252_),
    .B(_0300_),
    .C(_0406_),
    .D(_0460_),
    .X(_0465_));
 sky130_fd_sc_hd__or4_1 _1183_ (.A(_0049_),
    .B(_0389_),
    .C(_0414_),
    .D(_0459_),
    .X(_0466_));
 sky130_fd_sc_hd__or4_1 _1184_ (.A(_0060_),
    .B(_0228_),
    .C(_0446_),
    .D(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__or4_1 _1185_ (.A(_0132_),
    .B(_0334_),
    .C(_0465_),
    .D(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__o32a_1 _1186_ (.A1(net44),
    .A2(_0464_),
    .A3(_0468_),
    .B1(net154),
    .B2(net139),
    .X(_0009_));
 sky130_fd_sc_hd__or2_1 _1187_ (.A(_0157_),
    .B(_0174_),
    .X(_0469_));
 sky130_fd_sc_hd__or2_1 _1188_ (.A(_0081_),
    .B(_0225_),
    .X(_0470_));
 sky130_fd_sc_hd__or2_1 _1189_ (.A(_0082_),
    .B(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__or3_1 _1190_ (.A(_0113_),
    .B(_0164_),
    .C(_0166_),
    .X(_0472_));
 sky130_fd_sc_hd__or2_1 _1191_ (.A(_0185_),
    .B(_0187_),
    .X(_0473_));
 sky130_fd_sc_hd__or2_1 _1192_ (.A(_0107_),
    .B(_0250_),
    .X(_0474_));
 sky130_fd_sc_hd__or2_1 _1193_ (.A(_0058_),
    .B(_0122_),
    .X(_0475_));
 sky130_fd_sc_hd__or4_1 _1194_ (.A(_0246_),
    .B(_0457_),
    .C(_0471_),
    .D(_0472_),
    .X(_0476_));
 sky130_fd_sc_hd__or4_1 _1195_ (.A(_0045_),
    .B(_0128_),
    .C(_0260_),
    .D(_0373_),
    .X(_0477_));
 sky130_fd_sc_hd__or4_1 _1196_ (.A(_0696_),
    .B(_0074_),
    .C(_0181_),
    .D(_0201_),
    .X(_0478_));
 sky130_fd_sc_hd__or4_1 _1197_ (.A(_0051_),
    .B(_0170_),
    .C(_0194_),
    .D(_0210_),
    .X(_0479_));
 sky130_fd_sc_hd__or3_1 _1198_ (.A(_0299_),
    .B(_0478_),
    .C(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__or3_1 _1199_ (.A(_0476_),
    .B(_0477_),
    .C(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__or4_1 _1200_ (.A(_0109_),
    .B(_0277_),
    .C(_0474_),
    .D(_0475_),
    .X(_0482_));
 sky130_fd_sc_hd__or4_1 _1201_ (.A(_0032_),
    .B(_0036_),
    .C(_0104_),
    .D(_0105_),
    .X(_0483_));
 sky130_fd_sc_hd__or3_1 _1202_ (.A(_0204_),
    .B(_0312_),
    .C(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__or4_1 _1203_ (.A(_0272_),
    .B(_0365_),
    .C(_0460_),
    .D(_0473_),
    .X(_0485_));
 sky130_fd_sc_hd__or4_1 _1204_ (.A(_0469_),
    .B(_0482_),
    .C(_0484_),
    .D(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__o32a_1 _1205_ (.A1(net45),
    .A2(_0481_),
    .A3(_0486_),
    .B1(net142),
    .B2(net136),
    .X(_0010_));
 sky130_fd_sc_hd__or3_1 _1206_ (.A(_0135_),
    .B(_0141_),
    .C(_0430_),
    .X(_0487_));
 sky130_fd_sc_hd__or3_1 _1207_ (.A(_0057_),
    .B(_0058_),
    .C(_0164_),
    .X(_0488_));
 sky130_fd_sc_hd__or4_2 _1208_ (.A(_0136_),
    .B(_0250_),
    .C(_0252_),
    .D(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__or2_1 _1209_ (.A(_0072_),
    .B(_0075_),
    .X(_0490_));
 sky130_fd_sc_hd__or2_1 _1210_ (.A(net135),
    .B(_0118_),
    .X(_0491_));
 sky130_fd_sc_hd__or4_1 _1211_ (.A(_0469_),
    .B(_0470_),
    .C(_0487_),
    .D(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__or4_1 _1212_ (.A(_0040_),
    .B(_0123_),
    .C(_0212_),
    .D(_0236_),
    .X(_0493_));
 sky130_fd_sc_hd__or3_1 _1213_ (.A(_0288_),
    .B(_0291_),
    .C(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__or4_1 _1214_ (.A(_0049_),
    .B(_0102_),
    .C(_0270_),
    .D(_0282_),
    .X(_0495_));
 sky130_fd_sc_hd__or4_2 _1215_ (.A(_0235_),
    .B(_0492_),
    .C(_0494_),
    .D(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__or4_1 _1216_ (.A(_0189_),
    .B(_0371_),
    .C(_0428_),
    .D(_0490_),
    .X(_0497_));
 sky130_fd_sc_hd__or3_1 _1217_ (.A(_0705_),
    .B(_0711_),
    .C(_0301_),
    .X(_0498_));
 sky130_fd_sc_hd__or4_1 _1218_ (.A(_0068_),
    .B(_0268_),
    .C(_0307_),
    .D(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__or4_1 _1219_ (.A(_0166_),
    .B(_0489_),
    .C(_0497_),
    .D(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__o32a_1 _1220_ (.A1(net43),
    .A2(_0496_),
    .A3(_0500_),
    .B1(net152),
    .B2(net138),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _1221_ (.A(_0707_),
    .B(_0237_),
    .X(_0501_));
 sky130_fd_sc_hd__or2_1 _1222_ (.A(_0104_),
    .B(_0290_),
    .X(_0502_));
 sky130_fd_sc_hd__or3_1 _1223_ (.A(_0094_),
    .B(_0270_),
    .C(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__or4_1 _1224_ (.A(_0390_),
    .B(_0458_),
    .C(_0490_),
    .D(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__or4_1 _1225_ (.A(_0099_),
    .B(_0127_),
    .C(_0157_),
    .D(_0179_),
    .X(_0505_));
 sky130_fd_sc_hd__or4_1 _1226_ (.A(_0138_),
    .B(_0241_),
    .C(_0254_),
    .D(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__or4_1 _1227_ (.A(_0116_),
    .B(_0161_),
    .C(_0300_),
    .D(_0349_),
    .X(_0507_));
 sky130_fd_sc_hd__or4_1 _1228_ (.A(_0336_),
    .B(_0470_),
    .C(_0501_),
    .D(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__or3_1 _1229_ (.A(_0504_),
    .B(_0506_),
    .C(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__or3_1 _1230_ (.A(_0306_),
    .B(_0407_),
    .C(_0445_),
    .X(_0510_));
 sky130_fd_sc_hd__o32a_1 _1231_ (.A1(net43),
    .A2(_0509_),
    .A3(_0510_),
    .B1(net141),
    .B2(net138),
    .X(_0012_));
 sky130_fd_sc_hd__or4_1 _1232_ (.A(_0693_),
    .B(_0696_),
    .C(_0130_),
    .D(_0192_),
    .X(_0511_));
 sky130_fd_sc_hd__or4_2 _1233_ (.A(_0094_),
    .B(_0095_),
    .C(_0261_),
    .D(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__or2_1 _1234_ (.A(_0107_),
    .B(_0225_),
    .X(_0513_));
 sky130_fd_sc_hd__or2_2 _1235_ (.A(_0090_),
    .B(_0161_),
    .X(_0514_));
 sky130_fd_sc_hd__or4_1 _1236_ (.A(_0119_),
    .B(_0199_),
    .C(_0209_),
    .D(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__or2_1 _1237_ (.A(_0037_),
    .B(_0134_),
    .X(_0516_));
 sky130_fd_sc_hd__or4_1 _1238_ (.A(_0168_),
    .B(_0265_),
    .C(_0305_),
    .D(_0358_),
    .X(_0517_));
 sky130_fd_sc_hd__or4_1 _1239_ (.A(_0178_),
    .B(_0181_),
    .C(_0336_),
    .D(_0502_),
    .X(_0518_));
 sky130_fd_sc_hd__or4_1 _1240_ (.A(_0512_),
    .B(_0516_),
    .C(_0517_),
    .D(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__or4_1 _1241_ (.A(_0079_),
    .B(_0253_),
    .C(_0348_),
    .D(_0413_),
    .X(_0520_));
 sky130_fd_sc_hd__or4_1 _1242_ (.A(_0214_),
    .B(_0223_),
    .C(_0244_),
    .D(_0513_),
    .X(_0521_));
 sky130_fd_sc_hd__or4_1 _1243_ (.A(_0086_),
    .B(_0109_),
    .C(_0292_),
    .D(_0295_),
    .X(_0522_));
 sky130_fd_sc_hd__or4_1 _1244_ (.A(_0188_),
    .B(_0231_),
    .C(_0521_),
    .D(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__or3_1 _1245_ (.A(_0515_),
    .B(_0520_),
    .C(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__o32a_1 _1246_ (.A1(net44),
    .A2(_0519_),
    .A3(_0524_),
    .B1(net156),
    .B2(net139),
    .X(_0013_));
 sky130_fd_sc_hd__or3_2 _1247_ (.A(_0701_),
    .B(_0202_),
    .C(_0203_),
    .X(_0525_));
 sky130_fd_sc_hd__or3_1 _1248_ (.A(_0240_),
    .B(_0245_),
    .C(_0501_),
    .X(_0526_));
 sky130_fd_sc_hd__or4_1 _1249_ (.A(_0040_),
    .B(_0094_),
    .C(_0272_),
    .D(_0389_),
    .X(_0527_));
 sky130_fd_sc_hd__or4_1 _1250_ (.A(_0693_),
    .B(_0221_),
    .C(_0274_),
    .D(_0285_),
    .X(_0528_));
 sky130_fd_sc_hd__or4_1 _1251_ (.A(_0069_),
    .B(_0149_),
    .C(_0297_),
    .D(_0491_),
    .X(_0529_));
 sky130_fd_sc_hd__or4_1 _1252_ (.A(_0487_),
    .B(_0489_),
    .C(_0527_),
    .D(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__or4_1 _1253_ (.A(_0191_),
    .B(_0193_),
    .C(_0234_),
    .D(_0405_),
    .X(_0531_));
 sky130_fd_sc_hd__or4_1 _1254_ (.A(_0051_),
    .B(_0075_),
    .C(_0213_),
    .D(_0268_),
    .X(_0532_));
 sky130_fd_sc_hd__or4_1 _1255_ (.A(_0231_),
    .B(_0528_),
    .C(_0531_),
    .D(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__or4_1 _1256_ (.A(_0471_),
    .B(_0525_),
    .C(_0526_),
    .D(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__o32a_1 _1257_ (.A1(net45),
    .A2(_0530_),
    .A3(_0534_),
    .B1(net143),
    .B2(net137),
    .X(_0014_));
 sky130_fd_sc_hd__or3_1 _1258_ (.A(_0281_),
    .B(_0293_),
    .C(_0385_),
    .X(_0535_));
 sky130_fd_sc_hd__or4_1 _1259_ (.A(_0033_),
    .B(_0052_),
    .C(_0053_),
    .D(_0089_),
    .X(_0536_));
 sky130_fd_sc_hd__or3_1 _1260_ (.A(_0248_),
    .B(_0249_),
    .C(_0274_),
    .X(_0537_));
 sky130_fd_sc_hd__or4_1 _1261_ (.A(_0189_),
    .B(_0228_),
    .C(_0536_),
    .D(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__or3_1 _1262_ (.A(_0527_),
    .B(_0535_),
    .C(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__or2_1 _1263_ (.A(_0158_),
    .B(_0286_),
    .X(_0540_));
 sky130_fd_sc_hd__or4_1 _1264_ (.A(_0373_),
    .B(_0405_),
    .C(_0430_),
    .D(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__or4_1 _1265_ (.A(_0295_),
    .B(_0327_),
    .C(_0411_),
    .D(_0412_),
    .X(_0542_));
 sky130_fd_sc_hd__or4_1 _1266_ (.A(_0113_),
    .B(_0205_),
    .C(_0290_),
    .D(_0297_),
    .X(_0543_));
 sky130_fd_sc_hd__or2_1 _1267_ (.A(_0114_),
    .B(_0130_),
    .X(_0544_));
 sky130_fd_sc_hd__or4_1 _1268_ (.A(_0431_),
    .B(_0474_),
    .C(_0475_),
    .D(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__or4_1 _1269_ (.A(_0337_),
    .B(_0542_),
    .C(_0543_),
    .D(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__or3_1 _1270_ (.A(_0539_),
    .B(_0541_),
    .C(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__o22a_1 _1271_ (.A1(net137),
    .A2(net150),
    .B1(net42),
    .B2(_0547_),
    .X(_0015_));
 sky130_fd_sc_hd__or4_1 _1272_ (.A(_0215_),
    .B(_0248_),
    .C(_0251_),
    .D(_0283_),
    .X(_0548_));
 sky130_fd_sc_hd__or3_1 _1273_ (.A(_0100_),
    .B(_0178_),
    .C(_0181_),
    .X(_0549_));
 sky130_fd_sc_hd__or2_1 _1274_ (.A(_0125_),
    .B(_0229_),
    .X(_0550_));
 sky130_fd_sc_hd__or4_1 _1275_ (.A(_0267_),
    .B(_0275_),
    .C(_0285_),
    .D(_0471_),
    .X(_0551_));
 sky130_fd_sc_hd__or4_1 _1276_ (.A(_0391_),
    .B(_0409_),
    .C(_0449_),
    .D(_0548_),
    .X(_0552_));
 sky130_fd_sc_hd__or4_1 _1277_ (.A(_0135_),
    .B(_0172_),
    .C(_0232_),
    .D(_0247_),
    .X(_0553_));
 sky130_fd_sc_hd__or4_1 _1278_ (.A(_0369_),
    .B(_0429_),
    .C(_0491_),
    .D(_0550_),
    .X(_0554_));
 sky130_fd_sc_hd__or4_1 _1279_ (.A(_0130_),
    .B(_0140_),
    .C(_0166_),
    .D(_0203_),
    .X(_0555_));
 sky130_fd_sc_hd__or4_1 _1280_ (.A(_0069_),
    .B(_0074_),
    .C(_0093_),
    .D(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__or4_1 _1281_ (.A(_0370_),
    .B(_0553_),
    .C(_0554_),
    .D(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__or4_1 _1282_ (.A(_0549_),
    .B(_0551_),
    .C(_0552_),
    .D(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__o22a_1 _1283_ (.A1(net138),
    .A2(net164),
    .B1(net43),
    .B2(_0558_),
    .X(_0016_));
 sky130_fd_sc_hd__or3_1 _1284_ (.A(_0075_),
    .B(_0081_),
    .C(_0082_),
    .X(_0559_));
 sky130_fd_sc_hd__or3_1 _1285_ (.A(_0098_),
    .B(_0174_),
    .C(_0473_),
    .X(_0560_));
 sky130_fd_sc_hd__or2_1 _1286_ (.A(_0647_),
    .B(_0044_),
    .X(_0561_));
 sky130_fd_sc_hd__or4_1 _1287_ (.A(_0275_),
    .B(_0277_),
    .C(_0559_),
    .D(_0560_),
    .X(_0562_));
 sky130_fd_sc_hd__or4_1 _1288_ (.A(_0058_),
    .B(_0129_),
    .C(_0167_),
    .D(_0202_),
    .X(_0563_));
 sky130_fd_sc_hd__or4_1 _1289_ (.A(_0096_),
    .B(_0243_),
    .C(_0514_),
    .D(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__or4_1 _1290_ (.A(_0126_),
    .B(_0309_),
    .C(_0312_),
    .D(_0429_),
    .X(_0565_));
 sky130_fd_sc_hd__or3_1 _1291_ (.A(_0502_),
    .B(_0544_),
    .C(_0561_),
    .X(_0566_));
 sky130_fd_sc_hd__or4_1 _1292_ (.A(_0325_),
    .B(_0516_),
    .C(_0565_),
    .D(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__or4_1 _1293_ (.A(_0049_),
    .B(_0118_),
    .C(_0120_),
    .D(_0212_),
    .X(_0568_));
 sky130_fd_sc_hd__or3_1 _1294_ (.A(_0696_),
    .B(_0156_),
    .C(_0280_),
    .X(_0569_));
 sky130_fd_sc_hd__or4_1 _1295_ (.A(_0301_),
    .B(_0540_),
    .C(_0568_),
    .D(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__or4_1 _1296_ (.A(_0562_),
    .B(_0564_),
    .C(_0567_),
    .D(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__o22a_1 _1297_ (.A1(net136),
    .A2(net167),
    .B1(net42),
    .B2(_0571_),
    .X(_0017_));
 sky130_fd_sc_hd__or3_2 _1298_ (.A(_0137_),
    .B(_0140_),
    .C(_0142_),
    .X(_0572_));
 sky130_fd_sc_hd__or2_1 _1299_ (.A(_0113_),
    .B(_0214_),
    .X(_0573_));
 sky130_fd_sc_hd__or4_1 _1300_ (.A(_0088_),
    .B(_0125_),
    .C(_0134_),
    .D(_0225_),
    .X(_0574_));
 sky130_fd_sc_hd__or4_1 _1301_ (.A(_0076_),
    .B(_0090_),
    .C(_0181_),
    .D(_0264_),
    .X(_0575_));
 sky130_fd_sc_hd__or4_1 _1302_ (.A(_0101_),
    .B(_0262_),
    .C(_0574_),
    .D(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__or4_1 _1303_ (.A(_0180_),
    .B(_0288_),
    .C(_0305_),
    .D(_0308_),
    .X(_0577_));
 sky130_fd_sc_hd__or4_1 _1304_ (.A(_0165_),
    .B(_0171_),
    .C(_0219_),
    .D(_0250_),
    .X(_0578_));
 sky130_fd_sc_hd__or4_1 _1305_ (.A(_0158_),
    .B(_0576_),
    .C(_0577_),
    .D(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__or4_1 _1306_ (.A(_0503_),
    .B(_0572_),
    .C(_0573_),
    .D(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__or4_1 _1307_ (.A(_0054_),
    .B(_0072_),
    .C(_0074_),
    .D(_0394_),
    .X(_0581_));
 sky130_fd_sc_hd__or4_1 _1308_ (.A(_0195_),
    .B(_0393_),
    .C(_0501_),
    .D(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__o32a_1 _1309_ (.A1(net43),
    .A2(_0580_),
    .A3(_0582_),
    .B1(net145),
    .B2(net138),
    .X(_0018_));
 sky130_fd_sc_hd__or4_1 _1310_ (.A(_0106_),
    .B(_0273_),
    .C(_0310_),
    .D(_0332_),
    .X(_0583_));
 sky130_fd_sc_hd__or4_1 _1311_ (.A(_0114_),
    .B(_0197_),
    .C(_0232_),
    .D(_0245_),
    .X(_0584_));
 sky130_fd_sc_hd__or4_1 _1312_ (.A(_0085_),
    .B(_0089_),
    .C(_0229_),
    .D(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__or4_1 _1313_ (.A(_0056_),
    .B(_0243_),
    .C(_0583_),
    .D(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__or3_1 _1314_ (.A(_0175_),
    .B(_0354_),
    .C(_0430_),
    .X(_0587_));
 sky130_fd_sc_hd__or4_1 _1315_ (.A(_0299_),
    .B(_0387_),
    .C(_0424_),
    .D(_0513_),
    .X(_0588_));
 sky130_fd_sc_hd__or4_1 _1316_ (.A(_0043_),
    .B(_0044_),
    .C(_0209_),
    .D(_0327_),
    .X(_0589_));
 sky130_fd_sc_hd__or4_1 _1317_ (.A(_0083_),
    .B(_0351_),
    .C(_0588_),
    .D(_0589_),
    .X(_0590_));
 sky130_fd_sc_hd__or3_1 _1318_ (.A(_0586_),
    .B(_0587_),
    .C(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__o22a_1 _1319_ (.A1(net139),
    .A2(net158),
    .B1(net44),
    .B2(_0591_),
    .X(_0019_));
 sky130_fd_sc_hd__or4_1 _1320_ (.A(_0074_),
    .B(_0076_),
    .C(_0221_),
    .D(_0244_),
    .X(_0592_));
 sky130_fd_sc_hd__or4_1 _1321_ (.A(_0201_),
    .B(_0231_),
    .C(_0366_),
    .D(_0548_),
    .X(_0593_));
 sky130_fd_sc_hd__or2_1 _1322_ (.A(_0096_),
    .B(_0193_),
    .X(_0594_));
 sky130_fd_sc_hd__or4_1 _1323_ (.A(_0267_),
    .B(_0390_),
    .C(_0572_),
    .D(_0592_),
    .X(_0595_));
 sky130_fd_sc_hd__or4_1 _1324_ (.A(_0091_),
    .B(_0171_),
    .C(_0233_),
    .D(_0349_),
    .X(_0596_));
 sky130_fd_sc_hd__or4_1 _1325_ (.A(_0647_),
    .B(_0082_),
    .C(_0098_),
    .D(_0156_),
    .X(_0597_));
 sky130_fd_sc_hd__or4_1 _1326_ (.A(_0054_),
    .B(_0178_),
    .C(_0181_),
    .D(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__or4_1 _1327_ (.A(_0141_),
    .B(_0203_),
    .C(_0238_),
    .D(_0262_),
    .X(_0599_));
 sky130_fd_sc_hd__or4_1 _1328_ (.A(_0594_),
    .B(_0596_),
    .C(_0598_),
    .D(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__or3_1 _1329_ (.A(_0593_),
    .B(_0595_),
    .C(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__o22a_1 _1330_ (.A1(net138),
    .A2(net168),
    .B1(net43),
    .B2(_0601_),
    .X(_0020_));
 sky130_fd_sc_hd__or2_1 _1331_ (.A(_0647_),
    .B(_0251_),
    .X(_0602_));
 sky130_fd_sc_hd__or2_1 _1332_ (.A(_0095_),
    .B(_0264_),
    .X(_0603_));
 sky130_fd_sc_hd__or2_1 _1333_ (.A(_0065_),
    .B(_0258_),
    .X(_0604_));
 sky130_fd_sc_hd__or3_1 _1334_ (.A(_0087_),
    .B(_0109_),
    .C(_0277_),
    .X(_0605_));
 sky130_fd_sc_hd__or4_1 _1335_ (.A(_0710_),
    .B(_0080_),
    .C(_0123_),
    .D(_0187_),
    .X(_0606_));
 sky130_fd_sc_hd__or4_1 _1336_ (.A(_0573_),
    .B(_0602_),
    .C(_0604_),
    .D(_0605_),
    .X(_0607_));
 sky130_fd_sc_hd__or2_1 _1337_ (.A(_0514_),
    .B(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__or4_1 _1338_ (.A(_0097_),
    .B(_0156_),
    .C(_0416_),
    .D(_0603_),
    .X(_0609_));
 sky130_fd_sc_hd__or4_1 _1339_ (.A(_0200_),
    .B(_0385_),
    .C(_0404_),
    .D(_0412_),
    .X(_0610_));
 sky130_fd_sc_hd__or4_1 _1340_ (.A(_0338_),
    .B(_0516_),
    .C(_0609_),
    .D(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__or3_1 _1341_ (.A(_0244_),
    .B(_0245_),
    .C(_0294_),
    .X(_0612_));
 sky130_fd_sc_hd__or4_1 _1342_ (.A(_0194_),
    .B(_0205_),
    .C(_0357_),
    .D(_0488_),
    .X(_0613_));
 sky130_fd_sc_hd__or3_1 _1343_ (.A(_0157_),
    .B(_0266_),
    .C(_0297_),
    .X(_0614_));
 sky130_fd_sc_hd__or4_1 _1344_ (.A(_0078_),
    .B(_0606_),
    .C(_0613_),
    .D(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__or3_1 _1345_ (.A(_0611_),
    .B(_0612_),
    .C(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__o32a_1 _1346_ (.A1(net43),
    .A2(_0608_),
    .A3(_0616_),
    .B1(net170),
    .B2(net138),
    .X(_0021_));
 sky130_fd_sc_hd__or3_1 _1347_ (.A(_0129_),
    .B(_0193_),
    .C(_0525_),
    .X(_0617_));
 sky130_fd_sc_hd__or4_1 _1348_ (.A(_0091_),
    .B(_0333_),
    .C(_0372_),
    .D(_0432_),
    .X(_0618_));
 sky130_fd_sc_hd__or4_1 _1349_ (.A(_0278_),
    .B(_0286_),
    .C(_0472_),
    .D(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__or4_1 _1350_ (.A(_0072_),
    .B(_0074_),
    .C(_0365_),
    .D(_0561_),
    .X(_0620_));
 sky130_fd_sc_hd__or3_1 _1351_ (.A(_0408_),
    .B(_0617_),
    .C(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__or4_1 _1352_ (.A(_0107_),
    .B(_0141_),
    .C(_0142_),
    .D(_0217_),
    .X(_0622_));
 sky130_fd_sc_hd__or4_1 _1353_ (.A(_0081_),
    .B(_0160_),
    .C(_0196_),
    .D(_0292_),
    .X(_0623_));
 sky130_fd_sc_hd__or4_1 _1354_ (.A(_0175_),
    .B(_0367_),
    .C(_0622_),
    .D(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__or4_1 _1355_ (.A(_0331_),
    .B(_0619_),
    .C(_0621_),
    .D(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__o22a_1 _1356_ (.A1(net139),
    .A2(net169),
    .B1(net44),
    .B2(_0625_),
    .X(_0022_));
 sky130_fd_sc_hd__or4_1 _1357_ (.A(_0114_),
    .B(_0122_),
    .C(_0167_),
    .D(_0197_),
    .X(_0626_));
 sky130_fd_sc_hd__or4_1 _1358_ (.A(_0234_),
    .B(_0242_),
    .C(_0458_),
    .D(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__or4_1 _1359_ (.A(_0079_),
    .B(_0159_),
    .C(_0279_),
    .D(_0617_),
    .X(_0628_));
 sky130_fd_sc_hd__or4_1 _1360_ (.A(_0119_),
    .B(_0208_),
    .C(_0404_),
    .D(_0561_),
    .X(_0629_));
 sky130_fd_sc_hd__or4_1 _1361_ (.A(_0040_),
    .B(_0121_),
    .C(_0124_),
    .D(_0245_),
    .X(_0630_));
 sky130_fd_sc_hd__or4_1 _1362_ (.A(_0051_),
    .B(_0265_),
    .C(_0629_),
    .D(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__or4_1 _1363_ (.A(_0058_),
    .B(_0174_),
    .C(_0214_),
    .D(_0298_),
    .X(_0632_));
 sky130_fd_sc_hd__or4_1 _1364_ (.A(_0063_),
    .B(_0258_),
    .C(_0292_),
    .D(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__or3_1 _1365_ (.A(_0092_),
    .B(_0313_),
    .C(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__or3_1 _1366_ (.A(_0627_),
    .B(_0631_),
    .C(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__o32a_1 _1367_ (.A1(net42),
    .A2(_0628_),
    .A3(_0635_),
    .B1(net159),
    .B2(net136),
    .X(_0023_));
 sky130_fd_sc_hd__or3_1 _1368_ (.A(_0119_),
    .B(_0180_),
    .C(_0210_),
    .X(_0636_));
 sky130_fd_sc_hd__or4_1 _1369_ (.A(_0131_),
    .B(_0192_),
    .C(_0335_),
    .D(_0415_),
    .X(_0637_));
 sky130_fd_sc_hd__or4_1 _1370_ (.A(_0033_),
    .B(_0036_),
    .C(_0044_),
    .D(_0222_),
    .X(_0638_));
 sky130_fd_sc_hd__or4_1 _1371_ (.A(_0215_),
    .B(_0308_),
    .C(_0637_),
    .D(_0638_),
    .X(_0639_));
 sky130_fd_sc_hd__or4_1 _1372_ (.A(_0693_),
    .B(_0052_),
    .C(_0063_),
    .D(_0104_),
    .X(_0640_));
 sky130_fd_sc_hd__or4_1 _1373_ (.A(_0162_),
    .B(_0203_),
    .C(_0305_),
    .D(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__or3_1 _1374_ (.A(_0560_),
    .B(_0605_),
    .C(_0636_),
    .X(_0642_));
 sky130_fd_sc_hd__or4_1 _1375_ (.A(_0526_),
    .B(_0639_),
    .C(_0641_),
    .D(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__or4_1 _1376_ (.A(_0094_),
    .B(_0137_),
    .C(_0142_),
    .D(_0270_),
    .X(_0644_));
 sky130_fd_sc_hd__or4_1 _1377_ (.A(_0200_),
    .B(_0228_),
    .C(_0231_),
    .D(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__or2_1 _1378_ (.A(_0425_),
    .B(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__o32a_1 _1379_ (.A1(net43),
    .A2(_0643_),
    .A3(_0646_),
    .B1(net149),
    .B2(net139),
    .X(_0024_));
 sky130_fd_sc_hd__or3_1 _1380_ (.A(_0119_),
    .B(_0209_),
    .C(_0426_),
    .X(_0648_));
 sky130_fd_sc_hd__or4_1 _1381_ (.A(_0549_),
    .B(_0559_),
    .C(_0572_),
    .D(_0602_),
    .X(_0649_));
 sky130_fd_sc_hd__or3_1 _1382_ (.A(_0391_),
    .B(_0427_),
    .C(_0512_),
    .X(_0650_));
 sky130_fd_sc_hd__or4_1 _1383_ (.A(_0190_),
    .B(_0198_),
    .C(_0388_),
    .D(_0648_),
    .X(_0651_));
 sky130_fd_sc_hd__or3_1 _1384_ (.A(_0068_),
    .B(_0069_),
    .C(_0283_),
    .X(_0652_));
 sky130_fd_sc_hd__or4_1 _1385_ (.A(_0704_),
    .B(_0171_),
    .C(_0203_),
    .D(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__or4_1 _1386_ (.A(_0164_),
    .B(_0166_),
    .C(_0356_),
    .D(_0550_),
    .X(_0654_));
 sky130_fd_sc_hd__or4_1 _1387_ (.A(_0649_),
    .B(_0651_),
    .C(_0653_),
    .D(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__o32a_1 _1388_ (.A1(net43),
    .A2(_0650_),
    .A3(_0655_),
    .B1(net171),
    .B2(net139),
    .X(_0025_));
 sky130_fd_sc_hd__or4_1 _1389_ (.A(_0098_),
    .B(_0176_),
    .C(_0296_),
    .D(_0297_),
    .X(_0656_));
 sky130_fd_sc_hd__or4_1 _1390_ (.A(_0166_),
    .B(_0489_),
    .C(_0592_),
    .D(_0656_),
    .X(_0658_));
 sky130_fd_sc_hd__or3_1 _1391_ (.A(_0226_),
    .B(_0473_),
    .C(_0603_),
    .X(_0659_));
 sky130_fd_sc_hd__or3_1 _1392_ (.A(_0209_),
    .B(_0230_),
    .C(_0281_),
    .X(_0660_));
 sky130_fd_sc_hd__or4_1 _1393_ (.A(_0102_),
    .B(_0103_),
    .C(_0241_),
    .D(_0308_),
    .X(_0661_));
 sky130_fd_sc_hd__or4_1 _1394_ (.A(_0149_),
    .B(_0326_),
    .C(_0660_),
    .D(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__or4_1 _1395_ (.A(_0705_),
    .B(_0203_),
    .C(_0275_),
    .D(_0277_),
    .X(_0663_));
 sky130_fd_sc_hd__or4_1 _1396_ (.A(_0710_),
    .B(_0131_),
    .C(_0282_),
    .D(_0285_),
    .X(_0664_));
 sky130_fd_sc_hd__or4_1 _1397_ (.A(_0430_),
    .B(_0573_),
    .C(_0663_),
    .D(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__or4_1 _1398_ (.A(_0163_),
    .B(_0659_),
    .C(_0662_),
    .D(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__o32a_1 _1399_ (.A1(net42),
    .A2(_0658_),
    .A3(_0666_),
    .B1(net151),
    .B2(net137),
    .X(_0026_));
 sky130_fd_sc_hd__or4_1 _1400_ (.A(_0077_),
    .B(_0163_),
    .C(_0370_),
    .D(_0392_),
    .X(_0668_));
 sky130_fd_sc_hd__or4_1 _1401_ (.A(_0085_),
    .B(_0157_),
    .C(_0263_),
    .D(_0270_),
    .X(_0669_));
 sky130_fd_sc_hd__or4_1 _1402_ (.A(_0711_),
    .B(_0208_),
    .C(_0248_),
    .D(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__or3_1 _1403_ (.A(_0172_),
    .B(_0243_),
    .C(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__or4_1 _1404_ (.A(_0177_),
    .B(_0386_),
    .C(_0604_),
    .D(_0626_),
    .X(_0672_));
 sky130_fd_sc_hd__or4_1 _1405_ (.A(_0127_),
    .B(_0188_),
    .C(_0213_),
    .D(_0275_),
    .X(_0673_));
 sky130_fd_sc_hd__or4_1 _1406_ (.A(_0226_),
    .B(_0296_),
    .C(_0308_),
    .D(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__or4_1 _1407_ (.A(_0668_),
    .B(_0671_),
    .C(_0672_),
    .D(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__o22a_1 _1408_ (.A1(net136),
    .A2(net161),
    .B1(net42),
    .B2(_0675_),
    .X(_0027_));
 sky130_fd_sc_hd__or4_1 _1409_ (.A(_0201_),
    .B(_0231_),
    .C(_0273_),
    .D(_0296_),
    .X(_0676_));
 sky130_fd_sc_hd__or3_1 _1410_ (.A(_0077_),
    .B(_0370_),
    .C(_0676_),
    .X(_0678_));
 sky130_fd_sc_hd__or3_1 _1411_ (.A(_0115_),
    .B(_0130_),
    .C(_0131_),
    .X(_0679_));
 sky130_fd_sc_hd__or4_1 _1412_ (.A(_0040_),
    .B(_0350_),
    .C(_0389_),
    .D(_0525_),
    .X(_0680_));
 sky130_fd_sc_hd__or4_1 _1413_ (.A(_0182_),
    .B(_0226_),
    .C(_0278_),
    .D(_0491_),
    .X(_0681_));
 sky130_fd_sc_hd__or4_1 _1414_ (.A(_0265_),
    .B(_0268_),
    .C(_0679_),
    .D(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__or4_1 _1415_ (.A(_0636_),
    .B(_0678_),
    .C(_0680_),
    .D(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__o32a_1 _1416_ (.A1(_0173_),
    .A2(net42),
    .A3(_0683_),
    .B1(net146),
    .B2(net136),
    .X(_0028_));
 sky130_fd_sc_hd__or3_1 _1417_ (.A(_0191_),
    .B(_0273_),
    .C(_0296_),
    .X(_0684_));
 sky130_fd_sc_hd__or4_1 _1418_ (.A(_0083_),
    .B(_0194_),
    .C(_0283_),
    .D(_0291_),
    .X(_0685_));
 sky130_fd_sc_hd__or4_1 _1419_ (.A(net135),
    .B(_0696_),
    .C(_0159_),
    .D(_0370_),
    .X(_0686_));
 sky130_fd_sc_hd__or4_1 _1420_ (.A(_0183_),
    .B(_0684_),
    .C(_0685_),
    .D(_0686_),
    .X(_0688_));
 sky130_fd_sc_hd__or4_1 _1421_ (.A(_0072_),
    .B(_0201_),
    .C(_0216_),
    .D(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__o32a_1 _1422_ (.A1(_0173_),
    .A2(net42),
    .A3(_0689_),
    .B1(net155),
    .B2(net136),
    .X(_0029_));
 sky130_fd_sc_hd__or4_1 _1423_ (.A(_0108_),
    .B(_0247_),
    .C(_0269_),
    .D(_0299_),
    .X(_0690_));
 sky130_fd_sc_hd__or3_1 _1424_ (.A(_0184_),
    .B(_0207_),
    .C(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__o22a_1 _1425_ (.A1(net136),
    .A2(net153),
    .B1(net42),
    .B2(_0691_),
    .X(_0030_));
 sky130_fd_sc_hd__or2_1 _1426_ (.A(net136),
    .B(net172),
    .X(_0692_));
 sky130_fd_sc_hd__o31a_1 _1427_ (.A1(net135),
    .A2(_0207_),
    .A3(_0257_),
    .B1(_0692_),
    .X(_0031_));
 sky130_fd_sc_hd__dfxtp_1 _1428_ (.CLK(clknet_2_0__leaf_clk0),
    .D(_0000_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_1 _1429_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0001_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_1 _1430_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0002_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _1431_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0003_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _1432_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0004_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _1433_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0005_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _1434_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0006_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _1435_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0007_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _1436_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0008_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _1437_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0009_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _1438_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0010_),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_1 _1439_ (.CLK(clknet_2_0__leaf_clk0),
    .D(_0011_),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_1 _1440_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0012_),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_1 _1441_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0013_),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_1 _1442_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0014_),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_1 _1443_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0015_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_1 _1444_ (.CLK(clknet_2_0__leaf_clk0),
    .D(_0016_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_1 _1445_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0017_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_1 _1446_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0018_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_1 _1447_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0019_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_1 _1448_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0020_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_1 _1449_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0021_),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_1 _1450_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0022_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_1 _1451_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0023_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_1 _1452_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0024_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_1 _1453_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0025_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_1 _1454_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0026_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _1455_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0027_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_1 _1456_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0028_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _1457_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0029_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _1458_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0030_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _1459_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0031_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _1460_ (.CLK(clknet_2_1__leaf_clk0),
    .D(net1),
    .Q(\addr0_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1461_ (.CLK(clknet_2_1__leaf_clk0),
    .D(net2),
    .Q(\addr0_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1462_ (.CLK(clknet_2_1__leaf_clk0),
    .D(net3),
    .Q(\addr0_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1463_ (.CLK(clknet_2_1__leaf_clk0),
    .D(net4),
    .Q(\addr0_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1464_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net5),
    .Q(\addr0_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1465_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net6),
    .Q(\addr0_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1466_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net7),
    .Q(\addr0_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1467_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net8),
    .Q(\addr0_reg[7] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk0 (.A(clk0),
    .X(clknet_0_clk0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_345 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(addr0[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(addr0[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(addr0[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(addr0[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(addr0[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(addr0[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(addr0[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(addr0[7]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(cs0),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(dout0[0]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(dout0[10]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(dout0[11]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(dout0[12]));
 sky130_fd_sc_hd__clkbuf_4 output14 (.A(net14),
    .X(dout0[13]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(dout0[14]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(dout0[15]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(dout0[16]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(dout0[17]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(dout0[18]));
 sky130_fd_sc_hd__clkbuf_4 output20 (.A(net20),
    .X(dout0[19]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(dout0[1]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(dout0[20]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(dout0[21]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(dout0[22]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(dout0[23]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(dout0[24]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(dout0[25]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(dout0[26]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(dout0[27]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(dout0[28]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(dout0[29]));
 sky130_fd_sc_hd__clkbuf_4 output32 (.A(net32),
    .X(dout0[2]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(dout0[30]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(dout0[31]));
 sky130_fd_sc_hd__clkbuf_4 output35 (.A(net35),
    .X(dout0[3]));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net36),
    .X(dout0[4]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(dout0[5]));
 sky130_fd_sc_hd__clkbuf_4 output38 (.A(net38),
    .X(dout0[6]));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net39),
    .X(dout0[7]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(dout0[8]));
 sky130_fd_sc_hd__clkbuf_4 output41 (.A(net41),
    .X(dout0[9]));
 sky130_fd_sc_hd__buf_2 fanout42 (.A(net45),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 fanout45 (.A(_0304_),
    .X(net45));
 sky130_fd_sc_hd__buf_1 wire46 (.A(_0073_),
    .X(net46));
 sky130_fd_sc_hd__buf_2 fanout47 (.A(net48),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 fanout48 (.A(_0071_),
    .X(net48));
 sky130_fd_sc_hd__buf_2 fanout49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 fanout50 (.A(_0070_),
    .X(net50));
 sky130_fd_sc_hd__buf_2 fanout51 (.A(_0067_),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 fanout52 (.A(_0067_),
    .X(net52));
 sky130_fd_sc_hd__buf_2 fanout53 (.A(_0066_),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 fanout54 (.A(_0066_),
    .X(net54));
 sky130_fd_sc_hd__buf_2 fanout55 (.A(net57),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 wire57 (.A(_0062_),
    .X(net57));
 sky130_fd_sc_hd__buf_2 fanout58 (.A(_0061_),
    .X(net58));
 sky130_fd_sc_hd__buf_1 fanout59 (.A(_0061_),
    .X(net59));
 sky130_fd_sc_hd__buf_2 fanout60 (.A(_0048_),
    .X(net60));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout61 (.A(_0048_),
    .X(net61));
 sky130_fd_sc_hd__buf_2 fanout62 (.A(net65),
    .X(net62));
 sky130_fd_sc_hd__buf_1 fanout63 (.A(net64),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 max_cap64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 wire65 (.A(_0047_),
    .X(net65));
 sky130_fd_sc_hd__buf_2 fanout66 (.A(_0042_),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 fanout67 (.A(_0042_),
    .X(net67));
 sky130_fd_sc_hd__buf_2 fanout68 (.A(net70),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 fanout69 (.A(net71),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 wire70 (.A(_0041_),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 max_cap71 (.A(_0041_),
    .X(net71));
 sky130_fd_sc_hd__buf_2 fanout72 (.A(_0039_),
    .X(net72));
 sky130_fd_sc_hd__buf_1 fanout73 (.A(_0039_),
    .X(net73));
 sky130_fd_sc_hd__buf_2 fanout74 (.A(_0038_),
    .X(net74));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout75 (.A(_0038_),
    .X(net75));
 sky130_fd_sc_hd__buf_2 fanout76 (.A(_0035_),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 fanout77 (.A(_0035_),
    .X(net77));
 sky130_fd_sc_hd__buf_2 fanout78 (.A(_0034_),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 fanout79 (.A(_0034_),
    .X(net79));
 sky130_fd_sc_hd__buf_2 fanout80 (.A(net81),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 fanout81 (.A(_0713_),
    .X(net81));
 sky130_fd_sc_hd__buf_2 fanout82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 fanout83 (.A(_0712_),
    .X(net83));
 sky130_fd_sc_hd__buf_2 fanout84 (.A(net86),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 fanout85 (.A(net87),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 wire86 (.A(net88),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 max_cap87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 wire88 (.A(_0709_),
    .X(net88));
 sky130_fd_sc_hd__buf_2 fanout89 (.A(_0708_),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 fanout90 (.A(_0708_),
    .X(net90));
 sky130_fd_sc_hd__buf_2 fanout91 (.A(_0706_),
    .X(net91));
 sky130_fd_sc_hd__buf_1 fanout92 (.A(_0706_),
    .X(net92));
 sky130_fd_sc_hd__buf_2 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 fanout94 (.A(_0703_),
    .X(net94));
 sky130_fd_sc_hd__buf_2 fanout95 (.A(_0700_),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 fanout96 (.A(_0700_),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_4 fanout97 (.A(net100),
    .X(net97));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 max_cap99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 wire100 (.A(_0699_),
    .X(net100));
 sky130_fd_sc_hd__buf_2 fanout101 (.A(net103),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 fanout102 (.A(net104),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 max_cap103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 wire104 (.A(_0698_),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 fanout105 (.A(_0697_),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 fanout106 (.A(_0697_),
    .X(net106));
 sky130_fd_sc_hd__buf_2 fanout107 (.A(_0695_),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 fanout108 (.A(_0695_),
    .X(net108));
 sky130_fd_sc_hd__buf_2 fanout109 (.A(_0694_),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 fanout110 (.A(_0694_),
    .X(net110));
 sky130_fd_sc_hd__buf_2 fanout111 (.A(_0687_),
    .X(net111));
 sky130_fd_sc_hd__buf_1 fanout112 (.A(_0687_),
    .X(net112));
 sky130_fd_sc_hd__buf_2 fanout113 (.A(_0677_),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 fanout114 (.A(_0677_),
    .X(net114));
 sky130_fd_sc_hd__buf_2 fanout115 (.A(_0667_),
    .X(net115));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout116 (.A(_0667_),
    .X(net116));
 sky130_fd_sc_hd__buf_2 fanout117 (.A(_0657_),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 fanout118 (.A(_0657_),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 fanout119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout120 (.A(\addr0_reg[7] ),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 fanout121 (.A(\addr0_reg[6] ),
    .X(net121));
 sky130_fd_sc_hd__buf_1 fanout122 (.A(\addr0_reg[6] ),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 fanout123 (.A(\addr0_reg[5] ),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 fanout124 (.A(\addr0_reg[5] ),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 fanout125 (.A(\addr0_reg[4] ),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 fanout126 (.A(\addr0_reg[4] ),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 fanout127 (.A(\addr0_reg[3] ),
    .X(net127));
 sky130_fd_sc_hd__buf_1 fanout128 (.A(\addr0_reg[3] ),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 fanout129 (.A(\addr0_reg[2] ),
    .X(net129));
 sky130_fd_sc_hd__buf_1 fanout130 (.A(\addr0_reg[2] ),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 fanout131 (.A(\addr0_reg[1] ),
    .X(net131));
 sky130_fd_sc_hd__buf_1 fanout132 (.A(\addr0_reg[1] ),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 fanout133 (.A(\addr0_reg[0] ),
    .X(net133));
 sky130_fd_sc_hd__buf_1 fanout134 (.A(\addr0_reg[0] ),
    .X(net134));
 sky130_fd_sc_hd__buf_2 fanout135 (.A(_0647_),
    .X(net135));
 sky130_fd_sc_hd__buf_2 fanout136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 fanout137 (.A(net9),
    .X(net137));
 sky130_fd_sc_hd__buf_2 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__buf_2 fanout139 (.A(net9),
    .X(net139));
 sky130_fd_sc_hd__conb_1 cust_rom_140 (.LO(net140));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_0__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_1__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_2__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_3__leaf_clk0));
 sky130_fd_sc_hd__clkinv_4 clkload0 (.A(clknet_2_0__leaf_clk0));
 sky130_fd_sc_hd__bufinv_16 clkload1 (.A(clknet_2_1__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_8 clkload2 (.A(clknet_2_3__leaf_clk0));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net13),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net11),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net15),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net10),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net19),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net30),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net40),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net21),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net26),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net16),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net28),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net12),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net33),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net41),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net31),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net14),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net37),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net20),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net25),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net32),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net29),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net35),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net36),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net17),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net38),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net39),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net18),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net22),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net24),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net23),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net27),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net34),
    .X(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0060_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_0082_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_0130_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0132_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_0156_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0215_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_0216_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_0261_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_0267_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_0283_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_0283_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_0292_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_0292_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_0421_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_0441_));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_281 ();
 assign dout0[32] = net140;
endmodule
