* NGSPICE file created from cust_rom0.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

.subckt cust_rom0 addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7]
+ clk0 cs0 dout0[0] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[16]
+ dout0[17] dout0[18] dout0[19] dout0[1] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24]
+ dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[2] dout0[30] dout0[31] dout0[3]
+ dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] vccd1 vssd1
XTAP_TAPCELL_ROW_52_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1270_ net265 net187 net162 net151 vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0985_ net311 net229 vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__or2_2
XFILLER_0_22_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout127 _0220_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_2
Xfanout116 net117 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__buf_1
X_1468_ clknet_2_3__leaf_clk0 _0027_ vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__dfxtp_1
Xfanout105 _0238_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__buf_1
Xfanout149 _0200_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__buf_1
Xfanout138 _0210_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_1
X_1399_ net145 net78 _0265_ _0664_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0770_ net548 net542 net535 net555 vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__a22o_1
X_1322_ net314 net239 net128 net107 vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__or4_1
X_1253_ _0459_ _0474_ _0515_ _0525_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__or4_1
X_1184_ _0265_ _0411_ _0457_ _0458_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_19_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0968_ net501 net371 net364 net492 vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0899_ net405 net346 net517 vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout480 net481 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout491 net493 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_16_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0822_ net429 net421 net414 net436 vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0753_ net585 net577 net600 net592 vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__and4b_1
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1236_ net558 net648 net41 _0510_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__a22o_1
X_1305_ _0569_ _0574_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__or2_1
X_1167_ net125 net118 _0227_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__or3_2
X_1098_ net319 net316 net194 _0380_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1021_ net221 net218 net217 vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0805_ net263 net261 net259 vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0736_ net333 net330 net327 vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__or3_2
X_1219_ _0484_ _0486_ _0493_ _0494_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold30 net16 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_5 _0059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1004_ net199 net198 net112 net105 vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0719_ net600 net585 net578 net592 vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_12_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 dout0[29] sky130_fd_sc_hd__buf_2
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 dout0[19] sky130_fd_sc_hd__buf_2
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout309 net310 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_1
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0984_ net309 net232 vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout128 net129 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_1
Xfanout106 _0238_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__buf_1
X_1467_ clknet_2_3__leaf_clk0 _0026_ vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__dfxtp_1
Xfanout139 _0210_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_1
Xfanout117 _0227_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__buf_1
X_1398_ net223 net135 net134 net117 vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1321_ _0150_ _0294_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__or2_1
X_1252_ net172 net91 net85 vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__or3_1
X_1183_ net290 _0074_ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_19_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0967_ net466 net372 net365 net457 vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0898_ net500 net379 net346 net493 vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout481 net482 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_1
Xfanout470 net472 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_1
Xfanout492 net493 vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__buf_1
XFILLER_0_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0752_ net594 net602 net577 net587 vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0821_ net248 net246 net245 net242 vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1304_ _0485_ _0570_ _0571_ _0573_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__or4_1
X_1235_ _0503_ _0505_ _0507_ _0509_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1166_ _0441_ _0442_ _0443_ _0444_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__or4_1
X_1097_ net255 net236 net234 net139 vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_22_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1020_ net166 net164 net82 vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__or3_2
X_0735_ net557 net486 net478 net544 vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0804_ net545 net402 net397 net532 vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1149_ net322 net316 net315 vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__or3_1
X_1218_ net239 _0112_ _0428_ _0487_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold31 net32 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 net26 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 _0071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Left_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1003_ net112 net105 vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0718_ net614 net620 net626 net607 vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 dout0[2] sky130_fd_sc_hd__clkbuf_4
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 dout0[1] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_33_Left_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput10 net10 vssd1 vssd1 vccd1 vccd1 dout0[0] sky130_fd_sc_hd__buf_2
XFILLER_0_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0983_ _0077_ _0117_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout118 net120 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__buf_1
Xfanout129 net130 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_1
Xfanout107 net109 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__buf_1
X_1397_ _0386_ _0430_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__or2_1
X_1466_ clknet_2_3__leaf_clk0 _0025_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Left_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1320_ _0500_ _0516_ _0555_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__or3_1
X_1182_ net157 _0392_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__or2_1
X_1251_ net561 net634 net44 _0524_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_20_Left_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0897_ net433 net377 net344 net426 vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__a22o_1
X_0966_ net96 net93 net90 _0252_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__or4_1
X_1449_ clknet_2_3__leaf_clk0 _0008_ vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout471 net472 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_1
Xfanout482 _0706_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_1
Xfanout460 net462 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_1
Xfanout493 net494 vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_16_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0751_ net335 net334 _0714_ _0032_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__or4_2
X_0820_ net247 net244 vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__or2_1
X_1303_ net265 net253 _0180_ _0572_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1096_ _0075_ _0308_ _0374_ _0375_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__or4_1
X_1234_ _0126_ net177 _0415_ _0508_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__or4_1
X_1165_ net208 net206 net155 net148 vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__or4_1
X_0949_ net114 net113 net111 net108 vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout290 _0070_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_1
XFILLER_0_16_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0734_ net605 net611 net617 net623 vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0803_ net263 net261 vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1217_ _0489_ _0490_ _0491_ _0492_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__or4_1
X_1148_ net271 net270 net250 net247 vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__or4_1
X_1079_ net227 net197 _0197_ _0362_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__or4_2
XFILLER_0_47_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold10 net28 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 net37 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_7 _0094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1002_ net308 net232 net79 net71 vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__or4_1
XFILLER_0_32_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0717_ net592 net577 net585 net601 vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_35_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput11 net11 vssd1 vssd1 vccd1 vccd1 dout0[10] sky130_fd_sc_hd__buf_2
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 dout0[30] sky130_fd_sc_hd__buf_2
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 dout0[20] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0982_ _0035_ _0038_ _0062_ _0069_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__or4_1
Xfanout119 net120 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_1
Xfanout108 net109 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1465_ clknet_2_2__leaf_clk0 _0024_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__dfxtp_1
X_1396_ _0197_ _0310_ _0374_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout620 net621 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1181_ net279 net269 net263 vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__or3_1
X_1250_ _0517_ _0520_ _0523_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0896_ net448 net377 net344 net440 vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__a22o_1
X_0965_ net517 net366 vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__and2b_1
X_1448_ clknet_2_1__leaf_clk0 _0007_ vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1379_ net308 net231 _0239_ _0284_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__or4_1
XFILLER_0_52_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout472 net473 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_1
Xfanout461 net462 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_1
Xfanout494 net499 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__buf_1
Xfanout483 net484 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__buf_1
Xfanout450 net455 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_16_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0750_ net335 net334 net323 vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__or3_1
Xfanout90 net92 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_1
XFILLER_0_36_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1302_ net310 net211 net189 vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__or3_1
X_1233_ _0037_ net67 _0180_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1095_ _0056_ _0222_ _0376_ _0377_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1164_ net332 net289 net283 vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0948_ net508 net338 net410 vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_30_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0879_ net188 net184 vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout291 _0067_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__buf_1
Xfanout280 _0080_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0802_ net449 net401 net394 net441 vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0733_ net605 net611 net623 net617 vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__and4_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1216_ net66 net58 _0433_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1078_ net209 net202 net91 net69 vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__or4_1
X_1147_ net311 net229 net80 net76 vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold11 net15 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 net22 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_8 _0097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ net227 net225 net181 net180 vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0716_ cs0_reg vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput12 net12 vssd1 vssd1 vccd1 vccd1 dout0[11] sky130_fd_sc_hd__buf_2
Xoutput34 net34 vssd1 vssd1 vccd1 vccd1 dout0[3] sky130_fd_sc_hd__buf_2
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 dout0[21] sky130_fd_sc_hd__buf_2
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0981_ net76 net74 net73 net70 vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_14_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout109 net110 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__buf_1
XFILLER_0_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1464_ clknet_2_3__leaf_clk0 _0023_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__dfxtp_1
X_1395_ _0113_ _0316_ _0460_ _0565_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout621 net622 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_1
Xfanout610 addr0_reg\[3\] vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_5_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1180_ net149 net147 vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__or2_1
X_0964_ net489 net374 net368 net481 vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0895_ net590 net597 net574 net581 vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__and4b_1
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1447_ clknet_2_2__leaf_clk0 _0006_ vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1378_ _0408_ _0641_ _0642_ _0643_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout440 net441 vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_1
Xfanout473 net474 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__buf_1
Xfanout462 net463 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_1
Xfanout451 net452 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_1
Xfanout495 net496 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_1
Xfanout484 net485 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_1
XFILLER_0_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout91 net92 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__buf_1
Xfanout80 _0257_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__buf_1
XFILLER_0_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1232_ _0139_ _0282_ _0501_ _0506_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__or4_1
X_1301_ _0082_ net78 net69 _0563_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1094_ net185 net184 net182 vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__or3_2
X_1163_ net195 net193 net180 net178 vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__or4_1
X_0947_ net512 net429 net339 net436 vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0878_ net528 net360 net353 net519 vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload0 clknet_2_0__leaf_clk0 vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout281 net282 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_1
Xfanout292 _0067_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__buf_1
Xfanout270 _0084_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_1
XFILLER_0_24_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0801_ net433 net401 net394 net426 vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__a22o_1
X_0732_ net332 net329 vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1146_ net295 net293 _0315_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__or3_1
X_1215_ net159 net117 net101 _0306_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1077_ _0086_ _0214_ net60 _0304_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold12 net40 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 net17 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_9 _0103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1000_ net276 net271 net162 _0186_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__or4_1
XFILLER_0_32_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1129_ net227 _0201_ net147 net95 vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput35 net35 vssd1 vssd1 vccd1 vccd1 dout0[4] sky130_fd_sc_hd__buf_2
Xoutput13 net13 vssd1 vssd1 vccd1 vccd1 dout0[12] sky130_fd_sc_hd__buf_2
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 dout0[22] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0980_ net74 net71 vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1463_ clknet_2_2__leaf_clk0 _0022_ vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__dfxtp_1
X_1394_ net560 net650 net43 _0659_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout622 addr0_reg\[1\] vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__buf_1
Xfanout611 net612 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__buf_1
Xfanout600 net601 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_1
XFILLER_0_13_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0963_ net97 net94 vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_27_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0894_ net174 net173 net170 net168 vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1446_ clknet_2_1__leaf_clk0 _0005_ vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1377_ net219 net216 net95 net93 vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout474 _0709_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_1
Xfanout463 net464 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_1
Xfanout430 net431 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_1
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_1
Xfanout441 net442 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_1
Xfanout496 net497 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_1
Xfanout485 net490 vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout81 _0257_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__buf_1
Xfanout70 net71 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
Xfanout92 _0251_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_24_Left_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1231_ _0267_ _0271_ _0342_ _0496_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__or4_1
X_1300_ _0213_ net58 _0477_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1162_ net173 net95 net86 net69 vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_47_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1093_ net163 net82 net81 vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__or3_1
X_0946_ net535 net510 net340 net548 vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0877_ net434 net357 net350 net427 vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__a22o_1
X_1429_ _0191_ _0274_ _0275_ _0683_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_38_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload1 clknet_2_1__leaf_clk0 vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_18_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout282 _0073_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_2
Xfanout293 _0066_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__buf_1
Xfanout271 net272 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_1
Xfanout260 _0091_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_44_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0731_ net557 net503 net495 net544 vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__a22o_1
X_0800_ net525 net407 net399 net518 vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__a22o_1
X_1214_ net67 _0271_ _0341_ _0476_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__or4_1
X_1145_ net562 net651 net45 _0425_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1076_ _0708_ _0357_ _0358_ _0359_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__or4_1
X_0929_ net592 net585 net578 net600 vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_30_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold24 net11 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 net12 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1059_ net220 net216 vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_11_Left_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1128_ net271 _0408_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput36 net36 vssd1 vssd1 vccd1 vccd1 dout0[5] sky130_fd_sc_hd__clkbuf_4
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 dout0[23] sky130_fd_sc_hd__buf_2
Xoutput14 net14 vssd1 vssd1 vccd1 vccd1 dout0[13] sky130_fd_sc_hd__buf_2
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1462_ clknet_2_2__leaf_clk0 _0021_ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1393_ _0653_ _0657_ _0658_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout612 net616 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_1
Xfanout623 net624 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_1
Xfanout601 net602 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0962_ net476 net360 net353 net484 vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__a22o_1
X_0893_ net174 net169 vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__or2_1
X_1445_ clknet_2_3__leaf_clk0 _0004_ vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1376_ net328 net256 net130 net117 vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout464 net465 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_1
Xfanout453 net454 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__buf_1
Xfanout431 net432 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_1
Xfanout497 net498 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__clkbuf_1
Xfanout420 net425 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__clkbuf_1
Xfanout486 net488 vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_1
Xfanout475 net477 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__buf_1
Xfanout442 net447 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_1
Xfanout60 _0303_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_1
XFILLER_0_36_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout82 _0256_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__buf_1
Xfanout71 _0264_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_2
Xfanout93 _0249_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__buf_1
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1161_ net572 net659 net55 _0440_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__a22o_1
X_1092_ net267 _0091_ net175 net168 vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__or4_1
X_1230_ _0371_ _0409_ _0504_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_47_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0945_ net511 net461 net341 net471 vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0876_ net187 net185 vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1428_ net563 net636 net46 _0693_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_38_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1359_ net205 net204 net184 net182 vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_41_Left_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload2 clknet_2_3__leaf_clk0 vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_18_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout294 net295 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_1
Xfanout272 net274 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_2
Xfanout283 net285 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__buf_1
Xfanout261 _0089_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_1
Xfanout250 _0101_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_44_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0730_ net605 net611 net624 net621 vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1213_ net331 net326 _0076_ _0488_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1075_ net298 net294 net292 vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__or3_1
X_1144_ _0409_ _0419_ _0423_ _0424_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__or4_1
X_0859_ net458 net373 net366 net468 vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__a22o_1
X_0928_ net142 net140 net138 net135 vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__or4_2
Xhold14 net23 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 net20 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1058_ net252 net183 vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__or2_1
X_1127_ net276 net275 net268 net265 vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput15 net15 vssd1 vssd1 vccd1 vccd1 dout0[14] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput37 net37 vssd1 vssd1 vccd1 vccd1 dout0[6] sky130_fd_sc_hd__buf_2
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 dout0[24] sky130_fd_sc_hd__buf_2
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1461_ clknet_2_2__leaf_clk0 _0020_ vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1392_ _0554_ _0564_ _0577_ _0627_ vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout613 net616 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_1
Xfanout624 net629 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__buf_1
Xfanout602 net603 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_5_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0961_ net456 net359 net352 net467 vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0892_ net172 net170 vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1444_ clknet_2_1__leaf_clk0 _0003_ vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__dfxtp_1
X_1375_ net246 net213 net201 net150 vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_2_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout432 _0031_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__buf_1
Xfanout443 net444 vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_1
Xfanout410 _0050_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__buf_1
Xfanout421 net424 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_1
Xfanout498 net499 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_1
Xfanout454 net455 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_1
Xfanout487 net488 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_1
Xfanout476 net477 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_1
XFILLER_0_51_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout50 net52 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_1
Xfanout61 _0206_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_24_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout94 _0249_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_1
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout72 _0263_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__buf_1
Xfanout83 _0256_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_1
X_1160_ _0434_ _0438_ _0439_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__or3_1
X_1091_ net228 net214 net211 vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__or3_2
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0944_ net128 net125 net119 net116 vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_47_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0875_ net545 net356 net349 net532 vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__a22o_1
X_1427_ _0683_ _0692_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__or2_1
X_1358_ _0107_ _0213_ _0305_ _0432_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_38_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1289_ net289 net160 net80 _0559_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout240 net241 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_1
Xfanout273 net274 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_1
Xfanout284 net285 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_1
Xfanout295 net296 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_1
Xfanout251 net252 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_1
Xfanout262 _0089_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_1
X_1212_ net213 net171 net169 net142 vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_35_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1143_ net248 net242 _0158_ _0410_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__or4_1
X_1074_ net162 net160 net159 vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__or3_1
X_0927_ net143 net137 net136 vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0789_ net289 net282 vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__or2_1
X_0858_ _0143_ net200 vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__or2_1
Xhold26 net36 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 net29 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1126_ net59 _0406_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__or2_1
X_1057_ net332 net299 vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput38 net38 vssd1 vssd1 vccd1 vccd1 dout0[7] sky130_fd_sc_hd__clkbuf_4
Xoutput16 net16 vssd1 vssd1 vccd1 vccd1 dout0[15] sky130_fd_sc_hd__clkbuf_4
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 dout0[25] sky130_fd_sc_hd__buf_2
Xclkbuf_2_3__f_clk0 clknet_0_clk0 vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1109_ net312 net306 vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1391_ _0157_ _0292_ _0654_ _0656_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__or4_1
X_1460_ clknet_2_2__leaf_clk0 _0019_ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout625 net629 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_1
Xfanout614 net615 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_1
Xfanout603 net604 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_5_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0960_ net100 net99 vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__or2_1
X_0891_ net528 net374 net367 net521 vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__a22o_1
X_1443_ clknet_2_1__leaf_clk0 _0002_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__dfxtp_1
X_1374_ net64 net158 _0376_ _0487_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_2_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout422 net424 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_1
Xfanout411 net413 vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_1
Xfanout400 _0079_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_1
Xfanout455 _0712_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_1
Xfanout499 _0702_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_1
Xfanout444 net445 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_1
Xfanout488 net489 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_1
Xfanout477 net482 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_1
Xfanout433 net435 vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_1
Xfanout466 net467 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_1
Xfanout51 net52 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
Xfanout62 _0194_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__buf_1
Xfanout73 _0263_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout84 net85 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__buf_1
Xfanout95 net97 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__buf_1
X_1090_ _0140_ net61 vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0943_ net127 net116 vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__or2_1
X_0874_ net449 net356 net349 net441 vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1426_ _0133_ _0269_ _0687_ _0691_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__or4_1
X_1288_ _0714_ net195 net138 net72 vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__or4_1
X_1357_ _0098_ _0311_ _0620_ _0621_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout230 net231 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__buf_1
Xfanout241 _0109_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_2
Xfanout263 _0088_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_1
Xfanout252 _0097_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout285 _0072_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_2
Xfanout296 _0064_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_1
XFILLER_0_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1211_ _0153_ _0155_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__or2_1
X_1142_ _0290_ _0420_ _0421_ _0422_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1073_ net174 net171 net168 vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0857_ net476 net375 net367 net484 vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__a22o_1
X_0926_ net142 net138 vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold27 net39 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ net290 net281 net273 net75 vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__or4_1
X_0788_ net287 net285 _0073_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold16 net19 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1125_ net129 net126 net119 vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__or3_1
X_1056_ net260 net210 vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__or2_1
Xoutput39 net39 vssd1 vssd1 vccd1 vccd1 dout0[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 dout0[26] sky130_fd_sc_hd__buf_2
Xoutput17 net17 vssd1 vssd1 vccd1 vccd1 dout0[16] sky130_fd_sc_hd__buf_2
X_0909_ net491 net378 net345 net500 vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_15_Left_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1039_ net64 net129 net120 _0324_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__or4_1
X_1108_ net256 net114 vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_51_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1390_ _0044_ net237 net97 _0655_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout615 net616 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_1
Xfanout604 addr0_reg\[4\] vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_1
Xfanout626 net627 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0890_ net448 net370 net363 net440 vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__a22o_1
X_1442_ clknet_2_3__leaf_clk0 _0001_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__dfxtp_1
X_1373_ _0356_ _0627_ _0637_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout445 net446 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__buf_1
Xfanout423 net425 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_1
Xfanout412 net413 vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_1
Xfanout434 net435 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_1
Xfanout401 net402 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_18_Left_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout456 net457 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_1
Xfanout489 net490 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__clkbuf_1
Xfanout478 net480 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_1
Xfanout467 net468 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_1
XFILLER_0_36_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout74 net75 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__buf_1
Xfanout52 net54 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
Xfanout41 net42 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_1
Xfanout85 net86 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
Xfanout63 _0187_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_1
Xfanout96 net97 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__buf_1
XFILLER_0_51_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0942_ _0217_ net132 net124 _0224_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__or4_2
XFILLER_0_42_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0873_ net591 net597 net575 net582 vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__and4_1
XFILLER_0_27_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1425_ _0049_ _0056_ _0077_ _0215_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1287_ _0357_ _0433_ _0452_ _0473_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__or4_1
X_1356_ net221 net191 net122 net72 vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_46_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout286 _0072_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_1
Xfanout231 _0115_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_2
Xfanout264 net265 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_1
Xfanout220 _0125_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_1
Xfanout297 _0063_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_1
Xfanout275 _0081_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_2
Xfanout253 net255 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_3_Left_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout242 net243 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_1
XFILLER_0_49_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1072_ _0680_ net68 _0046_ _0225_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__or4_1
X_1210_ _0337_ _0485_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1141_ net67 _0411_ _0412_ _0413_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_35_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0787_ net287 net283 vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__or2_2
X_0856_ net492 net371 net364 net501 vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__a22o_1
X_0925_ net140 net138 net135 vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__or3_1
X_1408_ net303 net300 _0234_ net107 vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_45_Left_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold28 net34 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 net18 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__dlygate4sd3_1
X_1339_ net319 net318 net169 net107 vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1124_ net572 net656 net55 _0405_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__a22o_1
X_1055_ net201 net198 net130 net121 vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0839_ net222 _0125_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__or2_1
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 dout0[27] sky130_fd_sc_hd__buf_2
XFILLER_0_11_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0908_ net426 net378 net345 net433 vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__a22o_1
Xoutput18 net18 vssd1 vssd1 vccd1 vccd1 dout0[17] sky130_fd_sc_hd__buf_2
XFILLER_0_11_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1038_ net333 net324 net319 net312 vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__or4_1
X_1107_ net66 _0152_ _0156_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_32_Left_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout616 addr0_reg\[2\] vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__buf_1
Xfanout627 net628 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_1
Xfanout605 net610 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__buf_1
XFILLER_0_39_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1441_ clknet_2_2__leaf_clk0 _0000_ vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1372_ _0198_ _0333_ _0336_ _0502_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout446 net447 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_1
Xfanout424 net425 vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__clkbuf_1
Xfanout479 net480 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_1
Xfanout413 net418 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout402 net403 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_1
Xfanout435 net439 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_1
Xfanout457 net458 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_1
Xfanout468 net469 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout53 net54 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout75 _0261_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout64 _0187_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_1
Xfanout42 net49 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
Xfanout86 net87 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__buf_1
Xfanout97 _0248_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_51_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0941_ net118 net116 vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0872_ net591 net598 net575 net582 vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__nor4_1
X_1424_ net567 net645 net50 _0689_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__a22o_1
X_1355_ net335 net266 net218 vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_38_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1286_ _0554_ _0555_ _0556_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_46_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout232 _0115_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_1
Xfanout298 _0063_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_1
Xfanout210 _0134_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_1
Xfanout287 _0071_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_2
Xfanout221 net223 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_1
Xfanout243 net244 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_1
Xfanout254 net255 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_1
Xfanout265 _0088_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout276 net280 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_49_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1140_ net256 net253 net62 _0272_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__or4_1
X_1071_ net249 _0107_ _0354_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_43_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0924_ net389 net384 net409 vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_7_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0786_ net553 net412 net515 vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__o21ba_1
X_0855_ net591 net599 net584 net576 vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__nor4b_1
Xhold29 net38 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1338_ _0108_ _0222_ _0309_ _0416_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__or4_1
X_1407_ net564 net633 net47 _0673_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__a22o_1
Xhold18 net13 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__dlygate4sd3_1
X_1269_ _0156_ _0335_ _0339_ _0496_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_49_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1123_ _0394_ _0397_ _0404_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__or3_1
X_1054_ net166 net80 vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__or2_2
XFILLER_0_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0907_ _0192_ net155 vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__or2_1
X_0769_ _0051_ net309 _0053_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__or3_1
X_0838_ net527 net391 net387 net520 vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__a22o_1
Xoutput19 net19 vssd1 vssd1 vccd1 vccd1 dout0[18] sky130_fd_sc_hd__buf_2
XFILLER_0_3_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1106_ net214 _0386_ _0387_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__or3_1
X_1037_ _0696_ _0084_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout606 net610 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__buf_1
Xfanout628 net629 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_1
Xfanout617 net622 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__buf_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1371_ net560 net632 net43 _0636_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1440_ clknet_2_2__leaf_clk0 net9 vssd1 vssd1 vccd1 vccd1 cs0_reg sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout447 _0713_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__buf_1
Xfanout436 net437 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_1
Xfanout414 net417 vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__buf_1
Xfanout425 _0039_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_1
XFILLER_0_39_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout469 net474 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_1
Xfanout403 net404 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_1
Xfanout458 net459 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout54 net56 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__buf_1
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout98 net99 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__buf_1
Xfanout43 net44 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_1
Xfanout76 net77 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__buf_1
Xfanout65 _0166_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__buf_1
Xfanout87 _0255_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_1
XFILLER_0_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0940_ net374 net338 net516 vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0871_ _0150_ _0157_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__or2_1
X_1423_ _0683_ _0686_ _0687_ _0688_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__or4_1
X_1354_ net560 net644 net43 _0619_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__a22o_1
X_1285_ _0113_ net167 net163 vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_46_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout222 net223 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_1
Xfanout200 net201 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_1
Xfanout211 net213 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_1
Xfanout288 _0071_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_1
Xfanout233 _0114_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_1
Xfanout255 _0096_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__buf_1
Xfanout299 _0061_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout277 net280 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__buf_1
Xfanout266 net268 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_1
Xfanout244 _0104_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_21_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1070_ net301 net299 net267 net264 vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0923_ net538 net390 net385 net551 vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__a22o_1
X_0854_ net579 net588 net595 net603 vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__and4b_1
XFILLER_0_7_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0785_ net504 net419 net411 net496 vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1268_ _0388_ _0537_ _0538_ _0539_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__or4_1
X_1406_ _0661_ _0667_ _0672_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__or3_1
Xhold19 net33 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__dlygate4sd3_1
X_1337_ _0333_ _0502_ _0555_ _0603_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__or4_1
X_1199_ net228 net134 vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1122_ _0399_ _0400_ _0402_ _0403_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__or4_2
X_1053_ net239 net235 net79 net75 vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0837_ net551 net392 net386 net538 vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0906_ net456 net379 net348 net466 vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0768_ net311 net308 vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1105_ net224 net211 vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1036_ net209 net205 vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout618 net622 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_1
Xfanout607 net608 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__buf_1
Xfanout629 addr0_reg\[0\] vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__buf_1
XFILLER_0_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1019_ net163 net82 vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1370_ _0626_ _0628_ _0635_ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout404 net405 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_1
Xfanout415 net417 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_1
Xfanout437 net438 vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__buf_1
Xfanout459 net464 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout448 net449 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_1
Xfanout426 net428 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__buf_1
Xfanout55 net56 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__buf_1
Xfanout44 net45 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
Xfanout66 _0148_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__buf_1
Xfanout99 _0246_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout88 _0254_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__buf_1
Xfanout77 net78 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0870_ net195 net192 net189 _0155_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__or4_2
X_1422_ _0035_ _0038_ _0086_ _0093_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_50_Left_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1353_ _0273_ _0615_ _0618_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__or3_1
X_1284_ net254 _0099_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_46_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0999_ _0097_ net222 _0284_ _0285_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout234 _0114_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_1
Xfanout245 _0103_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_2
Xfanout223 _0124_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_1
Xfanout256 _0095_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout212 net213 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_1
Xfanout201 _0144_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_1
Xfanout267 net268 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_1
Xfanout289 _0070_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_1
Xfanout278 net280 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_32_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0922_ net518 net392 net386 net525 vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__a22o_1
X_0853_ net209 net207 net205 net204 vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__or4_2
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0784_ net487 net419 net411 net479 vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__a22o_1
X_1405_ _0407_ _0668_ _0669_ _0671_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1267_ net301 net276 net159 net103 vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__or4_1
Xinput1 addr0[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1198_ _0446_ _0472_ _0473_ _0474_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__or4_1
X_1336_ net91 net89 net84 vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire465 _0710_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1052_ net297 net181 _0310_ _0335_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__or4_1
X_1121_ net65 _0170_ _0247_ _0266_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_31_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0767_ net309 net308 vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0905_ net475 net380 net347 net483 vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__a22o_1
X_0836_ net227 net224 vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1319_ net563 net646 net46 _0587_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__a22o_1
XANTENNA_50 _0410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1104_ net210 net208 net206 vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__or3_1
X_1035_ _0100_ _0215_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0819_ net250 net245 vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout619 net620 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_1
Xfanout608 net609 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1018_ net237 net236 net115 net111 vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout438 net439 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_1
Xfanout416 net418 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_1
XFILLER_0_39_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout427 net428 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_1
Xfanout405 net408 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout449 net450 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_1
XFILLER_0_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout67 _0046_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_29_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout78 net79 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_24_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout56 _0281_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout89 _0254_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
Xfanout45 net48 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_1
XFILLER_0_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1421_ _0199_ _0206_ _0258_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1283_ _0194_ net153 vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__or2_1
X_1352_ _0556_ _0564_ _0603_ _0617_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_46_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0998_ net125 net118 vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout235 _0111_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_1
Xfanout279 net280 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_1
Xfanout224 net225 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_1
XFILLER_0_5_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout202 net203 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_1
Xfanout246 _0102_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_2
Xfanout268 _0087_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout257 net258 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__buf_1
Xfanout213 _0132_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_39_Left_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0921_ net445 net391 net385 net453 vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_23_Left_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0783_ net470 net420 net412 net460 vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__a22o_1
X_0852_ net210 net204 vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1335_ _0283_ _0599_ _0601_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__or3_1
X_1404_ _0090_ net233 net229 _0247_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__or4_1
Xinput2 addr0[1] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_1266_ net283 net282 net92 net87 vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__or4_1
X_1197_ net258 net255 net113 _0237_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_34_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1120_ _0106_ net152 net145 _0401_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__or4_1
X_1051_ net181 net179 vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0904_ net167 net165 net63 _0190_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0766_ net536 net422 net415 net549 vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__a22o_1
X_0835_ net387 net380 net515 vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1318_ _0576_ _0579_ _0580_ _0586_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__or4_1
X_1249_ _0447_ _0512_ _0521_ _0522_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__or4_1
XANTENNA_51 _0512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_40 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire274 _0083_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_1
XFILLER_0_40_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1103_ net571 net638 net54 _0385_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1034_ _0312_ _0314_ _0319_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Left_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0749_ net68 _0035_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0818_ net245 net242 vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_10_Left_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout609 net610 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1017_ net100 net98 net96 vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__or3_2
XFILLER_0_12_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout439 _0715_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_1
Xfanout417 net418 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout406 net408 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_1
Xfanout428 net432 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout68 _0033_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_24_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout79 _0260_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_2
Xfanout46 net47 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_1
XFILLER_0_35_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1420_ _0684_ _0685_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1351_ _0092_ _0268_ _0499_ _0616_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__or4_1
X_1282_ _0145_ _0548_ _0551_ _0552_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_46_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0997_ net325 net302 vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout236 _0111_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_1
Xfanout269 net270 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_1
Xfanout258 _0094_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__buf_1
Xfanout214 _0131_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_1
Xfanout225 _0122_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout203 _0143_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_1
Xfanout247 _0102_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0920_ _0199_ net61 vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__nor2_1
X_0782_ net297 net294 net293 net291 vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__or4_1
X_0851_ net207 net205 net204 vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1265_ net334 net68 net203 net66 vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__or4_1
X_1334_ _0059_ net260 net224 _0600_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1403_ _0098_ _0167_ _0258_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__or3_1
Xinput3 addr0[2] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1196_ net266 net262 net248 net242 vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__or4_1
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Left_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1050_ net307 net291 vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__or2_1
X_0834_ net597 net574 net581 net590 vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__nor4b_1
XTAP_TAPCELL_ROW_31_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0903_ net160 net157 vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0765_ net523 net422 net414 net530 vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_47_Left_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1248_ net62 _0339_ _0519_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__or3_1
X_1317_ _0578_ _0582_ _0583_ _0585_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1179_ net275 _0192_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_52 _0700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_30 _0586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1102_ _0371_ _0373_ _0383_ _0384_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1033_ _0075_ _0315_ _0316_ _0317_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__or4_1
X_0817_ net491 net404 net397 net500 vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__a22o_1
X_0748_ net333 net329 net327 net324 vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1016_ net631 net558 net41 _0302_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout429 net430 vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_1
Xfanout418 _0040_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__buf_1
Xfanout407 net408 vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout58 _0344_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_1
XFILLER_0_32_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout69 net71 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__buf_1
Xfanout47 net48 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_15_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1281_ _0065_ net272 net270 _0496_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__or4_1
X_1350_ net281 net251 net225 net99 vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0996_ _0212_ _0245_ net96 _0282_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__or4_1
Xfanout204 _0137_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_1
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout237 _0110_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_1
Xfanout215 _0131_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_1
Xfanout226 _0122_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__buf_1
Xfanout259 net260 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_1
Xfanout248 net249 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_1
XFILLER_0_49_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0850_ net476 net388 net383 net483 vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__a22o_1
X_0781_ net293 net292 vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1402_ _0150_ _0157_ _0181_ _0603_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1264_ net570 net641 net53 _0536_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__a22o_1
Xinput4 addr0[3] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_1333_ net311 net229 net148 net147 vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1195_ net137 net135 _0322_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0979_ net77 net72 vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_40_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout590 net591 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_1
X_0833_ net506 net390 net385 net498 vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__a22o_1
X_0902_ net485 net380 net347 net477 vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0764_ net421 net415 net410 vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__o21ba_1
X_1178_ net570 net657 net53 _0456_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1316_ _0123_ _0262_ _0584_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__or3_1
X_1247_ _0391_ _0458_ _0513_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_20 _0409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_31 _0591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_42 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 clknet_2_1__leaf_clk0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1101_ net301 net277 _0344_ _0372_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__or4_1
X_1032_ _0075_ _0317_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0747_ net330 net328 net325 vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__or3_1
X_0816_ net475 net406 net398 net483 vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1015_ _0092_ _0286_ _0295_ _0301_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout419 net420 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_1
Xfanout408 _0078_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout59 _0334_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_2
Xfanout48 net49 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_15_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1280_ _0044_ _0230_ _0272_ _0387_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0995_ net166 net83 vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__or2_1
Xfanout238 _0110_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_1
Xfanout216 _0129_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_1
Xfanout227 _0120_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_1
Xfanout205 net206 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_1
Xfanout249 net250 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0780_ net544 net505 net497 net557 vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__a22o_1
X_1401_ _0662_ _0663_ _0665_ _0666_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1194_ _0303_ _0334_ _0426_ _0470_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__or4_1
X_1263_ _0526_ _0532_ _0535_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__or3_1
X_1332_ net162 net160 _0457_ _0598_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__or4_1
Xinput5 addr0[4] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0978_ net72 net69 vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_40_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout580 addr0_reg\[7\] vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__buf_1
Xfanout591 net596 vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_31_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0763_ net613 net625 net618 net606 vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__or4b_1
XFILLER_0_43_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0832_ net603 net579 net588 net595 vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__and4b_1
X_0901_ net466 net379 net346 net456 vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__a22o_1
X_1315_ net192 _0155_ net149 net136 vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__or4_1
X_1177_ _0229_ _0374_ _0454_ _0455_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1246_ _0086_ _0149_ _0414_ _0518_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_32 _0644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_21 _0409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_10 _0164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1100_ _0378_ _0379_ _0381_ _0382_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__or4_1
X_1031_ net133 net132 net124 vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0746_ _0714_ net323 vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0815_ net456 net404 net397 net466 vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__a22o_1
X_1229_ _0105_ _0497_ _0502_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2__f_clk0 clknet_0_clk0 vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1014_ _0283_ _0298_ _0299_ _0300_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_14_Left_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0729_ net617 net623 net611 net605 vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__and4b_1
XFILLER_0_8_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout409 _0050_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__buf_1
XFILLER_0_29_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout49 net56 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_1
XFILLER_0_44_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0994_ _0244_ _0274_ _0276_ _0280_ cs0_reg vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__o41a_1
Xfanout239 _0109_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_1
Xfanout228 _0120_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_1
Xfanout217 _0129_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_1
Xfanout206 _0136_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_17_Left_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1400_ _0708_ net324 net278 net249 vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__or4_1
X_1331_ net328 net323 net219 net176 vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput6 addr0[5] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
X_1262_ _0036_ _0533_ _0534_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__or3_1
X_1193_ _0037_ _0173_ _0392_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__or3_1
XFILLER_0_52_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0977_ net500 net359 net352 net491 vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout592 net593 vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_1
Xfanout570 net571 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__buf_1
Xfanout581 net583 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0900_ _0185_ _0186_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0762_ net320 _0042_ net316 net312 vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__or4_1
X_0831_ net595 net579 net588 net603 vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1314_ net209 net207 _0305_ _0549_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1176_ _0445_ _0447_ _0450_ _0452_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1245_ net192 net189 net114 net112 vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_44_Left_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_11 _0175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_33 _0665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_22 _0411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1030_ net294 net292 vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0814_ net426 net401 net394 net433 vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__a22o_1
X_0745_ net554 net436 net429 net541 vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1228_ _0098_ _0498_ _0499_ _0500_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__or4_1
X_1159_ _0036_ _0389_ _0426_ _0430_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1013_ _0287_ _0294_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0728_ net540 net508 net515 vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0993_ _0275_ _0277_ _0278_ _0279_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout207 _0135_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__buf_1
Xfanout229 net231 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_1
Xfanout218 net219 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_1
XFILLER_0_49_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1261_ _0198_ net111 _0241_ _0448_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__or4_1
X_1330_ net563 net655 net46 _0597_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1192_ net567 net642 net50 _0469_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__a22o_1
Xinput7 addr0[6] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0976_ net467 net359 net352 net457 vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1459_ clknet_2_2__leaf_clk0 _0018_ vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout560 net561 vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_48_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout593 net594 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_1
Xfanout582 net583 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_1
Xfanout571 net573 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__buf_1
X_0830_ net240 net238 net236 net234 vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__or4_2
XFILLER_0_22_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0761_ net320 net313 vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1313_ _0049_ _0199_ _0395_ _0581_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__or4_1
X_1244_ net218 net170 net103 net84 vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__or4_1
X_1175_ _0291_ _0306_ _0453_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__or3_1
XANTENNA_12 _0205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_45 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _0431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_34 _0714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0959_ net427 net356 net349 net434 vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_53_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout390 net393 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0813_ net257 _0095_ net253 net251 vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__or4_1
X_0744_ net607 net627 net620 net614 vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_24_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1158_ _0322_ _0435_ _0436_ _0437_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__or4_1
X_1227_ net187 net182 vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__or2_1
X_1089_ net332 net98 vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1012_ _0138_ _0288_ _0291_ _0292_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0727_ net602 net577 net587 net594 vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_8_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0992_ _0181_ net63 _0190_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__or3_1
Xfanout219 _0128_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_1
Xfanout208 _0135_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_1
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1191_ _0466_ _0467_ _0468_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__or3_1
Xinput8 addr0[7] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
X_1260_ _0163_ _0262_ _0315_ _0413_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0975_ net79 net74 vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__or2_1
X_1389_ net301 net299 net284 net282 vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__or4_1
X_1458_ clknet_2_2__leaf_clk0 _0017_ vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout572 net573 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_48_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout550 net551 vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_1
Xfanout583 net584 vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout561 net562 vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__clkbuf_1
Xfanout594 net595 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_1
X_0760_ net318 net317 net313 vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1312_ net310 net302 net237 net143 vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__or4_1
X_1174_ net67 _0180_ _0451_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__or3_1
X_1243_ _0498_ _0514_ _0515_ _0516_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__or4_1
XANTENNA_13 _0238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_46 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_35 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0889_ net434 net369 net362 net427 vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0958_ net492 net356 net349 net501 vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__a22o_1
XANTENNA_24 _0431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout391 net392 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__clkbuf_1
Xfanout380 net382 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_1
XFILLER_0_33_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0743_ net626 net619 net608 net615 vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__and4bb_1
X_0812_ net258 net252 vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1226_ net287 net228 net216 net95 vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__or4_1
X_1157_ _0202_ _0242_ net88 net84 vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__or4_1
X_1088_ net113 _0239_ _0370_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__or3_2
XFILLER_0_15_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1011_ _0289_ _0293_ _0296_ _0297_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0726_ net609 net612 net623 net617 vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1209_ net62 net151 _0202_ net144 vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0991_ net167 net163 _0247_ _0253_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout209 _0134_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__buf_1
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1190_ _0113_ _0316_ _0460_ _0461_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__or4_1
Xinput9 cs0 vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0974_ net390 net354 net515 vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_14_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1457_ clknet_2_2__leaf_clk0 _0016_ vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1388_ _0287_ net59 _0377_ _0427_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__or4_1
Xfanout540 net543 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__buf_1
Xfanout551 net552 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__buf_1
Xfanout595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_1
Xfanout584 net589 vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_1
Xfanout562 net565 vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__buf_1
Xfanout573 _0629_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1311_ _0431_ _0451_ _0460_ _0511_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__or4_1
X_1173_ net185 net182 net146 net144 vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1242_ net142 _0322_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__or2_1
XANTENNA_36 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 _0454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_14 _0241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0957_ _0229_ _0231_ _0236_ _0243_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__or4_2
XFILLER_0_42_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0888_ net547 net369 net362 net534 vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_53_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout392 net393 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_1
Xfanout381 net382 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_1
Xfanout370 net371 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_1
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0742_ net553 net453 net445 net540 vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0811_ net256 net254 net251 vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__or3_1
X_1087_ net298 net293 net291 vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__or3_1
X_1156_ _0112_ _0228_ _0310_ _0343_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__or4_1
X_1225_ net156 net153 _0205_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_50_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1010_ net322 net289 net152 net150 vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_29_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0725_ net336 net334 vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__or2_1
X_1208_ net65 _0268_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1139_ _0038_ _0062_ _0259_ _0418_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_9_Left_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1 net10 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_35_Left_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0990_ _0140_ _0215_ _0259_ _0268_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0973_ net485 net360 net353 net477 vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1456_ clknet_2_1__leaf_clk0 _0015_ vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__dfxtp_1
X_1387_ _0537_ _0650_ _0652_ vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout530 net531 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_1
Xfanout541 net543 vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_1
Xfanout552 _0649_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_1
Xfanout585 net586 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_1
Xfanout574 net575 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_1
Xfanout596 addr0_reg\[5\] vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_1
Xfanout563 net564 vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__buf_1
XFILLER_0_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_38_Left_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1241_ net63 net161 vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__or2_1
X_1310_ net57 _0318_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_22_Left_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1172_ net278 net266 net261 net259 vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__or4_1
X_0956_ _0237_ net106 net104 net101 vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__or4_1
XANTENNA_26 _0462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 _0272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_48 _0088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0887_ net65 _0167_ _0170_ _0173_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__nor4_1
X_1439_ clknet_2_0__leaf_clk0 net8 vssd1 vssd1 vccd1 vccd1 addr0_reg\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_53_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout393 _0118_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_1
Xfanout382 _0121_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_1
Xfanout360 net361 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_1
Xfanout371 net372 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__buf_1
X_0810_ net533 net403 net396 net546 vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__a22o_1
X_0741_ net607 net619 net626 net615 vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1224_ net202 net199 net195 net190 vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_50_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1086_ net568 net658 net51 _0369_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__a22o_1
X_1155_ _0127_ _0295_ _0317_ _0358_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__or4_1
X_0939_ net509 net503 net495 net337 vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout190 net191 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_1
X_0724_ net554 net531 net521 net542 vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1207_ net570 net654 net53 _0483_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1069_ net572 net661 net55 _0353_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1138_ _0181_ _0307_ _0407_ _0417_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__or4_1
XFILLER_0_50_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 net24 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0972_ net88 net84 net82 net81 vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1455_ clknet_2_3__leaf_clk0 _0014_ vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__dfxtp_1
X_1386_ net268 net260 _0372_ _0651_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout542 net543 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__buf_1
Xfanout531 _0690_ vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__buf_1
Xfanout520 net521 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout586 net587 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_1
Xfanout553 net556 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__buf_1
Xfanout597 net599 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__buf_1
Xfanout575 net576 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_1
Xfanout564 net565 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1171_ _0106_ _0390_ _0448_ _0449_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__or4_1
X_1240_ _0123_ net211 vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_27 _0480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_16 _0272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0955_ net103 net102 vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__or2_1
XANTENNA_49 _0272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0886_ net179 net177 vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__or2_1
X_1438_ clknet_2_0__leaf_clk0 net7 vssd1 vssd1 vccd1 vccd1 addr0_reg\[6\] sky130_fd_sc_hd__dfxtp_1
X_1369_ _0273_ _0631_ _0633_ _0634_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_53_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout361 _0159_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_1
Xfanout383 net384 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_1
Xfanout350 net351 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_1
Xfanout372 net373 vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_1
Xfanout394 net395 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_1
X_0740_ net615 net628 net621 net609 vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__and4b_1
X_1154_ _0427_ _0428_ _0431_ _0433_ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__or4_1
X_1223_ net131 _0413_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_50_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1085_ _0365_ _0368_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0938_ net124 net122 vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0869_ net191 _0155_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__or2_2
XFILLER_0_2_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout191 _0154_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__buf_1
Xfanout180 _0169_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_1
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0723_ net608 net626 net619 net614 vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1206_ _0471_ _0475_ _0482_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1137_ net327 net257 net179 net123 vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1068_ _0345_ _0347_ _0352_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__or3_1
XFILLER_0_35_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold3 net27 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1471_ clknet_2_1__leaf_clk0 _0030_ vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_37_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0971_ net83 net81 vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__or2_1
X_1454_ clknet_2_2__leaf_clk0 _0013_ vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__dfxtp_1
X_1385_ net244 net147 net112 net110 vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout510 net512 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__buf_1
Xfanout543 _0660_ vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_1
Xfanout554 net556 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_1
Xfanout521 net524 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__buf_1
Xfanout532 net533 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_1
Xfanout565 net566 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_1
Xfanout587 net588 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_1
Xfanout576 net580 vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_1
Xfanout598 net599 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1170_ net306 net304 vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__or2_1
X_0954_ net509 net495 net337 net503 vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_17 _0312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_28 _0553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0885_ net533 net357 net350 net546 vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__a22o_1
XANTENNA_39 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1437_ clknet_2_0__leaf_clk0 net6 vssd1 vssd1 vccd1 vccd1 addr0_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1368_ _0117_ _0315_ _0316_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__or3_1
X_1299_ _0270_ _0566_ _0567_ _0568_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_53_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout340 net342 vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_1
Xfanout384 net387 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_1
Xfanout362 net363 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__buf_1
Xfanout395 net396 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_1
Xfanout373 net376 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_1
Xfanout351 net352 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__buf_1
XFILLER_0_24_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1084_ _0355_ _0356_ _0366_ _0367_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__or4_1
X_1222_ net102 net89 vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__or2_1
X_1153_ net100 net98 net93 vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_50_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0937_ net511 net451 net444 net341 vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__a22o_1
X_0799_ net278 net275 net272 net269 vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__or4_2
X_0868_ net519 net375 net367 net526 vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout181 _0168_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_1
Xfanout170 net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout192 net194 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_1
XFILLER_0_29_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0722_ net614 net627 net619 net607 vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1205_ _0479_ _0480_ _0481_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__or3_1
X_1067_ _0348_ _0349_ _0350_ _0351_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1136_ _0414_ _0415_ _0416_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4 net14 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1119_ net287 net276 net270 net216 vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_0_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1470_ clknet_2_2__leaf_clk0 _0029_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_46_Left_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0970_ net525 net381 net348 net518 vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__a22o_1
X_1453_ clknet_2_2__leaf_clk0 _0012_ vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1384_ _0139_ net141 net137 _0513_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout522 net523 vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__buf_1
Xfanout511 net513 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__buf_1
Xfanout555 net556 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_1
Xfanout544 _0660_ vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__buf_1
Xfanout577 net580 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__buf_1
Xfanout588 net589 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__buf_1
Xfanout599 net604 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__buf_1
Xfanout566 net573 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_1
XFILLER_0_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout533 net534 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_1
Xfanout500 net502 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_1
XFILLER_0_51_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_18 _0312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_29 _0560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0953_ net508 net479 net337 net487 vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0884_ net442 net358 net351 net450 vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__a22o_1
X_1436_ clknet_2_0__leaf_clk0 net5 vssd1 vssd1 vccd1 vccd1 addr0_reg\[4\] sky130_fd_sc_hd__dfxtp_1
X_1367_ net156 net153 _0458_ _0632_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_53_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1298_ _0038_ _0150_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout341 net342 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_1
Xfanout330 net331 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_1
Xfanout385 net386 vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_1
Xfanout374 net375 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_1
Xfanout363 net364 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_1
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__clkbuf_1
Xfanout352 net355 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_1
X_1221_ net143 net140 vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_9_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1083_ net283 net110 _0310_ _0339_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__or4_1
X_1152_ net100 net93 vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_50_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0936_ net529 net510 net339 net522 vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__a22o_1
X_0798_ net279 net273 vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0867_ net441 net369 net362 net449 vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1419_ _0059_ net257 net226 _0140_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__or4_1
XFILLER_0_53_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout193 net194 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_1
Xfanout182 _0165_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_1
Xfanout171 _0177_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_1
Xfanout160 _0188_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__buf_1
XFILLER_0_44_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0721_ net555 net548 net542 net535 vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_12_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1204_ _0704_ _0048_ _0085_ _0205_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1135_ net290 net286 net281 vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__or3_2
X_1066_ net271 _0123_ net196 _0346_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0919_ net149 net148 net146 net144 vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_3_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold5 net31 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1049_ net115 net104 net101 vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__or3_1
X_1118_ net336 net68 _0212_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_73 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1452_ clknet_2_1__leaf_clk0 _0011_ vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__dfxtp_1
X_1383_ net567 net637 net50 _0648_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout512 net513 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_1
Xfanout523 net524 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__clkbuf_1
Xfanout556 _0639_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__buf_1
Xfanout578 net579 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_1
Xfanout589 addr0_reg\[6\] vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_1
Xfanout567 net569 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_1
Xfanout545 net546 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__buf_1
Xfanout501 net502 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_16_Left_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout534 net539 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_1
XFILLER_0_51_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0952_ _0237_ net106 vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__or2_1
XANTENNA_19 _0352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0883_ net181 net180 vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1366_ net158 net111 net103 net101 vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__or4_1
X_1435_ clknet_2_0__leaf_clk0 net4 vssd1 vssd1 vccd1 vccd1 addr0_reg\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1297_ _0034_ _0047_ _0236_ net60 vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout320 net321 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_1
Xfanout331 _0703_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__buf_1
Xfanout342 net343 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_1
Xfanout375 net376 vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_1
Xfanout386 net387 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__buf_1
Xfanout353 net355 vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_1_Left_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout364 net365 vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__buf_1
Xfanout397 net400 vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_1
XFILLER_0_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1151_ net108 _0239_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__or2_1
X_1220_ net568 net643 net51 _0495_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1082_ _0054_ _0153_ _0262_ _0285_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_50_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0935_ net133 net132 net128 net125 vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__or4_1
X_0866_ _0151_ net193 vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0797_ net469 net407 net399 net459 vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_43_Left_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1418_ net230 _0117_ _0166_ _0268_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1349_ _0576_ _0611_ _0613_ _0614_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__or4_1
Xfanout183 _0165_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_1
Xfanout150 _0200_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout172 net173 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__buf_1
Xfanout161 _0188_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_1
Xfanout194 _0152_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0720_ net606 net612 net624 net618 vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__and4b_1
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1203_ net309 net150 _0476_ _0477_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1134_ net241 net233 _0186_ net157 vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__or4_1
X_1065_ _0074_ _0082_ _0340_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0849_ net494 net388 net383 net502 vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__a22o_1
X_0918_ net146 net144 vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__or2_2
XFILLER_0_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_1__f_clk0 clknet_0_clk0 vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6 net30 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1117_ net252 net235 net185 _0398_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1048_ net114 net102 vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1451_ clknet_2_3__leaf_clk0 _0010_ vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__dfxtp_1
X_1382_ _0472_ _0638_ _0640_ _0647_ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout513 net514 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_1
Xfanout524 _0695_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__buf_1
Xfanout502 net507 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__buf_1
XFILLER_0_13_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout535 net537 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__buf_1
Xfanout557 _0639_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__buf_1
Xfanout579 net580 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_1
Xfanout568 net569 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_1
Xfanout546 net547 vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__buf_1
XFILLER_0_47_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0951_ net522 net510 net339 net529 vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0882_ net361 net354 net409 vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_50_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1434_ clknet_2_0__leaf_clk0 net3 vssd1 vssd1 vccd1 vccd1 addr0_reg\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1296_ net63 net157 _0564_ _0565_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__or4_1
X_1365_ net272 net75 _0630_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_53_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout321 net322 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_1
Xfanout343 _0216_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__buf_1
Xfanout332 _0700_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout310 _0052_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout354 net355 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__buf_1
Xfanout365 net366 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_1
Xfanout376 _0141_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_1
Xfanout387 _0119_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_1
Xfanout398 net400 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_1
X_1150_ net319 net317 net312 net285 vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_9_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1081_ _0360_ _0361_ _0363_ _0364_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0934_ net130 net127 vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0865_ net533 net369 net362 net546 vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__a22o_1
X_0796_ net593 net516 net600 net586 vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__nor4b_1
X_1417_ _0244_ _0668_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1348_ _0198_ _0323_ _0336_ _0449_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__or4_1
X_1279_ net131 net105 _0497_ _0549_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout140 _0209_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_1
Xfanout195 _0151_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout184 _0164_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_1
Xfanout173 _0176_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout151 net152 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout162 _0185_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__buf_1
XFILLER_0_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1202_ _0338_ _0396_ _0416_ _0478_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__or4_1
X_1064_ net244 net62 net146 _0339_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__or4_1
X_1133_ net187 net186 net76 net70 vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0779_ net540 net470 net460 net553 vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__a22o_1
X_0848_ net459 net389 net384 net469 vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__a22o_1
X_0917_ net380 net347 net409 vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_3_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7 net25 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1047_ net570 net639 net53 _0332_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1116_ net164 _0192_ net134 net110 vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk0 clk0 vssd1 vssd1 vccd1 vccd1 clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1450_ clknet_2_1__leaf_clk0 _0009_ vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dfxtp_1
X_1381_ _0112_ _0644_ _0645_ _0646_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout536 net537 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_1
Xfanout514 _0699_ vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__buf_1
Xfanout503 net504 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_1
Xfanout525 net526 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__buf_1
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout547 net552 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_1
Xfanout569 net571 vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_1
Xfanout558 net559 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__buf_1
XFILLER_0_47_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0950_ net511 net443 net341 net451 vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0881_ net521 net360 net353 net528 vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1433_ clknet_2_0__leaf_clk0 net2 vssd1 vssd1 vccd1 vccd1 addr0_reg\[1\] sky130_fd_sc_hd__dfxtp_1
X_1295_ net303 net300 _0066_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__or3_1
X_1364_ net327 net323 net131 net105 vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout311 _0051_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout333 _0700_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_1
Xfanout300 _0061_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__buf_1
Xfanout322 _0041_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_1
Xfanout355 _0160_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_1
Xfanout399 net400 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_1
Xfanout388 net389 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_1
Xfanout344 net345 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_1
Xfanout377 net378 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_1
Xfanout366 net368 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__buf_1
XFILLER_0_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1080_ _0057_ net257 net61 net106 vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0933_ net511 net471 net461 net341 vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__a22o_1
X_0864_ net374 net367 net410 vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__o21ba_1
X_0795_ net277 net275 vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1416_ net567 net640 net50 _0682_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__a22o_1
X_1347_ _0190_ _0457_ _0612_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__or3_1
X_1278_ net335 net329 vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__or2_1
Xfanout130 _0219_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_2
Xfanout141 _0209_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_1
Xfanout163 net165 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout174 _0175_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_1
Xfanout196 _0147_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_1
Xfanout152 _0196_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_2
Xfanout185 _0162_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__buf_1
XFILLER_0_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1201_ net269 net220 net215 net94 vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__or4_1
X_1063_ _0341_ _0342_ _0343_ net58 vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__or4_1
X_1132_ net133 net122 vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0916_ net532 net378 net345 net545 vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__a22o_1
X_0847_ net431 net389 net384 net438 vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__a22o_1
X_0778_ net297 net296 vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold8 net35 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1115_ _0034_ _0370_ _0395_ _0396_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__or4_1
X_1046_ _0320_ _0328_ _0331_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_0_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1029_ net305 net299 vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_36_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1380_ _0065_ _0074_ _0099_ _0266_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout537 net538 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_1
Xfanout548 net550 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__buf_1
Xfanout504 net505 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_1
Xfanout515 net517 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__buf_1
Xfanout526 net527 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_1
XFILLER_0_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout559 net566 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0880_ net186 net183 vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__or2_1
X_1432_ clknet_2_0__leaf_clk0 net1 vssd1 vssd1 vccd1 vccd1 addr0_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1363_ _0446_ _0461_ _0514_ _0627_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__or4_1
XFILLER_0_53_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1294_ net131 net123 net122 vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__or3_1
XFILLER_0_53_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_52_Left_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout301 net303 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_1
Xfanout312 net314 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_1
Xfanout334 _0696_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__buf_1
Xfanout323 _0032_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout367 net368 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_1
Xfanout389 net393 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_1
Xfanout345 net346 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_1
Xfanout356 net358 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__buf_1
Xfanout378 net379 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_52_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0932_ net508 net486 net478 net338 vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0794_ net484 net406 net398 net475 vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__a22o_1
X_0863_ net203 net199 net198 net196 vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__or4_2
XFILLER_0_48_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1415_ _0678_ _0679_ _0681_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__or3_1
X_1346_ _0164_ net177 net127 net109 vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__or4_1
X_1277_ net218 _0170_ net176 net58 vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout120 net121 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_5_Left_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout131 _0218_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_1
Xfanout175 _0175_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout164 _0184_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout197 _0147_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_1
Xfanout153 net154 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_1
Xfanout186 _0162_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_1
Xfanout142 _0208_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_1
XFILLER_0_20_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1200_ net164 net80 vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1062_ _0214_ _0293_ _0338_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__or3_1
X_1131_ net329 net291 vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0915_ net149 net148 vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__or2_1
X_0777_ net541 net436 net429 net554 vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__a22o_1
X_0846_ _0127_ _0130_ net214 net212 vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1329_ _0470_ _0588_ _0594_ _0596_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__or4_1
Xhold9 net21 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1114_ net175 net92 net87 vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__or3_1
XFILLER_0_29_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1045_ net194 _0156_ _0329_ _0330_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__or4_1
X_0829_ net238 net233 vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_39_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_8_Left_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1028_ _0055_ net231 _0313_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_34_Left_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout549 net550 vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_1
Xfanout505 net506 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_1
Xfanout516 net517 vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__clkbuf_1
Xfanout538 net539 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_1
Xfanout527 net528 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1431_ net558 net649 _0252_ net41 vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__a22o_1
X_1293_ net250 net246 net90 net88 vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__or4_1
X_1362_ _0181_ _0603_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout313 net314 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_1
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout324 net326 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__buf_1
Xfanout368 _0142_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_1
Xfanout335 net336 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_1
Xfanout357 net358 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_1
Xfanout346 net348 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_1
Xfanout379 net382 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_52_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_37_Left_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0931_ net548 net510 net339 net535 vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__a22o_1
X_0862_ net202 net199 net196 vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_21_Left_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0793_ net501 net402 net395 net491 vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__a22o_1
X_1276_ net572 net660 net55 _0547_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1414_ _0108_ _0374_ _0668_ _0677_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1345_ _0704_ _0105_ _0179_ _0205_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout132 _0218_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_1
Xfanout110 _0235_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout143 _0208_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_1
Xfanout121 _0226_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__buf_1
Xfanout165 _0184_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__buf_1
Xfanout154 _0195_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout187 _0161_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__buf_1
Xfanout198 _0146_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_1
Xfanout176 _0172_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__buf_1
XFILLER_0_49_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1130_ net206 net140 vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__or2_1
X_1061_ net261 net207 net173 net90 vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__or4_1
XFILLER_0_50_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0845_ net483 net388 net383 net475 vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__a22o_1
X_0914_ net440 net377 net344 net448 vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0776_ net544 net486 net478 net557 vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1259_ _0221_ _0527_ _0529_ _0531_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_3_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1328_ _0163_ _0412_ _0432_ _0595_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1113_ net128 net118 net116 vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__or3_1
XFILLER_0_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1044_ _0307_ _0309_ _0311_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_0_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0828_ net443 net421 net414 net451 vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0759_ net318 net315 vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1027_ net113 net107 _0237_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_36_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout506 net507 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__buf_1
XFILLER_0_13_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout517 _0698_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout539 _0670_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__buf_1
Xfanout528 net531 vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__buf_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1430_ net563 net635 net46 _0694_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1292_ net559 net653 net42 _0562_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__a22o_1
X_1361_ _0622_ _0623_ _0625_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout314 net315 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__buf_1
Xfanout303 _0060_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__buf_1
Xfanout325 net326 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout336 _0680_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_1
Xfanout347 net348 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__buf_1
Xfanout369 net370 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__buf_1
Xfanout358 net359 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_1
XFILLER_0_32_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0930_ net509 net437 net430 net337 vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__a22o_1
X_0792_ net590 net597 net574 net581 vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__and4bb_1
X_0861_ net198 net196 vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__or2_1
X_1413_ _0371_ _0373_ _0676_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__or3_1
X_1275_ _0540_ _0543_ _0546_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__or3_1
X_1344_ net558 net652 net41 _0610_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__a22o_1
Xwire57 _0174_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout133 net134 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout111 _0234_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_1
Xfanout122 _0224_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__buf_1
Xfanout166 _0183_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_1
Xfanout144 _0204_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_1
Xfanout100 _0245_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__buf_1
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_1
Xfanout177 _0172_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__buf_1
Xfanout155 _0193_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_1
Xfanout188 _0161_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1060_ net60 _0314_ net59 _0337_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0775_ net307 net305 net304 net300 vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__or4_2
X_0844_ net473 net390 net385 net463 vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__a22o_1
X_0913_ net519 net381 net347 net526 vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1189_ _0708_ _0108_ _0236_ _0459_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__or4_1
X_1258_ net61 _0288_ _0429_ _0530_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__or4_1
X_1327_ _0055_ _0116_ _0123_ _0242_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_49_Left_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1043_ net60 _0304_ _0306_ _0308_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__or4_1
X_1112_ _0093_ _0388_ _0389_ _0393_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_0_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0758_ net452 net421 net414 net443 vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0827_ net460 net423 net416 net470 vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1026_ _0149_ net168 _0179_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__or3_2
XFILLER_0_47_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout529 net530 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__buf_1
Xfanout507 _0701_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__buf_1
Xfanout518 net519 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_1
XFILLER_0_6_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1009_ net336 net307 net305 net239 vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1360_ _0090_ net200 net197 _0624_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__or4_1
X_1291_ _0550_ _0553_ _0557_ _0561_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout337 net338 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_1
Xfanout304 _0060_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_1
Xfanout315 _0045_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_1
Xfanout348 _0182_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_1
Xfanout326 _0711_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_1
Xfanout359 net361 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_1
XFILLER_0_17_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0791_ net574 net581 net590 net598 vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0860_ net427 net370 net363 net434 vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1412_ net230 _0117_ _0548_ _0669_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__or4_1
X_1343_ _0602_ _0604_ _0609_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__or3_1
X_1274_ _0406_ _0512_ _0544_ _0545_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0989_ _0133_ _0158_ net57 _0207_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__or4bb_1
Xfanout101 net102 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__buf_1
Xfanout134 _0217_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout189 net190 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__buf_1
Xfanout156 _0193_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_1
Xfanout123 net124 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__buf_1
Xfanout167 _0183_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_1
Xfanout112 _0233_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__buf_1
Xfanout145 _0204_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_1
Xfanout178 _0171_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0912_ _0192_ net155 net154 net151 vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__or4_4
X_0774_ net543 net451 net443 net556 vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__a22o_1
X_0843_ _0128_ net217 vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_11_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1326_ _0355_ _0589_ _0591_ _0593_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__or4_1
X_1188_ _0312_ _0462_ _0463_ _0465_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__or4_1
X_1257_ net235 net208 net166 net98 vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1042_ _0321_ _0325_ _0326_ _0327_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__or4_1
X_1111_ _0116_ _0390_ _0391_ _0392_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_0_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0757_ net318 net316 vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__or2_1
X_0826_ net241 net236 vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1309_ net202 net66 _0525_ _0577_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1025_ _0169_ net178 net176 vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__or3_1
X_0809_ net518 net406 net398 net525 vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_1 _0033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout508 net514 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__buf_1
Xfanout519 net520 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__buf_1
X_1008_ net174 net172 net170 vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1290_ _0062_ _0138_ _0558_ _0560_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 _0058_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__buf_1
Xfanout327 net328 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_1
Xfanout316 _0043_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__buf_1
Xfanout338 net343 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__buf_1
Xfanout349 net351 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_1
XFILLER_0_17_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0790_ net290 net288 net286 net281 vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1273_ _0047_ net240 _0112_ _0375_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__or4_1
X_1342_ _0605_ _0606_ _0607_ _0608_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__or4_1
X_1411_ net294 net288 _0081_ net269 vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0988_ _0086_ _0093_ _0100_ _0108_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__or4_1
Xfanout102 _0241_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_2
Xfanout113 _0233_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__buf_1
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout124 _0223_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout168 net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_1
Xfanout135 _0211_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout146 _0203_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_1
Xfanout157 _0189_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__buf_1
Xfanout179 _0171_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Left_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0842_ net438 net392 net386 net431 vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0911_ net155 net151 vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__or2_1
X_0773_ net541 net529 net522 net554 vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1256_ _0106_ _0156_ _0528_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__or3_1
X_1325_ _0258_ _0267_ _0592_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1187_ net224 _0130_ net183 _0464_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1110_ _0186_ net161 vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__or2_1
X_1041_ _0137_ net65 _0167_ _0197_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0825_ net237 net235 vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0756_ net437 net423 net416 net430 vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1239_ net297 net241 vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__or2_1
X_1308_ net253 net251 net221 net217 vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1024_ net180 net178 vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_44_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Left_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0808_ net440 net401 net394 net448 vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_12_Left_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0739_ net553 net470 net460 net540 vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2 _0033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout509 net514 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_1
XFILLER_0_6_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1007_ net192 net189 net90 net88 vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout339 net340 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_1
Xfanout317 _0043_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_1
Xfanout306 _0058_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_1
Xfanout328 _0707_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1410_ _0229_ _0231_ _0674_ _0675_ vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1272_ _0708_ _0229_ _0289_ _0313_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__or4_1
X_1341_ _0054_ _0068_ _0126_ _0153_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0987_ _0269_ _0270_ _0273_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout125 net126 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_1
Xfanout114 _0232_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_2
Xfanout103 _0240_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_2
Xfanout136 _0211_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout147 _0203_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_1
Xfanout169 _0178_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_2
Xfanout158 net159 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0772_ net307 net305 vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__or2_1
X_0841_ net454 net388 net383 net446 vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0910_ net153 net152 vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1255_ net220 net219 net203 _0146_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__or4_1
X_1186_ net191 net164 net136 net94 vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__or4_1
X_1324_ net278 net172 net167 net123 vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Left_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1040_ net259 net225 _0322_ _0323_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0755_ net549 net423 net416 net536 vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__a22o_1
X_0824_ net495 net419 net411 net503 vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1169_ net298 net230 vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1238_ _0100_ net99 _0311_ _0511_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__or4_2
X_1307_ net59 _0359_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1023_ net76 net74 net73 vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_44_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0738_ net606 net613 net624 net618 vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0807_ net406 net398 net409 vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_3 _0055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1006_ net188 net184 net133 net123 vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 dout0[9] sky130_fd_sc_hd__buf_2
XFILLER_0_53_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout329 net331 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__buf_1
Xfanout307 _0057_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_1
Xfanout318 _0042_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_1
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1340_ net264 net233 _0168_ net154 vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1271_ _0130_ _0167_ _0541_ _0542_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0986_ _0049_ _0054_ _0272_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout126 net127 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_1
Xfanout104 _0240_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__buf_1
Xfanout115 _0232_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__buf_1
XFILLER_0_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout159 _0189_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout137 net139 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_1
X_1469_ clknet_2_3__leaf_clk0 _0028_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__dfxtp_1
Xfanout148 _0201_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_1
XFILLER_0_49_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0771_ net555 net541 net410 vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__o21ba_1
X_0840_ net228 net226 net221 net220 vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_11_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1323_ net284 net217 net215 _0590_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1185_ _0697_ _0099_ _0153_ _0230_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__or4_1
X_1254_ _0076_ _0139_ net141 net137 vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_19_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0969_ net545 net377 net344 net532 vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout490 _0705_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_1
XFILLER_0_28_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0754_ net529 net423 net416 net522 vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__a22o_1
X_0823_ net478 net419 net411 net486 vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1306_ net560 net647 net43 _0575_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__a22o_1
X_1099_ _0148_ net64 _0250_ _0267_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__or4_1
X_1168_ net324 _0033_ _0446_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__or3_1
X_1237_ net248 _0103_ net243 vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_0__f_clk0 clknet_0_clk0 vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1022_ net249 net246 net245 vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_44_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0737_ net625 net618 net606 net612 vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__and4b_1
XFILLER_0_24_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0806_ net266 net263 net262 net259 vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 _0057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xcust_rom0_630 vssd1 vssd1 vccd1 vccd1 cust_rom0_630/HI dout0[31] sky130_fd_sc_hd__conb_1
XFILLER_0_16_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1005_ net214 net212 net178 net176 vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__or4_1
XFILLER_0_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 dout0[28] sky130_fd_sc_hd__buf_2
XFILLER_0_53_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout308 _0053_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__buf_1
Xfanout319 net321 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__buf_1
.ends

