VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cust_rom
  CLASS BLOCK ;
  FOREIGN cust_rom ;
  ORIGIN 0.000 0.000 ;
  SIZE 142.880 BY 153.600 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 141.680 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 141.680 ;
    END
  END VPWR
  PIN addr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END addr0[7]
  PIN clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END clk0
  PIN cs0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 23.840 142.880 24.440 ;
    END
  END cs0
  PIN dout0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 68.040 142.880 68.640 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 81.640 142.880 82.240 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 108.840 142.880 109.440 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 87.030 149.600 87.310 153.600 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 64.640 142.880 65.240 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 57.840 142.880 58.440 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 78.240 142.880 78.840 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 47.640 142.880 48.240 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 98.640 142.880 99.240 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 77.370 149.600 77.650 153.600 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 71.440 142.880 72.040 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 95.240 142.880 95.840 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 105.440 142.880 106.040 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 119.040 142.880 119.640 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 115.640 142.880 116.240 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 88.440 142.880 89.040 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 54.440 142.880 55.040 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 51.040 142.880 51.640 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 40.840 142.880 41.440 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 37.440 142.880 38.040 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.470 149.600 93.750 153.600 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 27.240 142.880 27.840 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END dout0[31]
  PIN dout0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 149.600 16.470 153.600 ;
    END
  END dout0[32]
  PIN dout0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 67.710 149.600 67.990 153.600 ;
    END
  END dout0[3]
  PIN dout0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 99.910 149.600 100.190 153.600 ;
    END
  END dout0[4]
  PIN dout0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 91.840 142.880 92.440 ;
    END
  END dout0[5]
  PIN dout0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 106.350 149.600 106.630 153.600 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 109.570 149.600 109.850 153.600 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.880 44.240 142.880 44.840 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 70.930 149.600 71.210 153.600 ;
    END
  END dout0[9]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 137.270 141.525 ;
      LAYER li1 ;
        RECT 5.520 10.795 137.080 141.525 ;
      LAYER met1 ;
        RECT 2.830 10.640 137.470 141.680 ;
      LAYER met2 ;
        RECT 2.860 149.320 15.910 149.600 ;
        RECT 16.750 149.320 67.430 149.600 ;
        RECT 68.270 149.320 70.650 149.600 ;
        RECT 71.490 149.320 77.090 149.600 ;
        RECT 77.930 149.320 86.750 149.600 ;
        RECT 87.590 149.320 93.190 149.600 ;
        RECT 94.030 149.320 99.630 149.600 ;
        RECT 100.470 149.320 106.070 149.600 ;
        RECT 106.910 149.320 109.290 149.600 ;
        RECT 110.130 149.320 137.440 149.600 ;
        RECT 2.860 4.280 137.440 149.320 ;
        RECT 2.860 4.000 73.870 4.280 ;
        RECT 74.710 4.000 99.630 4.280 ;
        RECT 100.470 4.000 112.510 4.280 ;
        RECT 113.350 4.000 137.440 4.280 ;
      LAYER met3 ;
        RECT 2.110 130.240 138.880 141.605 ;
        RECT 4.400 128.840 138.880 130.240 ;
        RECT 2.110 126.840 138.880 128.840 ;
        RECT 4.400 125.440 138.880 126.840 ;
        RECT 2.110 123.440 138.880 125.440 ;
        RECT 4.400 122.040 138.880 123.440 ;
        RECT 2.110 120.040 138.880 122.040 ;
        RECT 4.400 118.640 138.480 120.040 ;
        RECT 2.110 116.640 138.880 118.640 ;
        RECT 2.110 115.240 138.480 116.640 ;
        RECT 2.110 109.840 138.880 115.240 ;
        RECT 4.400 108.440 138.480 109.840 ;
        RECT 2.110 106.440 138.880 108.440 ;
        RECT 2.110 105.040 138.480 106.440 ;
        RECT 2.110 99.640 138.880 105.040 ;
        RECT 2.110 98.240 138.480 99.640 ;
        RECT 2.110 96.240 138.880 98.240 ;
        RECT 2.110 94.840 138.480 96.240 ;
        RECT 2.110 92.840 138.880 94.840 ;
        RECT 2.110 91.440 138.480 92.840 ;
        RECT 2.110 89.440 138.880 91.440 ;
        RECT 2.110 88.040 138.480 89.440 ;
        RECT 2.110 82.640 138.880 88.040 ;
        RECT 2.110 81.240 138.480 82.640 ;
        RECT 2.110 79.240 138.880 81.240 ;
        RECT 2.110 77.840 138.480 79.240 ;
        RECT 2.110 72.440 138.880 77.840 ;
        RECT 2.110 71.040 138.480 72.440 ;
        RECT 2.110 69.040 138.880 71.040 ;
        RECT 2.110 67.640 138.480 69.040 ;
        RECT 2.110 65.640 138.880 67.640 ;
        RECT 2.110 64.240 138.480 65.640 ;
        RECT 2.110 58.840 138.880 64.240 ;
        RECT 2.110 57.440 138.480 58.840 ;
        RECT 2.110 55.440 138.880 57.440 ;
        RECT 2.110 54.040 138.480 55.440 ;
        RECT 2.110 52.040 138.880 54.040 ;
        RECT 2.110 50.640 138.480 52.040 ;
        RECT 2.110 48.640 138.880 50.640 ;
        RECT 2.110 47.240 138.480 48.640 ;
        RECT 2.110 45.240 138.880 47.240 ;
        RECT 4.400 43.840 138.480 45.240 ;
        RECT 2.110 41.840 138.880 43.840 ;
        RECT 4.400 40.440 138.480 41.840 ;
        RECT 2.110 38.440 138.880 40.440 ;
        RECT 2.110 37.040 138.480 38.440 ;
        RECT 2.110 31.640 138.880 37.040 ;
        RECT 4.400 30.240 138.880 31.640 ;
        RECT 2.110 28.240 138.880 30.240 ;
        RECT 4.400 26.840 138.480 28.240 ;
        RECT 2.110 24.840 138.880 26.840 ;
        RECT 2.110 23.440 138.480 24.840 ;
        RECT 2.110 10.715 138.880 23.440 ;
      LAYER met4 ;
        RECT 1.710 19.215 20.640 139.225 ;
        RECT 23.040 19.215 23.940 139.225 ;
        RECT 26.340 19.215 130.345 139.225 ;
      LAYER met5 ;
        RECT 1.500 51.900 128.220 101.100 ;
  END
END cust_rom
END LIBRARY

