VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MACRO rom_high
   CLASS BLOCK ;
   SIZE 102.91 BY 111.56 ;
   SYMMETRY X Y R90 ;
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 7.09 -7.1 7.47 ;
      END
   END clk0
   PIN cs0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  17.755 -7.48 18.135 -7.1 ;
      END
   END cs0
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  21.97 -7.48 22.35 -7.1 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  24.01 -7.48 24.39 -7.1 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 24.71 -7.1 25.09 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 25.455 -7.1 25.835 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 26.145 -7.1 26.525 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 23.24 -7.1 23.62 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 26.835 -7.1 27.215 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  -7.48 22.55 -7.1 22.93 ;
      END
   END addr0[7]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  52.895 -7.48 53.275 -7.1 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  54.435 -7.48 54.815 -7.1 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  55.975 -7.48 56.355 -7.1 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  57.515 -7.48 57.895 -7.1 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  59.055 -7.48 59.435 -7.1 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  60.595 -7.48 60.975 -7.1 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  61.355 -7.48 61.735 -7.1 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  63.675 -7.48 64.055 -7.1 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  65.215 -7.48 65.595 -7.1 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  66.755 -7.48 67.135 -7.1 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  68.295 -7.48 68.675 -7.1 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  69.835 -7.48 70.215 -7.1 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  71.375 -7.48 71.755 -7.1 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  72.915 -7.48 73.295 -7.1 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  74.455 -7.48 74.835 -7.1 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  75.905 -7.48 76.285 -7.1 ;
      END
   END dout0[15]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  -7.48 -7.48 110.39 -5.74 ;
         LAYER met3 ;
         RECT  -7.48 117.3 110.39 119.04 ;
         LAYER met4 ;
         RECT  108.65 -7.48 110.39 119.04 ;
         LAYER met4 ;
         RECT  -7.48 -7.48 -5.74 119.04 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  105.17 -4.0 106.91 115.56 ;
         LAYER met3 ;
         RECT  -4.0 -4.0 106.91 -2.26 ;
         LAYER met4 ;
         RECT  -4.0 -4.0 -2.26 115.56 ;
         LAYER met3 ;
         RECT  -4.0 113.82 106.91 115.56 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 102.29 110.94 ;
   LAYER  met2 ;
      RECT  0.62 0.62 102.29 110.94 ;
   LAYER  met3 ;
      RECT  0.62 0.62 102.29 110.94 ;
   LAYER  met4 ;
      RECT  0.62 0.62 102.29 110.94 ;
   END
END    rom_high
END    LIBRARY
