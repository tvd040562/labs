magic
tech sky130A
magscale 1 2
timestamp 1727310469
<< viali >>
rect 13093 17833 13127 17867
rect 14197 17833 14231 17867
rect 13369 17561 13403 17595
rect 14473 17561 14507 17595
rect 14749 17289 14783 17323
rect 11897 17153 11931 17187
rect 12164 17153 12198 17187
rect 13369 17153 13403 17187
rect 13636 17153 13670 17187
rect 15393 17153 15427 17187
rect 16497 17153 16531 17187
rect 16773 17153 16807 17187
rect 13277 16949 13311 16983
rect 14841 16949 14875 16983
rect 15853 16949 15887 16983
rect 16957 16949 16991 16983
rect 12541 16745 12575 16779
rect 17049 16745 17083 16779
rect 13737 16609 13771 16643
rect 15669 16609 15703 16643
rect 12725 16541 12759 16575
rect 13093 16541 13127 16575
rect 14289 16541 14323 16575
rect 14657 16541 14691 16575
rect 15577 16541 15611 16575
rect 12817 16473 12851 16507
rect 12909 16473 12943 16507
rect 13185 16473 13219 16507
rect 14473 16473 14507 16507
rect 14565 16473 14599 16507
rect 15914 16473 15948 16507
rect 14841 16405 14875 16439
rect 14933 16405 14967 16439
rect 13645 16201 13679 16235
rect 15945 16201 15979 16235
rect 10701 16133 10735 16167
rect 9965 16065 9999 16099
rect 10241 16065 10275 16099
rect 10885 16065 10919 16099
rect 12081 16065 12115 16099
rect 12265 16065 12299 16099
rect 12357 16065 12391 16099
rect 13093 16065 13127 16099
rect 13277 16065 13311 16099
rect 13369 16065 13403 16099
rect 13461 16065 13495 16099
rect 13921 16065 13955 16099
rect 14105 16065 14139 16099
rect 14197 16065 14231 16099
rect 14289 16065 14323 16099
rect 14565 16065 14599 16099
rect 14821 16065 14855 16099
rect 16773 16065 16807 16099
rect 10057 15997 10091 16031
rect 10517 15929 10551 15963
rect 12541 15929 12575 15963
rect 14473 15929 14507 15963
rect 10241 15861 10275 15895
rect 10425 15861 10459 15895
rect 12265 15861 12299 15895
rect 16957 15861 16991 15895
rect 5917 15657 5951 15691
rect 7849 15657 7883 15691
rect 8309 15657 8343 15691
rect 9137 15657 9171 15691
rect 9505 15657 9539 15691
rect 10425 15657 10459 15691
rect 10609 15657 10643 15691
rect 11345 15657 11379 15691
rect 12265 15657 12299 15691
rect 12633 15657 12667 15691
rect 11713 15589 11747 15623
rect 7941 15521 7975 15555
rect 10241 15521 10275 15555
rect 15669 15521 15703 15555
rect 5641 15453 5675 15487
rect 5825 15453 5859 15487
rect 5917 15453 5951 15487
rect 8125 15453 8159 15487
rect 9137 15453 9171 15487
rect 9321 15453 9355 15487
rect 10425 15453 10459 15487
rect 11345 15453 11379 15487
rect 11529 15453 11563 15487
rect 12541 15453 12575 15487
rect 12633 15453 12667 15487
rect 7849 15385 7883 15419
rect 10149 15385 10183 15419
rect 11805 15385 11839 15419
rect 11989 15385 12023 15419
rect 15914 15385 15948 15419
rect 6101 15317 6135 15351
rect 12173 15317 12207 15351
rect 17049 15317 17083 15351
rect 12357 15113 12391 15147
rect 13645 15113 13679 15147
rect 14565 15113 14599 15147
rect 15761 15113 15795 15147
rect 16957 15113 16991 15147
rect 11897 15045 11931 15079
rect 13185 15045 13219 15079
rect 15393 15045 15427 15079
rect 5641 14977 5675 15011
rect 5825 14977 5859 15011
rect 6561 14977 6595 15011
rect 6837 14977 6871 15011
rect 7205 14977 7239 15011
rect 7481 14977 7515 15011
rect 7849 14977 7883 15011
rect 8033 14977 8067 15011
rect 9321 14977 9355 15011
rect 9597 14977 9631 15011
rect 10977 14977 11011 15011
rect 11161 14977 11195 15011
rect 12081 14977 12115 15011
rect 12173 14977 12207 15011
rect 13461 14977 13495 15011
rect 13921 14977 13955 15011
rect 14105 14977 14139 15011
rect 14197 14977 14231 15011
rect 15209 14977 15243 15011
rect 15485 14977 15519 15011
rect 15577 14977 15611 15011
rect 15853 14977 15887 15011
rect 16497 14977 16531 15011
rect 16773 14977 16807 15011
rect 6653 14909 6687 14943
rect 7297 14909 7331 14943
rect 9505 14909 9539 14943
rect 13277 14909 13311 14943
rect 14289 14909 14323 14943
rect 9781 14841 9815 14875
rect 6009 14773 6043 14807
rect 6377 14773 6411 14807
rect 6561 14773 6595 14807
rect 7205 14773 7239 14807
rect 7665 14773 7699 14807
rect 8217 14773 8251 14807
rect 9321 14773 9355 14807
rect 11345 14773 11379 14807
rect 11989 14773 12023 14807
rect 13185 14773 13219 14807
rect 13737 14773 13771 14807
rect 14197 14773 14231 14807
rect 8493 14569 8527 14603
rect 11437 14569 11471 14603
rect 11805 14569 11839 14603
rect 12265 14569 12299 14603
rect 13461 14569 13495 14603
rect 12633 14501 12667 14535
rect 8401 14433 8435 14467
rect 11529 14433 11563 14467
rect 13553 14433 13587 14467
rect 15301 14433 15335 14467
rect 8217 14365 8251 14399
rect 8493 14365 8527 14399
rect 9137 14365 9171 14399
rect 9321 14365 9355 14399
rect 11437 14365 11471 14399
rect 12265 14365 12299 14399
rect 12449 14365 12483 14399
rect 13461 14365 13495 14399
rect 8953 14297 8987 14331
rect 15568 14297 15602 14331
rect 8677 14229 8711 14263
rect 13829 14229 13863 14263
rect 16681 14229 16715 14263
rect 3617 14025 3651 14059
rect 10149 14025 10183 14059
rect 11897 14025 11931 14059
rect 14381 14025 14415 14059
rect 15669 14025 15703 14059
rect 3249 13957 3283 13991
rect 7113 13957 7147 13991
rect 7481 13957 7515 13991
rect 8861 13957 8895 13991
rect 10425 13957 10459 13991
rect 3065 13889 3099 13923
rect 3341 13889 3375 13923
rect 3433 13889 3467 13923
rect 4353 13889 4387 13923
rect 4537 13889 4571 13923
rect 6837 13889 6871 13923
rect 7021 13889 7055 13923
rect 7205 13889 7239 13923
rect 7665 13889 7699 13923
rect 8401 13889 8435 13923
rect 8585 13889 8619 13923
rect 9137 13889 9171 13923
rect 9689 13889 9723 13923
rect 9965 13889 9999 13923
rect 10609 13889 10643 13923
rect 11529 13889 11563 13923
rect 13921 13889 13955 13923
rect 14197 13889 14231 13923
rect 14473 13889 14507 13923
rect 14657 13889 14691 13923
rect 15117 13889 15151 13923
rect 15301 13889 15335 13923
rect 15393 13889 15427 13923
rect 15485 13889 15519 13923
rect 15853 13889 15887 13923
rect 16497 13889 16531 13923
rect 16773 13889 16807 13923
rect 4721 13821 4755 13855
rect 7849 13821 7883 13855
rect 8769 13821 8803 13855
rect 9045 13821 9079 13855
rect 9873 13821 9907 13855
rect 10793 13821 10827 13855
rect 11621 13821 11655 13855
rect 14013 13821 14047 13855
rect 7389 13685 7423 13719
rect 9137 13685 9171 13719
rect 9321 13685 9355 13719
rect 9689 13685 9723 13719
rect 11529 13685 11563 13719
rect 13921 13685 13955 13719
rect 14473 13685 14507 13719
rect 14841 13685 14875 13719
rect 16957 13685 16991 13719
rect 4813 13481 4847 13515
rect 5457 13481 5491 13515
rect 6377 13481 6411 13515
rect 7021 13481 7055 13515
rect 8033 13481 8067 13515
rect 9781 13481 9815 13515
rect 9965 13481 9999 13515
rect 10517 13481 10551 13515
rect 10885 13481 10919 13515
rect 12541 13481 12575 13515
rect 13001 13481 13035 13515
rect 14105 13481 14139 13515
rect 3617 13413 3651 13447
rect 14565 13413 14599 13447
rect 10517 13345 10551 13379
rect 12633 13345 12667 13379
rect 14289 13345 14323 13379
rect 15669 13345 15703 13379
rect 3111 13277 3145 13311
rect 3433 13277 3467 13311
rect 3985 13277 4019 13311
rect 4261 13277 4295 13311
rect 4537 13277 4571 13311
rect 4629 13277 4663 13311
rect 4905 13277 4939 13311
rect 5273 13277 5307 13311
rect 5641 13277 5675 13311
rect 5825 13277 5859 13311
rect 6009 13277 6043 13311
rect 6469 13277 6503 13311
rect 6561 13277 6595 13311
rect 7021 13277 7055 13311
rect 7113 13277 7147 13311
rect 7389 13277 7423 13311
rect 7537 13277 7571 13311
rect 7665 13277 7699 13311
rect 7895 13277 7929 13311
rect 9597 13277 9631 13311
rect 9781 13277 9815 13311
rect 10701 13277 10735 13311
rect 12541 13277 12575 13311
rect 12817 13277 12851 13311
rect 14381 13277 14415 13311
rect 15025 13277 15059 13311
rect 15393 13277 15427 13311
rect 3249 13209 3283 13243
rect 3341 13209 3375 13243
rect 3801 13209 3835 13243
rect 4445 13209 4479 13243
rect 5089 13209 5123 13243
rect 5181 13209 5215 13243
rect 5917 13209 5951 13243
rect 6285 13209 6319 13243
rect 7297 13209 7331 13243
rect 7757 13209 7791 13243
rect 10425 13209 10459 13243
rect 14105 13209 14139 13243
rect 15209 13209 15243 13243
rect 15301 13209 15335 13243
rect 15914 13209 15948 13243
rect 4169 13141 4203 13175
rect 6193 13141 6227 13175
rect 6745 13141 6779 13175
rect 6837 13141 6871 13175
rect 15577 13141 15611 13175
rect 17049 13141 17083 13175
rect 3801 12937 3835 12971
rect 10609 12937 10643 12971
rect 12817 12937 12851 12971
rect 14657 12937 14691 12971
rect 15853 12937 15887 12971
rect 16957 12937 16991 12971
rect 3525 12869 3559 12903
rect 4813 12869 4847 12903
rect 12357 12869 12391 12903
rect 3249 12801 3283 12835
rect 3433 12801 3467 12835
rect 3617 12801 3651 12835
rect 4537 12801 4571 12835
rect 4721 12801 4755 12835
rect 4905 12801 4939 12835
rect 5549 12801 5583 12835
rect 5733 12801 5767 12835
rect 5825 12801 5859 12835
rect 5917 12801 5951 12835
rect 7113 12801 7147 12835
rect 7297 12801 7331 12835
rect 7389 12801 7423 12835
rect 7481 12801 7515 12835
rect 10793 12801 10827 12835
rect 10977 12801 11011 12835
rect 12633 12801 12667 12835
rect 12909 12801 12943 12835
rect 13001 12801 13035 12835
rect 14289 12801 14323 12835
rect 14473 12801 14507 12835
rect 16497 12801 16531 12835
rect 16773 12801 16807 12835
rect 12541 12733 12575 12767
rect 5089 12665 5123 12699
rect 13277 12665 13311 12699
rect 6101 12597 6135 12631
rect 7665 12597 7699 12631
rect 12357 12597 12391 12631
rect 12909 12597 12943 12631
rect 2973 12393 3007 12427
rect 6561 12393 6595 12427
rect 7205 12393 7239 12427
rect 7941 12393 7975 12427
rect 8769 12393 8803 12427
rect 9229 12393 9263 12427
rect 9597 12393 9631 12427
rect 10609 12393 10643 12427
rect 11161 12393 11195 12427
rect 11437 12393 11471 12427
rect 12541 12393 12575 12427
rect 10793 12325 10827 12359
rect 6469 12257 6503 12291
rect 9137 12257 9171 12291
rect 9689 12257 9723 12291
rect 10425 12257 10459 12291
rect 11621 12257 11655 12291
rect 12449 12257 12483 12291
rect 2421 12189 2455 12223
rect 2697 12189 2731 12223
rect 2789 12189 2823 12223
rect 3065 12189 3099 12223
rect 3249 12189 3283 12223
rect 3433 12189 3467 12223
rect 4261 12189 4295 12223
rect 4537 12189 4571 12223
rect 4629 12189 4663 12223
rect 4905 12189 4939 12223
rect 5273 12189 5307 12223
rect 6285 12189 6319 12223
rect 6561 12189 6595 12223
rect 6653 12189 6687 12223
rect 6929 12189 6963 12223
rect 7021 12189 7055 12223
rect 7297 12189 7331 12223
rect 7390 12189 7424 12223
rect 7762 12189 7796 12223
rect 8401 12189 8435 12223
rect 9321 12189 9355 12223
rect 9873 12189 9907 12223
rect 10609 12189 10643 12223
rect 11069 12189 11103 12223
rect 11161 12189 11195 12223
rect 11444 12189 11478 12223
rect 11713 12189 11747 12223
rect 12265 12189 12299 12223
rect 12541 12189 12575 12223
rect 15025 12189 15059 12223
rect 15301 12189 15335 12223
rect 15393 12189 15427 12223
rect 15669 12189 15703 12223
rect 2605 12121 2639 12155
rect 3341 12121 3375 12155
rect 4445 12121 4479 12155
rect 5089 12121 5123 12155
rect 5181 12121 5215 12155
rect 6837 12121 6871 12155
rect 7573 12121 7607 12155
rect 7665 12121 7699 12155
rect 8585 12121 8619 12155
rect 9045 12121 9079 12155
rect 9597 12121 9631 12155
rect 10333 12121 10367 12155
rect 10885 12121 10919 12155
rect 15209 12121 15243 12155
rect 15914 12121 15948 12155
rect 3617 12053 3651 12087
rect 4813 12053 4847 12087
rect 5457 12053 5491 12087
rect 6101 12053 6135 12087
rect 9505 12053 9539 12087
rect 10057 12053 10091 12087
rect 11345 12053 11379 12087
rect 11897 12053 11931 12087
rect 12725 12053 12759 12087
rect 15577 12053 15611 12087
rect 17049 12053 17083 12087
rect 3801 11849 3835 11883
rect 5089 11849 5123 11883
rect 6377 11849 6411 11883
rect 14197 11849 14231 11883
rect 15853 11849 15887 11883
rect 3433 11781 3467 11815
rect 4813 11781 4847 11815
rect 10609 11781 10643 11815
rect 13553 11781 13587 11815
rect 14473 11781 14507 11815
rect 3249 11713 3283 11747
rect 3525 11713 3559 11747
rect 3617 11713 3651 11747
rect 4537 11713 4571 11747
rect 4721 11713 4755 11747
rect 4905 11713 4939 11747
rect 6515 11713 6549 11747
rect 6653 11713 6687 11747
rect 6745 11713 6779 11747
rect 6928 11713 6962 11747
rect 7014 11713 7048 11747
rect 7665 11713 7699 11747
rect 8677 11713 8711 11747
rect 8861 11713 8895 11747
rect 9045 11713 9079 11747
rect 10517 11713 10551 11747
rect 10885 11713 10919 11747
rect 13369 11713 13403 11747
rect 13829 11713 13863 11747
rect 14749 11713 14783 11747
rect 15025 11713 15059 11747
rect 16497 11713 16531 11747
rect 16865 11713 16899 11747
rect 10793 11645 10827 11679
rect 13921 11645 13955 11679
rect 14565 11645 14599 11679
rect 15117 11645 15151 11679
rect 16681 11645 16715 11679
rect 7481 11577 7515 11611
rect 10885 11509 10919 11543
rect 11069 11509 11103 11543
rect 13737 11509 13771 11543
rect 13829 11509 13863 11543
rect 14473 11509 14507 11543
rect 14933 11509 14967 11543
rect 15025 11509 15059 11543
rect 15393 11509 15427 11543
rect 7021 11305 7055 11339
rect 8493 11305 8527 11339
rect 11529 11305 11563 11339
rect 12449 11305 12483 11339
rect 13093 11305 13127 11339
rect 13461 11305 13495 11339
rect 14105 11305 14139 11339
rect 14473 11305 14507 11339
rect 6009 11237 6043 11271
rect 7849 11237 7883 11271
rect 15669 11169 15703 11203
rect 4813 11101 4847 11135
rect 5089 11101 5123 11135
rect 5181 11101 5215 11135
rect 5457 11101 5491 11135
rect 5733 11101 5767 11135
rect 5825 11101 5859 11135
rect 7113 11101 7147 11135
rect 7297 11101 7331 11135
rect 7481 11101 7515 11135
rect 7689 11101 7723 11135
rect 7941 11101 7975 11135
rect 8309 11101 8343 11135
rect 9505 11101 9539 11135
rect 13093 11101 13127 11135
rect 13185 11101 13219 11135
rect 14105 11101 14139 11135
rect 14197 11101 14231 11135
rect 15025 11101 15059 11135
rect 15301 11101 15335 11135
rect 15393 11101 15427 11135
rect 4997 11033 5031 11067
rect 5641 11033 5675 11067
rect 7573 11033 7607 11067
rect 8125 11033 8159 11067
rect 8217 11033 8251 11067
rect 9137 11033 9171 11067
rect 9321 11033 9355 11067
rect 10241 11033 10275 11067
rect 12081 11033 12115 11067
rect 12265 11033 12299 11067
rect 15209 11033 15243 11067
rect 15914 11033 15948 11067
rect 5365 10965 5399 10999
rect 15577 10965 15611 10999
rect 17049 10965 17083 10999
rect 3341 10761 3375 10795
rect 5457 10761 5491 10795
rect 7389 10761 7423 10795
rect 10793 10761 10827 10795
rect 15853 10761 15887 10795
rect 16957 10761 16991 10795
rect 2973 10693 3007 10727
rect 3617 10693 3651 10727
rect 4261 10693 4295 10727
rect 7021 10693 7055 10727
rect 7665 10693 7699 10727
rect 8585 10693 8619 10727
rect 13277 10693 13311 10727
rect 2789 10625 2823 10659
rect 3065 10625 3099 10659
rect 3157 10625 3191 10659
rect 3433 10625 3467 10659
rect 3709 10625 3743 10659
rect 3801 10625 3835 10659
rect 4077 10625 4111 10659
rect 4445 10625 4479 10659
rect 4905 10625 4939 10659
rect 5089 10625 5123 10659
rect 5181 10625 5215 10659
rect 5273 10625 5307 10659
rect 6837 10625 6871 10659
rect 7113 10625 7147 10659
rect 7205 10625 7239 10659
rect 7481 10625 7515 10659
rect 7757 10625 7791 10659
rect 7895 10625 7929 10659
rect 10425 10625 10459 10659
rect 10517 10625 10551 10659
rect 11529 10625 11563 10659
rect 13553 10625 13587 10659
rect 16497 10625 16531 10659
rect 16773 10625 16807 10659
rect 10333 10557 10367 10591
rect 11621 10557 11655 10591
rect 13461 10557 13495 10591
rect 3985 10489 4019 10523
rect 11897 10489 11931 10523
rect 8033 10421 8067 10455
rect 10609 10421 10643 10455
rect 11529 10421 11563 10455
rect 13277 10421 13311 10455
rect 13737 10421 13771 10455
rect 2789 10217 2823 10251
rect 8217 10217 8251 10251
rect 8953 10217 8987 10251
rect 9505 10217 9539 10251
rect 11161 10217 11195 10251
rect 12265 10217 12299 10251
rect 13553 10217 13587 10251
rect 13737 10217 13771 10251
rect 14565 10217 14599 10251
rect 16957 10217 16991 10251
rect 4997 10149 5031 10183
rect 6561 10149 6595 10183
rect 7573 10149 7607 10183
rect 9413 10149 9447 10183
rect 5641 10081 5675 10115
rect 7665 10081 7699 10115
rect 9137 10081 9171 10115
rect 14657 10081 14691 10115
rect 2605 10013 2639 10047
rect 3801 10013 3835 10047
rect 4169 10013 4203 10047
rect 4445 10013 4479 10047
rect 4813 10013 4847 10047
rect 5917 10013 5951 10047
rect 6009 10013 6043 10047
rect 6193 10013 6227 10047
rect 6377 10013 6411 10047
rect 7021 10013 7055 10047
rect 7297 10013 7331 10047
rect 7389 10013 7423 10047
rect 8033 10013 8067 10047
rect 8401 10013 8435 10047
rect 9229 10013 9263 10047
rect 9689 10013 9723 10047
rect 12081 10013 12115 10047
rect 12817 10013 12851 10047
rect 13461 10013 13495 10047
rect 13553 10013 13587 10047
rect 14565 10013 14599 10047
rect 16405 10013 16439 10047
rect 16773 10013 16807 10047
rect 2145 9945 2179 9979
rect 2513 9945 2547 9979
rect 3985 9945 4019 9979
rect 4077 9945 4111 9979
rect 4629 9945 4663 9979
rect 4721 9945 4755 9979
rect 6285 9945 6319 9979
rect 6837 9945 6871 9979
rect 7205 9945 7239 9979
rect 7849 9945 7883 9979
rect 8953 9945 8987 9979
rect 9873 9945 9907 9979
rect 11345 9945 11379 9979
rect 11529 9945 11563 9979
rect 11897 9945 11931 9979
rect 13001 9945 13035 9979
rect 13277 9945 13311 9979
rect 2421 9877 2455 9911
rect 4353 9877 4387 9911
rect 6745 9877 6779 9911
rect 8585 9877 8619 9911
rect 13185 9877 13219 9911
rect 14933 9877 14967 9911
rect 16589 9877 16623 9911
rect 2421 9673 2455 9707
rect 2881 9673 2915 9707
rect 2513 9605 2547 9639
rect 6377 9605 6411 9639
rect 7573 9605 7607 9639
rect 7665 9605 7699 9639
rect 8217 9605 8251 9639
rect 8309 9605 8343 9639
rect 9229 9605 9263 9639
rect 9597 9605 9631 9639
rect 9873 9605 9907 9639
rect 11713 9605 11747 9639
rect 13829 9605 13863 9639
rect 2329 9537 2363 9571
rect 3065 9537 3099 9571
rect 6653 9537 6687 9571
rect 7389 9537 7423 9571
rect 7757 9537 7791 9571
rect 8033 9537 8067 9571
rect 8401 9537 8435 9571
rect 8677 9537 8711 9571
rect 8953 9537 8987 9571
rect 9413 9537 9447 9571
rect 10149 9537 10183 9571
rect 10885 9537 10919 9571
rect 11897 9537 11931 9571
rect 13645 9537 13679 9571
rect 14565 9537 14599 9571
rect 15117 9537 15151 9571
rect 15384 9537 15418 9571
rect 5457 9469 5491 9503
rect 5733 9469 5767 9503
rect 6469 9469 6503 9503
rect 8769 9469 8803 9503
rect 9965 9469 9999 9503
rect 10977 9469 11011 9503
rect 14657 9469 14691 9503
rect 6837 9401 6871 9435
rect 9137 9401 9171 9435
rect 10333 9401 10367 9435
rect 11253 9401 11287 9435
rect 6653 9333 6687 9367
rect 7941 9333 7975 9367
rect 8585 9333 8619 9367
rect 8677 9333 8711 9367
rect 9873 9333 9907 9367
rect 11069 9333 11103 9367
rect 11529 9333 11563 9367
rect 14013 9333 14047 9367
rect 14749 9333 14783 9367
rect 14933 9333 14967 9367
rect 16497 9333 16531 9367
rect 5457 9129 5491 9163
rect 8309 9129 8343 9163
rect 13369 9129 13403 9163
rect 13737 9129 13771 9163
rect 14105 9129 14139 9163
rect 14565 9129 14599 9163
rect 16129 9129 16163 9163
rect 3065 9061 3099 9095
rect 4445 9061 4479 9095
rect 7113 9061 7147 9095
rect 2973 8993 3007 9027
rect 4077 8993 4111 9027
rect 8309 8993 8343 9027
rect 13369 8993 13403 9027
rect 14197 8993 14231 9027
rect 16865 8993 16899 9027
rect 2237 8925 2271 8959
rect 3249 8925 3283 8959
rect 3341 8925 3375 8959
rect 3801 8925 3835 8959
rect 4905 8925 4939 8959
rect 5273 8925 5307 8959
rect 5549 8925 5583 8959
rect 5733 8925 5767 8959
rect 5917 8925 5951 8959
rect 6561 8925 6595 8959
rect 6837 8925 6871 8959
rect 6929 8925 6963 8959
rect 7481 8925 7515 8959
rect 7757 8925 7791 8959
rect 7849 8925 7883 8959
rect 8493 8925 8527 8959
rect 11253 8925 11287 8959
rect 13553 8925 13587 8959
rect 14105 8925 14139 8959
rect 14381 8925 14415 8959
rect 15577 8925 15611 8959
rect 15853 8925 15887 8959
rect 15945 8925 15979 8959
rect 16313 8925 16347 8959
rect 2329 8857 2363 8891
rect 2421 8857 2455 8891
rect 4261 8857 4295 8891
rect 5089 8857 5123 8891
rect 5181 8857 5215 8891
rect 5825 8857 5859 8891
rect 6745 8857 6779 8891
rect 7665 8857 7699 8891
rect 8217 8857 8251 8891
rect 11069 8857 11103 8891
rect 13277 8857 13311 8891
rect 15761 8857 15795 8891
rect 2789 8789 2823 8823
rect 3525 8789 3559 8823
rect 4169 8789 4203 8823
rect 6101 8789 6135 8823
rect 8033 8789 8067 8823
rect 8677 8789 8711 8823
rect 11437 8789 11471 8823
rect 2421 8585 2455 8619
rect 2789 8585 2823 8619
rect 8217 8585 8251 8619
rect 10701 8585 10735 8619
rect 11897 8585 11931 8619
rect 13001 8585 13035 8619
rect 13461 8585 13495 8619
rect 13921 8585 13955 8619
rect 16957 8585 16991 8619
rect 2237 8517 2271 8551
rect 2329 8517 2363 8551
rect 5089 8517 5123 8551
rect 7757 8517 7791 8551
rect 9505 8517 9539 8551
rect 9781 8517 9815 8551
rect 15393 8517 15427 8551
rect 3341 8449 3375 8483
rect 4813 8449 4847 8483
rect 4997 8449 5031 8483
rect 5181 8449 5215 8483
rect 7481 8449 7515 8483
rect 7665 8449 7699 8483
rect 7849 8449 7883 8483
rect 8309 8449 8343 8483
rect 9321 8449 9355 8483
rect 10057 8449 10091 8483
rect 10333 8449 10367 8483
rect 10517 8449 10551 8483
rect 11529 8449 11563 8483
rect 12541 8449 12575 8483
rect 12817 8449 12851 8483
rect 13093 8449 13127 8483
rect 13553 8449 13587 8483
rect 14013 8449 14047 8483
rect 14105 8449 14139 8483
rect 15209 8449 15243 8483
rect 15485 8449 15519 8483
rect 15577 8449 15611 8483
rect 15853 8449 15887 8483
rect 16773 8449 16807 8483
rect 2973 8381 3007 8415
rect 9689 8381 9723 8415
rect 9965 8381 9999 8415
rect 11621 8381 11655 8415
rect 12725 8381 12759 8415
rect 13185 8381 13219 8415
rect 13645 8381 13679 8415
rect 14289 8381 14323 8415
rect 16497 8381 16531 8415
rect 3525 8313 3559 8347
rect 5365 8313 5399 8347
rect 8033 8313 8067 8347
rect 14013 8313 14047 8347
rect 9781 8245 9815 8279
rect 10241 8245 10275 8279
rect 11529 8245 11563 8279
rect 12633 8245 12667 8279
rect 13093 8245 13127 8279
rect 13737 8245 13771 8279
rect 15761 8245 15795 8279
rect 3617 8041 3651 8075
rect 6009 8041 6043 8075
rect 6745 8041 6779 8075
rect 10977 8041 11011 8075
rect 11437 8041 11471 8075
rect 11713 8041 11747 8075
rect 13553 8041 13587 8075
rect 14565 8041 14599 8075
rect 15025 8041 15059 8075
rect 15393 8041 15427 8075
rect 17049 8041 17083 8075
rect 7849 7973 7883 8007
rect 8493 7973 8527 8007
rect 11253 7973 11287 8007
rect 14381 7973 14415 8007
rect 2237 7905 2271 7939
rect 4629 7905 4663 7939
rect 10885 7905 10919 7939
rect 13369 7905 13403 7939
rect 14473 7905 14507 7939
rect 15117 7905 15151 7939
rect 2053 7837 2087 7871
rect 2605 7837 2639 7871
rect 3433 7837 3467 7871
rect 3893 7837 3927 7871
rect 3985 7837 4019 7871
rect 4721 7837 4755 7871
rect 4905 7837 4939 7871
rect 4997 7837 5031 7871
rect 5089 7837 5123 7871
rect 5365 7837 5399 7871
rect 5549 7837 5583 7871
rect 5825 7837 5859 7871
rect 6101 7837 6135 7871
rect 6285 7837 6319 7871
rect 6561 7837 6595 7871
rect 7205 7837 7239 7871
rect 7353 7837 7387 7871
rect 7573 7837 7607 7871
rect 7709 7837 7743 7871
rect 7941 7837 7975 7871
rect 8125 7837 8159 7871
rect 8217 7837 8251 7871
rect 8309 7837 8343 7871
rect 10701 7837 10735 7871
rect 11069 7837 11103 7871
rect 11345 7837 11379 7871
rect 11437 7837 11471 7871
rect 13553 7837 13587 7871
rect 14197 7837 14231 7871
rect 14657 7837 14691 7871
rect 15025 7837 15059 7871
rect 15669 7837 15703 7871
rect 15925 7837 15959 7871
rect 2789 7769 2823 7803
rect 4445 7769 4479 7803
rect 7481 7769 7515 7803
rect 10793 7769 10827 7803
rect 13277 7769 13311 7803
rect 2697 7701 2731 7735
rect 4077 7701 4111 7735
rect 5273 7701 5307 7735
rect 9229 7701 9263 7735
rect 13737 7701 13771 7735
rect 14933 7701 14967 7735
rect 1777 7497 1811 7531
rect 3893 7497 3927 7531
rect 3985 7497 4019 7531
rect 9321 7497 9355 7531
rect 10057 7497 10091 7531
rect 10517 7497 10551 7531
rect 12541 7497 12575 7531
rect 15945 7497 15979 7531
rect 16313 7497 16347 7531
rect 16957 7497 16991 7531
rect 3249 7429 3283 7463
rect 3433 7429 3467 7463
rect 3617 7429 3651 7463
rect 4077 7429 4111 7463
rect 4353 7429 4387 7463
rect 4721 7429 4755 7463
rect 5273 7429 5307 7463
rect 9689 7429 9723 7463
rect 11529 7429 11563 7463
rect 12633 7429 12667 7463
rect 12817 7429 12851 7463
rect 1961 7361 1995 7395
rect 2237 7361 2271 7395
rect 2513 7361 2547 7395
rect 2697 7361 2731 7395
rect 3065 7361 3099 7395
rect 4445 7361 4479 7395
rect 4629 7361 4663 7395
rect 4813 7361 4847 7395
rect 5089 7361 5123 7395
rect 5365 7361 5399 7395
rect 5457 7361 5491 7395
rect 8861 7361 8895 7395
rect 9137 7361 9171 7395
rect 9873 7361 9907 7395
rect 10149 7361 10183 7395
rect 11805 7361 11839 7395
rect 12081 7361 12115 7395
rect 12357 7361 12391 7395
rect 16129 7361 16163 7395
rect 16497 7361 16531 7395
rect 16773 7361 16807 7395
rect 2789 7293 2823 7327
rect 8953 7293 8987 7327
rect 10241 7293 10275 7327
rect 11621 7293 11655 7327
rect 12173 7293 12207 7327
rect 4997 7225 5031 7259
rect 11989 7225 12023 7259
rect 5641 7157 5675 7191
rect 9137 7157 9171 7191
rect 10149 7157 10183 7191
rect 11621 7157 11655 7191
rect 12081 7157 12115 7191
rect 13001 7157 13035 7191
rect 2789 6953 2823 6987
rect 8953 6953 8987 6987
rect 11161 6953 11195 6987
rect 11621 6953 11655 6987
rect 12449 6953 12483 6987
rect 12909 6953 12943 6987
rect 14381 6953 14415 6987
rect 14841 6953 14875 6987
rect 7941 6885 7975 6919
rect 9413 6885 9447 6919
rect 6101 6817 6135 6851
rect 7021 6817 7055 6851
rect 9045 6817 9079 6851
rect 9873 6817 9907 6851
rect 11253 6817 11287 6851
rect 12541 6817 12575 6851
rect 13093 6817 13127 6851
rect 13185 6817 13219 6851
rect 13277 6817 13311 6851
rect 1409 6749 1443 6783
rect 4813 6749 4847 6783
rect 4997 6749 5031 6783
rect 5181 6749 5215 6783
rect 5457 6749 5491 6783
rect 5641 6749 5675 6783
rect 5917 6749 5951 6783
rect 7389 6749 7423 6783
rect 7573 6749 7607 6783
rect 7665 6749 7699 6783
rect 7757 6749 7791 6783
rect 8033 6749 8067 6783
rect 8309 6749 8343 6783
rect 8401 6749 8435 6783
rect 9229 6749 9263 6783
rect 11437 6749 11471 6783
rect 12725 6749 12759 6783
rect 14565 6749 14599 6783
rect 14657 6749 14691 6783
rect 15669 6749 15703 6783
rect 1676 6681 1710 6715
rect 5089 6681 5123 6715
rect 7205 6681 7239 6715
rect 8217 6681 8251 6715
rect 8953 6681 8987 6715
rect 9505 6681 9539 6715
rect 9689 6681 9723 6715
rect 11161 6681 11195 6715
rect 12449 6681 12483 6715
rect 13461 6681 13495 6715
rect 14381 6681 14415 6715
rect 15914 6681 15948 6715
rect 5365 6613 5399 6647
rect 8585 6613 8619 6647
rect 13369 6613 13403 6647
rect 17049 6613 17083 6647
rect 1593 6409 1627 6443
rect 4261 6409 4295 6443
rect 7941 6409 7975 6443
rect 13737 6409 13771 6443
rect 15761 6409 15795 6443
rect 5365 6341 5399 6375
rect 7573 6341 7607 6375
rect 15393 6341 15427 6375
rect 1409 6273 1443 6307
rect 1869 6273 1903 6307
rect 3065 6273 3099 6307
rect 3341 6273 3375 6307
rect 3525 6273 3559 6307
rect 4077 6273 4111 6307
rect 4169 6273 4203 6307
rect 4629 6273 4663 6307
rect 5089 6273 5123 6307
rect 5273 6273 5307 6307
rect 5462 6273 5496 6307
rect 7435 6273 7469 6307
rect 7661 6273 7695 6307
rect 7757 6273 7791 6307
rect 8033 6273 8067 6307
rect 8217 6273 8251 6307
rect 8309 6273 8343 6307
rect 8401 6273 8435 6307
rect 9321 6273 9355 6307
rect 9505 6273 9539 6307
rect 13369 6273 13403 6307
rect 13645 6273 13679 6307
rect 13921 6273 13955 6307
rect 14105 6273 14139 6307
rect 15209 6273 15243 6307
rect 15485 6273 15519 6307
rect 15577 6273 15611 6307
rect 15853 6273 15887 6307
rect 16497 6273 16531 6307
rect 16773 6273 16807 6307
rect 3617 6205 3651 6239
rect 4813 6205 4847 6239
rect 13461 6205 13495 6239
rect 3893 6137 3927 6171
rect 8585 6137 8619 6171
rect 13185 6137 13219 6171
rect 16957 6137 16991 6171
rect 1685 6069 1719 6103
rect 5089 6069 5123 6103
rect 9321 6069 9355 6103
rect 9689 6069 9723 6103
rect 13645 6069 13679 6103
rect 2789 5865 2823 5899
rect 4445 5865 4479 5899
rect 8493 5865 8527 5899
rect 10609 5865 10643 5899
rect 11621 5865 11655 5899
rect 14105 5865 14139 5899
rect 14565 5865 14599 5899
rect 17049 5865 17083 5899
rect 7481 5797 7515 5831
rect 4261 5729 4295 5763
rect 5825 5729 5859 5763
rect 6193 5729 6227 5763
rect 11437 5729 11471 5763
rect 14197 5729 14231 5763
rect 1409 5661 1443 5695
rect 1676 5661 1710 5695
rect 4077 5661 4111 5695
rect 5549 5661 5583 5695
rect 5922 5661 5956 5695
rect 6101 5661 6135 5695
rect 6278 5661 6312 5695
rect 6377 5661 6411 5695
rect 6561 5661 6595 5695
rect 7297 5661 7331 5695
rect 7665 5661 7699 5695
rect 7849 5661 7883 5695
rect 8033 5661 8067 5695
rect 8309 5661 8343 5695
rect 9321 5661 9355 5695
rect 10057 5661 10091 5695
rect 10701 5661 10735 5695
rect 10793 5661 10827 5695
rect 11621 5661 11655 5695
rect 13553 5661 13587 5695
rect 14381 5661 14415 5695
rect 15025 5661 15059 5695
rect 15209 5661 15243 5695
rect 15393 5661 15427 5695
rect 15669 5661 15703 5695
rect 3801 5593 3835 5627
rect 5733 5593 5767 5627
rect 5825 5593 5859 5627
rect 7113 5593 7147 5627
rect 7941 5593 7975 5627
rect 10241 5593 10275 5627
rect 10517 5593 10551 5627
rect 11345 5593 11379 5627
rect 13737 5593 13771 5627
rect 13921 5593 13955 5627
rect 14105 5593 14139 5627
rect 15301 5593 15335 5627
rect 15914 5593 15948 5627
rect 4169 5525 4203 5559
rect 6561 5525 6595 5559
rect 7021 5525 7055 5559
rect 8217 5525 8251 5559
rect 9505 5525 9539 5559
rect 10425 5525 10459 5559
rect 10977 5525 11011 5559
rect 11805 5525 11839 5559
rect 15577 5525 15611 5559
rect 2789 5321 2823 5355
rect 3249 5321 3283 5355
rect 8677 5321 8711 5355
rect 10241 5321 10275 5355
rect 12081 5321 12115 5355
rect 15853 5321 15887 5355
rect 16957 5321 16991 5355
rect 2973 5253 3007 5287
rect 5549 5253 5583 5287
rect 7389 5253 7423 5287
rect 7481 5253 7515 5287
rect 8125 5253 8159 5287
rect 12265 5253 12299 5287
rect 1665 5185 1699 5219
rect 3341 5185 3375 5219
rect 3617 5185 3651 5219
rect 3709 5185 3743 5219
rect 3985 5185 4019 5219
rect 4169 5185 4203 5219
rect 4721 5185 4755 5219
rect 4813 5185 4847 5219
rect 4905 5185 4939 5219
rect 5089 5185 5123 5219
rect 5273 5185 5307 5219
rect 5457 5185 5491 5219
rect 5646 5185 5680 5219
rect 5917 5185 5951 5219
rect 6101 5185 6135 5219
rect 6377 5185 6411 5219
rect 6561 5185 6595 5219
rect 6653 5185 6687 5219
rect 6745 5185 6779 5219
rect 7205 5185 7239 5219
rect 7573 5185 7607 5219
rect 7849 5185 7883 5219
rect 8033 5185 8067 5219
rect 8217 5185 8251 5219
rect 8493 5185 8527 5219
rect 8953 5185 8987 5219
rect 9045 5185 9079 5219
rect 9229 5185 9263 5219
rect 9505 5185 9539 5219
rect 9781 5185 9815 5219
rect 10057 5185 10091 5219
rect 12449 5185 12483 5219
rect 12541 5185 12575 5219
rect 12725 5185 12759 5219
rect 15485 5185 15519 5219
rect 16773 5185 16807 5219
rect 1409 5117 1443 5151
rect 3157 5117 3191 5151
rect 4537 5117 4571 5151
rect 5549 5117 5583 5151
rect 9965 5117 9999 5151
rect 16497 5117 16531 5151
rect 3065 5049 3099 5083
rect 4445 5049 4479 5083
rect 7757 5049 7791 5083
rect 8401 5049 8435 5083
rect 9413 5049 9447 5083
rect 15669 5049 15703 5083
rect 6929 4981 6963 5015
rect 9689 4981 9723 5015
rect 10057 4981 10091 5015
rect 12725 4981 12759 5015
rect 2789 4777 2823 4811
rect 3525 4777 3559 4811
rect 3985 4777 4019 4811
rect 4721 4777 4755 4811
rect 7389 4777 7423 4811
rect 9321 4777 9355 4811
rect 17049 4777 17083 4811
rect 4445 4709 4479 4743
rect 8125 4709 8159 4743
rect 9597 4709 9631 4743
rect 6653 4641 6687 4675
rect 1409 4573 1443 4607
rect 3341 4573 3375 4607
rect 4077 4573 4111 4607
rect 4261 4573 4295 4607
rect 7205 4573 7239 4607
rect 7573 4573 7607 4607
rect 7757 4573 7791 4607
rect 7849 4573 7883 4607
rect 7941 4573 7975 4607
rect 8217 4573 8251 4607
rect 9689 4573 9723 4607
rect 9781 4573 9815 4607
rect 10057 4573 10091 4607
rect 11069 4573 11103 4607
rect 13645 4573 13679 4607
rect 13737 4573 13771 4607
rect 13921 4573 13955 4607
rect 14933 4573 14967 4607
rect 15025 4573 15059 4607
rect 15209 4573 15243 4607
rect 15393 4573 15427 4607
rect 15669 4573 15703 4607
rect 1676 4505 1710 4539
rect 3801 4505 3835 4539
rect 4629 4505 4663 4539
rect 6837 4505 6871 4539
rect 15301 4505 15335 4539
rect 15914 4505 15948 4539
rect 8401 4437 8435 4471
rect 9965 4437 9999 4471
rect 11253 4437 11287 4471
rect 13829 4437 13863 4471
rect 14749 4437 14783 4471
rect 15577 4437 15611 4471
rect 1593 4233 1627 4267
rect 1685 4233 1719 4267
rect 7113 4233 7147 4267
rect 7665 4233 7699 4267
rect 9939 4233 9973 4267
rect 10333 4233 10367 4267
rect 14933 4233 14967 4267
rect 15853 4233 15887 4267
rect 7817 4165 7851 4199
rect 8033 4165 8067 4199
rect 10149 4165 10183 4199
rect 10885 4165 10919 4199
rect 11161 4165 11195 4199
rect 11345 4165 11379 4199
rect 11897 4165 11931 4199
rect 12081 4165 12115 4199
rect 13369 4165 13403 4199
rect 13737 4165 13771 4199
rect 14105 4165 14139 4199
rect 1409 4097 1443 4131
rect 1869 4097 1903 4131
rect 6377 4097 6411 4131
rect 6561 4097 6595 4131
rect 6837 4097 6871 4131
rect 7297 4097 7331 4131
rect 9229 4097 9263 4131
rect 9413 4097 9447 4131
rect 10425 4097 10459 4131
rect 10517 4097 10551 4131
rect 13553 4097 13587 4131
rect 13829 4097 13863 4131
rect 14013 4097 14047 4131
rect 14289 4097 14323 4131
rect 14749 4097 14783 4131
rect 15025 4097 15059 4131
rect 15117 4097 15151 4131
rect 15761 4097 15795 4131
rect 16497 4097 16531 4131
rect 7389 4029 7423 4063
rect 7481 4029 7515 4063
rect 9321 4029 9355 4063
rect 10701 4029 10735 4063
rect 10977 4029 11011 4063
rect 13185 4029 13219 4063
rect 13461 4029 13495 4063
rect 13645 4029 13679 4063
rect 14473 4029 14507 4063
rect 7021 3961 7055 3995
rect 13829 3961 13863 3995
rect 7849 3893 7883 3927
rect 9781 3893 9815 3927
rect 9965 3893 9999 3927
rect 10609 3893 10643 3927
rect 12265 3893 12299 3927
rect 14565 3893 14599 3927
rect 6653 3689 6687 3723
rect 7113 3689 7147 3723
rect 7757 3689 7791 3723
rect 9137 3689 9171 3723
rect 10977 3689 11011 3723
rect 12357 3689 12391 3723
rect 12541 3689 12575 3723
rect 16037 3689 16071 3723
rect 16221 3689 16255 3723
rect 6561 3621 6595 3655
rect 6745 3621 6779 3655
rect 7941 3621 7975 3655
rect 10609 3621 10643 3655
rect 11161 3621 11195 3655
rect 8401 3553 8435 3587
rect 12265 3553 12299 3587
rect 6653 3485 6687 3519
rect 7389 3485 7423 3519
rect 8217 3485 8251 3519
rect 8309 3485 8343 3519
rect 9505 3485 9539 3519
rect 11437 3485 11471 3519
rect 12081 3485 12115 3519
rect 12357 3485 12391 3519
rect 14657 3485 14691 3519
rect 16129 3485 16163 3519
rect 6377 3417 6411 3451
rect 7113 3417 7147 3451
rect 7757 3417 7791 3451
rect 9137 3417 9171 3451
rect 10977 3417 11011 3451
rect 11253 3417 11287 3451
rect 14902 3417 14936 3451
rect 7297 3349 7331 3383
rect 8033 3349 8067 3383
rect 8953 3349 8987 3383
rect 7757 3145 7791 3179
rect 9873 3145 9907 3179
rect 11345 3145 11379 3179
rect 6377 3009 6411 3043
rect 6633 3009 6667 3043
rect 8125 3009 8159 3043
rect 8217 3009 8251 3043
rect 8493 3009 8527 3043
rect 8760 3009 8794 3043
rect 9965 3009 9999 3043
rect 10232 3009 10266 3043
rect 14298 3009 14332 3043
rect 14565 3009 14599 3043
rect 8033 2941 8067 2975
rect 15209 2941 15243 2975
rect 7849 2805 7883 2839
rect 13185 2805 13219 2839
rect 14657 2805 14691 2839
rect 6101 2601 6135 2635
rect 9137 2601 9171 2635
rect 10425 2601 10459 2635
rect 14105 2601 14139 2635
rect 5917 2397 5951 2431
rect 9321 2397 9355 2431
rect 10609 2397 10643 2431
rect 13921 2397 13955 2431
rect 14289 2397 14323 2431
rect 14565 2397 14599 2431
rect 14749 2397 14783 2431
rect 13737 2261 13771 2295
<< metal1 >>
rect 1104 17978 17388 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 17388 17978
rect 1104 17904 17388 17926
rect 12894 17824 12900 17876
rect 12952 17864 12958 17876
rect 13081 17867 13139 17873
rect 13081 17864 13093 17867
rect 12952 17836 13093 17864
rect 12952 17824 12958 17836
rect 13081 17833 13093 17836
rect 13127 17833 13139 17867
rect 13081 17827 13139 17833
rect 13538 17824 13544 17876
rect 13596 17864 13602 17876
rect 14185 17867 14243 17873
rect 14185 17864 14197 17867
rect 13596 17836 14197 17864
rect 13596 17824 13602 17836
rect 14185 17833 14197 17836
rect 14231 17833 14243 17867
rect 14185 17827 14243 17833
rect 13262 17552 13268 17604
rect 13320 17592 13326 17604
rect 13357 17595 13415 17601
rect 13357 17592 13369 17595
rect 13320 17564 13369 17592
rect 13320 17552 13326 17564
rect 13357 17561 13369 17564
rect 13403 17561 13415 17595
rect 13357 17555 13415 17561
rect 14461 17595 14519 17601
rect 14461 17561 14473 17595
rect 14507 17592 14519 17595
rect 14734 17592 14740 17604
rect 14507 17564 14740 17592
rect 14507 17561 14519 17564
rect 14461 17555 14519 17561
rect 14734 17552 14740 17564
rect 14792 17552 14798 17604
rect 1104 17434 17388 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 17388 17434
rect 1104 17360 17388 17382
rect 14734 17280 14740 17332
rect 14792 17320 14798 17332
rect 14792 17292 15332 17320
rect 14792 17280 14798 17292
rect 15194 17252 15200 17264
rect 11900 17224 15200 17252
rect 11900 17193 11928 17224
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17153 11943 17187
rect 11885 17147 11943 17153
rect 12152 17187 12210 17193
rect 12152 17153 12164 17187
rect 12198 17184 12210 17187
rect 12526 17184 12532 17196
rect 12198 17156 12532 17184
rect 12198 17153 12210 17156
rect 12152 17147 12210 17153
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 13372 17193 13400 17224
rect 15194 17212 15200 17224
rect 15252 17212 15258 17264
rect 13630 17193 13636 17196
rect 13357 17187 13415 17193
rect 13357 17153 13369 17187
rect 13403 17153 13415 17187
rect 13357 17147 13415 17153
rect 13624 17147 13636 17193
rect 13630 17144 13636 17147
rect 13688 17144 13694 17196
rect 15304 17184 15332 17292
rect 15381 17187 15439 17193
rect 15381 17184 15393 17187
rect 15304 17156 15393 17184
rect 15381 17153 15393 17156
rect 15427 17153 15439 17187
rect 15381 17147 15439 17153
rect 16485 17187 16543 17193
rect 16485 17153 16497 17187
rect 16531 17184 16543 17187
rect 16758 17184 16764 17196
rect 16531 17156 16764 17184
rect 16531 17153 16543 17156
rect 16485 17147 16543 17153
rect 16758 17144 16764 17156
rect 16816 17144 16822 17196
rect 13262 16940 13268 16992
rect 13320 16940 13326 16992
rect 13998 16940 14004 16992
rect 14056 16980 14062 16992
rect 14829 16983 14887 16989
rect 14829 16980 14841 16983
rect 14056 16952 14841 16980
rect 14056 16940 14062 16952
rect 14829 16949 14841 16952
rect 14875 16949 14887 16983
rect 14829 16943 14887 16949
rect 15286 16940 15292 16992
rect 15344 16980 15350 16992
rect 15841 16983 15899 16989
rect 15841 16980 15853 16983
rect 15344 16952 15853 16980
rect 15344 16940 15350 16952
rect 15841 16949 15853 16952
rect 15887 16949 15899 16983
rect 15841 16943 15899 16949
rect 16482 16940 16488 16992
rect 16540 16980 16546 16992
rect 16945 16983 17003 16989
rect 16945 16980 16957 16983
rect 16540 16952 16957 16980
rect 16540 16940 16546 16952
rect 16945 16949 16957 16952
rect 16991 16949 17003 16983
rect 16945 16943 17003 16949
rect 1104 16890 17388 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 17388 16890
rect 1104 16816 17388 16838
rect 12526 16736 12532 16788
rect 12584 16736 12590 16788
rect 16758 16736 16764 16788
rect 16816 16776 16822 16788
rect 17037 16779 17095 16785
rect 17037 16776 17049 16779
rect 16816 16748 17049 16776
rect 16816 16736 16822 16748
rect 17037 16745 17049 16748
rect 17083 16745 17095 16779
rect 17037 16739 17095 16745
rect 13262 16600 13268 16652
rect 13320 16640 13326 16652
rect 13725 16643 13783 16649
rect 13725 16640 13737 16643
rect 13320 16612 13737 16640
rect 13320 16600 13326 16612
rect 13725 16609 13737 16612
rect 13771 16609 13783 16643
rect 13725 16603 13783 16609
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 15252 16612 15669 16640
rect 15252 16600 15258 16612
rect 15657 16609 15669 16612
rect 15703 16609 15715 16643
rect 15657 16603 15715 16609
rect 12713 16575 12771 16581
rect 12713 16541 12725 16575
rect 12759 16572 12771 16575
rect 12759 16544 13032 16572
rect 12759 16541 12771 16544
rect 12713 16535 12771 16541
rect 12802 16464 12808 16516
rect 12860 16464 12866 16516
rect 12897 16507 12955 16513
rect 12897 16473 12909 16507
rect 12943 16473 12955 16507
rect 13004 16504 13032 16544
rect 13078 16532 13084 16584
rect 13136 16532 13142 16584
rect 14277 16575 14335 16581
rect 14277 16541 14289 16575
rect 14323 16572 14335 16575
rect 14366 16572 14372 16584
rect 14323 16544 14372 16572
rect 14323 16541 14335 16544
rect 14277 16535 14335 16541
rect 14366 16532 14372 16544
rect 14424 16532 14430 16584
rect 14645 16575 14703 16581
rect 14645 16541 14657 16575
rect 14691 16572 14703 16575
rect 15286 16572 15292 16584
rect 14691 16544 15292 16572
rect 14691 16541 14703 16544
rect 14645 16535 14703 16541
rect 15286 16532 15292 16544
rect 15344 16532 15350 16584
rect 15562 16532 15568 16584
rect 15620 16532 15626 16584
rect 13173 16507 13231 16513
rect 13173 16504 13185 16507
rect 13004 16476 13185 16504
rect 12897 16467 12955 16473
rect 13173 16473 13185 16476
rect 13219 16473 13231 16507
rect 13173 16467 13231 16473
rect 12912 16436 12940 16467
rect 14090 16464 14096 16516
rect 14148 16504 14154 16516
rect 14461 16507 14519 16513
rect 14461 16504 14473 16507
rect 14148 16476 14473 16504
rect 14148 16464 14154 16476
rect 14461 16473 14473 16476
rect 14507 16473 14519 16507
rect 14461 16467 14519 16473
rect 14553 16507 14611 16513
rect 14553 16473 14565 16507
rect 14599 16473 14611 16507
rect 15902 16507 15960 16513
rect 15902 16504 15914 16507
rect 14553 16467 14611 16473
rect 14844 16476 15914 16504
rect 13262 16436 13268 16448
rect 12912 16408 13268 16436
rect 13262 16396 13268 16408
rect 13320 16396 13326 16448
rect 14182 16396 14188 16448
rect 14240 16436 14246 16448
rect 14568 16436 14596 16467
rect 14844 16445 14872 16476
rect 15902 16473 15914 16476
rect 15948 16473 15960 16507
rect 15902 16467 15960 16473
rect 14240 16408 14596 16436
rect 14829 16439 14887 16445
rect 14240 16396 14246 16408
rect 14829 16405 14841 16439
rect 14875 16405 14887 16439
rect 14829 16399 14887 16405
rect 14918 16396 14924 16448
rect 14976 16396 14982 16448
rect 1104 16346 17388 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 17388 16346
rect 1104 16272 17388 16294
rect 10244 16204 12296 16232
rect 10244 16108 10272 16204
rect 10689 16167 10747 16173
rect 10689 16133 10701 16167
rect 10735 16164 10747 16167
rect 11974 16164 11980 16176
rect 10735 16136 11980 16164
rect 10735 16133 10747 16136
rect 10689 16127 10747 16133
rect 11974 16124 11980 16136
rect 12032 16124 12038 16176
rect 8294 16056 8300 16108
rect 8352 16096 8358 16108
rect 9953 16099 10011 16105
rect 9953 16096 9965 16099
rect 8352 16068 9965 16096
rect 8352 16056 8358 16068
rect 9953 16065 9965 16068
rect 9999 16065 10011 16099
rect 9953 16059 10011 16065
rect 10226 16056 10232 16108
rect 10284 16056 10290 16108
rect 10873 16099 10931 16105
rect 10873 16065 10885 16099
rect 10919 16065 10931 16099
rect 10873 16059 10931 16065
rect 10042 15988 10048 16040
rect 10100 15988 10106 16040
rect 10505 15963 10563 15969
rect 10505 15960 10517 15963
rect 10244 15932 10517 15960
rect 10244 15901 10272 15932
rect 10505 15929 10517 15932
rect 10551 15929 10563 15963
rect 10888 15960 10916 16059
rect 10962 16056 10968 16108
rect 11020 16096 11026 16108
rect 12268 16105 12296 16204
rect 13630 16192 13636 16244
rect 13688 16192 13694 16244
rect 14918 16232 14924 16244
rect 14292 16204 14924 16232
rect 13998 16164 14004 16176
rect 13464 16136 14004 16164
rect 12069 16099 12127 16105
rect 12069 16096 12081 16099
rect 11020 16068 12081 16096
rect 11020 16056 11026 16068
rect 12069 16065 12081 16068
rect 12115 16065 12127 16099
rect 12069 16059 12127 16065
rect 12253 16099 12311 16105
rect 12253 16065 12265 16099
rect 12299 16065 12311 16099
rect 12253 16059 12311 16065
rect 12345 16099 12403 16105
rect 12345 16065 12357 16099
rect 12391 16096 12403 16099
rect 12434 16096 12440 16108
rect 12391 16068 12440 16096
rect 12391 16065 12403 16068
rect 12345 16059 12403 16065
rect 12434 16056 12440 16068
rect 12492 16056 12498 16108
rect 13081 16099 13139 16105
rect 13081 16096 13093 16099
rect 12544 16068 13093 16096
rect 11054 15960 11060 15972
rect 10888 15932 11060 15960
rect 10505 15923 10563 15929
rect 11054 15920 11060 15932
rect 11112 15960 11118 15972
rect 11882 15960 11888 15972
rect 11112 15932 11888 15960
rect 11112 15920 11118 15932
rect 11882 15920 11888 15932
rect 11940 15920 11946 15972
rect 12544 15969 12572 16068
rect 13081 16065 13093 16068
rect 13127 16065 13139 16099
rect 13081 16059 13139 16065
rect 13262 16056 13268 16108
rect 13320 16056 13326 16108
rect 13464 16105 13492 16136
rect 13998 16124 14004 16136
rect 14056 16124 14062 16176
rect 13357 16099 13415 16105
rect 13357 16065 13369 16099
rect 13403 16065 13415 16099
rect 13357 16059 13415 16065
rect 13449 16099 13507 16105
rect 13449 16065 13461 16099
rect 13495 16065 13507 16099
rect 13449 16059 13507 16065
rect 13909 16099 13967 16105
rect 13909 16065 13921 16099
rect 13955 16065 13967 16099
rect 13909 16059 13967 16065
rect 12529 15963 12587 15969
rect 12529 15929 12541 15963
rect 12575 15929 12587 15963
rect 13372 15960 13400 16059
rect 13924 16028 13952 16059
rect 14090 16056 14096 16108
rect 14148 16056 14154 16108
rect 14182 16056 14188 16108
rect 14240 16056 14246 16108
rect 14292 16105 14320 16204
rect 14918 16192 14924 16204
rect 14976 16192 14982 16244
rect 15562 16192 15568 16244
rect 15620 16232 15626 16244
rect 15933 16235 15991 16241
rect 15933 16232 15945 16235
rect 15620 16204 15945 16232
rect 15620 16192 15626 16204
rect 15933 16201 15945 16204
rect 15979 16201 15991 16235
rect 15933 16195 15991 16201
rect 15194 16164 15200 16176
rect 14568 16136 15200 16164
rect 14568 16105 14596 16136
rect 15194 16124 15200 16136
rect 15252 16124 15258 16176
rect 14277 16099 14335 16105
rect 14277 16065 14289 16099
rect 14323 16065 14335 16099
rect 14277 16059 14335 16065
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16065 14611 16099
rect 14809 16099 14867 16105
rect 14809 16096 14821 16099
rect 14553 16059 14611 16065
rect 14660 16068 14821 16096
rect 13998 16028 14004 16040
rect 13924 16000 14004 16028
rect 13998 15988 14004 16000
rect 14056 15988 14062 16040
rect 14108 16028 14136 16056
rect 14660 16028 14688 16068
rect 14809 16065 14821 16068
rect 14855 16065 14867 16099
rect 15948 16096 15976 16195
rect 16761 16099 16819 16105
rect 16761 16096 16773 16099
rect 15948 16068 16773 16096
rect 14809 16059 14867 16065
rect 16761 16065 16773 16068
rect 16807 16065 16819 16099
rect 16761 16059 16819 16065
rect 14108 16000 14228 16028
rect 14090 15960 14096 15972
rect 13372 15932 14096 15960
rect 12529 15923 12587 15929
rect 14090 15920 14096 15932
rect 14148 15920 14154 15972
rect 10229 15895 10287 15901
rect 10229 15861 10241 15895
rect 10275 15861 10287 15895
rect 10229 15855 10287 15861
rect 10413 15895 10471 15901
rect 10413 15861 10425 15895
rect 10459 15892 10471 15895
rect 11606 15892 11612 15904
rect 10459 15864 11612 15892
rect 10459 15861 10471 15864
rect 10413 15855 10471 15861
rect 11606 15852 11612 15864
rect 11664 15852 11670 15904
rect 12250 15852 12256 15904
rect 12308 15852 12314 15904
rect 14200 15892 14228 16000
rect 14476 16000 14688 16028
rect 14476 15969 14504 16000
rect 14461 15963 14519 15969
rect 14461 15929 14473 15963
rect 14507 15929 14519 15963
rect 14461 15923 14519 15929
rect 15470 15892 15476 15904
rect 14200 15864 15476 15892
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 16942 15852 16948 15904
rect 17000 15852 17006 15904
rect 1104 15802 17388 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 17388 15802
rect 1104 15728 17388 15750
rect 5905 15691 5963 15697
rect 5905 15657 5917 15691
rect 5951 15688 5963 15691
rect 6178 15688 6184 15700
rect 5951 15660 6184 15688
rect 5951 15657 5963 15660
rect 5905 15651 5963 15657
rect 6178 15648 6184 15660
rect 6236 15648 6242 15700
rect 7650 15648 7656 15700
rect 7708 15688 7714 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7708 15660 7849 15688
rect 7708 15648 7714 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 7837 15651 7895 15657
rect 8294 15648 8300 15700
rect 8352 15648 8358 15700
rect 9122 15648 9128 15700
rect 9180 15648 9186 15700
rect 9493 15691 9551 15697
rect 9493 15657 9505 15691
rect 9539 15688 9551 15691
rect 10226 15688 10232 15700
rect 9539 15660 10232 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 10226 15648 10232 15660
rect 10284 15648 10290 15700
rect 10413 15691 10471 15697
rect 10413 15657 10425 15691
rect 10459 15657 10471 15691
rect 10413 15651 10471 15657
rect 10597 15691 10655 15697
rect 10597 15657 10609 15691
rect 10643 15688 10655 15691
rect 10962 15688 10968 15700
rect 10643 15660 10968 15688
rect 10643 15657 10655 15660
rect 10597 15651 10655 15657
rect 7098 15620 7104 15632
rect 5644 15592 7104 15620
rect 5644 15493 5672 15592
rect 7098 15580 7104 15592
rect 7156 15620 7162 15632
rect 10428 15620 10456 15651
rect 10962 15648 10968 15660
rect 11020 15648 11026 15700
rect 11146 15648 11152 15700
rect 11204 15688 11210 15700
rect 11333 15691 11391 15697
rect 11333 15688 11345 15691
rect 11204 15660 11345 15688
rect 11204 15648 11210 15660
rect 11333 15657 11345 15660
rect 11379 15657 11391 15691
rect 11333 15651 11391 15657
rect 12250 15648 12256 15700
rect 12308 15648 12314 15700
rect 12621 15691 12679 15697
rect 12621 15657 12633 15691
rect 12667 15688 12679 15691
rect 12710 15688 12716 15700
rect 12667 15660 12716 15688
rect 12667 15657 12679 15660
rect 12621 15651 12679 15657
rect 12710 15648 12716 15660
rect 12768 15648 12774 15700
rect 14182 15648 14188 15700
rect 14240 15688 14246 15700
rect 15286 15688 15292 15700
rect 14240 15660 15292 15688
rect 14240 15648 14246 15660
rect 15286 15648 15292 15660
rect 15344 15648 15350 15700
rect 11054 15620 11060 15632
rect 7156 15592 10364 15620
rect 10428 15592 11060 15620
rect 7156 15580 7162 15592
rect 7926 15512 7932 15564
rect 7984 15512 7990 15564
rect 8036 15524 10180 15552
rect 5629 15487 5687 15493
rect 5629 15453 5641 15487
rect 5675 15453 5687 15487
rect 5629 15447 5687 15453
rect 5813 15487 5871 15493
rect 5813 15453 5825 15487
rect 5859 15453 5871 15487
rect 5813 15447 5871 15453
rect 5534 15376 5540 15428
rect 5592 15416 5598 15428
rect 5828 15416 5856 15447
rect 5902 15444 5908 15496
rect 5960 15444 5966 15496
rect 8036 15484 8064 15524
rect 6104 15456 8064 15484
rect 8113 15487 8171 15493
rect 6104 15416 6132 15456
rect 8113 15453 8125 15487
rect 8159 15484 8171 15487
rect 8294 15484 8300 15496
rect 8159 15456 8300 15484
rect 8159 15453 8171 15456
rect 8113 15447 8171 15453
rect 8294 15444 8300 15456
rect 8352 15444 8358 15496
rect 9122 15444 9128 15496
rect 9180 15444 9186 15496
rect 9309 15487 9367 15493
rect 9309 15453 9321 15487
rect 9355 15484 9367 15487
rect 9582 15484 9588 15496
rect 9355 15456 9588 15484
rect 9355 15453 9367 15456
rect 9309 15447 9367 15453
rect 9582 15444 9588 15456
rect 9640 15444 9646 15496
rect 10152 15484 10180 15524
rect 10226 15512 10232 15564
rect 10284 15512 10290 15564
rect 10336 15552 10364 15592
rect 11054 15580 11060 15592
rect 11112 15580 11118 15632
rect 11701 15623 11759 15629
rect 11701 15589 11713 15623
rect 11747 15620 11759 15623
rect 11747 15592 12434 15620
rect 11747 15589 11759 15592
rect 11701 15583 11759 15589
rect 12406 15552 12434 15592
rect 13262 15580 13268 15632
rect 13320 15620 13326 15632
rect 15102 15620 15108 15632
rect 13320 15592 15108 15620
rect 13320 15580 13326 15592
rect 15102 15580 15108 15592
rect 15160 15580 15166 15632
rect 10336 15524 11376 15552
rect 12406 15524 12664 15552
rect 10152 15456 10364 15484
rect 5592 15388 6132 15416
rect 5592 15376 5598 15388
rect 6822 15376 6828 15428
rect 6880 15416 6886 15428
rect 7837 15419 7895 15425
rect 7837 15416 7849 15419
rect 6880 15388 7849 15416
rect 6880 15376 6886 15388
rect 7837 15385 7849 15388
rect 7883 15385 7895 15419
rect 7837 15379 7895 15385
rect 10134 15376 10140 15428
rect 10192 15376 10198 15428
rect 10336 15416 10364 15456
rect 10410 15444 10416 15496
rect 10468 15444 10474 15496
rect 11348 15493 11376 15524
rect 11333 15487 11391 15493
rect 11333 15453 11345 15487
rect 11379 15453 11391 15487
rect 11333 15447 11391 15453
rect 11517 15487 11575 15493
rect 11517 15453 11529 15487
rect 11563 15484 11575 15487
rect 11698 15484 11704 15496
rect 11563 15456 11704 15484
rect 11563 15453 11575 15456
rect 11517 15447 11575 15453
rect 11054 15416 11060 15428
rect 10336 15388 11060 15416
rect 11054 15376 11060 15388
rect 11112 15376 11118 15428
rect 11348 15416 11376 15447
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 12636 15493 12664 15524
rect 15194 15512 15200 15564
rect 15252 15552 15258 15564
rect 15657 15555 15715 15561
rect 15657 15552 15669 15555
rect 15252 15524 15669 15552
rect 15252 15512 15258 15524
rect 15657 15521 15669 15524
rect 15703 15521 15715 15555
rect 15657 15515 15715 15521
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 12621 15487 12679 15493
rect 12621 15453 12633 15487
rect 12667 15453 12679 15487
rect 12621 15447 12679 15453
rect 11793 15419 11851 15425
rect 11793 15416 11805 15419
rect 11348 15388 11805 15416
rect 11793 15385 11805 15388
rect 11839 15385 11851 15419
rect 11793 15379 11851 15385
rect 11977 15419 12035 15425
rect 11977 15385 11989 15419
rect 12023 15385 12035 15419
rect 12544 15416 12572 15447
rect 14090 15416 14096 15428
rect 12544 15388 14096 15416
rect 11977 15379 12035 15385
rect 6089 15351 6147 15357
rect 6089 15317 6101 15351
rect 6135 15348 6147 15351
rect 9674 15348 9680 15360
rect 6135 15320 9680 15348
rect 6135 15317 6147 15320
rect 6089 15311 6147 15317
rect 9674 15308 9680 15320
rect 9732 15308 9738 15360
rect 11072 15348 11100 15376
rect 11992 15348 12020 15379
rect 14090 15376 14096 15388
rect 14148 15376 14154 15428
rect 15746 15376 15752 15428
rect 15804 15416 15810 15428
rect 15902 15419 15960 15425
rect 15902 15416 15914 15419
rect 15804 15388 15914 15416
rect 15804 15376 15810 15388
rect 15902 15385 15914 15388
rect 15948 15385 15960 15419
rect 15902 15379 15960 15385
rect 11072 15320 12020 15348
rect 12066 15308 12072 15360
rect 12124 15348 12130 15360
rect 12161 15351 12219 15357
rect 12161 15348 12173 15351
rect 12124 15320 12173 15348
rect 12124 15308 12130 15320
rect 12161 15317 12173 15320
rect 12207 15317 12219 15351
rect 12161 15311 12219 15317
rect 12802 15308 12808 15360
rect 12860 15348 12866 15360
rect 15654 15348 15660 15360
rect 12860 15320 15660 15348
rect 12860 15308 12866 15320
rect 15654 15308 15660 15320
rect 15712 15308 15718 15360
rect 17034 15308 17040 15360
rect 17092 15308 17098 15360
rect 1104 15258 17388 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 17388 15258
rect 1104 15184 17388 15206
rect 7558 15104 7564 15156
rect 7616 15144 7622 15156
rect 9122 15144 9128 15156
rect 7616 15116 9128 15144
rect 7616 15104 7622 15116
rect 9122 15104 9128 15116
rect 9180 15144 9186 15156
rect 9180 15116 9904 15144
rect 9180 15104 9186 15116
rect 6730 15076 6736 15088
rect 6472 15048 6736 15076
rect 5629 15011 5687 15017
rect 5629 14977 5641 15011
rect 5675 14977 5687 15011
rect 5629 14971 5687 14977
rect 5813 15011 5871 15017
rect 5813 14977 5825 15011
rect 5859 15008 5871 15011
rect 6472 15008 6500 15048
rect 6730 15036 6736 15048
rect 6788 15036 6794 15088
rect 7282 15076 7288 15088
rect 7116 15048 7288 15076
rect 5859 14980 6500 15008
rect 6549 15011 6607 15017
rect 5859 14977 5871 14980
rect 5813 14971 5871 14977
rect 6549 14977 6561 15011
rect 6595 15008 6607 15011
rect 6595 14980 6776 15008
rect 6595 14977 6607 14980
rect 6549 14971 6607 14977
rect 5644 14872 5672 14971
rect 5718 14900 5724 14952
rect 5776 14940 5782 14952
rect 6564 14940 6592 14971
rect 5776 14912 6592 14940
rect 5776 14900 5782 14912
rect 6638 14900 6644 14952
rect 6696 14900 6702 14952
rect 6748 14940 6776 14980
rect 6822 14968 6828 15020
rect 6880 14968 6886 15020
rect 7116 14940 7144 15048
rect 7282 15036 7288 15048
rect 7340 15036 7346 15088
rect 7193 15011 7251 15017
rect 7193 14977 7205 15011
rect 7239 15008 7251 15011
rect 7469 15011 7527 15017
rect 7239 14980 7420 15008
rect 7239 14977 7251 14980
rect 7193 14971 7251 14977
rect 6748 14912 7144 14940
rect 7282 14900 7288 14952
rect 7340 14900 7346 14952
rect 5902 14872 5908 14884
rect 5644 14844 5908 14872
rect 5902 14832 5908 14844
rect 5960 14872 5966 14884
rect 6656 14872 6684 14900
rect 7392 14872 7420 14980
rect 7469 14977 7481 15011
rect 7515 15008 7527 15011
rect 7558 15008 7564 15020
rect 7515 14980 7564 15008
rect 7515 14977 7527 14980
rect 7469 14971 7527 14977
rect 7558 14968 7564 14980
rect 7616 15008 7622 15020
rect 7616 14980 7793 15008
rect 7616 14968 7622 14980
rect 7765 14940 7793 14980
rect 7834 14968 7840 15020
rect 7892 14968 7898 15020
rect 8021 15011 8079 15017
rect 8021 14977 8033 15011
rect 8067 14977 8079 15011
rect 8021 14971 8079 14977
rect 8036 14940 8064 14971
rect 9122 14968 9128 15020
rect 9180 15008 9186 15020
rect 9309 15011 9367 15017
rect 9309 15008 9321 15011
rect 9180 14980 9321 15008
rect 9180 14968 9186 14980
rect 9309 14977 9321 14980
rect 9355 14977 9367 15011
rect 9309 14971 9367 14977
rect 9582 14968 9588 15020
rect 9640 14968 9646 15020
rect 9876 15008 9904 15116
rect 10410 15104 10416 15156
rect 10468 15144 10474 15156
rect 12345 15147 12403 15153
rect 10468 15116 12204 15144
rect 10468 15104 10474 15116
rect 11422 15036 11428 15088
rect 11480 15076 11486 15088
rect 11885 15079 11943 15085
rect 11885 15076 11897 15079
rect 11480 15048 11897 15076
rect 11480 15036 11486 15048
rect 11885 15045 11897 15048
rect 11931 15045 11943 15079
rect 11885 15039 11943 15045
rect 10965 15011 11023 15017
rect 10965 15008 10977 15011
rect 9876 14980 10977 15008
rect 10965 14977 10977 14980
rect 11011 14977 11023 15011
rect 10965 14971 11023 14977
rect 11146 14968 11152 15020
rect 11204 14968 11210 15020
rect 12066 14968 12072 15020
rect 12124 14968 12130 15020
rect 12176 15017 12204 15116
rect 12345 15113 12357 15147
rect 12391 15144 12403 15147
rect 13633 15147 13691 15153
rect 12391 15116 13216 15144
rect 12391 15113 12403 15116
rect 12345 15107 12403 15113
rect 13188 15085 13216 15116
rect 13633 15113 13645 15147
rect 13679 15113 13691 15147
rect 13633 15107 13691 15113
rect 14553 15147 14611 15153
rect 14553 15113 14565 15147
rect 14599 15113 14611 15147
rect 14553 15107 14611 15113
rect 13173 15079 13231 15085
rect 13173 15045 13185 15079
rect 13219 15045 13231 15079
rect 13648 15076 13676 15107
rect 13648 15048 14228 15076
rect 13173 15039 13231 15045
rect 12161 15011 12219 15017
rect 12161 14977 12173 15011
rect 12207 14977 12219 15011
rect 12161 14971 12219 14977
rect 13449 15011 13507 15017
rect 13449 14977 13461 15011
rect 13495 15008 13507 15011
rect 13538 15008 13544 15020
rect 13495 14980 13544 15008
rect 13495 14977 13507 14980
rect 13449 14971 13507 14977
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 13909 15011 13967 15017
rect 13909 14977 13921 15011
rect 13955 14977 13967 15011
rect 13909 14971 13967 14977
rect 7765 14912 8064 14940
rect 7466 14872 7472 14884
rect 5960 14844 6684 14872
rect 6932 14844 7472 14872
rect 5960 14832 5966 14844
rect 5994 14764 6000 14816
rect 6052 14764 6058 14816
rect 6362 14764 6368 14816
rect 6420 14764 6426 14816
rect 6546 14764 6552 14816
rect 6604 14804 6610 14816
rect 6932 14804 6960 14844
rect 7466 14832 7472 14844
rect 7524 14832 7530 14884
rect 7834 14872 7840 14884
rect 7576 14844 7840 14872
rect 6604 14776 6960 14804
rect 6604 14764 6610 14776
rect 7006 14764 7012 14816
rect 7064 14804 7070 14816
rect 7193 14807 7251 14813
rect 7193 14804 7205 14807
rect 7064 14776 7205 14804
rect 7064 14764 7070 14776
rect 7193 14773 7205 14776
rect 7239 14804 7251 14807
rect 7576 14804 7604 14844
rect 7834 14832 7840 14844
rect 7892 14832 7898 14884
rect 8036 14872 8064 14912
rect 8294 14900 8300 14952
rect 8352 14940 8358 14952
rect 9493 14943 9551 14949
rect 9493 14940 9505 14943
rect 8352 14912 9505 14940
rect 8352 14900 8358 14912
rect 9493 14909 9505 14912
rect 9539 14940 9551 14943
rect 9950 14940 9956 14952
rect 9539 14912 9956 14940
rect 9539 14909 9551 14912
rect 9493 14903 9551 14909
rect 9950 14900 9956 14912
rect 10008 14900 10014 14952
rect 12894 14900 12900 14952
rect 12952 14940 12958 14952
rect 13265 14943 13323 14949
rect 13265 14940 13277 14943
rect 12952 14912 13277 14940
rect 12952 14900 12958 14912
rect 13265 14909 13277 14912
rect 13311 14909 13323 14943
rect 13265 14903 13323 14909
rect 13354 14900 13360 14952
rect 13412 14940 13418 14952
rect 13924 14940 13952 14971
rect 14090 14968 14096 15020
rect 14148 14968 14154 15020
rect 14200 15017 14228 15048
rect 14185 15011 14243 15017
rect 14185 14977 14197 15011
rect 14231 14977 14243 15011
rect 14568 15008 14596 15107
rect 15746 15104 15752 15156
rect 15804 15104 15810 15156
rect 16942 15104 16948 15156
rect 17000 15104 17006 15156
rect 15378 15036 15384 15088
rect 15436 15036 15442 15088
rect 15197 15011 15255 15017
rect 15197 15008 15209 15011
rect 14568 14980 15209 15008
rect 14185 14971 14243 14977
rect 15197 14977 15209 14980
rect 15243 14977 15255 15011
rect 15197 14971 15255 14977
rect 15286 14968 15292 15020
rect 15344 15008 15350 15020
rect 15473 15011 15531 15017
rect 15473 15008 15485 15011
rect 15344 14980 15485 15008
rect 15344 14968 15350 14980
rect 15473 14977 15485 14980
rect 15519 14977 15531 15011
rect 15473 14971 15531 14977
rect 15565 15011 15623 15017
rect 15565 14977 15577 15011
rect 15611 15008 15623 15011
rect 15841 15011 15899 15017
rect 15841 15008 15853 15011
rect 15611 14980 15853 15008
rect 15611 14977 15623 14980
rect 15565 14971 15623 14977
rect 15841 14977 15853 14980
rect 15887 14977 15899 15011
rect 15841 14971 15899 14977
rect 16485 15011 16543 15017
rect 16485 14977 16497 15011
rect 16531 15008 16543 15011
rect 16761 15011 16819 15017
rect 16761 15008 16773 15011
rect 16531 14980 16773 15008
rect 16531 14977 16543 14980
rect 16485 14971 16543 14977
rect 16761 14977 16773 14980
rect 16807 15008 16819 15011
rect 17034 15008 17040 15020
rect 16807 14980 17040 15008
rect 16807 14977 16819 14980
rect 16761 14971 16819 14977
rect 17034 14968 17040 14980
rect 17092 14968 17098 15020
rect 13412 14912 13952 14940
rect 13412 14900 13418 14912
rect 14274 14900 14280 14952
rect 14332 14900 14338 14952
rect 9769 14875 9827 14881
rect 8036 14844 9674 14872
rect 7239 14776 7604 14804
rect 7653 14807 7711 14813
rect 7239 14773 7251 14776
rect 7193 14767 7251 14773
rect 7653 14773 7665 14807
rect 7699 14804 7711 14807
rect 8110 14804 8116 14816
rect 7699 14776 8116 14804
rect 7699 14773 7711 14776
rect 7653 14767 7711 14773
rect 8110 14764 8116 14776
rect 8168 14764 8174 14816
rect 8202 14764 8208 14816
rect 8260 14764 8266 14816
rect 8938 14764 8944 14816
rect 8996 14804 9002 14816
rect 9309 14807 9367 14813
rect 9309 14804 9321 14807
rect 8996 14776 9321 14804
rect 8996 14764 9002 14776
rect 9309 14773 9321 14776
rect 9355 14773 9367 14807
rect 9646 14804 9674 14844
rect 9769 14841 9781 14875
rect 9815 14872 9827 14875
rect 9815 14844 14228 14872
rect 9815 14841 9827 14844
rect 9769 14835 9827 14841
rect 11146 14804 11152 14816
rect 9646 14776 11152 14804
rect 9309 14767 9367 14773
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 11330 14764 11336 14816
rect 11388 14764 11394 14816
rect 11974 14764 11980 14816
rect 12032 14764 12038 14816
rect 13170 14764 13176 14816
rect 13228 14764 13234 14816
rect 13354 14764 13360 14816
rect 13412 14804 13418 14816
rect 14200 14813 14228 14844
rect 13725 14807 13783 14813
rect 13725 14804 13737 14807
rect 13412 14776 13737 14804
rect 13412 14764 13418 14776
rect 13725 14773 13737 14776
rect 13771 14773 13783 14807
rect 13725 14767 13783 14773
rect 14185 14807 14243 14813
rect 14185 14773 14197 14807
rect 14231 14773 14243 14807
rect 14185 14767 14243 14773
rect 1104 14714 17388 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 17388 14714
rect 1104 14640 17388 14662
rect 6178 14560 6184 14612
rect 6236 14600 6242 14612
rect 6822 14600 6828 14612
rect 6236 14572 6828 14600
rect 6236 14560 6242 14572
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 8478 14560 8484 14612
rect 8536 14560 8542 14612
rect 8754 14560 8760 14612
rect 8812 14600 8818 14612
rect 9582 14600 9588 14612
rect 8812 14572 9588 14600
rect 8812 14560 8818 14572
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 11422 14600 11428 14612
rect 9784 14572 11428 14600
rect 5994 14492 6000 14544
rect 6052 14532 6058 14544
rect 9784 14532 9812 14572
rect 11422 14560 11428 14572
rect 11480 14560 11486 14612
rect 11793 14603 11851 14609
rect 11793 14569 11805 14603
rect 11839 14600 11851 14603
rect 12253 14603 12311 14609
rect 12253 14600 12265 14603
rect 11839 14572 12265 14600
rect 11839 14569 11851 14572
rect 11793 14563 11851 14569
rect 12253 14569 12265 14572
rect 12299 14569 12311 14603
rect 13449 14603 13507 14609
rect 13449 14600 13461 14603
rect 12253 14563 12311 14569
rect 12406 14572 13461 14600
rect 6052 14504 9812 14532
rect 6052 14492 6058 14504
rect 11238 14492 11244 14544
rect 11296 14532 11302 14544
rect 11296 14504 11652 14532
rect 11296 14492 11302 14504
rect 8389 14467 8447 14473
rect 8389 14433 8401 14467
rect 8435 14464 8447 14467
rect 9398 14464 9404 14476
rect 8435 14436 9404 14464
rect 8435 14433 8447 14436
rect 8389 14427 8447 14433
rect 9398 14424 9404 14436
rect 9456 14424 9462 14476
rect 11330 14424 11336 14476
rect 11388 14464 11394 14476
rect 11517 14467 11575 14473
rect 11517 14464 11529 14467
rect 11388 14436 11529 14464
rect 11388 14424 11394 14436
rect 11517 14433 11529 14436
rect 11563 14433 11575 14467
rect 11517 14427 11575 14433
rect 3418 14356 3424 14408
rect 3476 14396 3482 14408
rect 7190 14396 7196 14408
rect 3476 14368 7196 14396
rect 3476 14356 3482 14368
rect 7190 14356 7196 14368
rect 7248 14356 7254 14408
rect 8202 14356 8208 14408
rect 8260 14356 8266 14408
rect 8294 14356 8300 14408
rect 8352 14396 8358 14408
rect 8481 14399 8539 14405
rect 8481 14396 8493 14399
rect 8352 14368 8493 14396
rect 8352 14356 8358 14368
rect 8481 14365 8493 14368
rect 8527 14365 8539 14399
rect 9125 14399 9183 14405
rect 9125 14396 9137 14399
rect 8481 14359 8539 14365
rect 8588 14368 9137 14396
rect 6638 14288 6644 14340
rect 6696 14328 6702 14340
rect 8386 14328 8392 14340
rect 6696 14300 8392 14328
rect 6696 14288 6702 14300
rect 8386 14288 8392 14300
rect 8444 14328 8450 14340
rect 8588 14328 8616 14368
rect 9125 14365 9137 14368
rect 9171 14365 9183 14399
rect 9125 14359 9183 14365
rect 9214 14356 9220 14408
rect 9272 14396 9278 14408
rect 9309 14399 9367 14405
rect 9309 14396 9321 14399
rect 9272 14368 9321 14396
rect 9272 14356 9278 14368
rect 9309 14365 9321 14368
rect 9355 14396 9367 14399
rect 11425 14399 11483 14405
rect 11425 14396 11437 14399
rect 9355 14368 11437 14396
rect 9355 14365 9367 14368
rect 9309 14359 9367 14365
rect 11425 14365 11437 14368
rect 11471 14365 11483 14399
rect 11624 14396 11652 14504
rect 12066 14492 12072 14544
rect 12124 14532 12130 14544
rect 12406 14532 12434 14572
rect 13449 14569 13461 14572
rect 13495 14569 13507 14603
rect 13449 14563 13507 14569
rect 12124 14504 12434 14532
rect 12621 14535 12679 14541
rect 12124 14492 12130 14504
rect 12621 14501 12633 14535
rect 12667 14532 12679 14535
rect 13078 14532 13084 14544
rect 12667 14504 13084 14532
rect 12667 14501 12679 14504
rect 12621 14495 12679 14501
rect 13078 14492 13084 14504
rect 13136 14492 13142 14544
rect 11790 14424 11796 14476
rect 11848 14464 11854 14476
rect 13541 14467 13599 14473
rect 13541 14464 13553 14467
rect 11848 14436 13553 14464
rect 11848 14424 11854 14436
rect 13541 14433 13553 14436
rect 13587 14433 13599 14467
rect 13541 14427 13599 14433
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 15289 14467 15347 14473
rect 15289 14464 15301 14467
rect 15252 14436 15301 14464
rect 15252 14424 15258 14436
rect 15289 14433 15301 14436
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 11624 14368 12265 14396
rect 11425 14359 11483 14365
rect 12253 14365 12265 14368
rect 12299 14365 12311 14399
rect 12253 14359 12311 14365
rect 12437 14399 12495 14405
rect 12437 14365 12449 14399
rect 12483 14396 12495 14399
rect 12986 14396 12992 14408
rect 12483 14368 12992 14396
rect 12483 14365 12495 14368
rect 12437 14359 12495 14365
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 13354 14356 13360 14408
rect 13412 14396 13418 14408
rect 13449 14399 13507 14405
rect 13449 14396 13461 14399
rect 13412 14368 13461 14396
rect 13412 14356 13418 14368
rect 13449 14365 13461 14368
rect 13495 14365 13507 14399
rect 13449 14359 13507 14365
rect 8444 14300 8616 14328
rect 8444 14288 8450 14300
rect 8938 14288 8944 14340
rect 8996 14288 9002 14340
rect 12894 14328 12900 14340
rect 9232 14300 12900 14328
rect 4614 14220 4620 14272
rect 4672 14260 4678 14272
rect 8294 14260 8300 14272
rect 4672 14232 8300 14260
rect 4672 14220 4678 14232
rect 8294 14220 8300 14232
rect 8352 14220 8358 14272
rect 8665 14263 8723 14269
rect 8665 14229 8677 14263
rect 8711 14260 8723 14263
rect 9232 14260 9260 14300
rect 12894 14288 12900 14300
rect 12952 14328 12958 14340
rect 14182 14328 14188 14340
rect 12952 14300 14188 14328
rect 12952 14288 12958 14300
rect 14182 14288 14188 14300
rect 14240 14288 14246 14340
rect 15556 14331 15614 14337
rect 15556 14297 15568 14331
rect 15602 14328 15614 14331
rect 15654 14328 15660 14340
rect 15602 14300 15660 14328
rect 15602 14297 15614 14300
rect 15556 14291 15614 14297
rect 15654 14288 15660 14300
rect 15712 14288 15718 14340
rect 8711 14232 9260 14260
rect 8711 14229 8723 14232
rect 8665 14223 8723 14229
rect 11054 14220 11060 14272
rect 11112 14260 11118 14272
rect 12066 14260 12072 14272
rect 11112 14232 12072 14260
rect 11112 14220 11118 14232
rect 12066 14220 12072 14232
rect 12124 14220 12130 14272
rect 13814 14220 13820 14272
rect 13872 14220 13878 14272
rect 16669 14263 16727 14269
rect 16669 14229 16681 14263
rect 16715 14260 16727 14263
rect 16758 14260 16764 14272
rect 16715 14232 16764 14260
rect 16715 14229 16727 14232
rect 16669 14223 16727 14229
rect 16758 14220 16764 14232
rect 16816 14220 16822 14272
rect 1104 14170 17388 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 17388 14170
rect 1104 14096 17388 14118
rect 3605 14059 3663 14065
rect 3605 14025 3617 14059
rect 3651 14056 3663 14059
rect 7006 14056 7012 14068
rect 3651 14028 7012 14056
rect 3651 14025 3663 14028
rect 3605 14019 3663 14025
rect 7006 14016 7012 14028
rect 7064 14056 7070 14068
rect 7064 14028 7512 14056
rect 7064 14016 7070 14028
rect 3237 13991 3295 13997
rect 3237 13957 3249 13991
rect 3283 13988 3295 13991
rect 3694 13988 3700 14000
rect 3283 13960 3700 13988
rect 3283 13957 3295 13960
rect 3237 13951 3295 13957
rect 3694 13948 3700 13960
rect 3752 13988 3758 14000
rect 7101 13991 7159 13997
rect 3752 13960 7052 13988
rect 3752 13948 3758 13960
rect 3053 13923 3111 13929
rect 3053 13889 3065 13923
rect 3099 13920 3111 13923
rect 3142 13920 3148 13932
rect 3099 13892 3148 13920
rect 3099 13889 3111 13892
rect 3053 13883 3111 13889
rect 3142 13880 3148 13892
rect 3200 13880 3206 13932
rect 3326 13880 3332 13932
rect 3384 13880 3390 13932
rect 3418 13880 3424 13932
rect 3476 13920 3482 13932
rect 3878 13920 3884 13932
rect 3476 13892 3884 13920
rect 3476 13880 3482 13892
rect 3878 13880 3884 13892
rect 3936 13880 3942 13932
rect 4154 13880 4160 13932
rect 4212 13920 4218 13932
rect 4341 13923 4399 13929
rect 4341 13920 4353 13923
rect 4212 13892 4353 13920
rect 4212 13880 4218 13892
rect 4341 13889 4353 13892
rect 4387 13889 4399 13923
rect 4341 13883 4399 13889
rect 4525 13923 4583 13929
rect 4525 13889 4537 13923
rect 4571 13920 4583 13923
rect 5902 13920 5908 13932
rect 4571 13892 5908 13920
rect 4571 13889 4583 13892
rect 4525 13883 4583 13889
rect 5902 13880 5908 13892
rect 5960 13880 5966 13932
rect 6822 13880 6828 13932
rect 6880 13880 6886 13932
rect 7024 13929 7052 13960
rect 7101 13957 7113 13991
rect 7147 13988 7159 13991
rect 7282 13988 7288 14000
rect 7147 13960 7288 13988
rect 7147 13957 7159 13960
rect 7101 13951 7159 13957
rect 7282 13948 7288 13960
rect 7340 13948 7346 14000
rect 7484 13997 7512 14028
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 10137 14059 10195 14065
rect 8260 14028 9168 14056
rect 8260 14016 8266 14028
rect 7469 13991 7527 13997
rect 7469 13957 7481 13991
rect 7515 13957 7527 13991
rect 7469 13951 7527 13957
rect 8018 13948 8024 14000
rect 8076 13988 8082 14000
rect 8849 13991 8907 13997
rect 8849 13988 8861 13991
rect 8076 13960 8861 13988
rect 8076 13948 8082 13960
rect 8849 13957 8861 13960
rect 8895 13957 8907 13991
rect 8849 13951 8907 13957
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13889 7067 13923
rect 7009 13883 7067 13889
rect 7190 13880 7196 13932
rect 7248 13880 7254 13932
rect 7653 13923 7711 13929
rect 7653 13889 7665 13923
rect 7699 13920 7711 13923
rect 8294 13920 8300 13932
rect 7699 13892 8300 13920
rect 7699 13889 7711 13892
rect 7653 13883 7711 13889
rect 8294 13880 8300 13892
rect 8352 13880 8358 13932
rect 8386 13880 8392 13932
rect 8444 13880 8450 13932
rect 9140 13929 9168 14028
rect 10137 14025 10149 14059
rect 10183 14056 10195 14059
rect 10226 14056 10232 14068
rect 10183 14028 10232 14056
rect 10183 14025 10195 14028
rect 10137 14019 10195 14025
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 11054 14016 11060 14068
rect 11112 14016 11118 14068
rect 11885 14059 11943 14065
rect 11885 14025 11897 14059
rect 11931 14056 11943 14059
rect 13262 14056 13268 14068
rect 11931 14028 13268 14056
rect 11931 14025 11943 14028
rect 11885 14019 11943 14025
rect 13262 14016 13268 14028
rect 13320 14016 13326 14068
rect 14369 14059 14427 14065
rect 14369 14025 14381 14059
rect 14415 14056 14427 14059
rect 14415 14028 14780 14056
rect 14415 14025 14427 14028
rect 14369 14019 14427 14025
rect 9398 13948 9404 14000
rect 9456 13988 9462 14000
rect 10413 13991 10471 13997
rect 9456 13960 9996 13988
rect 9456 13948 9462 13960
rect 8573 13923 8631 13929
rect 8573 13889 8585 13923
rect 8619 13889 8631 13923
rect 8573 13883 8631 13889
rect 9125 13923 9183 13929
rect 9125 13889 9137 13923
rect 9171 13889 9183 13923
rect 9125 13883 9183 13889
rect 4709 13855 4767 13861
rect 4709 13821 4721 13855
rect 4755 13852 4767 13855
rect 4755 13824 7793 13852
rect 4755 13821 4767 13824
rect 4709 13815 4767 13821
rect 5442 13744 5448 13796
rect 5500 13784 5506 13796
rect 7765 13784 7793 13824
rect 7834 13812 7840 13864
rect 7892 13812 7898 13864
rect 8588 13852 8616 13883
rect 9490 13880 9496 13932
rect 9548 13920 9554 13932
rect 9968 13929 9996 13960
rect 10413 13957 10425 13991
rect 10459 13988 10471 13991
rect 11072 13988 11100 14016
rect 10459 13960 11100 13988
rect 10459 13957 10471 13960
rect 10413 13951 10471 13957
rect 11606 13948 11612 14000
rect 11664 13988 11670 14000
rect 14752 13988 14780 14028
rect 15654 14016 15660 14068
rect 15712 14016 15718 14068
rect 11664 13960 14504 13988
rect 14752 13960 15148 13988
rect 11664 13948 11670 13960
rect 9677 13923 9735 13929
rect 9677 13920 9689 13923
rect 9548 13892 9689 13920
rect 9548 13880 9554 13892
rect 9677 13889 9689 13892
rect 9723 13889 9735 13923
rect 9677 13883 9735 13889
rect 9953 13923 10011 13929
rect 9953 13889 9965 13923
rect 9999 13920 10011 13923
rect 10134 13920 10140 13932
rect 9999 13892 10140 13920
rect 9999 13889 10011 13892
rect 9953 13883 10011 13889
rect 10134 13880 10140 13892
rect 10192 13880 10198 13932
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13889 10655 13923
rect 10597 13883 10655 13889
rect 8404 13824 8616 13852
rect 8202 13784 8208 13796
rect 5500 13756 7696 13784
rect 7765 13756 8208 13784
rect 5500 13744 5506 13756
rect 5994 13676 6000 13728
rect 6052 13716 6058 13728
rect 6822 13716 6828 13728
rect 6052 13688 6828 13716
rect 6052 13676 6058 13688
rect 6822 13676 6828 13688
rect 6880 13716 6886 13728
rect 7098 13716 7104 13728
rect 6880 13688 7104 13716
rect 6880 13676 6886 13688
rect 7098 13676 7104 13688
rect 7156 13676 7162 13728
rect 7377 13719 7435 13725
rect 7377 13685 7389 13719
rect 7423 13716 7435 13719
rect 7558 13716 7564 13728
rect 7423 13688 7564 13716
rect 7423 13685 7435 13688
rect 7377 13679 7435 13685
rect 7558 13676 7564 13688
rect 7616 13676 7622 13728
rect 7668 13716 7696 13756
rect 8202 13744 8208 13756
rect 8260 13744 8266 13796
rect 8404 13716 8432 13824
rect 8588 13784 8616 13824
rect 8754 13812 8760 13864
rect 8812 13812 8818 13864
rect 9033 13855 9091 13861
rect 9033 13821 9045 13855
rect 9079 13852 9091 13855
rect 9508 13852 9536 13880
rect 9079 13824 9536 13852
rect 9079 13821 9091 13824
rect 9033 13815 9091 13821
rect 9858 13812 9864 13864
rect 9916 13812 9922 13864
rect 10502 13784 10508 13796
rect 8588 13756 10508 13784
rect 10502 13744 10508 13756
rect 10560 13784 10566 13796
rect 10612 13784 10640 13883
rect 11054 13880 11060 13932
rect 11112 13920 11118 13932
rect 11517 13923 11575 13929
rect 11517 13920 11529 13923
rect 11112 13892 11529 13920
rect 11112 13880 11118 13892
rect 11517 13889 11529 13892
rect 11563 13889 11575 13923
rect 11517 13883 11575 13889
rect 13906 13880 13912 13932
rect 13964 13880 13970 13932
rect 14476 13929 14504 13960
rect 14185 13923 14243 13929
rect 14185 13920 14197 13923
rect 14108 13892 14197 13920
rect 10781 13855 10839 13861
rect 10781 13821 10793 13855
rect 10827 13852 10839 13855
rect 11606 13852 11612 13864
rect 10827 13824 11612 13852
rect 10827 13821 10839 13824
rect 10781 13815 10839 13821
rect 11606 13812 11612 13824
rect 11664 13812 11670 13864
rect 12434 13812 12440 13864
rect 12492 13852 12498 13864
rect 14001 13855 14059 13861
rect 14001 13852 14013 13855
rect 12492 13824 14013 13852
rect 12492 13812 12498 13824
rect 14001 13821 14013 13824
rect 14047 13821 14059 13855
rect 14001 13815 14059 13821
rect 10560 13756 10640 13784
rect 10560 13744 10566 13756
rect 12986 13744 12992 13796
rect 13044 13784 13050 13796
rect 14108 13784 14136 13892
rect 14185 13889 14197 13892
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13889 14519 13923
rect 14461 13883 14519 13889
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13920 14703 13923
rect 14734 13920 14740 13932
rect 14691 13892 14740 13920
rect 14691 13889 14703 13892
rect 14645 13883 14703 13889
rect 14734 13880 14740 13892
rect 14792 13880 14798 13932
rect 15120 13929 15148 13960
rect 15105 13923 15163 13929
rect 15105 13889 15117 13923
rect 15151 13889 15163 13923
rect 15105 13883 15163 13889
rect 15289 13923 15347 13929
rect 15289 13889 15301 13923
rect 15335 13889 15347 13923
rect 15289 13883 15347 13889
rect 15381 13923 15439 13929
rect 15381 13889 15393 13923
rect 15427 13889 15439 13923
rect 15381 13883 15439 13889
rect 15473 13923 15531 13929
rect 15473 13889 15485 13923
rect 15519 13920 15531 13923
rect 15841 13923 15899 13929
rect 15841 13920 15853 13923
rect 15519 13892 15853 13920
rect 15519 13889 15531 13892
rect 15473 13883 15531 13889
rect 15841 13889 15853 13892
rect 15887 13889 15899 13923
rect 15841 13883 15899 13889
rect 16485 13923 16543 13929
rect 16485 13889 16497 13923
rect 16531 13920 16543 13923
rect 16758 13920 16764 13932
rect 16531 13892 16764 13920
rect 16531 13889 16543 13892
rect 16485 13883 16543 13889
rect 15304 13852 15332 13883
rect 15120 13824 15332 13852
rect 15396 13852 15424 13883
rect 16758 13880 16764 13892
rect 16816 13880 16822 13932
rect 15746 13852 15752 13864
rect 15396 13824 15752 13852
rect 15120 13796 15148 13824
rect 15746 13812 15752 13824
rect 15804 13812 15810 13864
rect 13044 13756 14136 13784
rect 13044 13744 13050 13756
rect 15102 13744 15108 13796
rect 15160 13744 15166 13796
rect 7668 13688 8432 13716
rect 9125 13719 9183 13725
rect 9125 13685 9137 13719
rect 9171 13716 9183 13719
rect 9214 13716 9220 13728
rect 9171 13688 9220 13716
rect 9171 13685 9183 13688
rect 9125 13679 9183 13685
rect 9214 13676 9220 13688
rect 9272 13676 9278 13728
rect 9306 13676 9312 13728
rect 9364 13676 9370 13728
rect 9582 13676 9588 13728
rect 9640 13716 9646 13728
rect 9677 13719 9735 13725
rect 9677 13716 9689 13719
rect 9640 13688 9689 13716
rect 9640 13676 9646 13688
rect 9677 13685 9689 13688
rect 9723 13685 9735 13719
rect 9677 13679 9735 13685
rect 9766 13676 9772 13728
rect 9824 13716 9830 13728
rect 10870 13716 10876 13728
rect 9824 13688 10876 13716
rect 9824 13676 9830 13688
rect 10870 13676 10876 13688
rect 10928 13676 10934 13728
rect 11330 13676 11336 13728
rect 11388 13716 11394 13728
rect 11517 13719 11575 13725
rect 11517 13716 11529 13719
rect 11388 13688 11529 13716
rect 11388 13676 11394 13688
rect 11517 13685 11529 13688
rect 11563 13685 11575 13719
rect 11517 13679 11575 13685
rect 13814 13676 13820 13728
rect 13872 13716 13878 13728
rect 13909 13719 13967 13725
rect 13909 13716 13921 13719
rect 13872 13688 13921 13716
rect 13872 13676 13878 13688
rect 13909 13685 13921 13688
rect 13955 13716 13967 13719
rect 14461 13719 14519 13725
rect 14461 13716 14473 13719
rect 13955 13688 14473 13716
rect 13955 13685 13967 13688
rect 13909 13679 13967 13685
rect 14461 13685 14473 13688
rect 14507 13685 14519 13719
rect 14461 13679 14519 13685
rect 14829 13719 14887 13725
rect 14829 13685 14841 13719
rect 14875 13716 14887 13719
rect 15010 13716 15016 13728
rect 14875 13688 15016 13716
rect 14875 13685 14887 13688
rect 14829 13679 14887 13685
rect 15010 13676 15016 13688
rect 15068 13676 15074 13728
rect 16942 13676 16948 13728
rect 17000 13676 17006 13728
rect 1104 13626 17388 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 17388 13626
rect 1104 13552 17388 13574
rect 4706 13512 4712 13524
rect 4264 13484 4712 13512
rect 3605 13447 3663 13453
rect 3605 13413 3617 13447
rect 3651 13444 3663 13447
rect 4062 13444 4068 13456
rect 3651 13416 4068 13444
rect 3651 13413 3663 13416
rect 3605 13407 3663 13413
rect 4062 13404 4068 13416
rect 4120 13404 4126 13456
rect 3510 13376 3516 13388
rect 3344 13348 3516 13376
rect 3142 13317 3148 13320
rect 3099 13311 3148 13317
rect 3099 13277 3111 13311
rect 3145 13277 3148 13311
rect 3099 13271 3148 13277
rect 3142 13268 3148 13271
rect 3200 13308 3206 13320
rect 3344 13308 3372 13348
rect 3510 13336 3516 13348
rect 3568 13376 3574 13388
rect 4264 13376 4292 13484
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 4801 13515 4859 13521
rect 4801 13481 4813 13515
rect 4847 13512 4859 13515
rect 4847 13484 5396 13512
rect 4847 13481 4859 13484
rect 4801 13475 4859 13481
rect 4338 13404 4344 13456
rect 4396 13444 4402 13456
rect 5368 13444 5396 13484
rect 5442 13472 5448 13524
rect 5500 13472 5506 13524
rect 6365 13515 6423 13521
rect 6365 13481 6377 13515
rect 6411 13481 6423 13515
rect 6365 13475 6423 13481
rect 5534 13444 5540 13456
rect 4396 13416 5304 13444
rect 5368 13416 5540 13444
rect 4396 13404 4402 13416
rect 3568 13348 4292 13376
rect 3568 13336 3574 13348
rect 3200 13280 3372 13308
rect 3421 13311 3479 13317
rect 3200 13268 3206 13280
rect 3421 13277 3433 13311
rect 3467 13308 3479 13311
rect 3602 13308 3608 13320
rect 3467 13280 3608 13308
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 3602 13268 3608 13280
rect 3660 13268 3666 13320
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13308 4031 13311
rect 4062 13308 4068 13320
rect 4019 13280 4068 13308
rect 4019 13277 4031 13280
rect 3973 13271 4031 13277
rect 4062 13268 4068 13280
rect 4120 13268 4126 13320
rect 4264 13317 4292 13348
rect 5166 13336 5172 13388
rect 5224 13336 5230 13388
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13277 4307 13311
rect 4249 13271 4307 13277
rect 4338 13268 4344 13320
rect 4396 13308 4402 13320
rect 4525 13311 4583 13317
rect 4525 13308 4537 13311
rect 4396 13280 4537 13308
rect 4396 13268 4402 13280
rect 4525 13277 4537 13280
rect 4571 13277 4583 13311
rect 4525 13271 4583 13277
rect 4614 13268 4620 13320
rect 4672 13268 4678 13320
rect 4706 13268 4712 13320
rect 4764 13268 4770 13320
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13308 4951 13311
rect 5184 13308 5212 13336
rect 5276 13317 5304 13416
rect 5534 13404 5540 13416
rect 5592 13404 5598 13456
rect 5810 13444 5816 13456
rect 5736 13416 5816 13444
rect 4939 13280 5212 13308
rect 5261 13311 5319 13317
rect 4939 13277 4951 13280
rect 4893 13271 4951 13277
rect 5261 13277 5273 13311
rect 5307 13277 5319 13311
rect 5261 13271 5319 13277
rect 5629 13311 5687 13317
rect 5629 13277 5641 13311
rect 5675 13308 5687 13311
rect 5736 13308 5764 13416
rect 5810 13404 5816 13416
rect 5868 13404 5874 13456
rect 6270 13404 6276 13456
rect 6328 13444 6334 13456
rect 6380 13444 6408 13475
rect 7006 13472 7012 13524
rect 7064 13472 7070 13524
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 7834 13512 7840 13524
rect 7156 13484 7840 13512
rect 7156 13472 7162 13484
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 8018 13472 8024 13524
rect 8076 13472 8082 13524
rect 9766 13512 9772 13524
rect 8128 13484 9772 13512
rect 6328 13416 6408 13444
rect 6328 13404 6334 13416
rect 6914 13404 6920 13456
rect 6972 13444 6978 13456
rect 6972 13416 7696 13444
rect 6972 13404 6978 13416
rect 7282 13376 7288 13388
rect 5828 13348 7288 13376
rect 5828 13317 5856 13348
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 5675 13280 5764 13308
rect 5813 13311 5871 13317
rect 5675 13277 5687 13280
rect 5629 13271 5687 13277
rect 5813 13277 5825 13311
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 3234 13200 3240 13252
rect 3292 13200 3298 13252
rect 3329 13243 3387 13249
rect 3329 13209 3341 13243
rect 3375 13240 3387 13243
rect 3375 13212 3464 13240
rect 3375 13209 3387 13212
rect 3329 13203 3387 13209
rect 3436 13184 3464 13212
rect 3786 13200 3792 13252
rect 3844 13200 3850 13252
rect 4356 13240 4384 13268
rect 4080 13212 4384 13240
rect 4433 13243 4491 13249
rect 3418 13132 3424 13184
rect 3476 13172 3482 13184
rect 4080 13172 4108 13212
rect 4433 13209 4445 13243
rect 4479 13209 4491 13243
rect 4724 13240 4752 13268
rect 5077 13243 5135 13249
rect 5077 13240 5089 13243
rect 4724 13212 5089 13240
rect 4433 13203 4491 13209
rect 5077 13209 5089 13212
rect 5123 13209 5135 13243
rect 5077 13203 5135 13209
rect 5169 13243 5227 13249
rect 5169 13209 5181 13243
rect 5215 13240 5227 13243
rect 5644 13240 5672 13271
rect 5215 13212 5672 13240
rect 5215 13209 5227 13212
rect 5169 13203 5227 13209
rect 3476 13144 4108 13172
rect 3476 13132 3482 13144
rect 4154 13132 4160 13184
rect 4212 13132 4218 13184
rect 4448 13172 4476 13203
rect 4706 13172 4712 13184
rect 4448 13144 4712 13172
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 5350 13132 5356 13184
rect 5408 13172 5414 13184
rect 5828 13172 5856 13271
rect 5994 13268 6000 13320
rect 6052 13268 6058 13320
rect 6454 13268 6460 13320
rect 6512 13268 6518 13320
rect 6549 13311 6607 13317
rect 6549 13277 6561 13311
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 5905 13243 5963 13249
rect 5905 13209 5917 13243
rect 5951 13240 5963 13243
rect 6086 13240 6092 13252
rect 5951 13212 6092 13240
rect 5951 13209 5963 13212
rect 5905 13203 5963 13209
rect 6086 13200 6092 13212
rect 6144 13200 6150 13252
rect 6270 13200 6276 13252
rect 6328 13200 6334 13252
rect 6564 13240 6592 13271
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 7009 13311 7067 13317
rect 7009 13308 7021 13311
rect 6788 13280 7021 13308
rect 6788 13268 6794 13280
rect 7009 13277 7021 13280
rect 7055 13277 7067 13311
rect 7009 13271 7067 13277
rect 7101 13311 7159 13317
rect 7101 13277 7113 13311
rect 7147 13308 7159 13311
rect 7190 13308 7196 13320
rect 7147 13280 7196 13308
rect 7147 13277 7159 13280
rect 7101 13271 7159 13277
rect 7190 13268 7196 13280
rect 7248 13308 7254 13320
rect 7558 13317 7564 13320
rect 7377 13311 7435 13317
rect 7377 13308 7389 13311
rect 7248 13280 7389 13308
rect 7248 13268 7254 13280
rect 7377 13277 7389 13280
rect 7423 13277 7435 13311
rect 7377 13271 7435 13277
rect 7525 13311 7564 13317
rect 7525 13277 7537 13311
rect 7525 13271 7564 13277
rect 7558 13268 7564 13271
rect 7616 13268 7622 13320
rect 7668 13317 7696 13416
rect 7742 13336 7748 13388
rect 7800 13376 7806 13388
rect 7800 13348 7885 13376
rect 7800 13336 7806 13348
rect 7857 13317 7885 13348
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13277 7711 13311
rect 7857 13311 7941 13317
rect 7857 13280 7895 13311
rect 7653 13271 7711 13277
rect 7883 13277 7895 13280
rect 7929 13277 7941 13311
rect 7883 13271 7941 13277
rect 6638 13240 6644 13252
rect 6564 13212 6644 13240
rect 5408 13144 5856 13172
rect 6181 13175 6239 13181
rect 5408 13132 5414 13144
rect 6181 13141 6193 13175
rect 6227 13172 6239 13175
rect 6564 13172 6592 13212
rect 6638 13200 6644 13212
rect 6696 13200 6702 13252
rect 7285 13243 7343 13249
rect 7285 13240 7297 13243
rect 6748 13212 7297 13240
rect 6748 13181 6776 13212
rect 7285 13209 7297 13212
rect 7331 13209 7343 13243
rect 7285 13203 7343 13209
rect 7745 13243 7803 13249
rect 7745 13209 7757 13243
rect 7791 13240 7803 13243
rect 8018 13240 8024 13252
rect 7791 13212 8024 13240
rect 7791 13209 7803 13212
rect 7745 13203 7803 13209
rect 8018 13200 8024 13212
rect 8076 13200 8082 13252
rect 6227 13144 6592 13172
rect 6733 13175 6791 13181
rect 6227 13141 6239 13144
rect 6181 13135 6239 13141
rect 6733 13141 6745 13175
rect 6779 13141 6791 13175
rect 6733 13135 6791 13141
rect 6822 13132 6828 13184
rect 6880 13132 6886 13184
rect 7006 13132 7012 13184
rect 7064 13172 7070 13184
rect 8128 13172 8156 13484
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 9953 13515 10011 13521
rect 9953 13481 9965 13515
rect 9999 13512 10011 13515
rect 10042 13512 10048 13524
rect 9999 13484 10048 13512
rect 9999 13481 10011 13484
rect 9953 13475 10011 13481
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 10502 13472 10508 13524
rect 10560 13472 10566 13524
rect 10873 13515 10931 13521
rect 10873 13481 10885 13515
rect 10919 13512 10931 13515
rect 12434 13512 12440 13524
rect 10919 13484 12440 13512
rect 10919 13481 10931 13484
rect 10873 13475 10931 13481
rect 12434 13472 12440 13484
rect 12492 13472 12498 13524
rect 12529 13515 12587 13521
rect 12529 13481 12541 13515
rect 12575 13481 12587 13515
rect 12529 13475 12587 13481
rect 12544 13444 12572 13475
rect 12986 13472 12992 13524
rect 13044 13472 13050 13524
rect 13262 13472 13268 13524
rect 13320 13512 13326 13524
rect 14093 13515 14151 13521
rect 14093 13512 14105 13515
rect 13320 13484 14105 13512
rect 13320 13472 13326 13484
rect 14093 13481 14105 13484
rect 14139 13481 14151 13515
rect 14093 13475 14151 13481
rect 15194 13472 15200 13524
rect 15252 13512 15258 13524
rect 15252 13484 15700 13512
rect 15252 13472 15258 13484
rect 12406 13416 12572 13444
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 10042 13376 10048 13388
rect 9732 13348 10048 13376
rect 9732 13336 9738 13348
rect 10042 13336 10048 13348
rect 10100 13336 10106 13388
rect 10410 13336 10416 13388
rect 10468 13376 10474 13388
rect 10505 13379 10563 13385
rect 10505 13376 10517 13379
rect 10468 13348 10517 13376
rect 10468 13336 10474 13348
rect 10505 13345 10517 13348
rect 10551 13345 10563 13379
rect 10505 13339 10563 13345
rect 8202 13268 8208 13320
rect 8260 13308 8266 13320
rect 9582 13308 9588 13320
rect 8260 13280 9588 13308
rect 8260 13268 8266 13280
rect 9582 13268 9588 13280
rect 9640 13268 9646 13320
rect 9766 13268 9772 13320
rect 9824 13308 9830 13320
rect 10689 13311 10747 13317
rect 10689 13308 10701 13311
rect 9824 13280 10701 13308
rect 9824 13268 9830 13280
rect 10689 13277 10701 13280
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 10410 13200 10416 13252
rect 10468 13200 10474 13252
rect 12406 13240 12434 13416
rect 13998 13404 14004 13456
rect 14056 13444 14062 13456
rect 14553 13447 14611 13453
rect 14553 13444 14565 13447
rect 14056 13416 14565 13444
rect 14056 13404 14062 13416
rect 14553 13413 14565 13416
rect 14599 13413 14611 13447
rect 14553 13407 14611 13413
rect 15672 13388 15700 13484
rect 12618 13336 12624 13388
rect 12676 13336 12682 13388
rect 14274 13336 14280 13388
rect 14332 13336 14338 13388
rect 15654 13336 15660 13388
rect 15712 13336 15718 13388
rect 12526 13268 12532 13320
rect 12584 13268 12590 13320
rect 12802 13268 12808 13320
rect 12860 13268 12866 13320
rect 14369 13311 14427 13317
rect 14369 13277 14381 13311
rect 14415 13308 14427 13311
rect 14458 13308 14464 13320
rect 14415 13280 14464 13308
rect 14415 13277 14427 13280
rect 14369 13271 14427 13277
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 15010 13268 15016 13320
rect 15068 13268 15074 13320
rect 15378 13268 15384 13320
rect 15436 13268 15442 13320
rect 10520 13212 12434 13240
rect 12544 13240 12572 13268
rect 13262 13240 13268 13252
rect 12544 13212 13268 13240
rect 7064 13144 8156 13172
rect 7064 13132 7070 13144
rect 9214 13132 9220 13184
rect 9272 13172 9278 13184
rect 10520 13172 10548 13212
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 14090 13200 14096 13252
rect 14148 13200 14154 13252
rect 15194 13200 15200 13252
rect 15252 13200 15258 13252
rect 15286 13200 15292 13252
rect 15344 13200 15350 13252
rect 15902 13243 15960 13249
rect 15902 13209 15914 13243
rect 15948 13209 15960 13243
rect 15902 13203 15960 13209
rect 9272 13144 10548 13172
rect 9272 13132 9278 13144
rect 10686 13132 10692 13184
rect 10744 13172 10750 13184
rect 12894 13172 12900 13184
rect 10744 13144 12900 13172
rect 10744 13132 10750 13144
rect 12894 13132 12900 13144
rect 12952 13132 12958 13184
rect 15565 13175 15623 13181
rect 15565 13141 15577 13175
rect 15611 13172 15623 13175
rect 15917 13172 15945 13203
rect 15611 13144 15945 13172
rect 17037 13175 17095 13181
rect 15611 13141 15623 13144
rect 15565 13135 15623 13141
rect 17037 13141 17049 13175
rect 17083 13172 17095 13175
rect 17083 13144 17448 13172
rect 17083 13141 17095 13144
rect 17037 13135 17095 13141
rect 1104 13082 17388 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 17388 13082
rect 1104 13008 17388 13030
rect 3786 12928 3792 12980
rect 3844 12968 3850 12980
rect 4522 12968 4528 12980
rect 3844 12940 4528 12968
rect 3844 12928 3850 12940
rect 4522 12928 4528 12940
rect 4580 12928 4586 12980
rect 6086 12968 6092 12980
rect 5552 12940 6092 12968
rect 2866 12860 2872 12912
rect 2924 12900 2930 12912
rect 3513 12903 3571 12909
rect 3513 12900 3525 12903
rect 2924 12872 3525 12900
rect 2924 12860 2930 12872
rect 3513 12869 3525 12872
rect 3559 12869 3571 12903
rect 3513 12863 3571 12869
rect 4801 12903 4859 12909
rect 4801 12869 4813 12903
rect 4847 12900 4859 12903
rect 5350 12900 5356 12912
rect 4847 12872 5356 12900
rect 4847 12869 4859 12872
rect 4801 12863 4859 12869
rect 5350 12860 5356 12872
rect 5408 12860 5414 12912
rect 3050 12792 3056 12844
rect 3108 12832 3114 12844
rect 3237 12835 3295 12841
rect 3237 12832 3249 12835
rect 3108 12804 3249 12832
rect 3108 12792 3114 12804
rect 3237 12801 3249 12804
rect 3283 12801 3295 12835
rect 3237 12795 3295 12801
rect 3326 12792 3332 12844
rect 3384 12832 3390 12844
rect 3421 12835 3479 12841
rect 3421 12832 3433 12835
rect 3384 12804 3433 12832
rect 3384 12792 3390 12804
rect 3421 12801 3433 12804
rect 3467 12801 3479 12835
rect 3421 12795 3479 12801
rect 3602 12792 3608 12844
rect 3660 12792 3666 12844
rect 4525 12835 4583 12841
rect 4525 12801 4537 12835
rect 4571 12801 4583 12835
rect 4525 12795 4583 12801
rect 4540 12628 4568 12795
rect 4706 12792 4712 12844
rect 4764 12792 4770 12844
rect 4893 12835 4951 12841
rect 4893 12801 4905 12835
rect 4939 12801 4951 12835
rect 4893 12795 4951 12801
rect 4614 12724 4620 12776
rect 4672 12764 4678 12776
rect 4908 12764 4936 12795
rect 5166 12792 5172 12844
rect 5224 12832 5230 12844
rect 5552 12841 5580 12940
rect 6086 12928 6092 12940
rect 6144 12968 6150 12980
rect 6144 12940 7144 12968
rect 6144 12928 6150 12940
rect 6270 12860 6276 12912
rect 6328 12900 6334 12912
rect 7006 12900 7012 12912
rect 6328 12872 7012 12900
rect 6328 12860 6334 12872
rect 7006 12860 7012 12872
rect 7064 12860 7070 12912
rect 7116 12844 7144 12940
rect 7558 12928 7564 12980
rect 7616 12968 7622 12980
rect 8202 12968 8208 12980
rect 7616 12940 8208 12968
rect 7616 12928 7622 12940
rect 8202 12928 8208 12940
rect 8260 12928 8266 12980
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 10597 12971 10655 12977
rect 10597 12968 10609 12971
rect 10560 12940 10609 12968
rect 10560 12928 10566 12940
rect 10597 12937 10609 12940
rect 10643 12937 10655 12971
rect 12434 12968 12440 12980
rect 10597 12931 10655 12937
rect 11716 12940 12440 12968
rect 8754 12860 8760 12912
rect 8812 12900 8818 12912
rect 10686 12900 10692 12912
rect 8812 12872 10692 12900
rect 8812 12860 8818 12872
rect 10686 12860 10692 12872
rect 10744 12860 10750 12912
rect 5537 12835 5595 12841
rect 5537 12832 5549 12835
rect 5224 12804 5549 12832
rect 5224 12792 5230 12804
rect 5537 12801 5549 12804
rect 5583 12801 5595 12835
rect 5537 12795 5595 12801
rect 5721 12835 5779 12841
rect 5721 12801 5733 12835
rect 5767 12801 5779 12835
rect 5721 12795 5779 12801
rect 5626 12764 5632 12776
rect 4672 12736 4936 12764
rect 5092 12736 5632 12764
rect 4672 12724 4678 12736
rect 5092 12705 5120 12736
rect 5626 12724 5632 12736
rect 5684 12724 5690 12776
rect 5077 12699 5135 12705
rect 5077 12665 5089 12699
rect 5123 12665 5135 12699
rect 5736 12696 5764 12795
rect 5810 12792 5816 12844
rect 5868 12792 5874 12844
rect 5905 12835 5963 12841
rect 5905 12801 5917 12835
rect 5951 12801 5963 12835
rect 5905 12795 5963 12801
rect 5920 12764 5948 12795
rect 6086 12792 6092 12844
rect 6144 12832 6150 12844
rect 6454 12832 6460 12844
rect 6144 12804 6460 12832
rect 6144 12792 6150 12804
rect 6454 12792 6460 12804
rect 6512 12792 6518 12844
rect 7098 12792 7104 12844
rect 7156 12792 7162 12844
rect 7282 12792 7288 12844
rect 7340 12792 7346 12844
rect 7374 12792 7380 12844
rect 7432 12792 7438 12844
rect 7469 12835 7527 12841
rect 7469 12801 7481 12835
rect 7515 12832 7527 12835
rect 7834 12832 7840 12844
rect 7515 12804 7840 12832
rect 7515 12801 7527 12804
rect 7469 12795 7527 12801
rect 7834 12792 7840 12804
rect 7892 12792 7898 12844
rect 10502 12792 10508 12844
rect 10560 12832 10566 12844
rect 10781 12835 10839 12841
rect 10781 12832 10793 12835
rect 10560 12804 10793 12832
rect 10560 12792 10566 12804
rect 10781 12801 10793 12804
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 10870 12792 10876 12844
rect 10928 12832 10934 12844
rect 10965 12835 11023 12841
rect 10965 12832 10977 12835
rect 10928 12804 10977 12832
rect 10928 12792 10934 12804
rect 10965 12801 10977 12804
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 8018 12764 8024 12776
rect 5920 12736 8024 12764
rect 8018 12724 8024 12736
rect 8076 12724 8082 12776
rect 8938 12724 8944 12776
rect 8996 12764 9002 12776
rect 11716 12764 11744 12940
rect 12434 12928 12440 12940
rect 12492 12928 12498 12980
rect 12526 12928 12532 12980
rect 12584 12968 12590 12980
rect 12805 12971 12863 12977
rect 12584 12940 12756 12968
rect 12584 12928 12590 12940
rect 12342 12860 12348 12912
rect 12400 12860 12406 12912
rect 12728 12900 12756 12940
rect 12805 12937 12817 12971
rect 12851 12968 12863 12971
rect 14090 12968 14096 12980
rect 12851 12940 14096 12968
rect 12851 12937 12863 12940
rect 12805 12931 12863 12937
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 14366 12928 14372 12980
rect 14424 12968 14430 12980
rect 14645 12971 14703 12977
rect 14645 12968 14657 12971
rect 14424 12940 14657 12968
rect 14424 12928 14430 12940
rect 14645 12937 14657 12940
rect 14691 12937 14703 12971
rect 14645 12931 14703 12937
rect 15378 12928 15384 12980
rect 15436 12968 15442 12980
rect 15841 12971 15899 12977
rect 15841 12968 15853 12971
rect 15436 12940 15853 12968
rect 15436 12928 15442 12940
rect 15841 12937 15853 12940
rect 15887 12937 15899 12971
rect 15841 12931 15899 12937
rect 16942 12928 16948 12980
rect 17000 12928 17006 12980
rect 12728 12872 13032 12900
rect 12434 12792 12440 12844
rect 12492 12832 12498 12844
rect 12621 12835 12679 12841
rect 12621 12832 12633 12835
rect 12492 12804 12633 12832
rect 12492 12792 12498 12804
rect 12621 12801 12633 12804
rect 12667 12832 12679 12835
rect 12802 12832 12808 12844
rect 12667 12804 12808 12832
rect 12667 12801 12679 12804
rect 12621 12795 12679 12801
rect 12802 12792 12808 12804
rect 12860 12792 12866 12844
rect 12894 12792 12900 12844
rect 12952 12792 12958 12844
rect 13004 12841 13032 12872
rect 15562 12860 15568 12912
rect 15620 12900 15626 12912
rect 15746 12900 15752 12912
rect 15620 12872 15752 12900
rect 15620 12860 15626 12872
rect 15746 12860 15752 12872
rect 15804 12860 15810 12912
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 13078 12792 13084 12844
rect 13136 12832 13142 12844
rect 14277 12835 14335 12841
rect 14277 12832 14289 12835
rect 13136 12804 14289 12832
rect 13136 12792 13142 12804
rect 14277 12801 14289 12804
rect 14323 12801 14335 12835
rect 14277 12795 14335 12801
rect 14458 12792 14464 12844
rect 14516 12792 14522 12844
rect 16485 12835 16543 12841
rect 16485 12801 16497 12835
rect 16531 12832 16543 12835
rect 16761 12835 16819 12841
rect 16761 12832 16773 12835
rect 16531 12804 16773 12832
rect 16531 12801 16543 12804
rect 16485 12795 16543 12801
rect 16761 12801 16773 12804
rect 16807 12832 16819 12835
rect 17420 12832 17448 13144
rect 16807 12804 17448 12832
rect 16807 12801 16819 12804
rect 16761 12795 16819 12801
rect 8996 12736 11744 12764
rect 12529 12767 12587 12773
rect 8996 12724 9002 12736
rect 12529 12733 12541 12767
rect 12575 12764 12587 12767
rect 12575 12736 12940 12764
rect 12575 12733 12587 12736
rect 12529 12727 12587 12733
rect 7558 12696 7564 12708
rect 5736 12668 7564 12696
rect 5077 12659 5135 12665
rect 7558 12656 7564 12668
rect 7616 12656 7622 12708
rect 7926 12656 7932 12708
rect 7984 12696 7990 12708
rect 9214 12696 9220 12708
rect 7984 12668 9220 12696
rect 7984 12656 7990 12668
rect 9214 12656 9220 12668
rect 9272 12656 9278 12708
rect 11422 12656 11428 12708
rect 11480 12696 11486 12708
rect 12544 12696 12572 12727
rect 11480 12668 12572 12696
rect 11480 12656 11486 12668
rect 5994 12628 6000 12640
rect 4540 12600 6000 12628
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 6089 12631 6147 12637
rect 6089 12597 6101 12631
rect 6135 12628 6147 12631
rect 6270 12628 6276 12640
rect 6135 12600 6276 12628
rect 6135 12597 6147 12600
rect 6089 12591 6147 12597
rect 6270 12588 6276 12600
rect 6328 12588 6334 12640
rect 7653 12631 7711 12637
rect 7653 12597 7665 12631
rect 7699 12628 7711 12631
rect 12158 12628 12164 12640
rect 7699 12600 12164 12628
rect 7699 12597 7711 12600
rect 7653 12591 7711 12597
rect 12158 12588 12164 12600
rect 12216 12628 12222 12640
rect 12912 12637 12940 12736
rect 13262 12656 13268 12708
rect 13320 12656 13326 12708
rect 12345 12631 12403 12637
rect 12345 12628 12357 12631
rect 12216 12600 12357 12628
rect 12216 12588 12222 12600
rect 12345 12597 12357 12600
rect 12391 12597 12403 12631
rect 12345 12591 12403 12597
rect 12897 12631 12955 12637
rect 12897 12597 12909 12631
rect 12943 12597 12955 12631
rect 12897 12591 12955 12597
rect 1104 12538 17388 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 17388 12538
rect 1104 12464 17388 12486
rect 2961 12427 3019 12433
rect 2961 12393 2973 12427
rect 3007 12424 3019 12427
rect 5718 12424 5724 12436
rect 3007 12396 5724 12424
rect 3007 12393 3019 12396
rect 2961 12387 3019 12393
rect 5718 12384 5724 12396
rect 5776 12384 5782 12436
rect 6270 12384 6276 12436
rect 6328 12424 6334 12436
rect 6549 12427 6607 12433
rect 6549 12424 6561 12427
rect 6328 12396 6561 12424
rect 6328 12384 6334 12396
rect 6549 12393 6561 12396
rect 6595 12424 6607 12427
rect 7193 12427 7251 12433
rect 6595 12396 7144 12424
rect 6595 12393 6607 12396
rect 6549 12387 6607 12393
rect 4264 12328 5028 12356
rect 3878 12288 3884 12300
rect 3068 12260 3884 12288
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12189 2467 12223
rect 2409 12183 2467 12189
rect 2685 12223 2743 12229
rect 2685 12189 2697 12223
rect 2731 12189 2743 12223
rect 2685 12183 2743 12189
rect 2424 12084 2452 12183
rect 2590 12112 2596 12164
rect 2648 12112 2654 12164
rect 2700 12152 2728 12183
rect 2774 12180 2780 12232
rect 2832 12180 2838 12232
rect 3068 12229 3096 12260
rect 3878 12248 3884 12260
rect 3936 12288 3942 12300
rect 4264 12288 4292 12328
rect 3936 12260 4292 12288
rect 3936 12248 3942 12260
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12189 3111 12223
rect 3053 12183 3111 12189
rect 2866 12152 2872 12164
rect 2700 12124 2872 12152
rect 2866 12112 2872 12124
rect 2924 12152 2930 12164
rect 3068 12152 3096 12183
rect 3234 12180 3240 12232
rect 3292 12180 3298 12232
rect 3421 12223 3479 12229
rect 3421 12189 3433 12223
rect 3467 12220 3479 12223
rect 3602 12220 3608 12232
rect 3467 12192 3608 12220
rect 3467 12189 3479 12192
rect 3421 12183 3479 12189
rect 3602 12180 3608 12192
rect 3660 12180 3666 12232
rect 4264 12229 4292 12260
rect 4540 12260 4936 12288
rect 4540 12229 4568 12260
rect 4249 12223 4307 12229
rect 4249 12189 4261 12223
rect 4295 12189 4307 12223
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 4249 12183 4307 12189
rect 4356 12192 4537 12220
rect 4356 12164 4384 12192
rect 4525 12189 4537 12192
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 4614 12180 4620 12232
rect 4672 12180 4678 12232
rect 4908 12229 4936 12260
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12189 4951 12223
rect 5000 12220 5028 12328
rect 6362 12316 6368 12368
rect 6420 12356 6426 12368
rect 6420 12328 6500 12356
rect 6420 12316 6426 12328
rect 6472 12297 6500 12328
rect 6457 12291 6515 12297
rect 6457 12257 6469 12291
rect 6503 12257 6515 12291
rect 6822 12288 6828 12300
rect 6457 12251 6515 12257
rect 6564 12260 6828 12288
rect 6564 12229 6592 12260
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 7116 12288 7144 12396
rect 7193 12393 7205 12427
rect 7239 12424 7251 12427
rect 7650 12424 7656 12436
rect 7239 12396 7656 12424
rect 7239 12393 7251 12396
rect 7193 12387 7251 12393
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 7926 12384 7932 12436
rect 7984 12384 7990 12436
rect 8478 12384 8484 12436
rect 8536 12424 8542 12436
rect 8757 12427 8815 12433
rect 8757 12424 8769 12427
rect 8536 12396 8769 12424
rect 8536 12384 8542 12396
rect 8757 12393 8769 12396
rect 8803 12393 8815 12427
rect 8757 12387 8815 12393
rect 9214 12384 9220 12436
rect 9272 12384 9278 12436
rect 9585 12427 9643 12433
rect 9585 12424 9597 12427
rect 9324 12396 9597 12424
rect 7668 12356 7696 12384
rect 9324 12356 9352 12396
rect 9585 12393 9597 12396
rect 9631 12424 9643 12427
rect 10597 12427 10655 12433
rect 9631 12396 10548 12424
rect 9631 12393 9643 12396
rect 9585 12387 9643 12393
rect 7668 12328 9352 12356
rect 9398 12316 9404 12368
rect 9456 12356 9462 12368
rect 9456 12328 10456 12356
rect 9456 12316 9462 12328
rect 7116 12260 7880 12288
rect 5261 12223 5319 12229
rect 5261 12220 5273 12223
rect 5000 12192 5273 12220
rect 4893 12183 4951 12189
rect 5261 12189 5273 12192
rect 5307 12189 5319 12223
rect 5261 12183 5319 12189
rect 6273 12223 6331 12229
rect 6273 12189 6285 12223
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 6687 12192 6776 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 2924 12124 3096 12152
rect 3329 12155 3387 12161
rect 2924 12112 2930 12124
rect 3329 12121 3341 12155
rect 3375 12152 3387 12155
rect 4338 12152 4344 12164
rect 3375 12124 4344 12152
rect 3375 12121 3387 12124
rect 3329 12115 3387 12121
rect 3050 12084 3056 12096
rect 2424 12056 3056 12084
rect 3050 12044 3056 12056
rect 3108 12084 3114 12096
rect 3344 12084 3372 12115
rect 4338 12112 4344 12124
rect 4396 12112 4402 12164
rect 4430 12112 4436 12164
rect 4488 12112 4494 12164
rect 4706 12112 4712 12164
rect 4764 12152 4770 12164
rect 5074 12152 5080 12164
rect 4764 12124 5080 12152
rect 4764 12112 4770 12124
rect 5074 12112 5080 12124
rect 5132 12112 5138 12164
rect 5166 12112 5172 12164
rect 5224 12112 5230 12164
rect 6288 12152 6316 12183
rect 6362 12152 6368 12164
rect 6288 12124 6368 12152
rect 6362 12112 6368 12124
rect 6420 12112 6426 12164
rect 3108 12056 3372 12084
rect 3605 12087 3663 12093
rect 3108 12044 3114 12056
rect 3605 12053 3617 12087
rect 3651 12084 3663 12087
rect 4522 12084 4528 12096
rect 3651 12056 4528 12084
rect 3651 12053 3663 12056
rect 3605 12047 3663 12053
rect 4522 12044 4528 12056
rect 4580 12044 4586 12096
rect 4801 12087 4859 12093
rect 4801 12053 4813 12087
rect 4847 12084 4859 12087
rect 5258 12084 5264 12096
rect 4847 12056 5264 12084
rect 4847 12053 4859 12056
rect 4801 12047 4859 12053
rect 5258 12044 5264 12056
rect 5316 12044 5322 12096
rect 5445 12087 5503 12093
rect 5445 12053 5457 12087
rect 5491 12084 5503 12087
rect 5994 12084 6000 12096
rect 5491 12056 6000 12084
rect 5491 12053 5503 12056
rect 5445 12047 5503 12053
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6089 12087 6147 12093
rect 6089 12053 6101 12087
rect 6135 12084 6147 12087
rect 6454 12084 6460 12096
rect 6135 12056 6460 12084
rect 6135 12053 6147 12056
rect 6089 12047 6147 12053
rect 6454 12044 6460 12056
rect 6512 12044 6518 12096
rect 6748 12084 6776 12192
rect 6914 12180 6920 12232
rect 6972 12180 6978 12232
rect 7009 12223 7067 12229
rect 7009 12189 7021 12223
rect 7055 12220 7067 12223
rect 7098 12220 7104 12232
rect 7055 12192 7104 12220
rect 7055 12189 7067 12192
rect 7009 12183 7067 12189
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 7282 12180 7288 12232
rect 7340 12180 7346 12232
rect 7374 12180 7380 12232
rect 7432 12220 7438 12232
rect 7750 12223 7808 12229
rect 7432 12192 7477 12220
rect 7432 12180 7438 12192
rect 7750 12189 7762 12223
rect 7796 12189 7808 12223
rect 7750 12183 7808 12189
rect 6825 12155 6883 12161
rect 6825 12121 6837 12155
rect 6871 12152 6883 12155
rect 7190 12152 7196 12164
rect 6871 12124 7196 12152
rect 6871 12121 6883 12124
rect 6825 12115 6883 12121
rect 7190 12112 7196 12124
rect 7248 12152 7254 12164
rect 7561 12155 7619 12161
rect 7561 12152 7573 12155
rect 7248 12124 7573 12152
rect 7248 12112 7254 12124
rect 7561 12121 7573 12124
rect 7607 12121 7619 12155
rect 7561 12115 7619 12121
rect 7650 12112 7656 12164
rect 7708 12112 7714 12164
rect 7006 12084 7012 12096
rect 6748 12056 7012 12084
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 7765 12084 7793 12183
rect 7156 12056 7793 12084
rect 7852 12084 7880 12260
rect 8478 12248 8484 12300
rect 8536 12288 8542 12300
rect 9125 12291 9183 12297
rect 9125 12288 9137 12291
rect 8536 12260 9137 12288
rect 8536 12248 8542 12260
rect 9125 12257 9137 12260
rect 9171 12257 9183 12291
rect 9125 12251 9183 12257
rect 9214 12248 9220 12300
rect 9272 12288 9278 12300
rect 10428 12297 10456 12328
rect 9677 12291 9735 12297
rect 9677 12288 9689 12291
rect 9272 12260 9689 12288
rect 9272 12248 9278 12260
rect 9677 12257 9689 12260
rect 9723 12257 9735 12291
rect 9677 12251 9735 12257
rect 10413 12291 10471 12297
rect 10413 12257 10425 12291
rect 10459 12257 10471 12291
rect 10520 12288 10548 12396
rect 10597 12393 10609 12427
rect 10643 12424 10655 12427
rect 10686 12424 10692 12436
rect 10643 12396 10692 12424
rect 10643 12393 10655 12396
rect 10597 12387 10655 12393
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 10870 12384 10876 12436
rect 10928 12424 10934 12436
rect 11149 12427 11207 12433
rect 11149 12424 11161 12427
rect 10928 12396 11161 12424
rect 10928 12384 10934 12396
rect 11149 12393 11161 12396
rect 11195 12424 11207 12427
rect 11425 12427 11483 12433
rect 11425 12424 11437 12427
rect 11195 12396 11437 12424
rect 11195 12393 11207 12396
rect 11149 12387 11207 12393
rect 11425 12393 11437 12396
rect 11471 12393 11483 12427
rect 11425 12387 11483 12393
rect 12526 12384 12532 12436
rect 12584 12384 12590 12436
rect 10781 12359 10839 12365
rect 10781 12325 10793 12359
rect 10827 12356 10839 12359
rect 10962 12356 10968 12368
rect 10827 12328 10968 12356
rect 10827 12325 10839 12328
rect 10781 12319 10839 12325
rect 10962 12316 10968 12328
rect 11020 12316 11026 12368
rect 10520 12260 11376 12288
rect 10413 12251 10471 12257
rect 8386 12180 8392 12232
rect 8444 12180 8450 12232
rect 8938 12180 8944 12232
rect 8996 12220 9002 12232
rect 9309 12223 9367 12229
rect 9309 12220 9321 12223
rect 8996 12192 9321 12220
rect 8996 12180 9002 12192
rect 9309 12189 9321 12192
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 9416 12192 9720 12220
rect 8478 12112 8484 12164
rect 8536 12152 8542 12164
rect 8573 12155 8631 12161
rect 8573 12152 8585 12155
rect 8536 12124 8585 12152
rect 8536 12112 8542 12124
rect 8573 12121 8585 12124
rect 8619 12121 8631 12155
rect 8573 12115 8631 12121
rect 9030 12112 9036 12164
rect 9088 12112 9094 12164
rect 9416 12084 9444 12192
rect 9582 12112 9588 12164
rect 9640 12112 9646 12164
rect 9692 12152 9720 12192
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 9861 12223 9919 12229
rect 9861 12220 9873 12223
rect 9824 12192 9873 12220
rect 9824 12180 9830 12192
rect 9861 12189 9873 12192
rect 9907 12189 9919 12223
rect 9861 12183 9919 12189
rect 9968 12192 10456 12220
rect 9968 12152 9996 12192
rect 10321 12155 10379 12161
rect 10321 12152 10333 12155
rect 9692 12124 9996 12152
rect 10060 12124 10333 12152
rect 7852 12056 9444 12084
rect 9493 12087 9551 12093
rect 7156 12044 7162 12056
rect 9493 12053 9505 12087
rect 9539 12084 9551 12087
rect 9766 12084 9772 12096
rect 9539 12056 9772 12084
rect 9539 12053 9551 12056
rect 9493 12047 9551 12053
rect 9766 12044 9772 12056
rect 9824 12044 9830 12096
rect 10060 12093 10088 12124
rect 10321 12121 10333 12124
rect 10367 12121 10379 12155
rect 10428 12152 10456 12192
rect 10594 12180 10600 12232
rect 10652 12180 10658 12232
rect 11054 12180 11060 12232
rect 11112 12180 11118 12232
rect 11146 12180 11152 12232
rect 11204 12180 11210 12232
rect 11348 12220 11376 12260
rect 11514 12248 11520 12300
rect 11572 12288 11578 12300
rect 11609 12291 11667 12297
rect 11609 12288 11621 12291
rect 11572 12260 11621 12288
rect 11572 12248 11578 12260
rect 11609 12257 11621 12260
rect 11655 12288 11667 12291
rect 12158 12288 12164 12300
rect 11655 12260 12164 12288
rect 11655 12257 11667 12260
rect 11609 12251 11667 12257
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 12434 12248 12440 12300
rect 12492 12288 12498 12300
rect 13262 12288 13268 12300
rect 12492 12260 13268 12288
rect 12492 12248 12498 12260
rect 13262 12248 13268 12260
rect 13320 12248 13326 12300
rect 15562 12288 15568 12300
rect 15304 12260 15568 12288
rect 11422 12220 11428 12232
rect 11480 12229 11486 12232
rect 11348 12192 11428 12220
rect 11422 12180 11428 12192
rect 11480 12183 11490 12229
rect 11701 12223 11759 12229
rect 11701 12189 11713 12223
rect 11747 12189 11759 12223
rect 11701 12183 11759 12189
rect 11480 12180 11486 12183
rect 10873 12155 10931 12161
rect 10873 12152 10885 12155
rect 10428 12124 10885 12152
rect 10321 12115 10379 12121
rect 10873 12121 10885 12124
rect 10919 12121 10931 12155
rect 11716 12152 11744 12183
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 12253 12223 12311 12229
rect 12253 12220 12265 12223
rect 12124 12192 12265 12220
rect 12124 12180 12130 12192
rect 12253 12189 12265 12192
rect 12299 12189 12311 12223
rect 12253 12183 12311 12189
rect 12526 12180 12532 12232
rect 12584 12180 12590 12232
rect 15013 12223 15071 12229
rect 15013 12189 15025 12223
rect 15059 12220 15071 12223
rect 15102 12220 15108 12232
rect 15059 12192 15108 12220
rect 15059 12189 15071 12192
rect 15013 12183 15071 12189
rect 15102 12180 15108 12192
rect 15160 12180 15166 12232
rect 15304 12229 15332 12260
rect 15562 12248 15568 12260
rect 15620 12288 15626 12300
rect 15620 12260 15792 12288
rect 15620 12248 15626 12260
rect 15764 12232 15792 12260
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12189 15347 12223
rect 15289 12183 15347 12189
rect 15378 12180 15384 12232
rect 15436 12180 15442 12232
rect 15654 12180 15660 12232
rect 15712 12180 15718 12232
rect 15746 12180 15752 12232
rect 15804 12180 15810 12232
rect 14642 12152 14648 12164
rect 10873 12115 10931 12121
rect 11072 12124 11744 12152
rect 12406 12124 14648 12152
rect 10045 12087 10103 12093
rect 10045 12053 10057 12087
rect 10091 12053 10103 12087
rect 10045 12047 10103 12053
rect 10686 12044 10692 12096
rect 10744 12084 10750 12096
rect 11072 12084 11100 12124
rect 10744 12056 11100 12084
rect 10744 12044 10750 12056
rect 11330 12044 11336 12096
rect 11388 12044 11394 12096
rect 11885 12087 11943 12093
rect 11885 12053 11897 12087
rect 11931 12084 11943 12087
rect 12406 12084 12434 12124
rect 14642 12112 14648 12124
rect 14700 12112 14706 12164
rect 15197 12155 15255 12161
rect 15197 12121 15209 12155
rect 15243 12121 15255 12155
rect 15902 12155 15960 12161
rect 15902 12152 15914 12155
rect 15197 12115 15255 12121
rect 15580 12124 15914 12152
rect 11931 12056 12434 12084
rect 11931 12053 11943 12056
rect 11885 12047 11943 12053
rect 12710 12044 12716 12096
rect 12768 12044 12774 12096
rect 15212 12084 15240 12115
rect 15470 12084 15476 12096
rect 15212 12056 15476 12084
rect 15470 12044 15476 12056
rect 15528 12044 15534 12096
rect 15580 12093 15608 12124
rect 15902 12121 15914 12124
rect 15948 12121 15960 12155
rect 15902 12115 15960 12121
rect 15565 12087 15623 12093
rect 15565 12053 15577 12087
rect 15611 12053 15623 12087
rect 15565 12047 15623 12053
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 17037 12087 17095 12093
rect 17037 12084 17049 12087
rect 16632 12056 17049 12084
rect 16632 12044 16638 12056
rect 17037 12053 17049 12056
rect 17083 12053 17095 12087
rect 17037 12047 17095 12053
rect 1104 11994 17388 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 17388 11994
rect 1104 11920 17388 11942
rect 3234 11840 3240 11892
rect 3292 11840 3298 11892
rect 3786 11840 3792 11892
rect 3844 11840 3850 11892
rect 4614 11840 4620 11892
rect 4672 11880 4678 11892
rect 5077 11883 5135 11889
rect 4672 11852 4936 11880
rect 4672 11840 4678 11852
rect 3252 11812 3280 11840
rect 3421 11815 3479 11821
rect 3421 11812 3433 11815
rect 3252 11784 3433 11812
rect 3421 11781 3433 11784
rect 3467 11781 3479 11815
rect 3421 11775 3479 11781
rect 3878 11772 3884 11824
rect 3936 11812 3942 11824
rect 4801 11815 4859 11821
rect 4801 11812 4813 11815
rect 3936 11784 4813 11812
rect 3936 11772 3942 11784
rect 4801 11781 4813 11784
rect 4847 11781 4859 11815
rect 4801 11775 4859 11781
rect 3237 11747 3295 11753
rect 3237 11713 3249 11747
rect 3283 11744 3295 11747
rect 3326 11744 3332 11756
rect 3283 11716 3332 11744
rect 3283 11713 3295 11716
rect 3237 11707 3295 11713
rect 3326 11704 3332 11716
rect 3384 11704 3390 11756
rect 3510 11704 3516 11756
rect 3568 11704 3574 11756
rect 3602 11704 3608 11756
rect 3660 11704 3666 11756
rect 4338 11704 4344 11756
rect 4396 11744 4402 11756
rect 4525 11747 4583 11753
rect 4525 11744 4537 11747
rect 4396 11716 4537 11744
rect 4396 11704 4402 11716
rect 4525 11713 4537 11716
rect 4571 11744 4583 11747
rect 4614 11744 4620 11756
rect 4571 11716 4620 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 4908 11753 4936 11852
rect 5077 11849 5089 11883
rect 5123 11880 5135 11883
rect 5350 11880 5356 11892
rect 5123 11852 5356 11880
rect 5123 11849 5135 11852
rect 5077 11843 5135 11849
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 6270 11840 6276 11892
rect 6328 11880 6334 11892
rect 6365 11883 6423 11889
rect 6365 11880 6377 11883
rect 6328 11852 6377 11880
rect 6328 11840 6334 11852
rect 6365 11849 6377 11852
rect 6411 11849 6423 11883
rect 6365 11843 6423 11849
rect 6730 11840 6736 11892
rect 6788 11840 6794 11892
rect 7190 11880 7196 11892
rect 6840 11852 7196 11880
rect 6748 11812 6776 11840
rect 6518 11784 6776 11812
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11744 4767 11747
rect 4893 11747 4951 11753
rect 4755 11716 4844 11744
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 4816 11688 4844 11716
rect 4893 11713 4905 11747
rect 4939 11744 4951 11747
rect 5442 11744 5448 11756
rect 4939 11716 5448 11744
rect 4939 11713 4951 11716
rect 4893 11707 4951 11713
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 6518 11753 6546 11784
rect 6503 11747 6561 11753
rect 6503 11713 6515 11747
rect 6549 11713 6561 11747
rect 6503 11707 6561 11713
rect 6641 11747 6699 11753
rect 6641 11713 6653 11747
rect 6687 11713 6699 11747
rect 6641 11707 6699 11713
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11744 6791 11747
rect 6840 11744 6868 11852
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 7282 11840 7288 11892
rect 7340 11880 7346 11892
rect 12526 11880 12532 11892
rect 7340 11852 12532 11880
rect 7340 11840 7346 11852
rect 12526 11840 12532 11852
rect 12584 11880 12590 11892
rect 14185 11883 14243 11889
rect 12584 11852 13584 11880
rect 12584 11840 12590 11852
rect 7374 11812 7380 11824
rect 6931 11784 7380 11812
rect 6931 11753 6959 11784
rect 7374 11772 7380 11784
rect 7432 11772 7438 11824
rect 8110 11772 8116 11824
rect 8168 11812 8174 11824
rect 13556 11821 13584 11852
rect 14185 11849 14197 11883
rect 14231 11880 14243 11883
rect 14366 11880 14372 11892
rect 14231 11852 14372 11880
rect 14231 11849 14243 11852
rect 14185 11843 14243 11849
rect 14366 11840 14372 11852
rect 14424 11840 14430 11892
rect 15378 11840 15384 11892
rect 15436 11880 15442 11892
rect 15841 11883 15899 11889
rect 15841 11880 15853 11883
rect 15436 11852 15853 11880
rect 15436 11840 15442 11852
rect 15841 11849 15853 11852
rect 15887 11849 15899 11883
rect 15841 11843 15899 11849
rect 10597 11815 10655 11821
rect 10597 11812 10609 11815
rect 8168 11784 10609 11812
rect 8168 11772 8174 11784
rect 10597 11781 10609 11784
rect 10643 11812 10655 11815
rect 13541 11815 13599 11821
rect 10643 11784 11284 11812
rect 10643 11781 10655 11784
rect 10597 11775 10655 11781
rect 6779 11716 6868 11744
rect 6916 11747 6974 11753
rect 6779 11713 6791 11716
rect 6733 11707 6791 11713
rect 6916 11713 6928 11747
rect 6962 11713 6974 11747
rect 6916 11707 6974 11713
rect 7002 11747 7060 11753
rect 7002 11713 7014 11747
rect 7048 11713 7060 11747
rect 7002 11707 7060 11713
rect 4798 11636 4804 11688
rect 4856 11636 4862 11688
rect 5902 11636 5908 11688
rect 5960 11676 5966 11688
rect 6656 11676 6684 11707
rect 5960 11648 6684 11676
rect 7024 11676 7052 11707
rect 7098 11704 7104 11756
rect 7156 11744 7162 11756
rect 7653 11747 7711 11753
rect 7653 11744 7665 11747
rect 7156 11716 7665 11744
rect 7156 11704 7162 11716
rect 7653 11713 7665 11716
rect 7699 11713 7711 11747
rect 7653 11707 7711 11713
rect 8662 11704 8668 11756
rect 8720 11704 8726 11756
rect 8849 11747 8907 11753
rect 8849 11713 8861 11747
rect 8895 11744 8907 11747
rect 8938 11744 8944 11756
rect 8895 11716 8944 11744
rect 8895 11713 8907 11716
rect 8849 11707 8907 11713
rect 8938 11704 8944 11716
rect 8996 11704 9002 11756
rect 9030 11704 9036 11756
rect 9088 11704 9094 11756
rect 10502 11704 10508 11756
rect 10560 11704 10566 11756
rect 10873 11747 10931 11753
rect 10873 11744 10885 11747
rect 10612 11716 10885 11744
rect 7282 11676 7288 11688
rect 7024 11648 7288 11676
rect 5960 11636 5966 11648
rect 4430 11568 4436 11620
rect 4488 11608 4494 11620
rect 4816 11608 4844 11636
rect 4488 11580 4844 11608
rect 6656 11608 6684 11648
rect 7282 11636 7288 11648
rect 7340 11676 7346 11688
rect 7340 11648 7788 11676
rect 7340 11636 7346 11648
rect 7466 11608 7472 11620
rect 6656 11580 7472 11608
rect 4488 11568 4494 11580
rect 7466 11568 7472 11580
rect 7524 11608 7530 11620
rect 7650 11608 7656 11620
rect 7524 11580 7656 11608
rect 7524 11568 7530 11580
rect 7650 11568 7656 11580
rect 7708 11568 7714 11620
rect 7760 11608 7788 11648
rect 8478 11636 8484 11688
rect 8536 11676 8542 11688
rect 9674 11676 9680 11688
rect 8536 11648 9680 11676
rect 8536 11636 8542 11648
rect 9674 11636 9680 11648
rect 9732 11636 9738 11688
rect 10318 11636 10324 11688
rect 10376 11676 10382 11688
rect 10612 11676 10640 11716
rect 10873 11713 10885 11716
rect 10919 11713 10931 11747
rect 11256 11744 11284 11784
rect 13541 11781 13553 11815
rect 13587 11781 13599 11815
rect 13541 11775 13599 11781
rect 14458 11772 14464 11824
rect 14516 11772 14522 11824
rect 12250 11744 12256 11756
rect 11256 11716 12256 11744
rect 10873 11707 10931 11713
rect 12250 11704 12256 11716
rect 12308 11704 12314 11756
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11713 13415 11747
rect 13357 11707 13415 11713
rect 10376 11648 10640 11676
rect 10376 11636 10382 11648
rect 9030 11608 9036 11620
rect 7760 11580 9036 11608
rect 9030 11568 9036 11580
rect 9088 11568 9094 11620
rect 2590 11500 2596 11552
rect 2648 11540 2654 11552
rect 5902 11540 5908 11552
rect 2648 11512 5908 11540
rect 2648 11500 2654 11512
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 5994 11500 6000 11552
rect 6052 11540 6058 11552
rect 10134 11540 10140 11552
rect 6052 11512 10140 11540
rect 6052 11500 6058 11512
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 10612 11540 10640 11648
rect 10781 11679 10839 11685
rect 10781 11645 10793 11679
rect 10827 11676 10839 11679
rect 10962 11676 10968 11688
rect 10827 11648 10968 11676
rect 10827 11645 10839 11648
rect 10781 11639 10839 11645
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 11514 11608 11520 11620
rect 10888 11580 11520 11608
rect 10686 11540 10692 11552
rect 10612 11512 10692 11540
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 10888 11549 10916 11580
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 13372 11608 13400 11707
rect 13722 11704 13728 11756
rect 13780 11744 13786 11756
rect 13817 11747 13875 11753
rect 13817 11744 13829 11747
rect 13780 11716 13829 11744
rect 13780 11704 13786 11716
rect 13817 11713 13829 11716
rect 13863 11713 13875 11747
rect 13817 11707 13875 11713
rect 14366 11704 14372 11756
rect 14424 11744 14430 11756
rect 14737 11747 14795 11753
rect 14737 11744 14749 11747
rect 14424 11716 14749 11744
rect 14424 11704 14430 11716
rect 14737 11713 14749 11716
rect 14783 11713 14795 11747
rect 14737 11707 14795 11713
rect 15010 11704 15016 11756
rect 15068 11704 15074 11756
rect 16485 11747 16543 11753
rect 16485 11713 16497 11747
rect 16531 11744 16543 11747
rect 16574 11744 16580 11756
rect 16531 11716 16580 11744
rect 16531 11713 16543 11716
rect 16485 11707 16543 11713
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 16758 11704 16764 11756
rect 16816 11744 16822 11756
rect 16853 11747 16911 11753
rect 16853 11744 16865 11747
rect 16816 11716 16865 11744
rect 16816 11704 16822 11716
rect 16853 11713 16865 11716
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 13909 11679 13967 11685
rect 13909 11676 13921 11679
rect 13504 11648 13921 11676
rect 13504 11636 13510 11648
rect 13909 11645 13921 11648
rect 13955 11645 13967 11679
rect 13909 11639 13967 11645
rect 14458 11636 14464 11688
rect 14516 11676 14522 11688
rect 14553 11679 14611 11685
rect 14553 11676 14565 11679
rect 14516 11648 14565 11676
rect 14516 11636 14522 11648
rect 14553 11645 14565 11648
rect 14599 11676 14611 11679
rect 15105 11679 15163 11685
rect 15105 11676 15117 11679
rect 14599 11648 15117 11676
rect 14599 11645 14611 11648
rect 14553 11639 14611 11645
rect 15105 11645 15117 11648
rect 15151 11645 15163 11679
rect 15105 11639 15163 11645
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 16669 11679 16727 11685
rect 16669 11676 16681 11679
rect 15344 11648 16681 11676
rect 15344 11636 15350 11648
rect 16669 11645 16681 11648
rect 16715 11645 16727 11679
rect 16669 11639 16727 11645
rect 14090 11608 14096 11620
rect 13372 11580 14096 11608
rect 14090 11568 14096 11580
rect 14148 11568 14154 11620
rect 10873 11543 10931 11549
rect 10873 11509 10885 11543
rect 10919 11509 10931 11543
rect 10873 11503 10931 11509
rect 11057 11543 11115 11549
rect 11057 11509 11069 11543
rect 11103 11540 11115 11543
rect 11330 11540 11336 11552
rect 11103 11512 11336 11540
rect 11103 11509 11115 11512
rect 11057 11503 11115 11509
rect 11330 11500 11336 11512
rect 11388 11500 11394 11552
rect 13722 11500 13728 11552
rect 13780 11500 13786 11552
rect 13814 11500 13820 11552
rect 13872 11500 13878 11552
rect 13998 11500 14004 11552
rect 14056 11540 14062 11552
rect 14461 11543 14519 11549
rect 14461 11540 14473 11543
rect 14056 11512 14473 11540
rect 14056 11500 14062 11512
rect 14461 11509 14473 11512
rect 14507 11509 14519 11543
rect 14461 11503 14519 11509
rect 14918 11500 14924 11552
rect 14976 11500 14982 11552
rect 15010 11500 15016 11552
rect 15068 11500 15074 11552
rect 15102 11500 15108 11552
rect 15160 11540 15166 11552
rect 15381 11543 15439 11549
rect 15381 11540 15393 11543
rect 15160 11512 15393 11540
rect 15160 11500 15166 11512
rect 15381 11509 15393 11512
rect 15427 11509 15439 11543
rect 15381 11503 15439 11509
rect 1104 11450 17388 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 17388 11450
rect 1104 11376 17388 11398
rect 3602 11296 3608 11348
rect 3660 11336 3666 11348
rect 7009 11339 7067 11345
rect 7009 11336 7021 11339
rect 3660 11308 7021 11336
rect 3660 11296 3666 11308
rect 7009 11305 7021 11308
rect 7055 11336 7067 11339
rect 7374 11336 7380 11348
rect 7055 11308 7380 11336
rect 7055 11305 7067 11308
rect 7009 11299 7067 11305
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 7650 11296 7656 11348
rect 7708 11336 7714 11348
rect 8110 11336 8116 11348
rect 7708 11308 8116 11336
rect 7708 11296 7714 11308
rect 8110 11296 8116 11308
rect 8168 11296 8174 11348
rect 8481 11339 8539 11345
rect 8481 11305 8493 11339
rect 8527 11336 8539 11339
rect 10318 11336 10324 11348
rect 8527 11308 10324 11336
rect 8527 11305 8539 11308
rect 8481 11299 8539 11305
rect 10318 11296 10324 11308
rect 10376 11296 10382 11348
rect 10502 11296 10508 11348
rect 10560 11336 10566 11348
rect 11517 11339 11575 11345
rect 11517 11336 11529 11339
rect 10560 11308 11529 11336
rect 10560 11296 10566 11308
rect 11517 11305 11529 11308
rect 11563 11336 11575 11339
rect 12437 11339 12495 11345
rect 11563 11308 11652 11336
rect 11563 11305 11575 11308
rect 11517 11299 11575 11305
rect 5997 11271 6055 11277
rect 5997 11237 6009 11271
rect 6043 11268 6055 11271
rect 6178 11268 6184 11280
rect 6043 11240 6184 11268
rect 6043 11237 6055 11240
rect 5997 11231 6055 11237
rect 6178 11228 6184 11240
rect 6236 11268 6242 11280
rect 6454 11268 6460 11280
rect 6236 11240 6460 11268
rect 6236 11228 6242 11240
rect 6454 11228 6460 11240
rect 6512 11228 6518 11280
rect 7282 11228 7288 11280
rect 7340 11228 7346 11280
rect 7392 11268 7420 11296
rect 7837 11271 7895 11277
rect 7392 11240 7793 11268
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 7300 11200 7328 11228
rect 7558 11200 7564 11212
rect 3936 11172 5120 11200
rect 3936 11160 3942 11172
rect 4522 11092 4528 11144
rect 4580 11132 4586 11144
rect 5092 11141 5120 11172
rect 5736 11172 7328 11200
rect 7392 11172 7564 11200
rect 4801 11135 4859 11141
rect 4801 11132 4813 11135
rect 4580 11104 4813 11132
rect 4580 11092 4586 11104
rect 4801 11101 4813 11104
rect 4847 11101 4859 11135
rect 4801 11095 4859 11101
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11101 5135 11135
rect 5077 11095 5135 11101
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11132 5227 11135
rect 5258 11132 5264 11144
rect 5215 11104 5264 11132
rect 5215 11101 5227 11104
rect 5169 11095 5227 11101
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11132 5503 11135
rect 5534 11132 5540 11144
rect 5491 11104 5540 11132
rect 5491 11101 5503 11104
rect 5445 11095 5503 11101
rect 5534 11092 5540 11104
rect 5592 11092 5598 11144
rect 5736 11141 5764 11172
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11101 5779 11135
rect 5721 11095 5779 11101
rect 5813 11135 5871 11141
rect 5813 11101 5825 11135
rect 5859 11132 5871 11135
rect 6270 11132 6276 11144
rect 5859 11104 6276 11132
rect 5859 11101 5871 11104
rect 5813 11095 5871 11101
rect 6270 11092 6276 11104
rect 6328 11132 6334 11144
rect 6730 11132 6736 11144
rect 6328 11104 6736 11132
rect 6328 11092 6334 11104
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 6914 11092 6920 11144
rect 6972 11132 6978 11144
rect 7101 11135 7159 11141
rect 7101 11132 7113 11135
rect 6972 11104 7113 11132
rect 6972 11092 6978 11104
rect 7101 11101 7113 11104
rect 7147 11101 7159 11135
rect 7101 11095 7159 11101
rect 7285 11135 7343 11141
rect 7285 11101 7297 11135
rect 7331 11132 7343 11135
rect 7392 11132 7420 11172
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 7331 11104 7420 11132
rect 7331 11101 7343 11104
rect 7285 11095 7343 11101
rect 7466 11092 7472 11144
rect 7524 11092 7530 11144
rect 7677 11135 7735 11141
rect 7677 11101 7689 11135
rect 7723 11132 7735 11135
rect 7765 11132 7793 11240
rect 7837 11237 7849 11271
rect 7883 11237 7895 11271
rect 7837 11231 7895 11237
rect 7852 11200 7880 11231
rect 8018 11228 8024 11280
rect 8076 11268 8082 11280
rect 8076 11240 8432 11268
rect 8076 11228 8082 11240
rect 7852 11172 8064 11200
rect 7723 11104 7793 11132
rect 7929 11135 7987 11141
rect 7723 11101 7735 11104
rect 7677 11095 7735 11101
rect 7929 11101 7941 11135
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 4614 11024 4620 11076
rect 4672 11064 4678 11076
rect 4985 11067 5043 11073
rect 4985 11064 4997 11067
rect 4672 11036 4997 11064
rect 4672 11024 4678 11036
rect 4985 11033 4997 11036
rect 5031 11033 5043 11067
rect 4985 11027 5043 11033
rect 5626 11024 5632 11076
rect 5684 11024 5690 11076
rect 7561 11067 7619 11073
rect 7561 11033 7573 11067
rect 7607 11064 7619 11067
rect 7834 11064 7840 11076
rect 7607 11036 7840 11064
rect 7607 11033 7619 11036
rect 7561 11027 7619 11033
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 5350 10956 5356 11008
rect 5408 10956 5414 11008
rect 7098 10956 7104 11008
rect 7156 10996 7162 11008
rect 7944 10996 7972 11095
rect 7156 10968 7972 10996
rect 8036 10996 8064 11172
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11132 8355 11135
rect 8404 11132 8432 11240
rect 9766 11160 9772 11212
rect 9824 11200 9830 11212
rect 10502 11200 10508 11212
rect 9824 11172 10508 11200
rect 9824 11160 9830 11172
rect 10502 11160 10508 11172
rect 10560 11160 10566 11212
rect 11624 11200 11652 11308
rect 12437 11305 12449 11339
rect 12483 11336 12495 11339
rect 12526 11336 12532 11348
rect 12483 11308 12532 11336
rect 12483 11305 12495 11308
rect 12437 11299 12495 11305
rect 12526 11296 12532 11308
rect 12584 11336 12590 11348
rect 12802 11336 12808 11348
rect 12584 11308 12808 11336
rect 12584 11296 12590 11308
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 12894 11296 12900 11348
rect 12952 11336 12958 11348
rect 13081 11339 13139 11345
rect 13081 11336 13093 11339
rect 12952 11308 13093 11336
rect 12952 11296 12958 11308
rect 13081 11305 13093 11308
rect 13127 11305 13139 11339
rect 13081 11299 13139 11305
rect 13449 11339 13507 11345
rect 13449 11305 13461 11339
rect 13495 11336 13507 11339
rect 13814 11336 13820 11348
rect 13495 11308 13820 11336
rect 13495 11305 13507 11308
rect 13449 11299 13507 11305
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 13998 11296 14004 11348
rect 14056 11336 14062 11348
rect 14093 11339 14151 11345
rect 14093 11336 14105 11339
rect 14056 11308 14105 11336
rect 14056 11296 14062 11308
rect 14093 11305 14105 11308
rect 14139 11305 14151 11339
rect 14093 11299 14151 11305
rect 14461 11339 14519 11345
rect 14461 11305 14473 11339
rect 14507 11336 14519 11339
rect 15010 11336 15016 11348
rect 14507 11308 15016 11336
rect 14507 11305 14519 11308
rect 14461 11299 14519 11305
rect 15010 11296 15016 11308
rect 15068 11296 15074 11348
rect 12066 11228 12072 11280
rect 12124 11268 12130 11280
rect 13170 11268 13176 11280
rect 12124 11240 13176 11268
rect 12124 11228 12130 11240
rect 13170 11228 13176 11240
rect 13228 11228 13234 11280
rect 15194 11200 15200 11212
rect 11624 11172 15200 11200
rect 15194 11160 15200 11172
rect 15252 11200 15258 11212
rect 15654 11200 15660 11212
rect 15252 11172 15660 11200
rect 15252 11160 15258 11172
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 8343 11104 8432 11132
rect 9493 11135 9551 11141
rect 8343 11101 8355 11104
rect 8297 11095 8355 11101
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 12894 11132 12900 11144
rect 9539 11104 12900 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 12894 11092 12900 11104
rect 12952 11092 12958 11144
rect 13078 11092 13084 11144
rect 13136 11092 13142 11144
rect 13170 11092 13176 11144
rect 13228 11092 13234 11144
rect 13722 11092 13728 11144
rect 13780 11132 13786 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13780 11104 14105 11132
rect 13780 11092 13786 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 14185 11135 14243 11141
rect 14185 11101 14197 11135
rect 14231 11101 14243 11135
rect 14185 11095 14243 11101
rect 8110 11024 8116 11076
rect 8168 11024 8174 11076
rect 8205 11067 8263 11073
rect 8205 11033 8217 11067
rect 8251 11064 8263 11067
rect 8846 11064 8852 11076
rect 8251 11036 8852 11064
rect 8251 11033 8263 11036
rect 8205 11027 8263 11033
rect 8846 11024 8852 11036
rect 8904 11024 8910 11076
rect 9125 11067 9183 11073
rect 9125 11033 9137 11067
rect 9171 11033 9183 11067
rect 9125 11027 9183 11033
rect 9309 11067 9367 11073
rect 9309 11033 9321 11067
rect 9355 11064 9367 11067
rect 9398 11064 9404 11076
rect 9355 11036 9404 11064
rect 9355 11033 9367 11036
rect 9309 11027 9367 11033
rect 8938 10996 8944 11008
rect 8036 10968 8944 10996
rect 7156 10956 7162 10968
rect 8938 10956 8944 10968
rect 8996 10996 9002 11008
rect 9140 10996 9168 11027
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 10229 11067 10287 11073
rect 10229 11033 10241 11067
rect 10275 11064 10287 11067
rect 10318 11064 10324 11076
rect 10275 11036 10324 11064
rect 10275 11033 10287 11036
rect 10229 11027 10287 11033
rect 10318 11024 10324 11036
rect 10376 11024 10382 11076
rect 10594 11024 10600 11076
rect 10652 11064 10658 11076
rect 10652 11036 12020 11064
rect 10652 11024 10658 11036
rect 8996 10968 9168 10996
rect 11992 10996 12020 11036
rect 12066 11024 12072 11076
rect 12124 11024 12130 11076
rect 12250 11024 12256 11076
rect 12308 11024 12314 11076
rect 13814 11064 13820 11076
rect 12360 11036 13820 11064
rect 12360 10996 12388 11036
rect 13814 11024 13820 11036
rect 13872 11064 13878 11076
rect 14200 11064 14228 11095
rect 14918 11092 14924 11144
rect 14976 11132 14982 11144
rect 15013 11135 15071 11141
rect 15013 11132 15025 11135
rect 14976 11104 15025 11132
rect 14976 11092 14982 11104
rect 15013 11101 15025 11104
rect 15059 11101 15071 11135
rect 15013 11095 15071 11101
rect 15286 11092 15292 11144
rect 15344 11092 15350 11144
rect 15378 11092 15384 11144
rect 15436 11092 15442 11144
rect 13872 11036 14228 11064
rect 13872 11024 13878 11036
rect 15102 11024 15108 11076
rect 15160 11064 15166 11076
rect 15197 11067 15255 11073
rect 15197 11064 15209 11067
rect 15160 11036 15209 11064
rect 15160 11024 15166 11036
rect 15197 11033 15209 11036
rect 15243 11033 15255 11067
rect 15902 11067 15960 11073
rect 15902 11064 15914 11067
rect 15197 11027 15255 11033
rect 15580 11036 15914 11064
rect 11992 10968 12388 10996
rect 15212 10996 15240 11027
rect 15286 10996 15292 11008
rect 15212 10968 15292 10996
rect 8996 10956 9002 10968
rect 15286 10956 15292 10968
rect 15344 10956 15350 11008
rect 15580 11005 15608 11036
rect 15902 11033 15914 11036
rect 15948 11033 15960 11067
rect 15902 11027 15960 11033
rect 15565 10999 15623 11005
rect 15565 10965 15577 10999
rect 15611 10965 15623 10999
rect 15565 10959 15623 10965
rect 16574 10956 16580 11008
rect 16632 10996 16638 11008
rect 17037 10999 17095 11005
rect 17037 10996 17049 10999
rect 16632 10968 17049 10996
rect 16632 10956 16638 10968
rect 17037 10965 17049 10968
rect 17083 10965 17095 10999
rect 17037 10959 17095 10965
rect 1104 10906 17388 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 17388 10906
rect 1104 10832 17388 10854
rect 3329 10795 3387 10801
rect 3329 10761 3341 10795
rect 3375 10792 3387 10795
rect 3375 10764 4292 10792
rect 3375 10761 3387 10764
rect 3329 10755 3387 10761
rect 2961 10727 3019 10733
rect 2961 10693 2973 10727
rect 3007 10724 3019 10727
rect 3605 10727 3663 10733
rect 3605 10724 3617 10727
rect 3007 10696 3617 10724
rect 3007 10693 3019 10696
rect 2961 10687 3019 10693
rect 3605 10693 3617 10696
rect 3651 10724 3663 10727
rect 3878 10724 3884 10736
rect 3651 10696 3884 10724
rect 3651 10693 3663 10696
rect 3605 10687 3663 10693
rect 3878 10684 3884 10696
rect 3936 10684 3942 10736
rect 4264 10733 4292 10764
rect 4522 10752 4528 10804
rect 4580 10792 4586 10804
rect 5074 10792 5080 10804
rect 4580 10764 5080 10792
rect 4580 10752 4586 10764
rect 5074 10752 5080 10764
rect 5132 10752 5138 10804
rect 5445 10795 5503 10801
rect 5445 10761 5457 10795
rect 5491 10792 5503 10795
rect 7377 10795 7435 10801
rect 5491 10764 7328 10792
rect 5491 10761 5503 10764
rect 5445 10755 5503 10761
rect 4249 10727 4307 10733
rect 4249 10693 4261 10727
rect 4295 10724 4307 10727
rect 5350 10724 5356 10736
rect 4295 10696 5356 10724
rect 4295 10693 4307 10696
rect 4249 10687 4307 10693
rect 5350 10684 5356 10696
rect 5408 10684 5414 10736
rect 5534 10684 5540 10736
rect 5592 10724 5598 10736
rect 7009 10727 7067 10733
rect 7009 10724 7021 10727
rect 5592 10696 7021 10724
rect 5592 10684 5598 10696
rect 7009 10693 7021 10696
rect 7055 10693 7067 10727
rect 7300 10724 7328 10764
rect 7377 10761 7389 10795
rect 7423 10792 7435 10795
rect 7466 10792 7472 10804
rect 7423 10764 7472 10792
rect 7423 10761 7435 10764
rect 7377 10755 7435 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 7576 10764 9674 10792
rect 7576 10724 7604 10764
rect 7300 10696 7604 10724
rect 7009 10687 7067 10693
rect 2777 10659 2835 10665
rect 2777 10625 2789 10659
rect 2823 10656 2835 10659
rect 2866 10656 2872 10668
rect 2823 10628 2872 10656
rect 2823 10625 2835 10628
rect 2777 10619 2835 10625
rect 2866 10616 2872 10628
rect 2924 10616 2930 10668
rect 3050 10616 3056 10668
rect 3108 10616 3114 10668
rect 3145 10659 3203 10665
rect 3145 10625 3157 10659
rect 3191 10625 3203 10659
rect 3145 10619 3203 10625
rect 3160 10588 3188 10619
rect 3418 10616 3424 10668
rect 3476 10616 3482 10668
rect 3510 10616 3516 10668
rect 3568 10656 3574 10668
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 3568 10628 3709 10656
rect 3568 10616 3574 10628
rect 3697 10625 3709 10628
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 3789 10659 3847 10665
rect 3789 10625 3801 10659
rect 3835 10656 3847 10659
rect 3970 10656 3976 10668
rect 3835 10628 3976 10656
rect 3835 10625 3847 10628
rect 3789 10619 3847 10625
rect 3804 10588 3832 10619
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 4065 10659 4123 10665
rect 4065 10625 4077 10659
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 3160 10560 3832 10588
rect 3973 10523 4031 10529
rect 3973 10489 3985 10523
rect 4019 10520 4031 10523
rect 4080 10520 4108 10619
rect 4430 10616 4436 10668
rect 4488 10616 4494 10668
rect 4706 10616 4712 10668
rect 4764 10656 4770 10668
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4764 10628 4905 10656
rect 4764 10616 4770 10628
rect 4893 10625 4905 10628
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10625 5135 10659
rect 5077 10619 5135 10625
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10625 5227 10659
rect 5169 10619 5227 10625
rect 5092 10588 5120 10619
rect 4908 10560 5120 10588
rect 5184 10588 5212 10619
rect 5258 10616 5264 10668
rect 5316 10616 5322 10668
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10656 6883 10659
rect 6914 10656 6920 10668
rect 6871 10628 6920 10656
rect 6871 10625 6883 10628
rect 6825 10619 6883 10625
rect 6840 10588 6868 10619
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 5184 10560 6868 10588
rect 7024 10588 7052 10687
rect 7650 10684 7656 10736
rect 7708 10724 7714 10736
rect 8110 10724 8116 10736
rect 7708 10696 8116 10724
rect 7708 10684 7714 10696
rect 8110 10684 8116 10696
rect 8168 10684 8174 10736
rect 8570 10684 8576 10736
rect 8628 10684 8634 10736
rect 7098 10616 7104 10668
rect 7156 10616 7162 10668
rect 7193 10659 7251 10665
rect 7193 10625 7205 10659
rect 7239 10656 7251 10659
rect 7282 10656 7288 10668
rect 7239 10628 7288 10656
rect 7239 10625 7251 10628
rect 7193 10619 7251 10625
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 7374 10616 7380 10668
rect 7432 10656 7438 10668
rect 7469 10659 7527 10665
rect 7469 10656 7481 10659
rect 7432 10628 7481 10656
rect 7432 10616 7438 10628
rect 7469 10625 7481 10628
rect 7515 10625 7527 10659
rect 7469 10619 7527 10625
rect 7742 10616 7748 10668
rect 7800 10616 7806 10668
rect 7883 10659 7941 10665
rect 7883 10625 7895 10659
rect 7929 10656 7941 10659
rect 8018 10656 8024 10668
rect 7929 10628 8024 10656
rect 7929 10625 7941 10628
rect 7883 10619 7941 10625
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 9646 10656 9674 10764
rect 10594 10752 10600 10804
rect 10652 10792 10658 10804
rect 10781 10795 10839 10801
rect 10781 10792 10793 10795
rect 10652 10764 10793 10792
rect 10652 10752 10658 10764
rect 10781 10761 10793 10764
rect 10827 10761 10839 10795
rect 10781 10755 10839 10761
rect 15378 10752 15384 10804
rect 15436 10792 15442 10804
rect 15841 10795 15899 10801
rect 15841 10792 15853 10795
rect 15436 10764 15853 10792
rect 15436 10752 15442 10764
rect 15841 10761 15853 10764
rect 15887 10761 15899 10795
rect 15841 10755 15899 10761
rect 16945 10795 17003 10801
rect 16945 10761 16957 10795
rect 16991 10792 17003 10795
rect 17218 10792 17224 10804
rect 16991 10764 17224 10792
rect 16991 10761 17003 10764
rect 16945 10755 17003 10761
rect 17218 10752 17224 10764
rect 17276 10752 17282 10804
rect 10134 10684 10140 10736
rect 10192 10724 10198 10736
rect 10192 10696 10548 10724
rect 10192 10684 10198 10696
rect 9766 10656 9772 10668
rect 9646 10628 9772 10656
rect 9766 10616 9772 10628
rect 9824 10656 9830 10668
rect 10520 10665 10548 10696
rect 12710 10684 12716 10736
rect 12768 10724 12774 10736
rect 13265 10727 13323 10733
rect 13265 10724 13277 10727
rect 12768 10696 13277 10724
rect 12768 10684 12774 10696
rect 13265 10693 13277 10696
rect 13311 10693 13323 10727
rect 13265 10687 13323 10693
rect 10413 10659 10471 10665
rect 10413 10656 10425 10659
rect 9824 10628 10425 10656
rect 9824 10616 9830 10628
rect 10413 10625 10425 10628
rect 10459 10625 10471 10659
rect 10413 10619 10471 10625
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10625 10563 10659
rect 10505 10619 10563 10625
rect 7650 10588 7656 10600
rect 7024 10560 7656 10588
rect 4614 10520 4620 10532
rect 4019 10492 4620 10520
rect 4019 10489 4031 10492
rect 3973 10483 4031 10489
rect 4614 10480 4620 10492
rect 4672 10480 4678 10532
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 4908 10452 4936 10560
rect 7650 10548 7656 10560
rect 7708 10548 7714 10600
rect 10318 10548 10324 10600
rect 10376 10548 10382 10600
rect 10520 10588 10548 10619
rect 10686 10616 10692 10668
rect 10744 10656 10750 10668
rect 10962 10656 10968 10668
rect 10744 10628 10968 10656
rect 10744 10616 10750 10628
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 11517 10659 11575 10665
rect 11517 10625 11529 10659
rect 11563 10656 11575 10659
rect 12066 10656 12072 10668
rect 11563 10628 12072 10656
rect 11563 10625 11575 10628
rect 11517 10619 11575 10625
rect 11609 10591 11667 10597
rect 11609 10588 11621 10591
rect 10520 10560 11621 10588
rect 11609 10557 11621 10560
rect 11655 10557 11667 10591
rect 11609 10551 11667 10557
rect 8110 10480 8116 10532
rect 8168 10520 8174 10532
rect 11716 10520 11744 10628
rect 12066 10616 12072 10628
rect 12124 10616 12130 10668
rect 13538 10656 13544 10668
rect 12406 10628 13544 10656
rect 12406 10588 12434 10628
rect 13538 10616 13544 10628
rect 13596 10616 13602 10668
rect 16485 10659 16543 10665
rect 16485 10625 16497 10659
rect 16531 10656 16543 10659
rect 16574 10656 16580 10668
rect 16531 10628 16580 10656
rect 16531 10625 16543 10628
rect 16485 10619 16543 10625
rect 16574 10616 16580 10628
rect 16632 10616 16638 10668
rect 16666 10616 16672 10668
rect 16724 10656 16730 10668
rect 16761 10659 16819 10665
rect 16761 10656 16773 10659
rect 16724 10628 16773 10656
rect 16724 10616 16730 10628
rect 16761 10625 16773 10628
rect 16807 10625 16819 10659
rect 16761 10619 16819 10625
rect 8168 10492 11744 10520
rect 11808 10560 12434 10588
rect 8168 10480 8174 10492
rect 3568 10424 4936 10452
rect 3568 10412 3574 10424
rect 5074 10412 5080 10464
rect 5132 10452 5138 10464
rect 5718 10452 5724 10464
rect 5132 10424 5724 10452
rect 5132 10412 5138 10424
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 8021 10455 8079 10461
rect 8021 10421 8033 10455
rect 8067 10452 8079 10455
rect 8662 10452 8668 10464
rect 8067 10424 8668 10452
rect 8067 10421 8079 10424
rect 8021 10415 8079 10421
rect 8662 10412 8668 10424
rect 8720 10452 8726 10464
rect 9306 10452 9312 10464
rect 8720 10424 9312 10452
rect 8720 10412 8726 10424
rect 9306 10412 9312 10424
rect 9364 10412 9370 10464
rect 10594 10412 10600 10464
rect 10652 10412 10658 10464
rect 10870 10412 10876 10464
rect 10928 10452 10934 10464
rect 11517 10455 11575 10461
rect 11517 10452 11529 10455
rect 10928 10424 11529 10452
rect 10928 10412 10934 10424
rect 11517 10421 11529 10424
rect 11563 10452 11575 10455
rect 11808 10452 11836 10560
rect 13170 10548 13176 10600
rect 13228 10588 13234 10600
rect 13449 10591 13507 10597
rect 13449 10588 13461 10591
rect 13228 10560 13461 10588
rect 13228 10548 13234 10560
rect 13449 10557 13461 10560
rect 13495 10588 13507 10591
rect 13722 10588 13728 10600
rect 13495 10560 13728 10588
rect 13495 10557 13507 10560
rect 13449 10551 13507 10557
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 11885 10523 11943 10529
rect 11885 10489 11897 10523
rect 11931 10520 11943 10523
rect 14274 10520 14280 10532
rect 11931 10492 14280 10520
rect 11931 10489 11943 10492
rect 11885 10483 11943 10489
rect 14274 10480 14280 10492
rect 14332 10480 14338 10532
rect 11563 10424 11836 10452
rect 11563 10421 11575 10424
rect 11517 10415 11575 10421
rect 12802 10412 12808 10464
rect 12860 10452 12866 10464
rect 13265 10455 13323 10461
rect 13265 10452 13277 10455
rect 12860 10424 13277 10452
rect 12860 10412 12866 10424
rect 13265 10421 13277 10424
rect 13311 10421 13323 10455
rect 13265 10415 13323 10421
rect 13725 10455 13783 10461
rect 13725 10421 13737 10455
rect 13771 10452 13783 10455
rect 14550 10452 14556 10464
rect 13771 10424 14556 10452
rect 13771 10421 13783 10424
rect 13725 10415 13783 10421
rect 14550 10412 14556 10424
rect 14608 10412 14614 10464
rect 1104 10362 17388 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 17388 10362
rect 1104 10288 17388 10310
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 3418 10248 3424 10260
rect 2823 10220 3424 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 4120 10220 5672 10248
rect 4120 10208 4126 10220
rect 4706 10180 4712 10192
rect 3804 10152 4712 10180
rect 2222 10004 2228 10056
rect 2280 10044 2286 10056
rect 3804 10053 3832 10152
rect 4706 10140 4712 10152
rect 4764 10140 4770 10192
rect 4982 10140 4988 10192
rect 5040 10140 5046 10192
rect 5442 10112 5448 10124
rect 4448 10084 5448 10112
rect 2593 10047 2651 10053
rect 2593 10044 2605 10047
rect 2280 10016 2605 10044
rect 2280 10004 2286 10016
rect 2593 10013 2605 10016
rect 2639 10013 2651 10047
rect 2593 10007 2651 10013
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 4154 10004 4160 10056
rect 4212 10004 4218 10056
rect 4448 10053 4476 10084
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 5644 10121 5672 10220
rect 5736 10220 6776 10248
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10081 5687 10115
rect 5629 10075 5687 10081
rect 4433 10047 4491 10053
rect 4433 10013 4445 10047
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10044 4859 10047
rect 5534 10044 5540 10056
rect 4847 10016 5540 10044
rect 4847 10013 4859 10016
rect 4801 10007 4859 10013
rect 2130 9936 2136 9988
rect 2188 9936 2194 9988
rect 2314 9936 2320 9988
rect 2372 9976 2378 9988
rect 2501 9979 2559 9985
rect 2501 9976 2513 9979
rect 2372 9948 2513 9976
rect 2372 9936 2378 9948
rect 2501 9945 2513 9948
rect 2547 9945 2559 9979
rect 2501 9939 2559 9945
rect 3970 9936 3976 9988
rect 4028 9936 4034 9988
rect 4065 9979 4123 9985
rect 4065 9945 4077 9979
rect 4111 9976 4123 9979
rect 4448 9976 4476 10007
rect 5534 10004 5540 10016
rect 5592 10044 5598 10056
rect 5736 10044 5764 10220
rect 5902 10140 5908 10192
rect 5960 10140 5966 10192
rect 6549 10183 6607 10189
rect 6549 10149 6561 10183
rect 6595 10180 6607 10183
rect 6638 10180 6644 10192
rect 6595 10152 6644 10180
rect 6595 10149 6607 10152
rect 6549 10143 6607 10149
rect 6638 10140 6644 10152
rect 6696 10140 6702 10192
rect 6748 10180 6776 10220
rect 7098 10208 7104 10260
rect 7156 10248 7162 10260
rect 8205 10251 8263 10257
rect 8205 10248 8217 10251
rect 7156 10220 8217 10248
rect 7156 10208 7162 10220
rect 8205 10217 8217 10220
rect 8251 10217 8263 10251
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 8205 10211 8263 10217
rect 8772 10220 8953 10248
rect 8772 10192 8800 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 8941 10211 8999 10217
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 10962 10248 10968 10260
rect 9548 10220 10968 10248
rect 9548 10208 9554 10220
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 11054 10208 11060 10260
rect 11112 10248 11118 10260
rect 11149 10251 11207 10257
rect 11149 10248 11161 10251
rect 11112 10220 11161 10248
rect 11112 10208 11118 10220
rect 11149 10217 11161 10220
rect 11195 10217 11207 10251
rect 11149 10211 11207 10217
rect 12253 10251 12311 10257
rect 12253 10217 12265 10251
rect 12299 10248 12311 10251
rect 12618 10248 12624 10260
rect 12299 10220 12624 10248
rect 12299 10217 12311 10220
rect 12253 10211 12311 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 13541 10251 13599 10257
rect 13541 10248 13553 10251
rect 13464 10220 13553 10248
rect 7561 10183 7619 10189
rect 6748 10152 7420 10180
rect 5920 10112 5948 10140
rect 5920 10084 6224 10112
rect 6196 10056 6224 10084
rect 6270 10072 6276 10124
rect 6328 10112 6334 10124
rect 7392 10112 7420 10152
rect 7561 10149 7573 10183
rect 7607 10180 7619 10183
rect 8662 10180 8668 10192
rect 7607 10152 8668 10180
rect 7607 10149 7619 10152
rect 7561 10143 7619 10149
rect 8662 10140 8668 10152
rect 8720 10140 8726 10192
rect 8754 10140 8760 10192
rect 8812 10140 8818 10192
rect 9401 10183 9459 10189
rect 9401 10149 9413 10183
rect 9447 10180 9459 10183
rect 13464 10180 13492 10220
rect 13541 10217 13553 10220
rect 13587 10217 13599 10251
rect 13541 10211 13599 10217
rect 13725 10251 13783 10257
rect 13725 10217 13737 10251
rect 13771 10248 13783 10251
rect 13906 10248 13912 10260
rect 13771 10220 13912 10248
rect 13771 10217 13783 10220
rect 13725 10211 13783 10217
rect 13906 10208 13912 10220
rect 13964 10208 13970 10260
rect 14274 10208 14280 10260
rect 14332 10248 14338 10260
rect 14553 10251 14611 10257
rect 14553 10248 14565 10251
rect 14332 10220 14565 10248
rect 14332 10208 14338 10220
rect 14553 10217 14565 10220
rect 14599 10217 14611 10251
rect 14553 10211 14611 10217
rect 16942 10208 16948 10260
rect 17000 10208 17006 10260
rect 9447 10152 10824 10180
rect 9447 10149 9459 10152
rect 9401 10143 9459 10149
rect 7653 10115 7711 10121
rect 7653 10112 7665 10115
rect 6328 10084 6408 10112
rect 7392 10084 7665 10112
rect 6328 10072 6334 10084
rect 5592 10016 5764 10044
rect 5592 10004 5598 10016
rect 5902 10004 5908 10056
rect 5960 10004 5966 10056
rect 5997 10047 6055 10053
rect 5997 10013 6009 10047
rect 6043 10013 6055 10047
rect 5997 10007 6055 10013
rect 4111 9948 4476 9976
rect 4617 9979 4675 9985
rect 4111 9945 4123 9948
rect 4065 9939 4123 9945
rect 4617 9945 4629 9979
rect 4663 9945 4675 9979
rect 4617 9939 4675 9945
rect 2409 9911 2467 9917
rect 2409 9877 2421 9911
rect 2455 9908 2467 9911
rect 2682 9908 2688 9920
rect 2455 9880 2688 9908
rect 2455 9877 2467 9880
rect 2409 9871 2467 9877
rect 2682 9868 2688 9880
rect 2740 9868 2746 9920
rect 4338 9868 4344 9920
rect 4396 9868 4402 9920
rect 4632 9908 4660 9939
rect 4706 9936 4712 9988
rect 4764 9976 4770 9988
rect 4764 9948 5028 9976
rect 4764 9936 4770 9948
rect 4798 9908 4804 9920
rect 4632 9880 4804 9908
rect 4798 9868 4804 9880
rect 4856 9868 4862 9920
rect 5000 9908 5028 9948
rect 5442 9936 5448 9988
rect 5500 9976 5506 9988
rect 6012 9976 6040 10007
rect 6178 10004 6184 10056
rect 6236 10004 6242 10056
rect 6380 10053 6408 10084
rect 7653 10081 7665 10084
rect 7699 10112 7711 10115
rect 9125 10115 9183 10121
rect 7699 10084 8340 10112
rect 7699 10081 7711 10084
rect 7653 10075 7711 10081
rect 8312 10056 8340 10084
rect 9125 10081 9137 10115
rect 9171 10112 9183 10115
rect 9490 10112 9496 10124
rect 9171 10084 9496 10112
rect 9171 10081 9183 10084
rect 9125 10075 9183 10081
rect 9490 10072 9496 10084
rect 9548 10112 9554 10124
rect 10686 10112 10692 10124
rect 9548 10084 10692 10112
rect 9548 10072 9554 10084
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 6365 10047 6423 10053
rect 6365 10013 6377 10047
rect 6411 10013 6423 10047
rect 6365 10007 6423 10013
rect 5500 9948 6040 9976
rect 6273 9979 6331 9985
rect 5500 9936 5506 9948
rect 6273 9945 6285 9979
rect 6319 9945 6331 9979
rect 6273 9939 6331 9945
rect 5902 9908 5908 9920
rect 5000 9880 5908 9908
rect 5902 9868 5908 9880
rect 5960 9908 5966 9920
rect 6288 9908 6316 9939
rect 5960 9880 6316 9908
rect 6380 9908 6408 10007
rect 6454 10004 6460 10056
rect 6512 10044 6518 10056
rect 6512 10016 6960 10044
rect 6512 10004 6518 10016
rect 6822 9936 6828 9988
rect 6880 9936 6886 9988
rect 6454 9908 6460 9920
rect 6380 9880 6460 9908
rect 5960 9868 5966 9880
rect 6454 9868 6460 9880
rect 6512 9868 6518 9920
rect 6730 9868 6736 9920
rect 6788 9868 6794 9920
rect 6932 9908 6960 10016
rect 7006 10004 7012 10056
rect 7064 10004 7070 10056
rect 7098 10004 7104 10056
rect 7156 10044 7162 10056
rect 7285 10047 7343 10053
rect 7285 10044 7297 10047
rect 7156 10016 7297 10044
rect 7156 10004 7162 10016
rect 7285 10013 7297 10016
rect 7331 10013 7343 10047
rect 7285 10007 7343 10013
rect 7374 10004 7380 10056
rect 7432 10004 7438 10056
rect 7466 10004 7472 10056
rect 7524 10044 7530 10056
rect 8021 10047 8079 10053
rect 8021 10044 8033 10047
rect 7524 10016 8033 10044
rect 7524 10004 7530 10016
rect 8021 10013 8033 10016
rect 8067 10013 8079 10047
rect 8021 10007 8079 10013
rect 8294 10004 8300 10056
rect 8352 10004 8358 10056
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10044 8447 10047
rect 8478 10044 8484 10056
rect 8435 10016 8484 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 9214 10004 9220 10056
rect 9272 10004 9278 10056
rect 9306 10004 9312 10056
rect 9364 10044 9370 10056
rect 9677 10047 9735 10053
rect 9677 10044 9689 10047
rect 9364 10016 9689 10044
rect 9364 10004 9370 10016
rect 9677 10013 9689 10016
rect 9723 10013 9735 10047
rect 10796 10044 10824 10152
rect 13188 10152 13492 10180
rect 10962 10072 10968 10124
rect 11020 10112 11026 10124
rect 12158 10112 12164 10124
rect 11020 10084 12164 10112
rect 11020 10072 11026 10084
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 12710 10072 12716 10124
rect 12768 10112 12774 10124
rect 13188 10112 13216 10152
rect 12768 10084 13216 10112
rect 12768 10072 12774 10084
rect 14642 10072 14648 10124
rect 14700 10072 14706 10124
rect 12069 10047 12127 10053
rect 12069 10044 12081 10047
rect 10796 10016 11100 10044
rect 9677 10007 9735 10013
rect 7190 9936 7196 9988
rect 7248 9936 7254 9988
rect 7837 9979 7895 9985
rect 7300 9948 7788 9976
rect 7300 9908 7328 9948
rect 6932 9880 7328 9908
rect 7760 9908 7788 9948
rect 7837 9945 7849 9979
rect 7883 9976 7895 9979
rect 8110 9976 8116 9988
rect 7883 9948 8116 9976
rect 7883 9945 7895 9948
rect 7837 9939 7895 9945
rect 8110 9936 8116 9948
rect 8168 9936 8174 9988
rect 8941 9979 8999 9985
rect 8941 9976 8953 9979
rect 8220 9948 8953 9976
rect 8220 9908 8248 9948
rect 8941 9945 8953 9948
rect 8987 9945 8999 9979
rect 9861 9979 9919 9985
rect 9861 9976 9873 9979
rect 8941 9939 8999 9945
rect 9692 9948 9873 9976
rect 9692 9920 9720 9948
rect 9861 9945 9873 9948
rect 9907 9976 9919 9979
rect 10962 9976 10968 9988
rect 9907 9948 10968 9976
rect 9907 9945 9919 9948
rect 9861 9939 9919 9945
rect 10962 9936 10968 9948
rect 11020 9936 11026 9988
rect 7760 9880 8248 9908
rect 8573 9911 8631 9917
rect 8573 9877 8585 9911
rect 8619 9908 8631 9911
rect 8846 9908 8852 9920
rect 8619 9880 8852 9908
rect 8619 9877 8631 9880
rect 8573 9871 8631 9877
rect 8846 9868 8852 9880
rect 8904 9868 8910 9920
rect 9674 9868 9680 9920
rect 9732 9868 9738 9920
rect 11072 9908 11100 10016
rect 11532 10016 12081 10044
rect 11532 9988 11560 10016
rect 12069 10013 12081 10016
rect 12115 10013 12127 10047
rect 12069 10007 12127 10013
rect 12802 10004 12808 10056
rect 12860 10004 12866 10056
rect 13446 10004 13452 10056
rect 13504 10004 13510 10056
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10044 13599 10047
rect 13630 10044 13636 10056
rect 13587 10016 13636 10044
rect 13587 10013 13599 10016
rect 13541 10007 13599 10013
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 14550 10004 14556 10056
rect 14608 10004 14614 10056
rect 16390 10004 16396 10056
rect 16448 10004 16454 10056
rect 16574 10004 16580 10056
rect 16632 10044 16638 10056
rect 16761 10047 16819 10053
rect 16761 10044 16773 10047
rect 16632 10016 16773 10044
rect 16632 10004 16638 10016
rect 16761 10013 16773 10016
rect 16807 10013 16819 10047
rect 16761 10007 16819 10013
rect 11146 9936 11152 9988
rect 11204 9976 11210 9988
rect 11333 9979 11391 9985
rect 11333 9976 11345 9979
rect 11204 9948 11345 9976
rect 11204 9936 11210 9948
rect 11333 9945 11345 9948
rect 11379 9945 11391 9979
rect 11333 9939 11391 9945
rect 11514 9936 11520 9988
rect 11572 9936 11578 9988
rect 11882 9936 11888 9988
rect 11940 9936 11946 9988
rect 12986 9936 12992 9988
rect 13044 9936 13050 9988
rect 13262 9936 13268 9988
rect 13320 9936 13326 9988
rect 13078 9908 13084 9920
rect 11072 9880 13084 9908
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 13173 9911 13231 9917
rect 13173 9877 13185 9911
rect 13219 9908 13231 9911
rect 14090 9908 14096 9920
rect 13219 9880 14096 9908
rect 13219 9877 13231 9880
rect 13173 9871 13231 9877
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 14921 9911 14979 9917
rect 14921 9877 14933 9911
rect 14967 9908 14979 9911
rect 15010 9908 15016 9920
rect 14967 9880 15016 9908
rect 14967 9877 14979 9880
rect 14921 9871 14979 9877
rect 15010 9868 15016 9880
rect 15068 9868 15074 9920
rect 16482 9868 16488 9920
rect 16540 9908 16546 9920
rect 16577 9911 16635 9917
rect 16577 9908 16589 9911
rect 16540 9880 16589 9908
rect 16540 9868 16546 9880
rect 16577 9877 16589 9880
rect 16623 9877 16635 9911
rect 16577 9871 16635 9877
rect 1104 9818 17388 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 17388 9818
rect 1104 9744 17388 9766
rect 2130 9664 2136 9716
rect 2188 9704 2194 9716
rect 2409 9707 2467 9713
rect 2409 9704 2421 9707
rect 2188 9676 2421 9704
rect 2188 9664 2194 9676
rect 2409 9673 2421 9676
rect 2455 9673 2467 9707
rect 2409 9667 2467 9673
rect 2869 9707 2927 9713
rect 2869 9673 2881 9707
rect 2915 9704 2927 9707
rect 3510 9704 3516 9716
rect 2915 9676 3516 9704
rect 2915 9673 2927 9676
rect 2869 9667 2927 9673
rect 3510 9664 3516 9676
rect 3568 9664 3574 9716
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 4396 9676 6408 9704
rect 4396 9664 4402 9676
rect 2222 9596 2228 9648
rect 2280 9636 2286 9648
rect 2501 9639 2559 9645
rect 2501 9636 2513 9639
rect 2280 9608 2513 9636
rect 2280 9596 2286 9608
rect 2501 9605 2513 9608
rect 2547 9605 2559 9639
rect 2501 9599 2559 9605
rect 5718 9596 5724 9648
rect 5776 9636 5782 9648
rect 6270 9636 6276 9648
rect 5776 9608 6276 9636
rect 5776 9596 5782 9608
rect 6270 9596 6276 9608
rect 6328 9596 6334 9648
rect 6380 9645 6408 9676
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 7374 9704 7380 9716
rect 7156 9676 7380 9704
rect 7156 9664 7162 9676
rect 7374 9664 7380 9676
rect 7432 9664 7438 9716
rect 7484 9676 8616 9704
rect 6365 9639 6423 9645
rect 6365 9605 6377 9639
rect 6411 9636 6423 9639
rect 7484 9636 7512 9676
rect 6411 9608 6465 9636
rect 6748 9608 7512 9636
rect 6411 9605 6423 9608
rect 6365 9599 6423 9605
rect 2314 9528 2320 9580
rect 2372 9528 2378 9580
rect 2682 9528 2688 9580
rect 2740 9568 2746 9580
rect 3053 9571 3111 9577
rect 3053 9568 3065 9571
rect 2740 9540 3065 9568
rect 2740 9528 2746 9540
rect 3053 9537 3065 9540
rect 3099 9537 3111 9571
rect 6380 9568 6408 9599
rect 6380 9540 6592 9568
rect 3053 9531 3111 9537
rect 6564 9512 6592 9540
rect 6638 9528 6644 9580
rect 6696 9558 6702 9580
rect 6748 9558 6776 9608
rect 7558 9596 7564 9648
rect 7616 9596 7622 9648
rect 7650 9596 7656 9648
rect 7708 9596 7714 9648
rect 8205 9639 8263 9645
rect 8205 9605 8217 9639
rect 8251 9605 8263 9639
rect 8205 9599 8263 9605
rect 6696 9530 6776 9558
rect 6696 9528 6702 9530
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9537 7803 9571
rect 7745 9531 7803 9537
rect 3970 9460 3976 9512
rect 4028 9500 4034 9512
rect 5445 9503 5503 9509
rect 5445 9500 5457 9503
rect 4028 9472 5457 9500
rect 4028 9460 4034 9472
rect 5445 9469 5457 9472
rect 5491 9469 5503 9503
rect 5445 9463 5503 9469
rect 5718 9460 5724 9512
rect 5776 9460 5782 9512
rect 6457 9503 6515 9509
rect 6457 9469 6469 9503
rect 6503 9469 6515 9503
rect 6457 9463 6515 9469
rect 4614 9392 4620 9444
rect 4672 9432 4678 9444
rect 6472 9432 6500 9463
rect 6546 9460 6552 9512
rect 6604 9460 6610 9512
rect 6914 9460 6920 9512
rect 6972 9500 6978 9512
rect 7760 9500 7788 9531
rect 7926 9528 7932 9580
rect 7984 9568 7990 9580
rect 8021 9571 8079 9577
rect 8021 9568 8033 9571
rect 7984 9540 8033 9568
rect 7984 9528 7990 9540
rect 8021 9537 8033 9540
rect 8067 9537 8079 9571
rect 8021 9531 8079 9537
rect 8220 9500 8248 9599
rect 8294 9596 8300 9648
rect 8352 9596 8358 9648
rect 8588 9636 8616 9676
rect 8662 9664 8668 9716
rect 8720 9704 8726 9716
rect 12986 9704 12992 9716
rect 8720 9676 12992 9704
rect 8720 9664 8726 9676
rect 9214 9636 9220 9648
rect 8588 9608 9220 9636
rect 9214 9596 9220 9608
rect 9272 9596 9278 9648
rect 9585 9639 9643 9645
rect 9585 9605 9597 9639
rect 9631 9636 9643 9639
rect 9861 9639 9919 9645
rect 9861 9636 9873 9639
rect 9631 9608 9873 9636
rect 9631 9605 9643 9608
rect 9585 9599 9643 9605
rect 9861 9605 9873 9608
rect 9907 9636 9919 9639
rect 10410 9636 10416 9648
rect 9907 9608 10416 9636
rect 9907 9605 9919 9608
rect 9861 9599 9919 9605
rect 10410 9596 10416 9608
rect 10468 9596 10474 9648
rect 10962 9596 10968 9648
rect 11020 9596 11026 9648
rect 11716 9645 11744 9676
rect 12986 9664 12992 9676
rect 13044 9664 13050 9716
rect 11701 9639 11759 9645
rect 11701 9605 11713 9639
rect 11747 9605 11759 9639
rect 11701 9599 11759 9605
rect 12802 9596 12808 9648
rect 12860 9636 12866 9648
rect 13262 9636 13268 9648
rect 12860 9608 13268 9636
rect 12860 9596 12866 9608
rect 13262 9596 13268 9608
rect 13320 9636 13326 9648
rect 13817 9639 13875 9645
rect 13817 9636 13829 9639
rect 13320 9608 13829 9636
rect 13320 9596 13326 9608
rect 13817 9605 13829 9608
rect 13863 9605 13875 9639
rect 13817 9599 13875 9605
rect 8386 9528 8392 9580
rect 8444 9528 8450 9580
rect 8665 9571 8723 9577
rect 8665 9537 8677 9571
rect 8711 9568 8723 9571
rect 8846 9568 8852 9580
rect 8711 9540 8852 9568
rect 8711 9537 8723 9540
rect 8665 9531 8723 9537
rect 6972 9472 7144 9500
rect 6972 9460 6978 9472
rect 4672 9404 6500 9432
rect 6825 9435 6883 9441
rect 4672 9392 4678 9404
rect 5368 9376 5396 9404
rect 6825 9401 6837 9435
rect 6871 9432 6883 9435
rect 7006 9432 7012 9444
rect 6871 9404 7012 9432
rect 6871 9401 6883 9404
rect 6825 9395 6883 9401
rect 7006 9392 7012 9404
rect 7064 9392 7070 9444
rect 7116 9432 7144 9472
rect 7668 9472 7788 9500
rect 7820 9472 8248 9500
rect 7668 9432 7696 9472
rect 7116 9404 7696 9432
rect 5350 9324 5356 9376
rect 5408 9324 5414 9376
rect 6638 9324 6644 9376
rect 6696 9324 6702 9376
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 7820 9364 7848 9472
rect 8680 9432 8708 9531
rect 8846 9528 8852 9540
rect 8904 9528 8910 9580
rect 8938 9528 8944 9580
rect 8996 9528 9002 9580
rect 9122 9528 9128 9580
rect 9180 9528 9186 9580
rect 9401 9571 9459 9577
rect 9401 9568 9413 9571
rect 9232 9540 9413 9568
rect 8757 9503 8815 9509
rect 8757 9469 8769 9503
rect 8803 9500 8815 9503
rect 8803 9472 8984 9500
rect 8803 9469 8815 9472
rect 8757 9463 8815 9469
rect 8496 9404 8708 9432
rect 6788 9336 7848 9364
rect 7929 9367 7987 9373
rect 6788 9324 6794 9336
rect 7929 9333 7941 9367
rect 7975 9364 7987 9367
rect 8496 9364 8524 9404
rect 7975 9336 8524 9364
rect 7975 9333 7987 9336
rect 7929 9327 7987 9333
rect 8570 9324 8576 9376
rect 8628 9324 8634 9376
rect 8662 9324 8668 9376
rect 8720 9324 8726 9376
rect 8956 9364 8984 9472
rect 9140 9441 9168 9528
rect 9232 9512 9260 9540
rect 9401 9537 9413 9540
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 10134 9528 10140 9580
rect 10192 9528 10198 9580
rect 10873 9571 10931 9577
rect 10873 9568 10885 9571
rect 10336 9540 10885 9568
rect 9214 9460 9220 9512
rect 9272 9460 9278 9512
rect 9950 9460 9956 9512
rect 10008 9460 10014 9512
rect 9125 9435 9183 9441
rect 9125 9401 9137 9435
rect 9171 9401 9183 9435
rect 9125 9395 9183 9401
rect 9306 9392 9312 9444
rect 9364 9432 9370 9444
rect 10226 9432 10232 9444
rect 9364 9404 10232 9432
rect 9364 9392 9370 9404
rect 10226 9392 10232 9404
rect 10284 9392 10290 9444
rect 10336 9441 10364 9540
rect 10873 9537 10885 9540
rect 10919 9537 10931 9571
rect 10980 9568 11008 9596
rect 11885 9571 11943 9577
rect 11885 9568 11897 9571
rect 10980 9540 11897 9568
rect 10873 9531 10931 9537
rect 11885 9537 11897 9540
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 13170 9528 13176 9580
rect 13228 9568 13234 9580
rect 13633 9571 13691 9577
rect 13633 9568 13645 9571
rect 13228 9540 13645 9568
rect 13228 9528 13234 9540
rect 13633 9537 13645 9540
rect 13679 9537 13691 9571
rect 13633 9531 13691 9537
rect 13906 9528 13912 9580
rect 13964 9568 13970 9580
rect 14553 9571 14611 9577
rect 14553 9568 14565 9571
rect 13964 9540 14565 9568
rect 13964 9528 13970 9540
rect 14553 9537 14565 9540
rect 14599 9537 14611 9571
rect 14553 9531 14611 9537
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9568 15163 9571
rect 15194 9568 15200 9580
rect 15151 9540 15200 9568
rect 15151 9537 15163 9540
rect 15105 9531 15163 9537
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 15372 9571 15430 9577
rect 15372 9537 15384 9571
rect 15418 9568 15430 9571
rect 16114 9568 16120 9580
rect 15418 9540 16120 9568
rect 15418 9537 15430 9540
rect 15372 9531 15430 9537
rect 16114 9528 16120 9540
rect 16172 9528 16178 9580
rect 10778 9460 10784 9512
rect 10836 9500 10842 9512
rect 10965 9503 11023 9509
rect 10965 9500 10977 9503
rect 10836 9472 10977 9500
rect 10836 9460 10842 9472
rect 10965 9469 10977 9472
rect 11011 9469 11023 9503
rect 10965 9463 11023 9469
rect 11146 9460 11152 9512
rect 11204 9500 11210 9512
rect 14182 9500 14188 9512
rect 11204 9472 14188 9500
rect 11204 9460 11210 9472
rect 14182 9460 14188 9472
rect 14240 9460 14246 9512
rect 14642 9460 14648 9512
rect 14700 9460 14706 9512
rect 10321 9435 10379 9441
rect 10321 9401 10333 9435
rect 10367 9401 10379 9435
rect 10321 9395 10379 9401
rect 11238 9392 11244 9444
rect 11296 9392 11302 9444
rect 9324 9364 9352 9392
rect 8956 9336 9352 9364
rect 9766 9324 9772 9376
rect 9824 9364 9830 9376
rect 9861 9367 9919 9373
rect 9861 9364 9873 9367
rect 9824 9336 9873 9364
rect 9824 9324 9830 9336
rect 9861 9333 9873 9336
rect 9907 9333 9919 9367
rect 9861 9327 9919 9333
rect 10134 9324 10140 9376
rect 10192 9364 10198 9376
rect 10870 9364 10876 9376
rect 10192 9336 10876 9364
rect 10192 9324 10198 9336
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 11057 9367 11115 9373
rect 11057 9333 11069 9367
rect 11103 9364 11115 9367
rect 11422 9364 11428 9376
rect 11103 9336 11428 9364
rect 11103 9333 11115 9336
rect 11057 9327 11115 9333
rect 11422 9324 11428 9336
rect 11480 9364 11486 9376
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 11480 9336 11529 9364
rect 11480 9324 11486 9336
rect 11517 9333 11529 9336
rect 11563 9333 11575 9367
rect 11517 9327 11575 9333
rect 14001 9367 14059 9373
rect 14001 9333 14013 9367
rect 14047 9364 14059 9367
rect 14734 9364 14740 9376
rect 14047 9336 14740 9364
rect 14047 9333 14059 9336
rect 14001 9327 14059 9333
rect 14734 9324 14740 9336
rect 14792 9324 14798 9376
rect 14918 9324 14924 9376
rect 14976 9324 14982 9376
rect 16482 9324 16488 9376
rect 16540 9324 16546 9376
rect 1104 9274 17388 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 17388 9274
rect 1104 9200 17388 9222
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9160 5503 9163
rect 6178 9160 6184 9172
rect 5491 9132 6184 9160
rect 5491 9129 5503 9132
rect 5445 9123 5503 9129
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 6362 9120 6368 9172
rect 6420 9160 6426 9172
rect 6638 9160 6644 9172
rect 6420 9132 6644 9160
rect 6420 9120 6426 9132
rect 6638 9120 6644 9132
rect 6696 9160 6702 9172
rect 8297 9163 8355 9169
rect 8297 9160 8309 9163
rect 6696 9132 8309 9160
rect 6696 9120 6702 9132
rect 8297 9129 8309 9132
rect 8343 9160 8355 9163
rect 8754 9160 8760 9172
rect 8343 9132 8760 9160
rect 8343 9129 8355 9132
rect 8297 9123 8355 9129
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 9030 9120 9036 9172
rect 9088 9160 9094 9172
rect 9214 9160 9220 9172
rect 9088 9132 9220 9160
rect 9088 9120 9094 9132
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 13170 9160 13176 9172
rect 9646 9132 13176 9160
rect 3053 9095 3111 9101
rect 3053 9061 3065 9095
rect 3099 9092 3111 9095
rect 3970 9092 3976 9104
rect 3099 9064 3976 9092
rect 3099 9061 3111 9064
rect 3053 9055 3111 9061
rect 2682 8984 2688 9036
rect 2740 9024 2746 9036
rect 2961 9027 3019 9033
rect 2961 9024 2973 9027
rect 2740 8996 2973 9024
rect 2740 8984 2746 8996
rect 2961 8993 2973 8996
rect 3007 8993 3019 9027
rect 2961 8987 3019 8993
rect 2222 8916 2228 8968
rect 2280 8956 2286 8968
rect 3068 8956 3096 9055
rect 3970 9052 3976 9064
rect 4028 9052 4034 9104
rect 4433 9095 4491 9101
rect 4433 9061 4445 9095
rect 4479 9092 4491 9095
rect 7101 9095 7159 9101
rect 4479 9064 6868 9092
rect 4479 9061 4491 9064
rect 4433 9055 4491 9061
rect 3602 8984 3608 9036
rect 3660 9024 3666 9036
rect 4065 9027 4123 9033
rect 4065 9024 4077 9027
rect 3660 8996 4077 9024
rect 3660 8984 3666 8996
rect 4065 8993 4077 8996
rect 4111 8993 4123 9027
rect 5442 9024 5448 9036
rect 4065 8987 4123 8993
rect 4908 8996 5448 9024
rect 2280 8928 3096 8956
rect 2280 8916 2286 8928
rect 3234 8916 3240 8968
rect 3292 8916 3298 8968
rect 3326 8916 3332 8968
rect 3384 8916 3390 8968
rect 3418 8916 3424 8968
rect 3476 8956 3482 8968
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 3476 8928 3801 8956
rect 3476 8916 3482 8928
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 4798 8916 4804 8968
rect 4856 8956 4862 8968
rect 4908 8965 4936 8996
rect 5442 8984 5448 8996
rect 5500 9024 5506 9036
rect 5500 8996 5764 9024
rect 5500 8984 5506 8996
rect 4893 8959 4951 8965
rect 4893 8956 4905 8959
rect 4856 8928 4905 8956
rect 4856 8916 4862 8928
rect 4893 8925 4905 8928
rect 4939 8925 4951 8959
rect 4893 8919 4951 8925
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8925 5319 8959
rect 5261 8919 5319 8925
rect 5537 8959 5595 8965
rect 5537 8925 5549 8959
rect 5583 8956 5595 8959
rect 5626 8956 5632 8968
rect 5583 8928 5632 8956
rect 5583 8925 5595 8928
rect 5537 8919 5595 8925
rect 2130 8848 2136 8900
rect 2188 8888 2194 8900
rect 2317 8891 2375 8897
rect 2317 8888 2329 8891
rect 2188 8860 2329 8888
rect 2188 8848 2194 8860
rect 2317 8857 2329 8860
rect 2363 8857 2375 8891
rect 2317 8851 2375 8857
rect 2406 8848 2412 8900
rect 2464 8888 2470 8900
rect 2464 8860 3556 8888
rect 2464 8848 2470 8860
rect 2777 8823 2835 8829
rect 2777 8789 2789 8823
rect 2823 8820 2835 8823
rect 3050 8820 3056 8832
rect 2823 8792 3056 8820
rect 2823 8789 2835 8792
rect 2777 8783 2835 8789
rect 3050 8780 3056 8792
rect 3108 8780 3114 8832
rect 3528 8829 3556 8860
rect 3694 8848 3700 8900
rect 3752 8888 3758 8900
rect 4249 8891 4307 8897
rect 4249 8888 4261 8891
rect 3752 8860 4261 8888
rect 3752 8848 3758 8860
rect 4249 8857 4261 8860
rect 4295 8857 4307 8891
rect 4249 8851 4307 8857
rect 4614 8848 4620 8900
rect 4672 8888 4678 8900
rect 5077 8891 5135 8897
rect 5077 8888 5089 8891
rect 4672 8860 5089 8888
rect 4672 8848 4678 8860
rect 5077 8857 5089 8860
rect 5123 8857 5135 8891
rect 5077 8851 5135 8857
rect 5169 8891 5227 8897
rect 5169 8857 5181 8891
rect 5215 8857 5227 8891
rect 5276 8888 5304 8919
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 5736 8965 5764 8996
rect 5810 8984 5816 9036
rect 5868 9024 5874 9036
rect 6840 9024 6868 9064
rect 7101 9061 7113 9095
rect 7147 9092 7159 9095
rect 8938 9092 8944 9104
rect 7147 9064 8944 9092
rect 7147 9061 7159 9064
rect 7101 9055 7159 9061
rect 8938 9052 8944 9064
rect 8996 9052 9002 9104
rect 8018 9024 8024 9036
rect 5868 8996 6408 9024
rect 6840 8996 6960 9024
rect 5868 8984 5874 8996
rect 5721 8959 5779 8965
rect 5721 8925 5733 8959
rect 5767 8925 5779 8959
rect 5721 8919 5779 8925
rect 5902 8916 5908 8968
rect 5960 8916 5966 8968
rect 6270 8956 6276 8968
rect 6012 8928 6276 8956
rect 5442 8888 5448 8900
rect 5276 8860 5448 8888
rect 5169 8851 5227 8857
rect 3513 8823 3571 8829
rect 3513 8789 3525 8823
rect 3559 8820 3571 8823
rect 3878 8820 3884 8832
rect 3559 8792 3884 8820
rect 3559 8789 3571 8792
rect 3513 8783 3571 8789
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 4154 8780 4160 8832
rect 4212 8780 4218 8832
rect 5184 8820 5212 8851
rect 5442 8848 5448 8860
rect 5500 8848 5506 8900
rect 5813 8891 5871 8897
rect 5813 8857 5825 8891
rect 5859 8888 5871 8891
rect 6012 8888 6040 8928
rect 6270 8916 6276 8928
rect 6328 8916 6334 8968
rect 6380 8888 6408 8996
rect 6546 8916 6552 8968
rect 6604 8916 6610 8968
rect 6638 8916 6644 8968
rect 6696 8956 6702 8968
rect 6932 8965 6960 8996
rect 7852 8996 8024 9024
rect 6825 8959 6883 8965
rect 6825 8956 6837 8959
rect 6696 8928 6837 8956
rect 6696 8916 6702 8928
rect 6825 8925 6837 8928
rect 6871 8925 6883 8959
rect 6825 8919 6883 8925
rect 6917 8959 6975 8965
rect 6917 8925 6929 8959
rect 6963 8956 6975 8959
rect 7374 8956 7380 8968
rect 6963 8928 7380 8956
rect 6963 8925 6975 8928
rect 6917 8919 6975 8925
rect 7374 8916 7380 8928
rect 7432 8956 7438 8968
rect 7469 8959 7527 8965
rect 7469 8956 7481 8959
rect 7432 8928 7481 8956
rect 7432 8916 7438 8928
rect 7469 8925 7481 8928
rect 7515 8925 7527 8959
rect 7469 8919 7527 8925
rect 7558 8916 7564 8968
rect 7616 8956 7622 8968
rect 7852 8965 7880 8996
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 8294 8984 8300 9036
rect 8352 8984 8358 9036
rect 8386 8984 8392 9036
rect 8444 9024 8450 9036
rect 9646 9024 9674 9132
rect 13170 9120 13176 9132
rect 13228 9120 13234 9172
rect 13354 9120 13360 9172
rect 13412 9120 13418 9172
rect 13725 9163 13783 9169
rect 13725 9129 13737 9163
rect 13771 9160 13783 9163
rect 13906 9160 13912 9172
rect 13771 9132 13912 9160
rect 13771 9129 13783 9132
rect 13725 9123 13783 9129
rect 13906 9120 13912 9132
rect 13964 9120 13970 9172
rect 14090 9120 14096 9172
rect 14148 9120 14154 9172
rect 14553 9163 14611 9169
rect 14553 9129 14565 9163
rect 14599 9160 14611 9163
rect 14642 9160 14648 9172
rect 14599 9132 14648 9160
rect 14599 9129 14611 9132
rect 14553 9123 14611 9129
rect 14642 9120 14648 9132
rect 14700 9120 14706 9172
rect 16114 9120 16120 9172
rect 16172 9120 16178 9172
rect 11238 9052 11244 9104
rect 11296 9092 11302 9104
rect 11790 9092 11796 9104
rect 11296 9064 11796 9092
rect 11296 9052 11302 9064
rect 11790 9052 11796 9064
rect 11848 9052 11854 9104
rect 13262 9052 13268 9104
rect 13320 9092 13326 9104
rect 13538 9092 13544 9104
rect 13320 9064 13544 9092
rect 13320 9052 13326 9064
rect 13538 9052 13544 9064
rect 13596 9052 13602 9104
rect 8444 8996 9674 9024
rect 8444 8984 8450 8996
rect 9766 8984 9772 9036
rect 9824 9024 9830 9036
rect 10410 9024 10416 9036
rect 9824 8996 10416 9024
rect 9824 8984 9830 8996
rect 10410 8984 10416 8996
rect 10468 8984 10474 9036
rect 10686 8984 10692 9036
rect 10744 9024 10750 9036
rect 13357 9027 13415 9033
rect 13357 9024 13369 9027
rect 10744 8996 13369 9024
rect 10744 8984 10750 8996
rect 13357 8993 13369 8996
rect 13403 8993 13415 9027
rect 13357 8987 13415 8993
rect 14182 8984 14188 9036
rect 14240 8984 14246 9036
rect 15746 8984 15752 9036
rect 15804 9024 15810 9036
rect 15804 8996 15884 9024
rect 15804 8984 15810 8996
rect 7745 8959 7803 8965
rect 7745 8956 7757 8959
rect 7616 8928 7757 8956
rect 7616 8916 7622 8928
rect 7745 8925 7757 8928
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 7837 8959 7895 8965
rect 7837 8925 7849 8959
rect 7883 8925 7895 8959
rect 8478 8956 8484 8968
rect 7837 8919 7895 8925
rect 7944 8928 8484 8956
rect 5859 8860 6040 8888
rect 6104 8860 6408 8888
rect 5859 8857 5871 8860
rect 5813 8851 5871 8857
rect 5902 8820 5908 8832
rect 5184 8792 5908 8820
rect 5902 8780 5908 8792
rect 5960 8780 5966 8832
rect 6104 8829 6132 8860
rect 6730 8848 6736 8900
rect 6788 8848 6794 8900
rect 7282 8848 7288 8900
rect 7340 8888 7346 8900
rect 7650 8888 7656 8900
rect 7340 8860 7656 8888
rect 7340 8848 7346 8860
rect 7650 8848 7656 8860
rect 7708 8848 7714 8900
rect 6089 8823 6147 8829
rect 6089 8789 6101 8823
rect 6135 8789 6147 8823
rect 6089 8783 6147 8789
rect 6178 8780 6184 8832
rect 6236 8820 6242 8832
rect 7944 8820 7972 8928
rect 8478 8916 8484 8928
rect 8536 8916 8542 8968
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 11241 8959 11299 8965
rect 11241 8956 11253 8959
rect 8628 8928 11253 8956
rect 8628 8916 8634 8928
rect 11241 8925 11253 8928
rect 11287 8956 11299 8959
rect 11514 8956 11520 8968
rect 11287 8928 11520 8956
rect 11287 8925 11299 8928
rect 11241 8919 11299 8925
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 12526 8916 12532 8968
rect 12584 8956 12590 8968
rect 12584 8928 13400 8956
rect 12584 8916 12590 8928
rect 8205 8891 8263 8897
rect 8205 8857 8217 8891
rect 8251 8888 8263 8891
rect 8251 8860 8616 8888
rect 8251 8857 8263 8860
rect 8205 8851 8263 8857
rect 8588 8832 8616 8860
rect 8846 8848 8852 8900
rect 8904 8888 8910 8900
rect 9582 8888 9588 8900
rect 8904 8860 9588 8888
rect 8904 8848 8910 8860
rect 9582 8848 9588 8860
rect 9640 8888 9646 8900
rect 11057 8891 11115 8897
rect 11057 8888 11069 8891
rect 9640 8860 11069 8888
rect 9640 8848 9646 8860
rect 11057 8857 11069 8860
rect 11103 8857 11115 8891
rect 11057 8851 11115 8857
rect 12986 8848 12992 8900
rect 13044 8888 13050 8900
rect 13265 8891 13323 8897
rect 13265 8888 13277 8891
rect 13044 8860 13277 8888
rect 13044 8848 13050 8860
rect 13265 8857 13277 8860
rect 13311 8857 13323 8891
rect 13372 8888 13400 8928
rect 13538 8916 13544 8968
rect 13596 8916 13602 8968
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13688 8928 14105 8956
rect 13688 8916 13694 8928
rect 14093 8925 14105 8928
rect 14139 8925 14151 8959
rect 14093 8919 14151 8925
rect 14369 8959 14427 8965
rect 14369 8925 14381 8959
rect 14415 8956 14427 8959
rect 14550 8956 14556 8968
rect 14415 8928 14556 8956
rect 14415 8925 14427 8928
rect 14369 8919 14427 8925
rect 14550 8916 14556 8928
rect 14608 8916 14614 8968
rect 14918 8916 14924 8968
rect 14976 8956 14982 8968
rect 15856 8965 15884 8996
rect 16482 8984 16488 9036
rect 16540 9024 16546 9036
rect 16853 9027 16911 9033
rect 16853 9024 16865 9027
rect 16540 8996 16865 9024
rect 16540 8984 16546 8996
rect 16853 8993 16865 8996
rect 16899 8993 16911 9027
rect 16853 8987 16911 8993
rect 15565 8959 15623 8965
rect 15565 8956 15577 8959
rect 14976 8928 15577 8956
rect 14976 8916 14982 8928
rect 15565 8925 15577 8928
rect 15611 8925 15623 8959
rect 15565 8919 15623 8925
rect 15841 8959 15899 8965
rect 15841 8925 15853 8959
rect 15887 8925 15899 8959
rect 15841 8919 15899 8925
rect 15933 8959 15991 8965
rect 15933 8925 15945 8959
rect 15979 8956 15991 8959
rect 16301 8959 16359 8965
rect 16301 8956 16313 8959
rect 15979 8928 16313 8956
rect 15979 8925 15991 8928
rect 15933 8919 15991 8925
rect 16301 8925 16313 8928
rect 16347 8925 16359 8959
rect 16301 8919 16359 8925
rect 14182 8888 14188 8900
rect 13372 8860 14188 8888
rect 13265 8851 13323 8857
rect 14182 8848 14188 8860
rect 14240 8848 14246 8900
rect 15286 8848 15292 8900
rect 15344 8888 15350 8900
rect 15749 8891 15807 8897
rect 15749 8888 15761 8891
rect 15344 8860 15761 8888
rect 15344 8848 15350 8860
rect 15749 8857 15761 8860
rect 15795 8857 15807 8891
rect 15749 8851 15807 8857
rect 6236 8792 7972 8820
rect 8021 8823 8079 8829
rect 6236 8780 6242 8792
rect 8021 8789 8033 8823
rect 8067 8820 8079 8823
rect 8294 8820 8300 8832
rect 8067 8792 8300 8820
rect 8067 8789 8079 8792
rect 8021 8783 8079 8789
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 8570 8780 8576 8832
rect 8628 8780 8634 8832
rect 8665 8823 8723 8829
rect 8665 8789 8677 8823
rect 8711 8820 8723 8823
rect 9766 8820 9772 8832
rect 8711 8792 9772 8820
rect 8711 8789 8723 8792
rect 8665 8783 8723 8789
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 10042 8780 10048 8832
rect 10100 8820 10106 8832
rect 10962 8820 10968 8832
rect 10100 8792 10968 8820
rect 10100 8780 10106 8792
rect 10962 8780 10968 8792
rect 11020 8780 11026 8832
rect 11425 8823 11483 8829
rect 11425 8789 11437 8823
rect 11471 8820 11483 8823
rect 11790 8820 11796 8832
rect 11471 8792 11796 8820
rect 11471 8789 11483 8792
rect 11425 8783 11483 8789
rect 11790 8780 11796 8792
rect 11848 8780 11854 8832
rect 11882 8780 11888 8832
rect 11940 8820 11946 8832
rect 14366 8820 14372 8832
rect 11940 8792 14372 8820
rect 11940 8780 11946 8792
rect 14366 8780 14372 8792
rect 14424 8780 14430 8832
rect 1104 8730 17388 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 17388 8730
rect 1104 8656 17388 8678
rect 2406 8576 2412 8628
rect 2464 8576 2470 8628
rect 2777 8619 2835 8625
rect 2777 8585 2789 8619
rect 2823 8616 2835 8619
rect 2866 8616 2872 8628
rect 2823 8588 2872 8616
rect 2823 8585 2835 8588
rect 2777 8579 2835 8585
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 2958 8576 2964 8628
rect 3016 8616 3022 8628
rect 6730 8616 6736 8628
rect 3016 8588 6736 8616
rect 3016 8576 3022 8588
rect 6730 8576 6736 8588
rect 6788 8576 6794 8628
rect 7834 8576 7840 8628
rect 7892 8616 7898 8628
rect 8205 8619 8263 8625
rect 8205 8616 8217 8619
rect 7892 8588 8217 8616
rect 7892 8576 7898 8588
rect 8205 8585 8217 8588
rect 8251 8585 8263 8619
rect 8205 8579 8263 8585
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 9030 8616 9036 8628
rect 8352 8588 9036 8616
rect 8352 8576 8358 8588
rect 9030 8576 9036 8588
rect 9088 8576 9094 8628
rect 9858 8576 9864 8628
rect 9916 8616 9922 8628
rect 10686 8616 10692 8628
rect 9916 8588 10692 8616
rect 9916 8576 9922 8588
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 11882 8576 11888 8628
rect 11940 8576 11946 8628
rect 12986 8576 12992 8628
rect 13044 8576 13050 8628
rect 13446 8576 13452 8628
rect 13504 8576 13510 8628
rect 13909 8619 13967 8625
rect 13909 8585 13921 8619
rect 13955 8585 13967 8619
rect 13909 8579 13967 8585
rect 2222 8508 2228 8560
rect 2280 8508 2286 8560
rect 2317 8551 2375 8557
rect 2317 8517 2329 8551
rect 2363 8548 2375 8551
rect 2682 8548 2688 8560
rect 2363 8520 2688 8548
rect 2363 8517 2375 8520
rect 2317 8511 2375 8517
rect 2682 8508 2688 8520
rect 2740 8508 2746 8560
rect 3510 8508 3516 8560
rect 3568 8548 3574 8560
rect 5077 8551 5135 8557
rect 5077 8548 5089 8551
rect 3568 8520 5089 8548
rect 3568 8508 3574 8520
rect 5077 8517 5089 8520
rect 5123 8517 5135 8551
rect 5077 8511 5135 8517
rect 5534 8508 5540 8560
rect 5592 8548 5598 8560
rect 6638 8548 6644 8560
rect 5592 8520 6644 8548
rect 5592 8508 5598 8520
rect 6638 8508 6644 8520
rect 6696 8508 6702 8560
rect 3050 8440 3056 8492
rect 3108 8480 3114 8492
rect 3329 8483 3387 8489
rect 3329 8480 3341 8483
rect 3108 8452 3341 8480
rect 3108 8440 3114 8452
rect 3329 8449 3341 8452
rect 3375 8449 3387 8483
rect 3329 8443 3387 8449
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8381 3019 8415
rect 4816 8412 4844 8443
rect 4982 8440 4988 8492
rect 5040 8440 5046 8492
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 6748 8480 6776 8576
rect 7374 8508 7380 8560
rect 7432 8548 7438 8560
rect 7745 8551 7803 8557
rect 7745 8548 7757 8551
rect 7432 8520 7757 8548
rect 7432 8508 7438 8520
rect 7745 8517 7757 8520
rect 7791 8517 7803 8551
rect 7745 8511 7803 8517
rect 9493 8551 9551 8557
rect 9493 8517 9505 8551
rect 9539 8548 9551 8551
rect 9582 8548 9588 8560
rect 9539 8520 9588 8548
rect 9539 8517 9551 8520
rect 9493 8511 9551 8517
rect 9582 8508 9588 8520
rect 9640 8508 9646 8560
rect 9766 8508 9772 8560
rect 9824 8508 9830 8560
rect 10594 8548 10600 8560
rect 10060 8520 10600 8548
rect 7469 8483 7527 8489
rect 7469 8480 7481 8483
rect 5215 8452 5764 8480
rect 6748 8452 7481 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 5258 8412 5264 8424
rect 4816 8384 5264 8412
rect 2961 8375 3019 8381
rect 2130 8304 2136 8356
rect 2188 8344 2194 8356
rect 2976 8344 3004 8375
rect 5258 8372 5264 8384
rect 5316 8372 5322 8424
rect 3513 8347 3571 8353
rect 3513 8344 3525 8347
rect 2188 8316 3525 8344
rect 2188 8304 2194 8316
rect 3513 8313 3525 8316
rect 3559 8344 3571 8347
rect 4062 8344 4068 8356
rect 3559 8316 4068 8344
rect 3559 8313 3571 8316
rect 3513 8307 3571 8313
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 5350 8304 5356 8356
rect 5408 8304 5414 8356
rect 5736 8344 5764 8452
rect 7469 8449 7481 8452
rect 7515 8480 7527 8483
rect 7558 8480 7564 8492
rect 7515 8452 7564 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 7650 8440 7656 8492
rect 7708 8440 7714 8492
rect 7834 8440 7840 8492
rect 7892 8480 7898 8492
rect 8018 8480 8024 8492
rect 7892 8452 8024 8480
rect 7892 8440 7898 8452
rect 8018 8440 8024 8452
rect 8076 8440 8082 8492
rect 8294 8440 8300 8492
rect 8352 8440 8358 8492
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8480 9367 8483
rect 9398 8480 9404 8492
rect 9355 8452 9404 8480
rect 9355 8449 9367 8452
rect 9309 8443 9367 8449
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 10060 8489 10088 8520
rect 10594 8508 10600 8520
rect 10652 8508 10658 8560
rect 11054 8508 11060 8560
rect 11112 8548 11118 8560
rect 11112 8520 13676 8548
rect 11112 8508 11118 8520
rect 10045 8483 10103 8489
rect 10045 8480 10057 8483
rect 9600 8452 10057 8480
rect 5810 8372 5816 8424
rect 5868 8412 5874 8424
rect 9600 8412 9628 8452
rect 10045 8449 10057 8452
rect 10091 8449 10103 8483
rect 10045 8443 10103 8449
rect 10226 8440 10232 8492
rect 10284 8480 10290 8492
rect 10321 8483 10379 8489
rect 10321 8480 10333 8483
rect 10284 8452 10333 8480
rect 10284 8440 10290 8452
rect 10321 8449 10333 8452
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 10410 8440 10416 8492
rect 10468 8480 10474 8492
rect 10505 8483 10563 8489
rect 10505 8480 10517 8483
rect 10468 8452 10517 8480
rect 10468 8440 10474 8452
rect 10505 8449 10517 8452
rect 10551 8480 10563 8483
rect 10686 8480 10692 8492
rect 10551 8452 10692 8480
rect 10551 8449 10563 8452
rect 10505 8443 10563 8449
rect 10686 8440 10692 8452
rect 10744 8440 10750 8492
rect 11514 8440 11520 8492
rect 11572 8440 11578 8492
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8480 12863 8483
rect 12894 8480 12900 8492
rect 12851 8452 12900 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 13078 8440 13084 8492
rect 13136 8440 13142 8492
rect 13538 8440 13544 8492
rect 13596 8440 13602 8492
rect 13648 8480 13676 8520
rect 13924 8480 13952 8579
rect 15286 8576 15292 8628
rect 15344 8616 15350 8628
rect 15470 8616 15476 8628
rect 15344 8588 15476 8616
rect 15344 8576 15350 8588
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 16942 8576 16948 8628
rect 17000 8576 17006 8628
rect 15304 8548 15332 8576
rect 15381 8551 15439 8557
rect 15381 8548 15393 8551
rect 15304 8520 15393 8548
rect 15381 8517 15393 8520
rect 15427 8517 15439 8551
rect 15746 8548 15752 8560
rect 15381 8511 15439 8517
rect 15488 8520 15752 8548
rect 14001 8483 14059 8489
rect 14001 8480 14013 8483
rect 13648 8452 13768 8480
rect 13924 8452 14013 8480
rect 5868 8384 9628 8412
rect 9677 8415 9735 8421
rect 5868 8372 5874 8384
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 9950 8412 9956 8424
rect 9723 8384 9956 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 10962 8372 10968 8424
rect 11020 8412 11026 8424
rect 11609 8415 11667 8421
rect 11609 8412 11621 8415
rect 11020 8384 11621 8412
rect 11020 8372 11026 8384
rect 11609 8381 11621 8384
rect 11655 8381 11667 8415
rect 11609 8375 11667 8381
rect 11698 8372 11704 8424
rect 11756 8412 11762 8424
rect 12618 8412 12624 8424
rect 11756 8384 12624 8412
rect 11756 8372 11762 8384
rect 12618 8372 12624 8384
rect 12676 8372 12682 8424
rect 12713 8415 12771 8421
rect 12713 8381 12725 8415
rect 12759 8381 12771 8415
rect 12713 8375 12771 8381
rect 6178 8344 6184 8356
rect 5736 8316 6184 8344
rect 6178 8304 6184 8316
rect 6236 8344 6242 8356
rect 6914 8344 6920 8356
rect 6236 8316 6920 8344
rect 6236 8304 6242 8316
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 7558 8304 7564 8356
rect 7616 8344 7622 8356
rect 7926 8344 7932 8356
rect 7616 8316 7932 8344
rect 7616 8304 7622 8316
rect 7926 8304 7932 8316
rect 7984 8304 7990 8356
rect 8021 8347 8079 8353
rect 8021 8313 8033 8347
rect 8067 8344 8079 8347
rect 11146 8344 11152 8356
rect 8067 8316 11152 8344
rect 8067 8313 8079 8316
rect 8021 8307 8079 8313
rect 11146 8304 11152 8316
rect 11204 8344 11210 8356
rect 12728 8344 12756 8375
rect 12986 8372 12992 8424
rect 13044 8412 13050 8424
rect 13173 8415 13231 8421
rect 13173 8412 13185 8415
rect 13044 8384 13185 8412
rect 13044 8372 13050 8384
rect 13173 8381 13185 8384
rect 13219 8381 13231 8415
rect 13173 8375 13231 8381
rect 13262 8372 13268 8424
rect 13320 8412 13326 8424
rect 13446 8412 13452 8424
rect 13320 8384 13452 8412
rect 13320 8372 13326 8384
rect 13446 8372 13452 8384
rect 13504 8412 13510 8424
rect 13633 8415 13691 8421
rect 13633 8412 13645 8415
rect 13504 8384 13645 8412
rect 13504 8372 13510 8384
rect 13633 8381 13645 8384
rect 13679 8381 13691 8415
rect 13740 8412 13768 8452
rect 14001 8449 14013 8452
rect 14047 8449 14059 8483
rect 14001 8443 14059 8449
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8480 14151 8483
rect 14550 8480 14556 8492
rect 14139 8452 14556 8480
rect 14139 8449 14151 8452
rect 14093 8443 14151 8449
rect 14550 8440 14556 8452
rect 14608 8440 14614 8492
rect 15194 8440 15200 8492
rect 15252 8440 15258 8492
rect 15286 8440 15292 8492
rect 15344 8480 15350 8492
rect 15488 8489 15516 8520
rect 15746 8508 15752 8520
rect 15804 8508 15810 8560
rect 15473 8483 15531 8489
rect 15473 8480 15485 8483
rect 15344 8452 15485 8480
rect 15344 8440 15350 8452
rect 15473 8449 15485 8452
rect 15519 8449 15531 8483
rect 15473 8443 15531 8449
rect 15565 8483 15623 8489
rect 15565 8449 15577 8483
rect 15611 8480 15623 8483
rect 15841 8483 15899 8489
rect 15841 8480 15853 8483
rect 15611 8452 15853 8480
rect 15611 8449 15623 8452
rect 15565 8443 15623 8449
rect 15841 8449 15853 8452
rect 15887 8449 15899 8483
rect 15841 8443 15899 8449
rect 16761 8483 16819 8489
rect 16761 8449 16773 8483
rect 16807 8480 16819 8483
rect 16850 8480 16856 8492
rect 16807 8452 16856 8480
rect 16807 8449 16819 8452
rect 16761 8443 16819 8449
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 14277 8415 14335 8421
rect 14277 8412 14289 8415
rect 13740 8384 14289 8412
rect 13633 8375 13691 8381
rect 14277 8381 14289 8384
rect 14323 8381 14335 8415
rect 14277 8375 14335 8381
rect 16485 8415 16543 8421
rect 16485 8381 16497 8415
rect 16531 8412 16543 8415
rect 17034 8412 17040 8424
rect 16531 8384 17040 8412
rect 16531 8381 16543 8384
rect 16485 8375 16543 8381
rect 17034 8372 17040 8384
rect 17092 8372 17098 8424
rect 11204 8316 13124 8344
rect 11204 8304 11210 8316
rect 3786 8236 3792 8288
rect 3844 8276 3850 8288
rect 4154 8276 4160 8288
rect 3844 8248 4160 8276
rect 3844 8236 3850 8248
rect 4154 8236 4160 8248
rect 4212 8236 4218 8288
rect 5074 8236 5080 8288
rect 5132 8276 5138 8288
rect 5902 8276 5908 8288
rect 5132 8248 5908 8276
rect 5132 8236 5138 8248
rect 5902 8236 5908 8248
rect 5960 8236 5966 8288
rect 8570 8236 8576 8288
rect 8628 8276 8634 8288
rect 9306 8276 9312 8288
rect 8628 8248 9312 8276
rect 8628 8236 8634 8248
rect 9306 8236 9312 8248
rect 9364 8236 9370 8288
rect 9766 8236 9772 8288
rect 9824 8276 9830 8288
rect 10134 8276 10140 8288
rect 9824 8248 10140 8276
rect 9824 8236 9830 8248
rect 10134 8236 10140 8248
rect 10192 8236 10198 8288
rect 10229 8279 10287 8285
rect 10229 8245 10241 8279
rect 10275 8276 10287 8279
rect 10594 8276 10600 8288
rect 10275 8248 10600 8276
rect 10275 8245 10287 8248
rect 10229 8239 10287 8245
rect 10594 8236 10600 8248
rect 10652 8236 10658 8288
rect 11330 8236 11336 8288
rect 11388 8276 11394 8288
rect 11517 8279 11575 8285
rect 11517 8276 11529 8279
rect 11388 8248 11529 8276
rect 11388 8236 11394 8248
rect 11517 8245 11529 8248
rect 11563 8276 11575 8279
rect 11882 8276 11888 8288
rect 11563 8248 11888 8276
rect 11563 8245 11575 8248
rect 11517 8239 11575 8245
rect 11882 8236 11888 8248
rect 11940 8236 11946 8288
rect 12618 8236 12624 8288
rect 12676 8276 12682 8288
rect 12986 8276 12992 8288
rect 12676 8248 12992 8276
rect 12676 8236 12682 8248
rect 12986 8236 12992 8248
rect 13044 8236 13050 8288
rect 13096 8285 13124 8316
rect 13998 8304 14004 8356
rect 14056 8304 14062 8356
rect 13081 8279 13139 8285
rect 13081 8245 13093 8279
rect 13127 8245 13139 8279
rect 13081 8239 13139 8245
rect 13725 8279 13783 8285
rect 13725 8245 13737 8279
rect 13771 8276 13783 8279
rect 13814 8276 13820 8288
rect 13771 8248 13820 8276
rect 13771 8245 13783 8248
rect 13725 8239 13783 8245
rect 13814 8236 13820 8248
rect 13872 8236 13878 8288
rect 15746 8236 15752 8288
rect 15804 8236 15810 8288
rect 1104 8186 17388 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 17388 8186
rect 1104 8112 17388 8134
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 3602 8072 3608 8084
rect 2832 8044 3608 8072
rect 2832 8032 2838 8044
rect 3602 8032 3608 8044
rect 3660 8072 3666 8084
rect 5997 8075 6055 8081
rect 3660 8044 4016 8072
rect 3660 8032 3666 8044
rect 2682 7964 2688 8016
rect 2740 8004 2746 8016
rect 3694 8004 3700 8016
rect 2740 7976 3700 8004
rect 2740 7964 2746 7976
rect 3694 7964 3700 7976
rect 3752 7964 3758 8016
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7936 2283 7939
rect 2958 7936 2964 7948
rect 2271 7908 2964 7936
rect 2271 7905 2283 7908
rect 2225 7899 2283 7905
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 2038 7828 2044 7880
rect 2096 7828 2102 7880
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 2639 7840 2912 7868
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 2774 7760 2780 7812
rect 2832 7760 2838 7812
rect 2884 7800 2912 7840
rect 3142 7828 3148 7880
rect 3200 7868 3206 7880
rect 3421 7871 3479 7877
rect 3421 7868 3433 7871
rect 3200 7840 3433 7868
rect 3200 7828 3206 7840
rect 3421 7837 3433 7840
rect 3467 7837 3479 7871
rect 3421 7831 3479 7837
rect 3878 7828 3884 7880
rect 3936 7828 3942 7880
rect 3988 7877 4016 8044
rect 4816 8044 5948 8072
rect 4062 7896 4068 7948
rect 4120 7936 4126 7948
rect 4617 7939 4675 7945
rect 4617 7936 4629 7939
rect 4120 7908 4629 7936
rect 4120 7896 4126 7908
rect 4617 7905 4629 7908
rect 4663 7905 4675 7939
rect 4816 7936 4844 8044
rect 5350 7964 5356 8016
rect 5408 8004 5414 8016
rect 5534 8004 5540 8016
rect 5408 7976 5540 8004
rect 5408 7964 5414 7976
rect 5534 7964 5540 7976
rect 5592 7964 5598 8016
rect 5810 7964 5816 8016
rect 5868 7964 5874 8016
rect 5920 8004 5948 8044
rect 5997 8041 6009 8075
rect 6043 8072 6055 8075
rect 6086 8072 6092 8084
rect 6043 8044 6092 8072
rect 6043 8041 6055 8044
rect 5997 8035 6055 8041
rect 6086 8032 6092 8044
rect 6144 8032 6150 8084
rect 6733 8075 6791 8081
rect 6733 8041 6745 8075
rect 6779 8072 6791 8075
rect 9766 8072 9772 8084
rect 6779 8044 9772 8072
rect 6779 8041 6791 8044
rect 6733 8035 6791 8041
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 10965 8075 11023 8081
rect 10965 8072 10977 8075
rect 9968 8044 10977 8072
rect 6270 8004 6276 8016
rect 5920 7976 6276 8004
rect 6270 7964 6276 7976
rect 6328 7964 6334 8016
rect 6638 7964 6644 8016
rect 6696 8004 6702 8016
rect 7837 8007 7895 8013
rect 6696 7976 7788 8004
rect 6696 7964 6702 7976
rect 5626 7936 5632 7948
rect 4617 7899 4675 7905
rect 4724 7908 4844 7936
rect 5000 7908 5632 7936
rect 4724 7877 4752 7908
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7837 4767 7871
rect 4709 7831 4767 7837
rect 4798 7828 4804 7880
rect 4856 7868 4862 7880
rect 5000 7877 5028 7908
rect 5626 7896 5632 7908
rect 5684 7936 5690 7948
rect 5828 7936 5856 7964
rect 7466 7936 7472 7948
rect 5684 7908 6316 7936
rect 5684 7896 5690 7908
rect 4893 7871 4951 7877
rect 4893 7868 4905 7871
rect 4856 7840 4905 7868
rect 4856 7828 4862 7840
rect 4893 7837 4905 7840
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 5074 7828 5080 7880
rect 5132 7828 5138 7880
rect 5350 7828 5356 7880
rect 5408 7828 5414 7880
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7868 5595 7871
rect 5813 7871 5871 7877
rect 5583 7840 5764 7868
rect 5583 7837 5595 7840
rect 5537 7831 5595 7837
rect 2958 7800 2964 7812
rect 2884 7772 2964 7800
rect 2958 7760 2964 7772
rect 3016 7760 3022 7812
rect 4430 7760 4436 7812
rect 4488 7800 4494 7812
rect 5092 7800 5120 7828
rect 5626 7800 5632 7812
rect 4488 7772 5120 7800
rect 5276 7772 5632 7800
rect 4488 7760 4494 7772
rect 2682 7692 2688 7744
rect 2740 7732 2746 7744
rect 2866 7732 2872 7744
rect 2740 7704 2872 7732
rect 2740 7692 2746 7704
rect 2866 7692 2872 7704
rect 2924 7692 2930 7744
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 5276 7741 5304 7772
rect 5626 7760 5632 7772
rect 5684 7760 5690 7812
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 4028 7704 4077 7732
rect 4028 7692 4034 7704
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 4065 7695 4123 7701
rect 5261 7735 5319 7741
rect 5261 7701 5273 7735
rect 5307 7701 5319 7735
rect 5261 7695 5319 7701
rect 5350 7692 5356 7744
rect 5408 7732 5414 7744
rect 5736 7732 5764 7840
rect 5813 7837 5825 7871
rect 5859 7868 5871 7871
rect 5902 7868 5908 7880
rect 5859 7840 5908 7868
rect 5859 7837 5871 7840
rect 5813 7831 5871 7837
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7868 6147 7871
rect 6178 7868 6184 7880
rect 6135 7840 6184 7868
rect 6135 7837 6147 7840
rect 6089 7831 6147 7837
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 6288 7877 6316 7908
rect 7208 7908 7472 7936
rect 7208 7877 7236 7908
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 7760 7936 7788 7976
rect 7837 7973 7849 8007
rect 7883 8004 7895 8007
rect 8386 8004 8392 8016
rect 7883 7976 8392 8004
rect 7883 7973 7895 7976
rect 7837 7967 7895 7973
rect 8386 7964 8392 7976
rect 8444 7964 8450 8016
rect 8481 8007 8539 8013
rect 8481 7973 8493 8007
rect 8527 8004 8539 8007
rect 9968 8004 9996 8044
rect 10965 8041 10977 8044
rect 11011 8072 11023 8075
rect 11330 8072 11336 8084
rect 11011 8044 11336 8072
rect 11011 8041 11023 8044
rect 10965 8035 11023 8041
rect 11330 8032 11336 8044
rect 11388 8032 11394 8084
rect 11422 8032 11428 8084
rect 11480 8032 11486 8084
rect 11514 8032 11520 8084
rect 11572 8072 11578 8084
rect 11701 8075 11759 8081
rect 11701 8072 11713 8075
rect 11572 8044 11713 8072
rect 11572 8032 11578 8044
rect 11701 8041 11713 8044
rect 11747 8041 11759 8075
rect 11701 8035 11759 8041
rect 13541 8075 13599 8081
rect 13541 8041 13553 8075
rect 13587 8072 13599 8075
rect 13814 8072 13820 8084
rect 13587 8044 13820 8072
rect 13587 8041 13599 8044
rect 13541 8035 13599 8041
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 14553 8075 14611 8081
rect 14553 8041 14565 8075
rect 14599 8072 14611 8075
rect 14642 8072 14648 8084
rect 14599 8044 14648 8072
rect 14599 8041 14611 8044
rect 14553 8035 14611 8041
rect 14642 8032 14648 8044
rect 14700 8032 14706 8084
rect 15010 8032 15016 8084
rect 15068 8032 15074 8084
rect 15194 8032 15200 8084
rect 15252 8072 15258 8084
rect 15381 8075 15439 8081
rect 15381 8072 15393 8075
rect 15252 8044 15393 8072
rect 15252 8032 15258 8044
rect 15381 8041 15393 8044
rect 15427 8041 15439 8075
rect 15381 8035 15439 8041
rect 17034 8032 17040 8084
rect 17092 8032 17098 8084
rect 8527 7976 9812 8004
rect 8527 7973 8539 7976
rect 8481 7967 8539 7973
rect 9784 7948 9812 7976
rect 9876 7976 9996 8004
rect 7714 7908 7972 7936
rect 7374 7877 7380 7880
rect 6273 7871 6331 7877
rect 6273 7837 6285 7871
rect 6319 7837 6331 7871
rect 6273 7831 6331 7837
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 7193 7871 7251 7877
rect 7193 7837 7205 7871
rect 7239 7837 7251 7871
rect 7193 7831 7251 7837
rect 7341 7871 7380 7877
rect 7341 7837 7353 7871
rect 7341 7831 7380 7837
rect 5920 7800 5948 7828
rect 6564 7800 6592 7831
rect 7374 7828 7380 7831
rect 7432 7828 7438 7880
rect 7558 7828 7564 7880
rect 7616 7828 7622 7880
rect 7714 7877 7742 7908
rect 7944 7880 7972 7908
rect 9766 7896 9772 7948
rect 9824 7896 9830 7948
rect 7697 7871 7755 7877
rect 7697 7837 7709 7871
rect 7743 7837 7755 7871
rect 7697 7831 7755 7837
rect 7926 7828 7932 7880
rect 7984 7828 7990 7880
rect 8018 7828 8024 7880
rect 8076 7868 8082 7880
rect 8113 7871 8171 7877
rect 8113 7868 8125 7871
rect 8076 7840 8125 7868
rect 8076 7828 8082 7840
rect 8113 7837 8125 7840
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 8202 7828 8208 7880
rect 8260 7828 8266 7880
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 5920 7772 6592 7800
rect 7469 7803 7527 7809
rect 7469 7769 7481 7803
rect 7515 7800 7527 7803
rect 8312 7800 8340 7831
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 9876 7868 9904 7976
rect 10502 7964 10508 8016
rect 10560 8004 10566 8016
rect 11241 8007 11299 8013
rect 10560 7976 11192 8004
rect 10560 7964 10566 7976
rect 9950 7896 9956 7948
rect 10008 7936 10014 7948
rect 10873 7939 10931 7945
rect 10873 7936 10885 7939
rect 10008 7908 10885 7936
rect 10008 7896 10014 7908
rect 10873 7905 10885 7908
rect 10919 7905 10931 7939
rect 11164 7936 11192 7976
rect 11241 7973 11253 8007
rect 11287 8004 11299 8007
rect 14369 8007 14427 8013
rect 14369 8004 14381 8007
rect 11287 7976 14381 8004
rect 11287 7973 11299 7976
rect 11241 7967 11299 7973
rect 14369 7973 14381 7976
rect 14415 8004 14427 8007
rect 14415 7976 15148 8004
rect 14415 7973 14427 7976
rect 14369 7967 14427 7973
rect 11514 7936 11520 7948
rect 11164 7908 11520 7936
rect 10873 7899 10931 7905
rect 11514 7896 11520 7908
rect 11572 7936 11578 7948
rect 11572 7908 12434 7936
rect 11572 7896 11578 7908
rect 8536 7840 9904 7868
rect 8536 7828 8542 7840
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 10689 7871 10747 7877
rect 10689 7868 10701 7871
rect 10376 7840 10701 7868
rect 10376 7828 10382 7840
rect 10689 7837 10701 7840
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 11054 7828 11060 7880
rect 11112 7828 11118 7880
rect 11330 7828 11336 7880
rect 11388 7828 11394 7880
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7837 11483 7871
rect 12406 7868 12434 7908
rect 12894 7896 12900 7948
rect 12952 7936 12958 7948
rect 15120 7945 15148 7976
rect 13357 7939 13415 7945
rect 13357 7936 13369 7939
rect 12952 7908 13369 7936
rect 12952 7896 12958 7908
rect 13357 7905 13369 7908
rect 13403 7905 13415 7939
rect 14461 7939 14519 7945
rect 14461 7936 14473 7939
rect 13357 7899 13415 7905
rect 13464 7908 14473 7936
rect 13464 7868 13492 7908
rect 14461 7905 14473 7908
rect 14507 7905 14519 7939
rect 14461 7899 14519 7905
rect 15105 7939 15163 7945
rect 15105 7905 15117 7939
rect 15151 7905 15163 7939
rect 15105 7899 15163 7905
rect 12406 7840 13492 7868
rect 11425 7831 11483 7837
rect 7515 7772 8340 7800
rect 7515 7769 7527 7772
rect 7469 7763 7527 7769
rect 6546 7732 6552 7744
rect 5408 7704 6552 7732
rect 5408 7692 5414 7704
rect 6546 7692 6552 7704
rect 6604 7732 6610 7744
rect 7484 7732 7512 7763
rect 8036 7744 8064 7772
rect 8662 7760 8668 7812
rect 8720 7800 8726 7812
rect 8720 7772 9674 7800
rect 8720 7760 8726 7772
rect 6604 7704 7512 7732
rect 6604 7692 6610 7704
rect 8018 7692 8024 7744
rect 8076 7692 8082 7744
rect 9214 7692 9220 7744
rect 9272 7692 9278 7744
rect 9646 7732 9674 7772
rect 10042 7760 10048 7812
rect 10100 7800 10106 7812
rect 10781 7803 10839 7809
rect 10781 7800 10793 7803
rect 10100 7772 10793 7800
rect 10100 7760 10106 7772
rect 10781 7769 10793 7772
rect 10827 7800 10839 7803
rect 11440 7800 11468 7831
rect 13538 7828 13544 7880
rect 13596 7828 13602 7880
rect 14185 7871 14243 7877
rect 14185 7868 14197 7871
rect 13740 7840 14197 7868
rect 10827 7772 11468 7800
rect 10827 7769 10839 7772
rect 10781 7763 10839 7769
rect 13262 7760 13268 7812
rect 13320 7760 13326 7812
rect 10134 7732 10140 7744
rect 9646 7704 10140 7732
rect 10134 7692 10140 7704
rect 10192 7692 10198 7744
rect 10594 7692 10600 7744
rect 10652 7732 10658 7744
rect 12802 7732 12808 7744
rect 10652 7704 12808 7732
rect 10652 7692 10658 7704
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 13740 7741 13768 7840
rect 14185 7837 14197 7840
rect 14231 7837 14243 7871
rect 14185 7831 14243 7837
rect 14645 7871 14703 7877
rect 14645 7837 14657 7871
rect 14691 7837 14703 7871
rect 14645 7831 14703 7837
rect 14660 7800 14688 7831
rect 15010 7828 15016 7880
rect 15068 7828 15074 7880
rect 15654 7828 15660 7880
rect 15712 7828 15718 7880
rect 15746 7828 15752 7880
rect 15804 7868 15810 7880
rect 15913 7871 15971 7877
rect 15913 7868 15925 7871
rect 15804 7840 15925 7868
rect 15804 7828 15810 7840
rect 15913 7837 15925 7840
rect 15959 7837 15971 7871
rect 15913 7831 15971 7837
rect 15562 7800 15568 7812
rect 14660 7772 15568 7800
rect 15562 7760 15568 7772
rect 15620 7760 15626 7812
rect 13725 7735 13783 7741
rect 13725 7701 13737 7735
rect 13771 7701 13783 7735
rect 13725 7695 13783 7701
rect 14734 7692 14740 7744
rect 14792 7732 14798 7744
rect 14921 7735 14979 7741
rect 14921 7732 14933 7735
rect 14792 7704 14933 7732
rect 14792 7692 14798 7704
rect 14921 7701 14933 7704
rect 14967 7701 14979 7735
rect 14921 7695 14979 7701
rect 1104 7642 17388 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 17388 7642
rect 1104 7568 17388 7590
rect 1765 7531 1823 7537
rect 1765 7497 1777 7531
rect 1811 7528 1823 7531
rect 2590 7528 2596 7540
rect 1811 7500 2596 7528
rect 1811 7497 1823 7500
rect 1765 7491 1823 7497
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 2866 7488 2872 7540
rect 2924 7528 2930 7540
rect 3510 7528 3516 7540
rect 2924 7500 3516 7528
rect 2924 7488 2930 7500
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 3878 7488 3884 7540
rect 3936 7488 3942 7540
rect 3970 7488 3976 7540
rect 4028 7488 4034 7540
rect 4798 7488 4804 7540
rect 4856 7488 4862 7540
rect 4982 7488 4988 7540
rect 5040 7528 5046 7540
rect 5442 7528 5448 7540
rect 5040 7500 5448 7528
rect 5040 7488 5046 7500
rect 2774 7460 2780 7472
rect 1964 7432 2780 7460
rect 1964 7401 1992 7432
rect 2774 7420 2780 7432
rect 2832 7460 2838 7472
rect 3142 7460 3148 7472
rect 2832 7432 3148 7460
rect 2832 7420 2838 7432
rect 3142 7420 3148 7432
rect 3200 7420 3206 7472
rect 3237 7463 3295 7469
rect 3237 7429 3249 7463
rect 3283 7460 3295 7463
rect 3326 7460 3332 7472
rect 3283 7432 3332 7460
rect 3283 7429 3295 7432
rect 3237 7423 3295 7429
rect 3326 7420 3332 7432
rect 3384 7420 3390 7472
rect 3418 7420 3424 7472
rect 3476 7420 3482 7472
rect 3602 7420 3608 7472
rect 3660 7420 3666 7472
rect 4062 7420 4068 7472
rect 4120 7420 4126 7472
rect 4341 7463 4399 7469
rect 4341 7429 4353 7463
rect 4387 7460 4399 7463
rect 4709 7463 4767 7469
rect 4709 7460 4721 7463
rect 4387 7432 4721 7460
rect 4387 7429 4399 7432
rect 4341 7423 4399 7429
rect 4709 7429 4721 7432
rect 4755 7460 4767 7463
rect 4816 7460 4844 7488
rect 5276 7469 5304 7500
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 9122 7488 9128 7540
rect 9180 7488 9186 7540
rect 9306 7488 9312 7540
rect 9364 7488 9370 7540
rect 10042 7488 10048 7540
rect 10100 7488 10106 7540
rect 10505 7531 10563 7537
rect 10505 7497 10517 7531
rect 10551 7528 10563 7531
rect 11330 7528 11336 7540
rect 10551 7500 11336 7528
rect 10551 7497 10563 7500
rect 10505 7491 10563 7497
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 12529 7531 12587 7537
rect 12529 7497 12541 7531
rect 12575 7528 12587 7531
rect 12575 7500 12664 7528
rect 12575 7497 12587 7500
rect 12529 7491 12587 7497
rect 5261 7463 5319 7469
rect 4755 7432 5212 7460
rect 4755 7429 4767 7432
rect 4709 7423 4767 7429
rect 1949 7395 2007 7401
rect 1949 7361 1961 7395
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 2038 7352 2044 7404
rect 2096 7392 2102 7404
rect 2225 7395 2283 7401
rect 2225 7392 2237 7395
rect 2096 7364 2237 7392
rect 2096 7352 2102 7364
rect 2225 7361 2237 7364
rect 2271 7361 2283 7395
rect 2225 7355 2283 7361
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 2590 7392 2596 7404
rect 2547 7364 2596 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2240 7324 2268 7355
rect 2590 7352 2596 7364
rect 2648 7352 2654 7404
rect 2682 7352 2688 7404
rect 2740 7352 2746 7404
rect 2958 7352 2964 7404
rect 3016 7392 3022 7404
rect 3053 7395 3111 7401
rect 3053 7392 3065 7395
rect 3016 7364 3065 7392
rect 3016 7352 3022 7364
rect 3053 7361 3065 7364
rect 3099 7392 3111 7395
rect 3436 7392 3464 7420
rect 3099 7364 3464 7392
rect 3099 7361 3111 7364
rect 3053 7355 3111 7361
rect 4430 7352 4436 7404
rect 4488 7352 4494 7404
rect 4614 7352 4620 7404
rect 4672 7352 4678 7404
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 2777 7327 2835 7333
rect 2240 7296 2360 7324
rect 2332 7256 2360 7296
rect 2777 7293 2789 7327
rect 2823 7324 2835 7327
rect 4062 7324 4068 7336
rect 2823 7296 4068 7324
rect 2823 7293 2835 7296
rect 2777 7287 2835 7293
rect 4062 7284 4068 7296
rect 4120 7284 4126 7336
rect 3786 7256 3792 7268
rect 2332 7228 3792 7256
rect 3786 7216 3792 7228
rect 3844 7216 3850 7268
rect 4632 7188 4660 7352
rect 4816 7324 4844 7355
rect 5074 7352 5080 7404
rect 5132 7352 5138 7404
rect 5184 7392 5212 7432
rect 5261 7429 5273 7463
rect 5307 7429 5319 7463
rect 6086 7460 6092 7472
rect 5261 7423 5319 7429
rect 5460 7432 6092 7460
rect 5460 7404 5488 7432
rect 6086 7420 6092 7432
rect 6144 7420 6150 7472
rect 9140 7460 9168 7488
rect 9677 7463 9735 7469
rect 9140 7432 9352 7460
rect 9324 7404 9352 7432
rect 9677 7429 9689 7463
rect 9723 7460 9735 7463
rect 9766 7460 9772 7472
rect 9723 7432 9772 7460
rect 9723 7429 9735 7432
rect 9677 7423 9735 7429
rect 9766 7420 9772 7432
rect 9824 7460 9830 7472
rect 10226 7460 10232 7472
rect 9824 7432 10232 7460
rect 9824 7420 9830 7432
rect 10226 7420 10232 7432
rect 10284 7420 10290 7472
rect 11238 7420 11244 7472
rect 11296 7460 11302 7472
rect 12636 7469 12664 7500
rect 15562 7488 15568 7540
rect 15620 7528 15626 7540
rect 15930 7528 15936 7540
rect 15620 7500 15936 7528
rect 15620 7488 15626 7500
rect 15930 7488 15936 7500
rect 15988 7488 15994 7540
rect 16298 7488 16304 7540
rect 16356 7488 16362 7540
rect 16942 7488 16948 7540
rect 17000 7488 17006 7540
rect 11517 7463 11575 7469
rect 11517 7460 11529 7463
rect 11296 7432 11529 7460
rect 11296 7420 11302 7432
rect 11517 7429 11529 7432
rect 11563 7460 11575 7463
rect 12621 7463 12679 7469
rect 11563 7432 12296 7460
rect 11563 7429 11575 7432
rect 11517 7423 11575 7429
rect 5353 7395 5411 7401
rect 5353 7392 5365 7395
rect 5184 7364 5365 7392
rect 5353 7361 5365 7364
rect 5399 7361 5411 7395
rect 5353 7355 5411 7361
rect 5442 7352 5448 7404
rect 5500 7352 5506 7404
rect 5626 7352 5632 7404
rect 5684 7392 5690 7404
rect 8386 7392 8392 7404
rect 5684 7364 8392 7392
rect 5684 7352 5690 7364
rect 8386 7352 8392 7364
rect 8444 7352 8450 7404
rect 8846 7352 8852 7404
rect 8904 7352 8910 7404
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 9306 7352 9312 7404
rect 9364 7352 9370 7404
rect 9858 7352 9864 7404
rect 9916 7352 9922 7404
rect 10134 7352 10140 7404
rect 10192 7352 10198 7404
rect 11790 7352 11796 7404
rect 11848 7352 11854 7404
rect 12066 7352 12072 7404
rect 12124 7352 12130 7404
rect 5534 7324 5540 7336
rect 4816 7296 5540 7324
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 7466 7284 7472 7336
rect 7524 7324 7530 7336
rect 8938 7324 8944 7336
rect 7524 7296 8944 7324
rect 7524 7284 7530 7296
rect 8938 7284 8944 7296
rect 8996 7284 9002 7336
rect 9140 7324 9168 7352
rect 10229 7327 10287 7333
rect 10229 7324 10241 7327
rect 9140 7296 10241 7324
rect 10229 7293 10241 7296
rect 10275 7293 10287 7327
rect 10229 7287 10287 7293
rect 11422 7284 11428 7336
rect 11480 7324 11486 7336
rect 11609 7327 11667 7333
rect 11609 7324 11621 7327
rect 11480 7296 11621 7324
rect 11480 7284 11486 7296
rect 11609 7293 11621 7296
rect 11655 7293 11667 7327
rect 11609 7287 11667 7293
rect 12161 7327 12219 7333
rect 12161 7293 12173 7327
rect 12207 7293 12219 7327
rect 12268 7324 12296 7432
rect 12621 7429 12633 7463
rect 12667 7429 12679 7463
rect 12621 7423 12679 7429
rect 12802 7420 12808 7472
rect 12860 7420 12866 7472
rect 12342 7352 12348 7404
rect 12400 7352 12406 7404
rect 16114 7352 16120 7404
rect 16172 7352 16178 7404
rect 16482 7352 16488 7404
rect 16540 7352 16546 7404
rect 16761 7395 16819 7401
rect 16761 7361 16773 7395
rect 16807 7392 16819 7395
rect 17034 7392 17040 7404
rect 16807 7364 17040 7392
rect 16807 7361 16819 7364
rect 16761 7355 16819 7361
rect 17034 7352 17040 7364
rect 17092 7352 17098 7404
rect 14366 7324 14372 7336
rect 12268 7296 14372 7324
rect 12161 7287 12219 7293
rect 4985 7259 5043 7265
rect 4985 7225 4997 7259
rect 5031 7256 5043 7259
rect 9398 7256 9404 7268
rect 5031 7228 9404 7256
rect 5031 7225 5043 7228
rect 4985 7219 5043 7225
rect 9398 7216 9404 7228
rect 9456 7256 9462 7268
rect 11977 7259 12035 7265
rect 9456 7228 10180 7256
rect 9456 7216 9462 7228
rect 5350 7188 5356 7200
rect 4632 7160 5356 7188
rect 5350 7148 5356 7160
rect 5408 7148 5414 7200
rect 5629 7191 5687 7197
rect 5629 7157 5641 7191
rect 5675 7188 5687 7191
rect 8662 7188 8668 7200
rect 5675 7160 8668 7188
rect 5675 7157 5687 7160
rect 5629 7151 5687 7157
rect 8662 7148 8668 7160
rect 8720 7148 8726 7200
rect 9125 7191 9183 7197
rect 9125 7157 9137 7191
rect 9171 7188 9183 7191
rect 9306 7188 9312 7200
rect 9171 7160 9312 7188
rect 9171 7157 9183 7160
rect 9125 7151 9183 7157
rect 9306 7148 9312 7160
rect 9364 7148 9370 7200
rect 10152 7197 10180 7228
rect 11977 7225 11989 7259
rect 12023 7256 12035 7259
rect 12176 7256 12204 7287
rect 14366 7284 14372 7296
rect 14424 7284 14430 7336
rect 12023 7228 12204 7256
rect 12023 7225 12035 7228
rect 11977 7219 12035 7225
rect 12526 7216 12532 7268
rect 12584 7256 12590 7268
rect 13078 7256 13084 7268
rect 12584 7228 13084 7256
rect 12584 7216 12590 7228
rect 13078 7216 13084 7228
rect 13136 7216 13142 7268
rect 10137 7191 10195 7197
rect 10137 7157 10149 7191
rect 10183 7157 10195 7191
rect 10137 7151 10195 7157
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 11606 7188 11612 7200
rect 11112 7160 11612 7188
rect 11112 7148 11118 7160
rect 11606 7148 11612 7160
rect 11664 7148 11670 7200
rect 11882 7148 11888 7200
rect 11940 7188 11946 7200
rect 12069 7191 12127 7197
rect 12069 7188 12081 7191
rect 11940 7160 12081 7188
rect 11940 7148 11946 7160
rect 12069 7157 12081 7160
rect 12115 7157 12127 7191
rect 12069 7151 12127 7157
rect 12986 7148 12992 7200
rect 13044 7148 13050 7200
rect 1104 7098 17388 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 17388 7098
rect 1104 7024 17388 7046
rect 2777 6987 2835 6993
rect 2777 6953 2789 6987
rect 2823 6984 2835 6987
rect 3326 6984 3332 6996
rect 2823 6956 3332 6984
rect 2823 6953 2835 6956
rect 2777 6947 2835 6953
rect 3326 6944 3332 6956
rect 3384 6944 3390 6996
rect 6086 6944 6092 6996
rect 6144 6984 6150 6996
rect 7558 6984 7564 6996
rect 6144 6956 7564 6984
rect 6144 6944 6150 6956
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 7668 6956 8432 6984
rect 7098 6876 7104 6928
rect 7156 6916 7162 6928
rect 7668 6916 7696 6956
rect 8404 6928 8432 6956
rect 8754 6944 8760 6996
rect 8812 6984 8818 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8812 6956 8953 6984
rect 8812 6944 8818 6956
rect 8941 6953 8953 6956
rect 8987 6953 8999 6987
rect 8941 6947 8999 6953
rect 9582 6944 9588 6996
rect 9640 6984 9646 6996
rect 9950 6984 9956 6996
rect 9640 6956 9956 6984
rect 9640 6944 9646 6956
rect 9950 6944 9956 6956
rect 10008 6944 10014 6996
rect 11146 6944 11152 6996
rect 11204 6944 11210 6996
rect 11609 6987 11667 6993
rect 11609 6953 11621 6987
rect 11655 6984 11667 6987
rect 12066 6984 12072 6996
rect 11655 6956 12072 6984
rect 11655 6953 11667 6956
rect 11609 6947 11667 6953
rect 12066 6944 12072 6956
rect 12124 6944 12130 6996
rect 12437 6987 12495 6993
rect 12437 6953 12449 6987
rect 12483 6953 12495 6987
rect 12437 6947 12495 6953
rect 12897 6987 12955 6993
rect 12897 6953 12909 6987
rect 12943 6984 12955 6987
rect 12943 6956 13308 6984
rect 12943 6953 12955 6956
rect 12897 6947 12955 6953
rect 7156 6888 7696 6916
rect 7156 6876 7162 6888
rect 6089 6851 6147 6857
rect 5644 6820 6040 6848
rect 1394 6740 1400 6792
rect 1452 6740 1458 6792
rect 4062 6740 4068 6792
rect 4120 6780 4126 6792
rect 4798 6780 4804 6792
rect 4120 6752 4804 6780
rect 4120 6740 4126 6752
rect 4798 6740 4804 6752
rect 4856 6740 4862 6792
rect 4982 6740 4988 6792
rect 5040 6740 5046 6792
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6780 5227 6783
rect 5350 6780 5356 6792
rect 5215 6752 5356 6780
rect 5215 6749 5227 6752
rect 5169 6743 5227 6749
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 5644 6789 5672 6820
rect 5445 6783 5503 6789
rect 5445 6749 5457 6783
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6749 5687 6783
rect 5629 6743 5687 6749
rect 1670 6721 1676 6724
rect 1664 6675 1676 6721
rect 1670 6672 1676 6675
rect 1728 6672 1734 6724
rect 4706 6672 4712 6724
rect 4764 6712 4770 6724
rect 5077 6715 5135 6721
rect 5077 6712 5089 6715
rect 4764 6684 5089 6712
rect 4764 6672 4770 6684
rect 5077 6681 5089 6684
rect 5123 6681 5135 6715
rect 5460 6712 5488 6743
rect 5902 6740 5908 6792
rect 5960 6740 5966 6792
rect 6012 6780 6040 6820
rect 6089 6817 6101 6851
rect 6135 6848 6147 6851
rect 6362 6848 6368 6860
rect 6135 6820 6368 6848
rect 6135 6817 6147 6820
rect 6089 6811 6147 6817
rect 6362 6808 6368 6820
rect 6420 6808 6426 6860
rect 7009 6851 7067 6857
rect 7009 6817 7021 6851
rect 7055 6848 7067 6851
rect 7190 6848 7196 6860
rect 7055 6820 7196 6848
rect 7055 6817 7067 6820
rect 7009 6811 7067 6817
rect 7190 6808 7196 6820
rect 7248 6808 7254 6860
rect 7300 6820 7604 6848
rect 7300 6792 7328 6820
rect 7576 6792 7604 6820
rect 7282 6780 7288 6792
rect 6012 6752 7288 6780
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6749 7435 6783
rect 7377 6743 7435 6749
rect 6270 6712 6276 6724
rect 5460 6684 6276 6712
rect 5077 6675 5135 6681
rect 6270 6672 6276 6684
rect 6328 6672 6334 6724
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 7392 6712 7420 6743
rect 7558 6740 7564 6792
rect 7616 6740 7622 6792
rect 7668 6789 7696 6888
rect 7929 6919 7987 6925
rect 7929 6885 7941 6919
rect 7975 6885 7987 6919
rect 7929 6879 7987 6885
rect 7944 6848 7972 6879
rect 8386 6876 8392 6928
rect 8444 6876 8450 6928
rect 9398 6876 9404 6928
rect 9456 6876 9462 6928
rect 11164 6916 11192 6944
rect 12452 6916 12480 6947
rect 11164 6888 12480 6916
rect 9033 6851 9091 6857
rect 9033 6848 9045 6851
rect 7944 6820 9045 6848
rect 9033 6817 9045 6820
rect 9079 6848 9091 6851
rect 9861 6851 9919 6857
rect 9079 6820 9674 6848
rect 9079 6817 9091 6820
rect 9033 6811 9091 6817
rect 7653 6783 7711 6789
rect 7653 6749 7665 6783
rect 7699 6749 7711 6783
rect 7653 6743 7711 6749
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6780 7803 6783
rect 7834 6780 7840 6792
rect 7791 6752 7840 6780
rect 7791 6749 7803 6752
rect 7745 6743 7803 6749
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 8018 6740 8024 6792
rect 8076 6740 8082 6792
rect 8297 6783 8355 6789
rect 8297 6780 8309 6783
rect 8128 6752 8309 6780
rect 7248 6684 7420 6712
rect 7248 6672 7254 6684
rect 5353 6647 5411 6653
rect 5353 6613 5365 6647
rect 5399 6644 5411 6647
rect 5626 6644 5632 6656
rect 5399 6616 5632 6644
rect 5399 6613 5411 6616
rect 5353 6607 5411 6613
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 7392 6644 7420 6684
rect 7926 6672 7932 6724
rect 7984 6712 7990 6724
rect 8128 6712 8156 6752
rect 8297 6749 8309 6752
rect 8343 6749 8355 6783
rect 8297 6743 8355 6749
rect 8386 6740 8392 6792
rect 8444 6740 8450 6792
rect 8846 6740 8852 6792
rect 8904 6780 8910 6792
rect 9217 6783 9275 6789
rect 9217 6780 9229 6783
rect 8904 6752 9229 6780
rect 8904 6740 8910 6752
rect 9217 6749 9229 6752
rect 9263 6749 9275 6783
rect 9646 6780 9674 6820
rect 9861 6817 9873 6851
rect 9907 6848 9919 6851
rect 10134 6848 10140 6860
rect 9907 6820 10140 6848
rect 9907 6817 9919 6820
rect 9861 6811 9919 6817
rect 10134 6808 10140 6820
rect 10192 6848 10198 6860
rect 10962 6848 10968 6860
rect 10192 6820 10968 6848
rect 10192 6808 10198 6820
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 11238 6808 11244 6860
rect 11296 6808 11302 6860
rect 12250 6808 12256 6860
rect 12308 6848 12314 6860
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 12308 6820 12541 6848
rect 12308 6808 12314 6820
rect 12529 6817 12541 6820
rect 12575 6817 12587 6851
rect 12529 6811 12587 6817
rect 12894 6808 12900 6860
rect 12952 6848 12958 6860
rect 13081 6851 13139 6857
rect 13081 6848 13093 6851
rect 12952 6820 13093 6848
rect 12952 6808 12958 6820
rect 13081 6817 13093 6820
rect 13127 6817 13139 6851
rect 13081 6811 13139 6817
rect 13170 6808 13176 6860
rect 13228 6808 13234 6860
rect 13280 6857 13308 6956
rect 14090 6944 14096 6996
rect 14148 6984 14154 6996
rect 14369 6987 14427 6993
rect 14369 6984 14381 6987
rect 14148 6956 14381 6984
rect 14148 6944 14154 6956
rect 14369 6953 14381 6956
rect 14415 6953 14427 6987
rect 14369 6947 14427 6953
rect 14829 6987 14887 6993
rect 14829 6953 14841 6987
rect 14875 6984 14887 6987
rect 15010 6984 15016 6996
rect 14875 6956 15016 6984
rect 14875 6953 14887 6956
rect 14829 6947 14887 6953
rect 15010 6944 15016 6956
rect 15068 6944 15074 6996
rect 13265 6851 13323 6857
rect 13265 6817 13277 6851
rect 13311 6848 13323 6851
rect 13906 6848 13912 6860
rect 13311 6820 13912 6848
rect 13311 6817 13323 6820
rect 13265 6811 13323 6817
rect 13906 6808 13912 6820
rect 13964 6808 13970 6860
rect 11330 6780 11336 6792
rect 9646 6752 11336 6780
rect 9217 6743 9275 6749
rect 11330 6740 11336 6752
rect 11388 6740 11394 6792
rect 11422 6740 11428 6792
rect 11480 6740 11486 6792
rect 12713 6783 12771 6789
rect 12713 6749 12725 6783
rect 12759 6749 12771 6783
rect 14553 6783 14611 6789
rect 14553 6780 14565 6783
rect 12452 6724 12572 6746
rect 12713 6743 12771 6749
rect 13280 6752 14565 6780
rect 7984 6684 8156 6712
rect 8205 6715 8263 6721
rect 7984 6672 7990 6684
rect 8205 6681 8217 6715
rect 8251 6681 8263 6715
rect 8205 6675 8263 6681
rect 8220 6644 8248 6675
rect 8938 6672 8944 6724
rect 8996 6672 9002 6724
rect 9493 6715 9551 6721
rect 9493 6681 9505 6715
rect 9539 6712 9551 6715
rect 9582 6712 9588 6724
rect 9539 6684 9588 6712
rect 9539 6681 9551 6684
rect 9493 6675 9551 6681
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 9677 6715 9735 6721
rect 9677 6681 9689 6715
rect 9723 6712 9735 6715
rect 9766 6712 9772 6724
rect 9723 6684 9772 6712
rect 9723 6681 9735 6684
rect 9677 6675 9735 6681
rect 9766 6672 9772 6684
rect 9824 6672 9830 6724
rect 11146 6672 11152 6724
rect 11204 6672 11210 6724
rect 12452 6721 12532 6724
rect 12437 6718 12532 6721
rect 12437 6715 12495 6718
rect 12437 6681 12449 6715
rect 12483 6681 12495 6715
rect 12437 6675 12495 6681
rect 12526 6672 12532 6718
rect 12584 6672 12590 6724
rect 12618 6672 12624 6724
rect 12676 6712 12682 6724
rect 12728 6712 12756 6743
rect 12676 6684 12756 6712
rect 12820 6684 13032 6712
rect 12676 6672 12682 6684
rect 7392 6616 8248 6644
rect 8573 6647 8631 6653
rect 8573 6613 8585 6647
rect 8619 6644 8631 6647
rect 9858 6644 9864 6656
rect 8619 6616 9864 6644
rect 8619 6613 8631 6616
rect 8573 6607 8631 6613
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 12158 6604 12164 6656
rect 12216 6644 12222 6656
rect 12820 6644 12848 6684
rect 12216 6616 12848 6644
rect 13004 6644 13032 6684
rect 13280 6644 13308 6752
rect 14553 6749 14565 6752
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 14645 6783 14703 6789
rect 14645 6749 14657 6783
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 13449 6715 13507 6721
rect 13449 6681 13461 6715
rect 13495 6712 13507 6715
rect 13630 6712 13636 6724
rect 13495 6684 13636 6712
rect 13495 6681 13507 6684
rect 13449 6675 13507 6681
rect 13630 6672 13636 6684
rect 13688 6672 13694 6724
rect 14366 6672 14372 6724
rect 14424 6672 14430 6724
rect 13004 6616 13308 6644
rect 12216 6604 12222 6616
rect 13354 6604 13360 6656
rect 13412 6604 13418 6656
rect 13814 6604 13820 6656
rect 13872 6644 13878 6656
rect 14182 6644 14188 6656
rect 13872 6616 14188 6644
rect 13872 6604 13878 6616
rect 14182 6604 14188 6616
rect 14240 6644 14246 6656
rect 14660 6644 14688 6743
rect 15654 6740 15660 6792
rect 15712 6740 15718 6792
rect 15746 6672 15752 6724
rect 15804 6712 15810 6724
rect 15902 6715 15960 6721
rect 15902 6712 15914 6715
rect 15804 6684 15914 6712
rect 15804 6672 15810 6684
rect 15902 6681 15914 6684
rect 15948 6681 15960 6715
rect 15902 6675 15960 6681
rect 14240 6616 14688 6644
rect 14240 6604 14246 6616
rect 16482 6604 16488 6656
rect 16540 6644 16546 6656
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 16540 6616 17049 6644
rect 16540 6604 16546 6616
rect 17037 6613 17049 6616
rect 17083 6613 17095 6647
rect 17037 6607 17095 6613
rect 1104 6554 17388 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 17388 6554
rect 1104 6480 17388 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1670 6440 1676 6452
rect 1627 6412 1676 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 3786 6400 3792 6452
rect 3844 6440 3850 6452
rect 4249 6443 4307 6449
rect 4249 6440 4261 6443
rect 3844 6412 4261 6440
rect 3844 6400 3850 6412
rect 4249 6409 4261 6412
rect 4295 6409 4307 6443
rect 4249 6403 4307 6409
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 7742 6440 7748 6452
rect 6328 6412 7748 6440
rect 6328 6400 6334 6412
rect 7742 6400 7748 6412
rect 7800 6400 7806 6452
rect 7929 6443 7987 6449
rect 7929 6409 7941 6443
rect 7975 6440 7987 6443
rect 8846 6440 8852 6452
rect 7975 6412 8852 6440
rect 7975 6409 7987 6412
rect 7929 6403 7987 6409
rect 8846 6400 8852 6412
rect 8904 6400 8910 6452
rect 8938 6400 8944 6452
rect 8996 6440 9002 6452
rect 9306 6440 9312 6452
rect 8996 6412 9312 6440
rect 8996 6400 9002 6412
rect 9306 6400 9312 6412
rect 9364 6440 9370 6452
rect 9582 6440 9588 6452
rect 9364 6412 9588 6440
rect 9364 6400 9370 6412
rect 9582 6400 9588 6412
rect 9640 6400 9646 6452
rect 11330 6400 11336 6452
rect 11388 6440 11394 6452
rect 12618 6440 12624 6452
rect 11388 6412 12624 6440
rect 11388 6400 11394 6412
rect 12618 6400 12624 6412
rect 12676 6400 12682 6452
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 13630 6440 13636 6452
rect 12768 6412 13636 6440
rect 12768 6400 12774 6412
rect 13630 6400 13636 6412
rect 13688 6400 13694 6452
rect 13722 6400 13728 6452
rect 13780 6400 13786 6452
rect 15470 6440 15476 6452
rect 15396 6412 15476 6440
rect 3694 6372 3700 6384
rect 3068 6344 3700 6372
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 900 6276 1409 6304
rect 900 6264 906 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 1854 6264 1860 6316
rect 1912 6264 1918 6316
rect 3068 6313 3096 6344
rect 3694 6332 3700 6344
rect 3752 6372 3758 6384
rect 3752 6344 4200 6372
rect 3752 6332 3758 6344
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6273 3111 6307
rect 3053 6267 3111 6273
rect 3329 6307 3387 6313
rect 3329 6273 3341 6307
rect 3375 6304 3387 6307
rect 3418 6304 3424 6316
rect 3375 6276 3424 6304
rect 3375 6273 3387 6276
rect 3329 6267 3387 6273
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6304 3571 6307
rect 3878 6304 3884 6316
rect 3559 6276 3884 6304
rect 3559 6273 3571 6276
rect 3513 6267 3571 6273
rect 2866 6196 2872 6248
rect 2924 6236 2930 6248
rect 3528 6236 3556 6267
rect 3878 6264 3884 6276
rect 3936 6304 3942 6316
rect 4172 6313 4200 6344
rect 4798 6332 4804 6384
rect 4856 6372 4862 6384
rect 5353 6375 5411 6381
rect 5353 6372 5365 6375
rect 4856 6344 5365 6372
rect 4856 6332 4862 6344
rect 5353 6341 5365 6344
rect 5399 6372 5411 6375
rect 7190 6372 7196 6384
rect 5399 6344 7196 6372
rect 5399 6341 5411 6344
rect 5353 6335 5411 6341
rect 7190 6332 7196 6344
rect 7248 6332 7254 6384
rect 7558 6332 7564 6384
rect 7616 6332 7622 6384
rect 7834 6332 7840 6384
rect 7892 6372 7898 6384
rect 7892 6344 8064 6372
rect 7892 6332 7898 6344
rect 4065 6307 4123 6313
rect 4065 6304 4077 6307
rect 3936 6276 4077 6304
rect 3936 6264 3942 6276
rect 4065 6273 4077 6276
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6273 4215 6307
rect 4157 6267 4215 6273
rect 4614 6264 4620 6316
rect 4672 6264 4678 6316
rect 4706 6264 4712 6316
rect 4764 6304 4770 6316
rect 5077 6307 5135 6313
rect 5077 6304 5089 6307
rect 4764 6276 5089 6304
rect 4764 6264 4770 6276
rect 5077 6273 5089 6276
rect 5123 6273 5135 6307
rect 5077 6267 5135 6273
rect 2924 6208 3556 6236
rect 2924 6196 2930 6208
rect 3602 6196 3608 6248
rect 3660 6196 3666 6248
rect 3970 6196 3976 6248
rect 4028 6236 4034 6248
rect 4798 6236 4804 6248
rect 4028 6208 4804 6236
rect 4028 6196 4034 6208
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 5092 6236 5120 6267
rect 5258 6264 5264 6316
rect 5316 6264 5322 6316
rect 5442 6264 5448 6316
rect 5500 6313 5506 6316
rect 5500 6304 5508 6313
rect 7098 6304 7104 6316
rect 5500 6276 5545 6304
rect 5644 6276 7104 6304
rect 5500 6267 5508 6276
rect 5500 6264 5506 6267
rect 5644 6236 5672 6276
rect 7098 6264 7104 6276
rect 7156 6304 7162 6316
rect 7423 6310 7481 6313
rect 7300 6307 7481 6310
rect 7300 6304 7435 6307
rect 7156 6282 7435 6304
rect 7156 6276 7328 6282
rect 7412 6276 7435 6282
rect 7156 6264 7162 6276
rect 7423 6273 7435 6276
rect 7469 6273 7481 6307
rect 7423 6267 7481 6273
rect 7649 6307 7707 6313
rect 7649 6273 7661 6307
rect 7695 6273 7707 6307
rect 7649 6270 7707 6273
rect 7576 6267 7707 6270
rect 5092 6208 5672 6236
rect 5994 6196 6000 6248
rect 6052 6236 6058 6248
rect 7282 6236 7288 6248
rect 6052 6208 7288 6236
rect 6052 6196 6058 6208
rect 7282 6196 7288 6208
rect 7340 6196 7346 6248
rect 7576 6242 7696 6267
rect 7742 6264 7748 6316
rect 7800 6264 7806 6316
rect 8036 6313 8064 6344
rect 8754 6332 8760 6384
rect 8812 6372 8818 6384
rect 12066 6372 12072 6384
rect 8812 6344 12072 6372
rect 8812 6332 8818 6344
rect 12066 6332 12072 6344
rect 12124 6332 12130 6384
rect 12986 6332 12992 6384
rect 13044 6372 13050 6384
rect 15396 6381 15424 6412
rect 15470 6400 15476 6412
rect 15528 6400 15534 6452
rect 15746 6400 15752 6452
rect 15804 6400 15810 6452
rect 15381 6375 15439 6381
rect 13044 6344 15240 6372
rect 13044 6332 13050 6344
rect 8021 6307 8079 6313
rect 8021 6273 8033 6307
rect 8067 6273 8079 6307
rect 8021 6267 8079 6273
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 7576 6236 7604 6242
rect 7412 6208 7604 6236
rect 7760 6236 7788 6264
rect 7834 6236 7840 6248
rect 7760 6208 7840 6236
rect 3786 6128 3792 6180
rect 3844 6168 3850 6180
rect 3881 6171 3939 6177
rect 3881 6168 3893 6171
rect 3844 6140 3893 6168
rect 3844 6128 3850 6140
rect 3881 6137 3893 6140
rect 3927 6137 3939 6171
rect 3881 6131 3939 6137
rect 7190 6128 7196 6180
rect 7248 6168 7254 6180
rect 7412 6168 7440 6208
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 7248 6140 7440 6168
rect 7248 6128 7254 6140
rect 7558 6128 7564 6180
rect 7616 6168 7622 6180
rect 8220 6168 8248 6267
rect 8294 6264 8300 6316
rect 8352 6264 8358 6316
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6304 8447 6307
rect 8478 6304 8484 6316
rect 8435 6276 8484 6304
rect 8435 6273 8447 6276
rect 8389 6267 8447 6273
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 9306 6264 9312 6316
rect 9364 6264 9370 6316
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6304 9551 6307
rect 9858 6304 9864 6316
rect 9539 6276 9864 6304
rect 9539 6273 9551 6276
rect 9493 6267 9551 6273
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 13354 6304 13360 6316
rect 10100 6276 13360 6304
rect 10100 6264 10106 6276
rect 13354 6264 13360 6276
rect 13412 6264 13418 6316
rect 13630 6264 13636 6316
rect 13688 6264 13694 6316
rect 15212 6313 15240 6344
rect 15381 6341 15393 6375
rect 15427 6341 15439 6375
rect 15381 6335 15439 6341
rect 13909 6307 13967 6313
rect 13909 6273 13921 6307
rect 13955 6273 13967 6307
rect 13909 6267 13967 6273
rect 14093 6307 14151 6313
rect 14093 6273 14105 6307
rect 14139 6273 14151 6307
rect 14093 6267 14151 6273
rect 15197 6307 15255 6313
rect 15197 6273 15209 6307
rect 15243 6273 15255 6307
rect 15197 6267 15255 6273
rect 8846 6196 8852 6248
rect 8904 6236 8910 6248
rect 13449 6239 13507 6245
rect 13449 6236 13461 6239
rect 8904 6208 13461 6236
rect 8904 6196 8910 6208
rect 13449 6205 13461 6208
rect 13495 6236 13507 6239
rect 13924 6236 13952 6267
rect 13495 6208 13952 6236
rect 13495 6205 13507 6208
rect 13449 6199 13507 6205
rect 7616 6140 8248 6168
rect 8573 6171 8631 6177
rect 7616 6128 7622 6140
rect 8573 6137 8585 6171
rect 8619 6168 8631 6171
rect 10042 6168 10048 6180
rect 8619 6140 10048 6168
rect 8619 6137 8631 6140
rect 8573 6131 8631 6137
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 11422 6128 11428 6180
rect 11480 6168 11486 6180
rect 12894 6168 12900 6180
rect 11480 6140 12900 6168
rect 11480 6128 11486 6140
rect 12894 6128 12900 6140
rect 12952 6168 12958 6180
rect 13173 6171 13231 6177
rect 13173 6168 13185 6171
rect 12952 6140 13185 6168
rect 12952 6128 12958 6140
rect 13173 6137 13185 6140
rect 13219 6137 13231 6171
rect 13173 6131 13231 6137
rect 13722 6128 13728 6180
rect 13780 6168 13786 6180
rect 14108 6168 14136 6267
rect 15286 6264 15292 6316
rect 15344 6304 15350 6316
rect 15473 6307 15531 6313
rect 15473 6304 15485 6307
rect 15344 6276 15485 6304
rect 15344 6264 15350 6276
rect 15473 6273 15485 6276
rect 15519 6273 15531 6307
rect 15473 6267 15531 6273
rect 15565 6307 15623 6313
rect 15565 6273 15577 6307
rect 15611 6304 15623 6307
rect 15841 6307 15899 6313
rect 15841 6304 15853 6307
rect 15611 6276 15853 6304
rect 15611 6273 15623 6276
rect 15565 6267 15623 6273
rect 15841 6273 15853 6276
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 16482 6264 16488 6316
rect 16540 6264 16546 6316
rect 16758 6264 16764 6316
rect 16816 6264 16822 6316
rect 13780 6140 14136 6168
rect 13780 6128 13786 6140
rect 16942 6128 16948 6180
rect 17000 6128 17006 6180
rect 1670 6060 1676 6112
rect 1728 6060 1734 6112
rect 5077 6103 5135 6109
rect 5077 6069 5089 6103
rect 5123 6100 5135 6103
rect 6362 6100 6368 6112
rect 5123 6072 6368 6100
rect 5123 6069 5135 6072
rect 5077 6063 5135 6069
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 7466 6100 7472 6112
rect 7340 6072 7472 6100
rect 7340 6060 7346 6072
rect 7466 6060 7472 6072
rect 7524 6100 7530 6112
rect 8386 6100 8392 6112
rect 7524 6072 8392 6100
rect 7524 6060 7530 6072
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 8662 6060 8668 6112
rect 8720 6100 8726 6112
rect 9309 6103 9367 6109
rect 9309 6100 9321 6103
rect 8720 6072 9321 6100
rect 8720 6060 8726 6072
rect 9309 6069 9321 6072
rect 9355 6069 9367 6103
rect 9309 6063 9367 6069
rect 9677 6103 9735 6109
rect 9677 6069 9689 6103
rect 9723 6100 9735 6103
rect 11606 6100 11612 6112
rect 9723 6072 11612 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 13630 6060 13636 6112
rect 13688 6060 13694 6112
rect 1104 6010 17388 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 17388 6010
rect 1104 5936 17388 5958
rect 2774 5856 2780 5908
rect 2832 5856 2838 5908
rect 4433 5899 4491 5905
rect 4433 5865 4445 5899
rect 4479 5896 4491 5899
rect 4706 5896 4712 5908
rect 4479 5868 4712 5896
rect 4479 5865 4491 5868
rect 4433 5859 4491 5865
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 7374 5896 7380 5908
rect 5465 5868 7380 5896
rect 3602 5788 3608 5840
rect 3660 5828 3666 5840
rect 5465 5828 5493 5868
rect 7374 5856 7380 5868
rect 7432 5896 7438 5908
rect 8294 5896 8300 5908
rect 7432 5868 8300 5896
rect 7432 5856 7438 5868
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 8478 5856 8484 5908
rect 8536 5856 8542 5908
rect 9030 5856 9036 5908
rect 9088 5896 9094 5908
rect 9582 5896 9588 5908
rect 9088 5868 9588 5896
rect 9088 5856 9094 5868
rect 9582 5856 9588 5868
rect 9640 5856 9646 5908
rect 10594 5856 10600 5908
rect 10652 5856 10658 5908
rect 11606 5856 11612 5908
rect 11664 5896 11670 5908
rect 12342 5896 12348 5908
rect 11664 5868 12348 5896
rect 11664 5856 11670 5868
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 13722 5856 13728 5908
rect 13780 5896 13786 5908
rect 14093 5899 14151 5905
rect 14093 5896 14105 5899
rect 13780 5868 14105 5896
rect 13780 5856 13786 5868
rect 14093 5865 14105 5868
rect 14139 5865 14151 5899
rect 14093 5859 14151 5865
rect 14458 5856 14464 5908
rect 14516 5896 14522 5908
rect 14553 5899 14611 5905
rect 14553 5896 14565 5899
rect 14516 5868 14565 5896
rect 14516 5856 14522 5868
rect 14553 5865 14565 5868
rect 14599 5865 14611 5899
rect 14553 5859 14611 5865
rect 16850 5856 16856 5908
rect 16908 5896 16914 5908
rect 17037 5899 17095 5905
rect 17037 5896 17049 5899
rect 16908 5868 17049 5896
rect 16908 5856 16914 5868
rect 17037 5865 17049 5868
rect 17083 5865 17095 5899
rect 17037 5859 17095 5865
rect 3660 5800 5493 5828
rect 3660 5788 3666 5800
rect 3786 5720 3792 5772
rect 3844 5760 3850 5772
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 3844 5732 4261 5760
rect 3844 5720 3850 5732
rect 4249 5729 4261 5732
rect 4295 5729 4307 5763
rect 4249 5723 4307 5729
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 1670 5701 1676 5704
rect 1664 5692 1676 5701
rect 1631 5664 1676 5692
rect 1664 5655 1676 5664
rect 1670 5652 1676 5655
rect 1728 5652 1734 5704
rect 3418 5652 3424 5704
rect 3476 5692 3482 5704
rect 3970 5692 3976 5704
rect 3476 5664 3976 5692
rect 3476 5652 3482 5664
rect 3970 5652 3976 5664
rect 4028 5692 4034 5704
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 4028 5664 4077 5692
rect 4028 5652 4034 5664
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 5465 5692 5493 5800
rect 5718 5788 5724 5840
rect 5776 5828 5782 5840
rect 6638 5828 6644 5840
rect 5776 5800 6644 5828
rect 5776 5788 5782 5800
rect 6638 5788 6644 5800
rect 6696 5828 6702 5840
rect 7469 5831 7527 5837
rect 6696 5800 6960 5828
rect 6696 5788 6702 5800
rect 5813 5763 5871 5769
rect 5813 5729 5825 5763
rect 5859 5760 5871 5763
rect 6181 5763 6239 5769
rect 5859 5732 6132 5760
rect 5859 5729 5871 5732
rect 5813 5723 5871 5729
rect 5537 5695 5595 5701
rect 5537 5692 5549 5695
rect 5465 5664 5549 5692
rect 4065 5655 4123 5661
rect 5537 5661 5549 5664
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 5626 5652 5632 5704
rect 5684 5692 5690 5704
rect 6104 5701 6132 5732
rect 6181 5729 6193 5763
rect 6227 5760 6239 5763
rect 6454 5760 6460 5772
rect 6227 5732 6460 5760
rect 6227 5729 6239 5732
rect 6181 5723 6239 5729
rect 6454 5720 6460 5732
rect 6512 5720 6518 5772
rect 6270 5701 6276 5704
rect 5910 5695 5968 5701
rect 5910 5692 5922 5695
rect 5684 5664 5922 5692
rect 5684 5652 5690 5664
rect 5910 5661 5922 5664
rect 5956 5661 5968 5695
rect 5910 5655 5968 5661
rect 6089 5695 6147 5701
rect 6089 5661 6101 5695
rect 6135 5661 6147 5695
rect 6266 5692 6276 5701
rect 6231 5664 6276 5692
rect 6089 5655 6147 5661
rect 6266 5655 6276 5664
rect 6270 5652 6276 5655
rect 6328 5652 6334 5704
rect 6362 5652 6368 5704
rect 6420 5652 6426 5704
rect 6546 5652 6552 5704
rect 6604 5652 6610 5704
rect 6932 5692 6960 5800
rect 7469 5797 7481 5831
rect 7515 5828 7527 5831
rect 7558 5828 7564 5840
rect 7515 5800 7564 5828
rect 7515 5797 7527 5800
rect 7469 5791 7527 5797
rect 7558 5788 7564 5800
rect 7616 5788 7622 5840
rect 7834 5788 7840 5840
rect 7892 5828 7898 5840
rect 8496 5828 8524 5856
rect 7892 5800 8524 5828
rect 7892 5788 7898 5800
rect 7374 5720 7380 5772
rect 7432 5760 7438 5772
rect 7576 5760 7604 5788
rect 7432 5732 7880 5760
rect 7432 5720 7438 5732
rect 7285 5695 7343 5701
rect 7285 5692 7297 5695
rect 6932 5664 7297 5692
rect 7285 5661 7297 5664
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 7650 5652 7656 5704
rect 7708 5652 7714 5704
rect 7852 5701 7880 5732
rect 7837 5695 7895 5701
rect 7837 5661 7849 5695
rect 7883 5661 7895 5695
rect 7944 5692 7972 5800
rect 9398 5788 9404 5840
rect 9456 5828 9462 5840
rect 9456 5800 11468 5828
rect 9456 5788 9462 5800
rect 11440 5769 11468 5800
rect 15286 5788 15292 5840
rect 15344 5828 15350 5840
rect 15344 5800 15608 5828
rect 15344 5788 15350 5800
rect 11425 5763 11483 5769
rect 9646 5732 11376 5760
rect 8021 5695 8079 5701
rect 8021 5692 8033 5695
rect 7944 5664 8033 5692
rect 7837 5655 7895 5661
rect 8021 5661 8033 5664
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 8202 5652 8208 5704
rect 8260 5652 8266 5704
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5692 8355 5695
rect 8386 5692 8392 5704
rect 8343 5664 8392 5692
rect 8343 5661 8355 5664
rect 8297 5655 8355 5661
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 9306 5652 9312 5704
rect 9364 5652 9370 5704
rect 3326 5584 3332 5636
rect 3384 5624 3390 5636
rect 3789 5627 3847 5633
rect 3789 5624 3801 5627
rect 3384 5596 3801 5624
rect 3384 5584 3390 5596
rect 3789 5593 3801 5596
rect 3835 5624 3847 5627
rect 3878 5624 3884 5636
rect 3835 5596 3884 5624
rect 3835 5593 3847 5596
rect 3789 5587 3847 5593
rect 3878 5584 3884 5596
rect 3936 5584 3942 5636
rect 5718 5584 5724 5636
rect 5776 5584 5782 5636
rect 5813 5627 5871 5633
rect 5813 5593 5825 5627
rect 5859 5593 5871 5627
rect 6730 5624 6736 5636
rect 5813 5587 5871 5593
rect 6564 5596 6736 5624
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 4062 5556 4068 5568
rect 3752 5528 4068 5556
rect 3752 5516 3758 5528
rect 4062 5516 4068 5528
rect 4120 5556 4126 5568
rect 4157 5559 4215 5565
rect 4157 5556 4169 5559
rect 4120 5528 4169 5556
rect 4120 5516 4126 5528
rect 4157 5525 4169 5528
rect 4203 5525 4215 5559
rect 4157 5519 4215 5525
rect 4614 5516 4620 5568
rect 4672 5556 4678 5568
rect 5828 5556 5856 5587
rect 6086 5556 6092 5568
rect 4672 5528 6092 5556
rect 4672 5516 4678 5528
rect 6086 5516 6092 5528
rect 6144 5516 6150 5568
rect 6564 5565 6592 5596
rect 6730 5584 6736 5596
rect 6788 5584 6794 5636
rect 7098 5584 7104 5636
rect 7156 5584 7162 5636
rect 7929 5627 7987 5633
rect 7929 5593 7941 5627
rect 7975 5624 7987 5627
rect 8220 5624 8248 5652
rect 9646 5624 9674 5732
rect 10045 5695 10103 5701
rect 10045 5661 10057 5695
rect 10091 5692 10103 5695
rect 10410 5692 10416 5704
rect 10091 5664 10416 5692
rect 10091 5661 10103 5664
rect 10045 5655 10103 5661
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 10689 5695 10747 5701
rect 10689 5661 10701 5695
rect 10735 5661 10747 5695
rect 10689 5655 10747 5661
rect 10781 5695 10839 5701
rect 10781 5661 10793 5695
rect 10827 5692 10839 5695
rect 10870 5692 10876 5704
rect 10827 5664 10876 5692
rect 10827 5661 10839 5664
rect 10781 5655 10839 5661
rect 7975 5596 8248 5624
rect 8312 5596 9674 5624
rect 7975 5593 7987 5596
rect 7929 5587 7987 5593
rect 6549 5559 6607 5565
rect 6549 5525 6561 5559
rect 6595 5525 6607 5559
rect 6549 5519 6607 5525
rect 7009 5559 7067 5565
rect 7009 5525 7021 5559
rect 7055 5556 7067 5559
rect 7944 5556 7972 5587
rect 7055 5528 7972 5556
rect 8205 5559 8263 5565
rect 7055 5525 7067 5528
rect 7009 5519 7067 5525
rect 8205 5525 8217 5559
rect 8251 5556 8263 5559
rect 8312 5556 8340 5596
rect 10226 5584 10232 5636
rect 10284 5584 10290 5636
rect 10502 5584 10508 5636
rect 10560 5584 10566 5636
rect 10704 5624 10732 5655
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 11348 5692 11376 5732
rect 11425 5729 11437 5763
rect 11471 5729 11483 5763
rect 11425 5723 11483 5729
rect 12342 5720 12348 5772
rect 12400 5760 12406 5772
rect 12400 5732 13676 5760
rect 12400 5720 12406 5732
rect 13648 5704 13676 5732
rect 14182 5720 14188 5772
rect 14240 5720 14246 5772
rect 15470 5760 15476 5772
rect 15212 5732 15476 5760
rect 11348 5664 11468 5692
rect 11054 5624 11060 5636
rect 10704 5596 11060 5624
rect 11054 5584 11060 5596
rect 11112 5584 11118 5636
rect 11333 5627 11391 5633
rect 11333 5593 11345 5627
rect 11379 5593 11391 5627
rect 11440 5624 11468 5664
rect 11514 5652 11520 5704
rect 11572 5692 11578 5704
rect 11609 5695 11667 5701
rect 11609 5692 11621 5695
rect 11572 5664 11621 5692
rect 11572 5652 11578 5664
rect 11609 5661 11621 5664
rect 11655 5661 11667 5695
rect 11609 5655 11667 5661
rect 13538 5652 13544 5704
rect 13596 5652 13602 5704
rect 13630 5652 13636 5704
rect 13688 5692 13694 5704
rect 15212 5701 15240 5732
rect 15470 5720 15476 5732
rect 15528 5720 15534 5772
rect 14369 5695 14427 5701
rect 14369 5692 14381 5695
rect 13688 5664 14381 5692
rect 13688 5652 13694 5664
rect 14369 5661 14381 5664
rect 14415 5661 14427 5695
rect 14369 5655 14427 5661
rect 15013 5695 15071 5701
rect 15013 5661 15025 5695
rect 15059 5661 15071 5695
rect 15013 5655 15071 5661
rect 15197 5695 15255 5701
rect 15197 5661 15209 5695
rect 15243 5661 15255 5695
rect 15197 5655 15255 5661
rect 15381 5695 15439 5701
rect 15381 5661 15393 5695
rect 15427 5692 15439 5695
rect 15580 5692 15608 5800
rect 15427 5664 15608 5692
rect 15427 5661 15439 5664
rect 15381 5655 15439 5661
rect 12618 5624 12624 5636
rect 11440 5596 12624 5624
rect 11333 5587 11391 5593
rect 8251 5528 8340 5556
rect 8251 5525 8263 5528
rect 8205 5519 8263 5525
rect 9030 5516 9036 5568
rect 9088 5556 9094 5568
rect 9493 5559 9551 5565
rect 9493 5556 9505 5559
rect 9088 5528 9505 5556
rect 9088 5516 9094 5528
rect 9493 5525 9505 5528
rect 9539 5525 9551 5559
rect 9493 5519 9551 5525
rect 10413 5559 10471 5565
rect 10413 5525 10425 5559
rect 10459 5556 10471 5559
rect 10594 5556 10600 5568
rect 10459 5528 10600 5556
rect 10459 5525 10471 5528
rect 10413 5519 10471 5525
rect 10594 5516 10600 5528
rect 10652 5516 10658 5568
rect 10965 5559 11023 5565
rect 10965 5525 10977 5559
rect 11011 5556 11023 5559
rect 11348 5556 11376 5587
rect 12618 5584 12624 5596
rect 12676 5584 12682 5636
rect 13354 5584 13360 5636
rect 13412 5624 13418 5636
rect 13725 5627 13783 5633
rect 13725 5624 13737 5627
rect 13412 5596 13737 5624
rect 13412 5584 13418 5596
rect 13725 5593 13737 5596
rect 13771 5593 13783 5627
rect 13725 5587 13783 5593
rect 13909 5627 13967 5633
rect 13909 5593 13921 5627
rect 13955 5624 13967 5627
rect 14090 5624 14096 5636
rect 13955 5596 14096 5624
rect 13955 5593 13967 5596
rect 13909 5587 13967 5593
rect 14090 5584 14096 5596
rect 14148 5584 14154 5636
rect 15028 5624 15056 5655
rect 15654 5652 15660 5704
rect 15712 5652 15718 5704
rect 14200 5596 15056 5624
rect 11011 5528 11376 5556
rect 11793 5559 11851 5565
rect 11011 5525 11023 5528
rect 10965 5519 11023 5525
rect 11793 5525 11805 5559
rect 11839 5556 11851 5559
rect 14200 5556 14228 5596
rect 15286 5584 15292 5636
rect 15344 5584 15350 5636
rect 15902 5627 15960 5633
rect 15902 5624 15914 5627
rect 15580 5596 15914 5624
rect 15580 5565 15608 5596
rect 15902 5593 15914 5596
rect 15948 5593 15960 5627
rect 15902 5587 15960 5593
rect 11839 5528 14228 5556
rect 15565 5559 15623 5565
rect 11839 5525 11851 5528
rect 11793 5519 11851 5525
rect 15565 5525 15577 5559
rect 15611 5525 15623 5559
rect 15565 5519 15623 5525
rect 1104 5466 17388 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 17388 5466
rect 1104 5392 17388 5414
rect 2777 5355 2835 5361
rect 2777 5321 2789 5355
rect 2823 5352 2835 5355
rect 3050 5352 3056 5364
rect 2823 5324 3056 5352
rect 2823 5321 2835 5324
rect 2777 5315 2835 5321
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 3237 5355 3295 5361
rect 3237 5321 3249 5355
rect 3283 5352 3295 5355
rect 3283 5324 8616 5352
rect 3283 5321 3295 5324
rect 3237 5315 3295 5321
rect 2961 5287 3019 5293
rect 2961 5253 2973 5287
rect 3007 5284 3019 5287
rect 3786 5284 3792 5296
rect 3007 5256 3792 5284
rect 3007 5253 3019 5256
rect 2961 5247 3019 5253
rect 1486 5176 1492 5228
rect 1544 5216 1550 5228
rect 1653 5219 1711 5225
rect 1653 5216 1665 5219
rect 1544 5188 1665 5216
rect 1544 5176 1550 5188
rect 1653 5185 1665 5188
rect 1699 5185 1711 5219
rect 1653 5179 1711 5185
rect 3326 5176 3332 5228
rect 3384 5176 3390 5228
rect 3620 5225 3648 5256
rect 3786 5244 3792 5256
rect 3844 5244 3850 5296
rect 5537 5287 5595 5293
rect 5537 5284 5549 5287
rect 4172 5256 5549 5284
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5185 3663 5219
rect 3605 5179 3663 5185
rect 1394 5108 1400 5160
rect 1452 5108 1458 5160
rect 3145 5151 3203 5157
rect 3145 5117 3157 5151
rect 3191 5148 3203 5151
rect 3418 5148 3424 5160
rect 3191 5120 3424 5148
rect 3191 5117 3203 5120
rect 3145 5111 3203 5117
rect 3418 5108 3424 5120
rect 3476 5108 3482 5160
rect 3620 5148 3648 5179
rect 3694 5176 3700 5228
rect 3752 5176 3758 5228
rect 3970 5176 3976 5228
rect 4028 5176 4034 5228
rect 4172 5225 4200 5256
rect 5537 5253 5549 5256
rect 5583 5284 5595 5287
rect 5583 5256 6776 5284
rect 5583 5253 5595 5256
rect 5537 5247 5595 5253
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 4246 5176 4252 5228
rect 4304 5216 4310 5228
rect 4709 5219 4767 5225
rect 4709 5216 4721 5219
rect 4304 5188 4721 5216
rect 4304 5176 4310 5188
rect 4709 5185 4721 5188
rect 4755 5185 4767 5219
rect 4709 5179 4767 5185
rect 4798 5176 4804 5228
rect 4856 5176 4862 5228
rect 4890 5176 4896 5228
rect 4948 5176 4954 5228
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5216 5135 5219
rect 5166 5216 5172 5228
rect 5123 5188 5172 5216
rect 5123 5185 5135 5188
rect 5077 5179 5135 5185
rect 5166 5176 5172 5188
rect 5224 5216 5230 5228
rect 5261 5219 5319 5225
rect 5261 5216 5273 5219
rect 5224 5188 5273 5216
rect 5224 5176 5230 5188
rect 5261 5185 5273 5188
rect 5307 5185 5319 5219
rect 5261 5179 5319 5185
rect 5350 5176 5356 5228
rect 5408 5216 5414 5228
rect 5445 5219 5503 5225
rect 5445 5216 5457 5219
rect 5408 5188 5457 5216
rect 5408 5176 5414 5188
rect 5445 5185 5457 5188
rect 5491 5185 5503 5219
rect 5445 5179 5503 5185
rect 5626 5176 5632 5228
rect 5684 5225 5690 5228
rect 5684 5216 5692 5225
rect 5684 5188 5729 5216
rect 5684 5179 5692 5188
rect 5684 5176 5690 5179
rect 5810 5176 5816 5228
rect 5868 5216 5874 5228
rect 5905 5219 5963 5225
rect 5905 5216 5917 5219
rect 5868 5188 5917 5216
rect 5868 5176 5874 5188
rect 5905 5185 5917 5188
rect 5951 5185 5963 5219
rect 5905 5179 5963 5185
rect 6089 5219 6147 5225
rect 6089 5185 6101 5219
rect 6135 5185 6147 5219
rect 6089 5179 6147 5185
rect 4525 5151 4583 5157
rect 4525 5148 4537 5151
rect 3620 5120 4537 5148
rect 4525 5117 4537 5120
rect 4571 5117 4583 5151
rect 4525 5111 4583 5117
rect 5537 5151 5595 5157
rect 5537 5117 5549 5151
rect 5583 5148 5595 5151
rect 5994 5148 6000 5160
rect 5583 5120 6000 5148
rect 5583 5117 5595 5120
rect 5537 5111 5595 5117
rect 5994 5108 6000 5120
rect 6052 5108 6058 5160
rect 3053 5083 3111 5089
rect 3053 5049 3065 5083
rect 3099 5080 3111 5083
rect 3694 5080 3700 5092
rect 3099 5052 3700 5080
rect 3099 5049 3111 5052
rect 3053 5043 3111 5049
rect 3694 5040 3700 5052
rect 3752 5040 3758 5092
rect 3878 5040 3884 5092
rect 3936 5080 3942 5092
rect 4062 5080 4068 5092
rect 3936 5052 4068 5080
rect 3936 5040 3942 5052
rect 4062 5040 4068 5052
rect 4120 5080 4126 5092
rect 4433 5083 4491 5089
rect 4433 5080 4445 5083
rect 4120 5052 4445 5080
rect 4120 5040 4126 5052
rect 4433 5049 4445 5052
rect 4479 5049 4491 5083
rect 4433 5043 4491 5049
rect 6104 5024 6132 5179
rect 6362 5176 6368 5228
rect 6420 5176 6426 5228
rect 6546 5176 6552 5228
rect 6604 5176 6610 5228
rect 6748 5225 6776 5256
rect 7374 5244 7380 5296
rect 7432 5244 7438 5296
rect 7469 5287 7527 5293
rect 7469 5253 7481 5287
rect 7515 5284 7527 5287
rect 7515 5256 7696 5284
rect 7515 5253 7527 5256
rect 7469 5247 7527 5253
rect 7668 5228 7696 5256
rect 7926 5244 7932 5296
rect 7984 5284 7990 5296
rect 8113 5287 8171 5293
rect 8113 5284 8125 5287
rect 7984 5256 8125 5284
rect 7984 5244 7990 5256
rect 8113 5253 8125 5256
rect 8159 5253 8171 5287
rect 8113 5247 8171 5253
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5216 6791 5219
rect 7098 5216 7104 5228
rect 6779 5188 7104 5216
rect 6779 5185 6791 5188
rect 6733 5179 6791 5185
rect 6454 5108 6460 5160
rect 6512 5148 6518 5160
rect 6656 5148 6684 5179
rect 7098 5176 7104 5188
rect 7156 5216 7162 5228
rect 7193 5219 7251 5225
rect 7193 5216 7205 5219
rect 7156 5188 7205 5216
rect 7156 5176 7162 5188
rect 7193 5185 7205 5188
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 7558 5176 7564 5228
rect 7616 5176 7622 5228
rect 7650 5176 7656 5228
rect 7708 5216 7714 5228
rect 7834 5216 7840 5228
rect 7708 5188 7840 5216
rect 7708 5176 7714 5188
rect 7834 5176 7840 5188
rect 7892 5176 7898 5228
rect 8018 5176 8024 5228
rect 8076 5176 8082 5228
rect 6512 5120 6684 5148
rect 8128 5148 8156 5247
rect 8202 5176 8208 5228
rect 8260 5176 8266 5228
rect 8478 5176 8484 5228
rect 8536 5176 8542 5228
rect 8588 5216 8616 5324
rect 8662 5312 8668 5364
rect 8720 5312 8726 5364
rect 10229 5355 10287 5361
rect 10229 5321 10241 5355
rect 10275 5352 10287 5355
rect 10502 5352 10508 5364
rect 10275 5324 10508 5352
rect 10275 5321 10287 5324
rect 10229 5315 10287 5321
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 11974 5312 11980 5364
rect 12032 5352 12038 5364
rect 12069 5355 12127 5361
rect 12069 5352 12081 5355
rect 12032 5324 12081 5352
rect 12032 5312 12038 5324
rect 12069 5321 12081 5324
rect 12115 5321 12127 5355
rect 12342 5352 12348 5364
rect 12069 5315 12127 5321
rect 12176 5324 12348 5352
rect 10318 5284 10324 5296
rect 8956 5256 9536 5284
rect 8956 5225 8984 5256
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8588 5188 8953 5216
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 9030 5176 9036 5228
rect 9088 5176 9094 5228
rect 9122 5176 9128 5228
rect 9180 5216 9186 5228
rect 9508 5225 9536 5256
rect 9600 5256 10324 5284
rect 9217 5219 9275 5225
rect 9217 5216 9229 5219
rect 9180 5188 9229 5216
rect 9180 5176 9186 5188
rect 9217 5185 9229 5188
rect 9263 5185 9275 5219
rect 9217 5179 9275 5185
rect 9493 5219 9551 5225
rect 9493 5185 9505 5219
rect 9539 5185 9551 5219
rect 9493 5179 9551 5185
rect 9048 5148 9076 5176
rect 8128 5120 9076 5148
rect 6512 5108 6518 5120
rect 7745 5083 7803 5089
rect 7745 5049 7757 5083
rect 7791 5080 7803 5083
rect 8389 5083 8447 5089
rect 7791 5052 8340 5080
rect 7791 5049 7803 5052
rect 7745 5043 7803 5049
rect 6086 4972 6092 5024
rect 6144 4972 6150 5024
rect 6917 5015 6975 5021
rect 6917 4981 6929 5015
rect 6963 5012 6975 5015
rect 8018 5012 8024 5024
rect 6963 4984 8024 5012
rect 6963 4981 6975 4984
rect 6917 4975 6975 4981
rect 8018 4972 8024 4984
rect 8076 4972 8082 5024
rect 8312 5012 8340 5052
rect 8389 5049 8401 5083
rect 8435 5080 8447 5083
rect 9232 5080 9260 5179
rect 9600 5148 9628 5256
rect 10318 5244 10324 5256
rect 10376 5244 10382 5296
rect 12176 5284 12204 5324
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 15286 5312 15292 5364
rect 15344 5352 15350 5364
rect 15841 5355 15899 5361
rect 15841 5352 15853 5355
rect 15344 5324 15853 5352
rect 15344 5312 15350 5324
rect 15841 5321 15853 5324
rect 15887 5321 15899 5355
rect 15841 5315 15899 5321
rect 16942 5312 16948 5364
rect 17000 5312 17006 5364
rect 11716 5256 12204 5284
rect 9674 5176 9680 5228
rect 9732 5176 9738 5228
rect 9766 5176 9772 5228
rect 9824 5176 9830 5228
rect 10045 5219 10103 5225
rect 10045 5185 10057 5219
rect 10091 5216 10103 5219
rect 10134 5216 10140 5228
rect 10091 5188 10140 5216
rect 10091 5185 10103 5188
rect 10045 5179 10103 5185
rect 10134 5176 10140 5188
rect 10192 5176 10198 5228
rect 8435 5052 9260 5080
rect 9324 5120 9628 5148
rect 9692 5148 9720 5176
rect 9953 5151 10011 5157
rect 9953 5148 9965 5151
rect 9692 5120 9965 5148
rect 8435 5049 8447 5052
rect 8389 5043 8447 5049
rect 9324 5012 9352 5120
rect 9953 5117 9965 5120
rect 9999 5148 10011 5151
rect 11716 5148 11744 5256
rect 12250 5244 12256 5296
rect 12308 5244 12314 5296
rect 12360 5256 12572 5284
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 12360 5216 12388 5256
rect 11848 5188 12388 5216
rect 11848 5176 11854 5188
rect 12434 5176 12440 5228
rect 12492 5176 12498 5228
rect 12544 5225 12572 5256
rect 12529 5219 12587 5225
rect 12529 5185 12541 5219
rect 12575 5185 12587 5219
rect 12529 5179 12587 5185
rect 12710 5176 12716 5228
rect 12768 5176 12774 5228
rect 15286 5176 15292 5228
rect 15344 5216 15350 5228
rect 15473 5219 15531 5225
rect 15473 5216 15485 5219
rect 15344 5188 15485 5216
rect 15344 5176 15350 5188
rect 15473 5185 15485 5188
rect 15519 5185 15531 5219
rect 15473 5179 15531 5185
rect 15746 5176 15752 5228
rect 15804 5216 15810 5228
rect 16761 5219 16819 5225
rect 16761 5216 16773 5219
rect 15804 5188 16773 5216
rect 15804 5176 15810 5188
rect 16761 5185 16773 5188
rect 16807 5185 16819 5219
rect 16761 5179 16819 5185
rect 13262 5148 13268 5160
rect 9999 5120 11744 5148
rect 12406 5120 13268 5148
rect 9999 5117 10011 5120
rect 9953 5111 10011 5117
rect 9401 5083 9459 5089
rect 9401 5049 9413 5083
rect 9447 5080 9459 5083
rect 12406 5080 12434 5120
rect 13262 5108 13268 5120
rect 13320 5108 13326 5160
rect 16485 5151 16543 5157
rect 16485 5117 16497 5151
rect 16531 5148 16543 5151
rect 16850 5148 16856 5160
rect 16531 5120 16856 5148
rect 16531 5117 16543 5120
rect 16485 5111 16543 5117
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 9447 5052 12434 5080
rect 9447 5049 9459 5052
rect 9401 5043 9459 5049
rect 15470 5040 15476 5092
rect 15528 5080 15534 5092
rect 15657 5083 15715 5089
rect 15657 5080 15669 5083
rect 15528 5052 15669 5080
rect 15528 5040 15534 5052
rect 15657 5049 15669 5052
rect 15703 5049 15715 5083
rect 15657 5043 15715 5049
rect 8312 4984 9352 5012
rect 9674 4972 9680 5024
rect 9732 4972 9738 5024
rect 10042 4972 10048 5024
rect 10100 4972 10106 5024
rect 12713 5015 12771 5021
rect 12713 4981 12725 5015
rect 12759 5012 12771 5015
rect 13722 5012 13728 5024
rect 12759 4984 13728 5012
rect 12759 4981 12771 4984
rect 12713 4975 12771 4981
rect 13722 4972 13728 4984
rect 13780 4972 13786 5024
rect 1104 4922 17388 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 17388 4922
rect 1104 4848 17388 4870
rect 2777 4811 2835 4817
rect 2777 4777 2789 4811
rect 2823 4808 2835 4811
rect 3234 4808 3240 4820
rect 2823 4780 3240 4808
rect 2823 4777 2835 4780
rect 2777 4771 2835 4777
rect 3234 4768 3240 4780
rect 3292 4768 3298 4820
rect 3513 4811 3571 4817
rect 3513 4777 3525 4811
rect 3559 4808 3571 4811
rect 3786 4808 3792 4820
rect 3559 4780 3792 4808
rect 3559 4777 3571 4780
rect 3513 4771 3571 4777
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 3970 4768 3976 4820
rect 4028 4768 4034 4820
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 4709 4811 4767 4817
rect 4709 4808 4721 4811
rect 4120 4780 4721 4808
rect 4120 4768 4126 4780
rect 4709 4777 4721 4780
rect 4755 4808 4767 4811
rect 4890 4808 4896 4820
rect 4755 4780 4896 4808
rect 4755 4777 4767 4780
rect 4709 4771 4767 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 5350 4768 5356 4820
rect 5408 4808 5414 4820
rect 6546 4808 6552 4820
rect 5408 4780 6552 4808
rect 5408 4768 5414 4780
rect 6546 4768 6552 4780
rect 6604 4808 6610 4820
rect 7377 4811 7435 4817
rect 7377 4808 7389 4811
rect 6604 4780 7389 4808
rect 6604 4768 6610 4780
rect 7377 4777 7389 4780
rect 7423 4777 7435 4811
rect 7377 4771 7435 4777
rect 9309 4811 9367 4817
rect 9309 4777 9321 4811
rect 9355 4808 9367 4811
rect 9766 4808 9772 4820
rect 9355 4780 9772 4808
rect 9355 4777 9367 4780
rect 9309 4771 9367 4777
rect 3252 4672 3280 4768
rect 3804 4672 3832 4768
rect 4433 4743 4491 4749
rect 4433 4709 4445 4743
rect 4479 4740 4491 4743
rect 5902 4740 5908 4752
rect 4479 4712 5908 4740
rect 4479 4709 4491 4712
rect 4433 4703 4491 4709
rect 5902 4700 5908 4712
rect 5960 4740 5966 4752
rect 6730 4740 6736 4752
rect 5960 4712 6736 4740
rect 5960 4700 5966 4712
rect 6730 4700 6736 4712
rect 6788 4700 6794 4752
rect 7098 4700 7104 4752
rect 7156 4740 7162 4752
rect 7156 4712 7328 4740
rect 7156 4700 7162 4712
rect 3252 4644 3556 4672
rect 3804 4644 4292 4672
rect 1394 4564 1400 4616
rect 1452 4564 1458 4616
rect 3050 4564 3056 4616
rect 3108 4604 3114 4616
rect 3329 4607 3387 4613
rect 3329 4604 3341 4607
rect 3108 4576 3341 4604
rect 3108 4564 3114 4576
rect 3329 4573 3341 4576
rect 3375 4573 3387 4607
rect 3528 4604 3556 4644
rect 3528 4576 3924 4604
rect 3329 4567 3387 4573
rect 1670 4545 1676 4548
rect 1664 4499 1676 4545
rect 1670 4496 1676 4499
rect 1728 4496 1734 4548
rect 3694 4496 3700 4548
rect 3752 4536 3758 4548
rect 3789 4539 3847 4545
rect 3789 4536 3801 4539
rect 3752 4508 3801 4536
rect 3752 4496 3758 4508
rect 3789 4505 3801 4508
rect 3835 4505 3847 4539
rect 3896 4536 3924 4576
rect 4062 4564 4068 4616
rect 4120 4564 4126 4616
rect 4264 4613 4292 4644
rect 6454 4632 6460 4684
rect 6512 4672 6518 4684
rect 6641 4675 6699 4681
rect 6641 4672 6653 4675
rect 6512 4644 6653 4672
rect 6512 4632 6518 4644
rect 6641 4641 6653 4644
rect 6687 4641 6699 4675
rect 6641 4635 6699 4641
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 6880 4644 7236 4672
rect 6880 4632 6886 4644
rect 7208 4613 7236 4644
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 7193 4607 7251 4613
rect 7193 4573 7205 4607
rect 7239 4573 7251 4607
rect 7300 4604 7328 4712
rect 7392 4672 7420 4771
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 16574 4808 16580 4820
rect 15028 4780 16580 4808
rect 8113 4743 8171 4749
rect 8113 4709 8125 4743
rect 8159 4740 8171 4743
rect 9490 4740 9496 4752
rect 8159 4712 9496 4740
rect 8159 4709 8171 4712
rect 8113 4703 8171 4709
rect 9490 4700 9496 4712
rect 9548 4700 9554 4752
rect 9585 4743 9643 4749
rect 9585 4709 9597 4743
rect 9631 4740 9643 4743
rect 10686 4740 10692 4752
rect 9631 4712 10692 4740
rect 9631 4709 9643 4712
rect 9585 4703 9643 4709
rect 10686 4700 10692 4712
rect 10744 4700 10750 4752
rect 7392 4644 7788 4672
rect 7760 4613 7788 4644
rect 8018 4632 8024 4684
rect 8076 4672 8082 4684
rect 8570 4672 8576 4684
rect 8076 4644 8576 4672
rect 8076 4632 8082 4644
rect 8570 4632 8576 4644
rect 8628 4672 8634 4684
rect 15028 4672 15056 4780
rect 16574 4768 16580 4780
rect 16632 4768 16638 4820
rect 16758 4768 16764 4820
rect 16816 4808 16822 4820
rect 17037 4811 17095 4817
rect 17037 4808 17049 4811
rect 16816 4780 17049 4808
rect 16816 4768 16822 4780
rect 17037 4777 17049 4780
rect 17083 4777 17095 4811
rect 17037 4771 17095 4777
rect 15470 4672 15476 4684
rect 8628 4644 9628 4672
rect 8628 4632 8634 4644
rect 7561 4607 7619 4613
rect 7561 4604 7573 4607
rect 7300 4576 7573 4604
rect 7193 4567 7251 4573
rect 7561 4573 7573 4576
rect 7607 4573 7619 4607
rect 7561 4567 7619 4573
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 7834 4564 7840 4616
rect 7892 4564 7898 4616
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 4617 4539 4675 4545
rect 4617 4536 4629 4539
rect 3896 4508 4629 4536
rect 3789 4499 3847 4505
rect 4617 4505 4629 4508
rect 4663 4505 4675 4539
rect 4617 4499 4675 4505
rect 6825 4539 6883 4545
rect 6825 4505 6837 4539
rect 6871 4536 6883 4539
rect 7650 4536 7656 4548
rect 6871 4508 7656 4536
rect 6871 4505 6883 4508
rect 6825 4499 6883 4505
rect 7650 4496 7656 4508
rect 7708 4496 7714 4548
rect 7944 4536 7972 4567
rect 8110 4564 8116 4616
rect 8168 4604 8174 4616
rect 8205 4607 8263 4613
rect 8205 4604 8217 4607
rect 8168 4576 8217 4604
rect 8168 4564 8174 4576
rect 8205 4573 8217 4576
rect 8251 4573 8263 4607
rect 9600 4604 9628 4644
rect 14936 4644 15056 4672
rect 15212 4644 15476 4672
rect 9677 4607 9735 4613
rect 9677 4604 9689 4607
rect 9600 4576 9689 4604
rect 8205 4567 8263 4573
rect 9677 4573 9689 4576
rect 9723 4573 9735 4607
rect 9677 4567 9735 4573
rect 9769 4607 9827 4613
rect 9769 4573 9781 4607
rect 9815 4604 9827 4607
rect 9950 4604 9956 4616
rect 9815 4576 9956 4604
rect 9815 4573 9827 4576
rect 9769 4567 9827 4573
rect 9950 4564 9956 4576
rect 10008 4564 10014 4616
rect 10045 4607 10103 4613
rect 10045 4573 10057 4607
rect 10091 4573 10103 4607
rect 10045 4567 10103 4573
rect 10060 4536 10088 4567
rect 10870 4564 10876 4616
rect 10928 4604 10934 4616
rect 11057 4607 11115 4613
rect 11057 4604 11069 4607
rect 10928 4576 11069 4604
rect 10928 4564 10934 4576
rect 11057 4573 11069 4576
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 13446 4564 13452 4616
rect 13504 4604 13510 4616
rect 13633 4607 13691 4613
rect 13633 4604 13645 4607
rect 13504 4576 13645 4604
rect 13504 4564 13510 4576
rect 13633 4573 13645 4576
rect 13679 4573 13691 4607
rect 13633 4567 13691 4573
rect 13722 4564 13728 4616
rect 13780 4564 13786 4616
rect 13909 4607 13967 4613
rect 13909 4573 13921 4607
rect 13955 4604 13967 4607
rect 13998 4604 14004 4616
rect 13955 4576 14004 4604
rect 13955 4573 13967 4576
rect 13909 4567 13967 4573
rect 13998 4564 14004 4576
rect 14056 4564 14062 4616
rect 14936 4613 14964 4644
rect 15212 4613 15240 4644
rect 15470 4632 15476 4644
rect 15528 4632 15534 4684
rect 14921 4607 14979 4613
rect 14921 4573 14933 4607
rect 14967 4573 14979 4607
rect 14921 4567 14979 4573
rect 15013 4607 15071 4613
rect 15013 4573 15025 4607
rect 15059 4573 15071 4607
rect 15013 4567 15071 4573
rect 15197 4607 15255 4613
rect 15197 4573 15209 4607
rect 15243 4573 15255 4607
rect 15197 4567 15255 4573
rect 15028 4536 15056 4567
rect 15378 4564 15384 4616
rect 15436 4564 15442 4616
rect 15654 4564 15660 4616
rect 15712 4564 15718 4616
rect 7852 4508 7972 4536
rect 9692 4508 10088 4536
rect 13832 4508 15056 4536
rect 15289 4539 15347 4545
rect 5626 4428 5632 4480
rect 5684 4468 5690 4480
rect 6362 4468 6368 4480
rect 5684 4440 6368 4468
rect 5684 4428 5690 4440
rect 6362 4428 6368 4440
rect 6420 4468 6426 4480
rect 7852 4468 7880 4508
rect 9692 4480 9720 4508
rect 8389 4471 8447 4477
rect 8389 4468 8401 4471
rect 6420 4440 8401 4468
rect 6420 4428 6426 4440
rect 8389 4437 8401 4440
rect 8435 4437 8447 4471
rect 8389 4431 8447 4437
rect 9674 4428 9680 4480
rect 9732 4428 9738 4480
rect 9953 4471 10011 4477
rect 9953 4437 9965 4471
rect 9999 4468 10011 4471
rect 10134 4468 10140 4480
rect 9999 4440 10140 4468
rect 9999 4437 10011 4440
rect 9953 4431 10011 4437
rect 10134 4428 10140 4440
rect 10192 4468 10198 4480
rect 11146 4468 11152 4480
rect 10192 4440 11152 4468
rect 10192 4428 10198 4440
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 11241 4471 11299 4477
rect 11241 4437 11253 4471
rect 11287 4468 11299 4471
rect 13538 4468 13544 4480
rect 11287 4440 13544 4468
rect 11287 4437 11299 4440
rect 11241 4431 11299 4437
rect 13538 4428 13544 4440
rect 13596 4428 13602 4480
rect 13832 4477 13860 4508
rect 15289 4505 15301 4539
rect 15335 4505 15347 4539
rect 15902 4539 15960 4545
rect 15902 4536 15914 4539
rect 15289 4499 15347 4505
rect 15580 4508 15914 4536
rect 13817 4471 13875 4477
rect 13817 4437 13829 4471
rect 13863 4437 13875 4471
rect 13817 4431 13875 4437
rect 14737 4471 14795 4477
rect 14737 4437 14749 4471
rect 14783 4468 14795 4471
rect 15194 4468 15200 4480
rect 14783 4440 15200 4468
rect 14783 4437 14795 4440
rect 14737 4431 14795 4437
rect 15194 4428 15200 4440
rect 15252 4468 15258 4480
rect 15304 4468 15332 4499
rect 15580 4477 15608 4508
rect 15902 4505 15914 4508
rect 15948 4505 15960 4539
rect 15902 4499 15960 4505
rect 15252 4440 15332 4468
rect 15565 4471 15623 4477
rect 15252 4428 15258 4440
rect 15565 4437 15577 4471
rect 15611 4437 15623 4471
rect 15565 4431 15623 4437
rect 1104 4378 17388 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 17388 4378
rect 1104 4304 17388 4326
rect 1486 4224 1492 4276
rect 1544 4264 1550 4276
rect 1581 4267 1639 4273
rect 1581 4264 1593 4267
rect 1544 4236 1593 4264
rect 1544 4224 1550 4236
rect 1581 4233 1593 4236
rect 1627 4233 1639 4267
rect 1581 4227 1639 4233
rect 1670 4224 1676 4276
rect 1728 4224 1734 4276
rect 6086 4224 6092 4276
rect 6144 4264 6150 4276
rect 7101 4267 7159 4273
rect 7101 4264 7113 4267
rect 6144 4236 7113 4264
rect 6144 4224 6150 4236
rect 7101 4233 7113 4236
rect 7147 4233 7159 4267
rect 7101 4227 7159 4233
rect 7650 4224 7656 4276
rect 7708 4224 7714 4276
rect 9674 4224 9680 4276
rect 9732 4264 9738 4276
rect 9927 4267 9985 4273
rect 9927 4264 9939 4267
rect 9732 4236 9939 4264
rect 9732 4224 9738 4236
rect 9927 4233 9939 4236
rect 9973 4264 9985 4267
rect 10321 4267 10379 4273
rect 10321 4264 10333 4267
rect 9973 4236 10333 4264
rect 9973 4233 9985 4236
rect 9927 4227 9985 4233
rect 10321 4233 10333 4236
rect 10367 4264 10379 4267
rect 10962 4264 10968 4276
rect 10367 4236 10968 4264
rect 10367 4233 10379 4236
rect 10321 4227 10379 4233
rect 10962 4224 10968 4236
rect 11020 4224 11026 4276
rect 14921 4267 14979 4273
rect 14921 4264 14933 4267
rect 14200 4236 14933 4264
rect 7466 4156 7472 4208
rect 7524 4196 7530 4208
rect 7805 4199 7863 4205
rect 7805 4196 7817 4199
rect 7524 4168 7817 4196
rect 7524 4156 7530 4168
rect 7805 4165 7817 4168
rect 7851 4165 7863 4199
rect 7805 4159 7863 4165
rect 8021 4199 8079 4205
rect 8021 4165 8033 4199
rect 8067 4196 8079 4199
rect 8202 4196 8208 4208
rect 8067 4168 8208 4196
rect 8067 4165 8079 4168
rect 8021 4159 8079 4165
rect 8202 4156 8208 4168
rect 8260 4156 8266 4208
rect 10134 4156 10140 4208
rect 10192 4156 10198 4208
rect 10870 4156 10876 4208
rect 10928 4156 10934 4208
rect 11149 4199 11207 4205
rect 11149 4196 11161 4199
rect 10980 4168 11161 4196
rect 1302 4088 1308 4140
rect 1360 4128 1366 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 1360 4100 1409 4128
rect 1360 4088 1366 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 1854 4088 1860 4140
rect 1912 4088 1918 4140
rect 6362 4088 6368 4140
rect 6420 4088 6426 4140
rect 6546 4088 6552 4140
rect 6604 4088 6610 4140
rect 6730 4088 6736 4140
rect 6788 4128 6794 4140
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6788 4100 6837 4128
rect 6788 4088 6794 4100
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 7285 4131 7343 4137
rect 7285 4097 7297 4131
rect 7331 4128 7343 4131
rect 7331 4100 7880 4128
rect 7331 4097 7343 4100
rect 7285 4091 7343 4097
rect 7852 4072 7880 4100
rect 9122 4088 9128 4140
rect 9180 4128 9186 4140
rect 9217 4131 9275 4137
rect 9217 4128 9229 4131
rect 9180 4100 9229 4128
rect 9180 4088 9186 4100
rect 9217 4097 9229 4100
rect 9263 4097 9275 4131
rect 9217 4091 9275 4097
rect 9398 4088 9404 4140
rect 9456 4088 9462 4140
rect 9490 4088 9496 4140
rect 9548 4128 9554 4140
rect 10318 4128 10324 4140
rect 9548 4100 10324 4128
rect 9548 4088 9554 4100
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 10413 4131 10471 4137
rect 10413 4097 10425 4131
rect 10459 4097 10471 4131
rect 10413 4091 10471 4097
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 10594 4128 10600 4140
rect 10551 4100 10600 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 7190 4020 7196 4072
rect 7248 4060 7254 4072
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 7248 4032 7389 4060
rect 7248 4020 7254 4032
rect 7377 4029 7389 4032
rect 7423 4029 7435 4063
rect 7377 4023 7435 4029
rect 7466 4020 7472 4072
rect 7524 4020 7530 4072
rect 7834 4020 7840 4072
rect 7892 4020 7898 4072
rect 9309 4063 9367 4069
rect 9309 4029 9321 4063
rect 9355 4060 9367 4063
rect 10428 4060 10456 4091
rect 10594 4088 10600 4100
rect 10652 4128 10658 4140
rect 10980 4128 11008 4168
rect 11149 4165 11161 4168
rect 11195 4165 11207 4199
rect 11333 4199 11391 4205
rect 11333 4196 11345 4199
rect 11149 4159 11207 4165
rect 11256 4168 11345 4196
rect 10652 4100 11008 4128
rect 10652 4088 10658 4100
rect 9355 4032 10456 4060
rect 9355 4029 9367 4032
rect 9309 4023 9367 4029
rect 10686 4020 10692 4072
rect 10744 4020 10750 4072
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 10965 4063 11023 4069
rect 10965 4060 10977 4063
rect 10836 4032 10977 4060
rect 10836 4020 10842 4032
rect 10965 4029 10977 4032
rect 11011 4029 11023 4063
rect 10965 4023 11023 4029
rect 7009 3995 7067 4001
rect 7009 3961 7021 3995
rect 7055 3992 7067 3995
rect 11256 3992 11284 4168
rect 11333 4165 11345 4168
rect 11379 4196 11391 4199
rect 11885 4199 11943 4205
rect 11885 4196 11897 4199
rect 11379 4168 11897 4196
rect 11379 4165 11391 4168
rect 11333 4159 11391 4165
rect 11885 4165 11897 4168
rect 11931 4165 11943 4199
rect 11885 4159 11943 4165
rect 12066 4156 12072 4208
rect 12124 4156 12130 4208
rect 13357 4199 13415 4205
rect 13357 4165 13369 4199
rect 13403 4196 13415 4199
rect 13630 4196 13636 4208
rect 13403 4168 13636 4196
rect 13403 4165 13415 4168
rect 13357 4159 13415 4165
rect 13630 4156 13636 4168
rect 13688 4156 13694 4208
rect 13725 4199 13783 4205
rect 13725 4165 13737 4199
rect 13771 4196 13783 4199
rect 14090 4196 14096 4208
rect 13771 4168 14096 4196
rect 13771 4165 13783 4168
rect 13725 4159 13783 4165
rect 14090 4156 14096 4168
rect 14148 4156 14154 4208
rect 13538 4088 13544 4140
rect 13596 4088 13602 4140
rect 13814 4088 13820 4140
rect 13872 4088 13878 4140
rect 13998 4088 14004 4140
rect 14056 4088 14062 4140
rect 13173 4063 13231 4069
rect 13173 4029 13185 4063
rect 13219 4060 13231 4063
rect 13354 4060 13360 4072
rect 13219 4032 13360 4060
rect 13219 4029 13231 4032
rect 13173 4023 13231 4029
rect 13354 4020 13360 4032
rect 13412 4020 13418 4072
rect 13449 4063 13507 4069
rect 13449 4029 13461 4063
rect 13495 4029 13507 4063
rect 13449 4023 13507 4029
rect 13633 4063 13691 4069
rect 13633 4029 13645 4063
rect 13679 4060 13691 4063
rect 14200 4060 14228 4236
rect 14921 4233 14933 4236
rect 14967 4264 14979 4267
rect 15194 4264 15200 4276
rect 14967 4236 15200 4264
rect 14967 4233 14979 4236
rect 14921 4227 14979 4233
rect 15194 4224 15200 4236
rect 15252 4224 15258 4276
rect 15378 4224 15384 4276
rect 15436 4264 15442 4276
rect 15841 4267 15899 4273
rect 15841 4264 15853 4267
rect 15436 4236 15853 4264
rect 15436 4224 15442 4236
rect 15841 4233 15853 4236
rect 15887 4233 15899 4267
rect 15841 4227 15899 4233
rect 14277 4131 14335 4137
rect 14277 4097 14289 4131
rect 14323 4128 14335 4131
rect 14734 4128 14740 4140
rect 14323 4100 14740 4128
rect 14323 4097 14335 4100
rect 14277 4091 14335 4097
rect 14734 4088 14740 4100
rect 14792 4088 14798 4140
rect 15013 4131 15071 4137
rect 15013 4097 15025 4131
rect 15059 4128 15071 4131
rect 15105 4131 15163 4137
rect 15105 4128 15117 4131
rect 15059 4100 15117 4128
rect 15059 4097 15071 4100
rect 15013 4091 15071 4097
rect 15105 4097 15117 4100
rect 15151 4097 15163 4131
rect 15105 4091 15163 4097
rect 15746 4088 15752 4140
rect 15804 4088 15810 4140
rect 16485 4131 16543 4137
rect 16485 4097 16497 4131
rect 16531 4128 16543 4131
rect 16758 4128 16764 4140
rect 16531 4100 16764 4128
rect 16531 4097 16543 4100
rect 16485 4091 16543 4097
rect 16758 4088 16764 4100
rect 16816 4088 16822 4140
rect 13679 4032 14228 4060
rect 14461 4063 14519 4069
rect 13679 4029 13691 4032
rect 13633 4023 13691 4029
rect 14461 4029 14473 4063
rect 14507 4060 14519 4063
rect 15286 4060 15292 4072
rect 14507 4032 15292 4060
rect 14507 4029 14519 4032
rect 14461 4023 14519 4029
rect 7055 3964 11284 3992
rect 13464 3992 13492 4023
rect 15286 4020 15292 4032
rect 15344 4020 15350 4072
rect 13817 3995 13875 4001
rect 13817 3992 13829 3995
rect 13464 3964 13829 3992
rect 7055 3961 7067 3964
rect 7009 3955 7067 3961
rect 13817 3961 13829 3964
rect 13863 3961 13875 3995
rect 13817 3955 13875 3961
rect 7834 3884 7840 3936
rect 7892 3884 7898 3936
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 9490 3924 9496 3936
rect 8996 3896 9496 3924
rect 8996 3884 9002 3896
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 9769 3927 9827 3933
rect 9769 3893 9781 3927
rect 9815 3924 9827 3927
rect 9858 3924 9864 3936
rect 9815 3896 9864 3924
rect 9815 3893 9827 3896
rect 9769 3887 9827 3893
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 9950 3884 9956 3936
rect 10008 3884 10014 3936
rect 10318 3884 10324 3936
rect 10376 3924 10382 3936
rect 10597 3927 10655 3933
rect 10597 3924 10609 3927
rect 10376 3896 10609 3924
rect 10376 3884 10382 3896
rect 10597 3893 10609 3896
rect 10643 3893 10655 3927
rect 10597 3887 10655 3893
rect 12253 3927 12311 3933
rect 12253 3893 12265 3927
rect 12299 3924 12311 3927
rect 13998 3924 14004 3936
rect 12299 3896 14004 3924
rect 12299 3893 12311 3896
rect 12253 3887 12311 3893
rect 13998 3884 14004 3896
rect 14056 3884 14062 3936
rect 14550 3884 14556 3936
rect 14608 3884 14614 3936
rect 1104 3834 17388 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 17388 3834
rect 1104 3760 17388 3782
rect 6641 3723 6699 3729
rect 6641 3689 6653 3723
rect 6687 3720 6699 3723
rect 6822 3720 6828 3732
rect 6687 3692 6828 3720
rect 6687 3689 6699 3692
rect 6641 3683 6699 3689
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7101 3723 7159 3729
rect 7101 3689 7113 3723
rect 7147 3720 7159 3723
rect 7466 3720 7472 3732
rect 7147 3692 7472 3720
rect 7147 3689 7159 3692
rect 7101 3683 7159 3689
rect 7466 3680 7472 3692
rect 7524 3680 7530 3732
rect 7745 3723 7803 3729
rect 7745 3689 7757 3723
rect 7791 3720 7803 3723
rect 7834 3720 7840 3732
rect 7791 3692 7840 3720
rect 7791 3689 7803 3692
rect 7745 3683 7803 3689
rect 6549 3655 6607 3661
rect 6549 3621 6561 3655
rect 6595 3652 6607 3655
rect 6733 3655 6791 3661
rect 6733 3652 6745 3655
rect 6595 3624 6745 3652
rect 6595 3621 6607 3624
rect 6549 3615 6607 3621
rect 6733 3621 6745 3624
rect 6779 3652 6791 3655
rect 7760 3652 7788 3683
rect 7834 3680 7840 3692
rect 7892 3720 7898 3732
rect 7892 3692 8432 3720
rect 7892 3680 7898 3692
rect 6779 3624 7788 3652
rect 7929 3655 7987 3661
rect 6779 3621 6791 3624
rect 6733 3615 6791 3621
rect 7929 3621 7941 3655
rect 7975 3652 7987 3655
rect 8110 3652 8116 3664
rect 7975 3624 8116 3652
rect 7975 3621 7987 3624
rect 7929 3615 7987 3621
rect 8110 3612 8116 3624
rect 8168 3612 8174 3664
rect 8202 3612 8208 3664
rect 8260 3652 8266 3664
rect 8260 3624 8340 3652
rect 8260 3612 8266 3624
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3516 6699 3519
rect 7377 3519 7435 3525
rect 7377 3516 7389 3519
rect 6687 3488 7389 3516
rect 6687 3485 6699 3488
rect 6641 3479 6699 3485
rect 7377 3485 7389 3488
rect 7423 3516 7435 3519
rect 7466 3516 7472 3528
rect 7423 3488 7472 3516
rect 7423 3485 7435 3488
rect 7377 3479 7435 3485
rect 7466 3476 7472 3488
rect 7524 3516 7530 3528
rect 8018 3516 8024 3528
rect 7524 3488 8024 3516
rect 7524 3476 7530 3488
rect 8018 3476 8024 3488
rect 8076 3516 8082 3528
rect 8312 3525 8340 3624
rect 8404 3593 8432 3692
rect 9122 3680 9128 3732
rect 9180 3680 9186 3732
rect 10962 3680 10968 3732
rect 11020 3680 11026 3732
rect 12342 3680 12348 3732
rect 12400 3680 12406 3732
rect 12526 3680 12532 3732
rect 12584 3680 12590 3732
rect 15746 3680 15752 3732
rect 15804 3720 15810 3732
rect 16025 3723 16083 3729
rect 16025 3720 16037 3723
rect 15804 3692 16037 3720
rect 15804 3680 15810 3692
rect 16025 3689 16037 3692
rect 16071 3689 16083 3723
rect 16025 3683 16083 3689
rect 16209 3723 16267 3729
rect 16209 3689 16221 3723
rect 16255 3720 16267 3723
rect 16482 3720 16488 3732
rect 16255 3692 16488 3720
rect 16255 3689 16267 3692
rect 16209 3683 16267 3689
rect 16482 3680 16488 3692
rect 16540 3680 16546 3732
rect 8389 3587 8447 3593
rect 8389 3553 8401 3587
rect 8435 3584 8447 3587
rect 9140 3584 9168 3680
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 10597 3655 10655 3661
rect 10597 3652 10609 3655
rect 10008 3624 10609 3652
rect 10008 3612 10014 3624
rect 10597 3621 10609 3624
rect 10643 3621 10655 3655
rect 10597 3615 10655 3621
rect 11149 3655 11207 3661
rect 11149 3621 11161 3655
rect 11195 3621 11207 3655
rect 11149 3615 11207 3621
rect 8435 3556 9168 3584
rect 11164 3584 11192 3615
rect 12250 3584 12256 3596
rect 11164 3556 12256 3584
rect 8435 3553 8447 3556
rect 8389 3547 8447 3553
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 8076 3488 8217 3516
rect 8076 3476 8082 3488
rect 8205 3485 8217 3488
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 8297 3519 8355 3525
rect 8297 3485 8309 3519
rect 8343 3516 8355 3519
rect 9398 3516 9404 3528
rect 8343 3488 9404 3516
rect 8343 3485 8355 3488
rect 8297 3479 8355 3485
rect 6365 3451 6423 3457
rect 6365 3417 6377 3451
rect 6411 3448 6423 3451
rect 7101 3451 7159 3457
rect 7101 3448 7113 3451
rect 6411 3420 7113 3448
rect 6411 3417 6423 3420
rect 6365 3411 6423 3417
rect 7101 3417 7113 3420
rect 7147 3448 7159 3451
rect 7190 3448 7196 3460
rect 7147 3420 7196 3448
rect 7147 3417 7159 3420
rect 7101 3411 7159 3417
rect 7190 3408 7196 3420
rect 7248 3448 7254 3460
rect 7745 3451 7803 3457
rect 7745 3448 7757 3451
rect 7248 3420 7757 3448
rect 7248 3408 7254 3420
rect 7745 3417 7757 3420
rect 7791 3448 7803 3451
rect 8110 3448 8116 3460
rect 7791 3420 8116 3448
rect 7791 3417 7803 3420
rect 7745 3411 7803 3417
rect 8110 3408 8116 3420
rect 8168 3408 8174 3460
rect 8220 3448 8248 3479
rect 9398 3476 9404 3488
rect 9456 3516 9462 3528
rect 9493 3519 9551 3525
rect 9493 3516 9505 3519
rect 9456 3488 9505 3516
rect 9456 3476 9462 3488
rect 9493 3485 9505 3488
rect 9539 3516 9551 3519
rect 9539 3488 11008 3516
rect 9539 3485 9551 3488
rect 9493 3479 9551 3485
rect 9125 3451 9183 3457
rect 9125 3448 9137 3451
rect 8220 3420 9137 3448
rect 9125 3417 9137 3420
rect 9171 3448 9183 3451
rect 9950 3448 9956 3460
rect 9171 3420 9956 3448
rect 9171 3417 9183 3420
rect 9125 3411 9183 3417
rect 9950 3408 9956 3420
rect 10008 3408 10014 3460
rect 10980 3457 11008 3488
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 11425 3519 11483 3525
rect 11425 3516 11437 3519
rect 11204 3488 11437 3516
rect 11204 3476 11210 3488
rect 11425 3485 11437 3488
rect 11471 3485 11483 3519
rect 11425 3479 11483 3485
rect 12066 3476 12072 3528
rect 12124 3476 12130 3528
rect 12345 3519 12403 3525
rect 12345 3485 12357 3519
rect 12391 3485 12403 3519
rect 12345 3479 12403 3485
rect 10965 3451 11023 3457
rect 10965 3417 10977 3451
rect 11011 3448 11023 3451
rect 11241 3451 11299 3457
rect 11241 3448 11253 3451
rect 11011 3420 11253 3448
rect 11011 3417 11023 3420
rect 10965 3411 11023 3417
rect 11241 3417 11253 3420
rect 11287 3417 11299 3451
rect 11241 3411 11299 3417
rect 7282 3340 7288 3392
rect 7340 3340 7346 3392
rect 7558 3340 7564 3392
rect 7616 3380 7622 3392
rect 8021 3383 8079 3389
rect 8021 3380 8033 3383
rect 7616 3352 8033 3380
rect 7616 3340 7622 3352
rect 8021 3349 8033 3352
rect 8067 3349 8079 3383
rect 8021 3343 8079 3349
rect 8941 3383 8999 3389
rect 8941 3349 8953 3383
rect 8987 3380 8999 3383
rect 9306 3380 9312 3392
rect 8987 3352 9312 3380
rect 8987 3349 8999 3352
rect 8941 3343 8999 3349
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9490 3340 9496 3392
rect 9548 3380 9554 3392
rect 12360 3380 12388 3479
rect 14642 3476 14648 3528
rect 14700 3516 14706 3528
rect 15654 3516 15660 3528
rect 14700 3488 15660 3516
rect 14700 3476 14706 3488
rect 15654 3476 15660 3488
rect 15712 3476 15718 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 16117 3519 16175 3525
rect 16117 3516 16129 3519
rect 15988 3488 16129 3516
rect 15988 3476 15994 3488
rect 16117 3485 16129 3488
rect 16163 3485 16175 3519
rect 16117 3479 16175 3485
rect 14550 3408 14556 3460
rect 14608 3448 14614 3460
rect 14890 3451 14948 3457
rect 14890 3448 14902 3451
rect 14608 3420 14902 3448
rect 14608 3408 14614 3420
rect 14890 3417 14902 3420
rect 14936 3417 14948 3451
rect 14890 3411 14948 3417
rect 9548 3352 12388 3380
rect 9548 3340 9554 3352
rect 1104 3290 17388 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 17388 3290
rect 1104 3216 17388 3238
rect 7745 3179 7803 3185
rect 7745 3145 7757 3179
rect 7791 3176 7803 3179
rect 7834 3176 7840 3188
rect 7791 3148 7840 3176
rect 7791 3145 7803 3148
rect 7745 3139 7803 3145
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 9861 3179 9919 3185
rect 9861 3145 9873 3179
rect 9907 3176 9919 3179
rect 9950 3176 9956 3188
rect 9907 3148 9956 3176
rect 9907 3145 9919 3148
rect 9861 3139 9919 3145
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 11146 3136 11152 3188
rect 11204 3176 11210 3188
rect 11333 3179 11391 3185
rect 11333 3176 11345 3179
rect 11204 3148 11345 3176
rect 11204 3136 11210 3148
rect 11333 3145 11345 3148
rect 11379 3145 11391 3179
rect 11333 3139 11391 3145
rect 1394 3068 1400 3120
rect 1452 3108 1458 3120
rect 9214 3108 9220 3120
rect 1452 3080 9220 3108
rect 1452 3068 1458 3080
rect 6380 3049 6408 3080
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 6621 3043 6679 3049
rect 6621 3040 6633 3043
rect 6512 3012 6633 3040
rect 6512 3000 6518 3012
rect 6621 3009 6633 3012
rect 6667 3009 6679 3043
rect 6621 3003 6679 3009
rect 7834 3000 7840 3052
rect 7892 3040 7898 3052
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 7892 3012 8125 3040
rect 7892 3000 7898 3012
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 8113 3003 8171 3009
rect 8202 3000 8208 3052
rect 8260 3000 8266 3052
rect 8496 3049 8524 3080
rect 9214 3068 9220 3080
rect 9272 3108 9278 3120
rect 14642 3108 14648 3120
rect 9272 3080 14648 3108
rect 9272 3068 9278 3080
rect 8481 3043 8539 3049
rect 8481 3009 8493 3043
rect 8527 3009 8539 3043
rect 8481 3003 8539 3009
rect 8748 3043 8806 3049
rect 8748 3009 8760 3043
rect 8794 3040 8806 3043
rect 9122 3040 9128 3052
rect 8794 3012 9128 3040
rect 8794 3009 8806 3012
rect 8748 3003 8806 3009
rect 9122 3000 9128 3012
rect 9180 3000 9186 3052
rect 9968 3049 9996 3080
rect 10226 3049 10232 3052
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3009 10011 3043
rect 9953 3003 10011 3009
rect 10220 3003 10232 3049
rect 10226 3000 10232 3003
rect 10284 3000 10290 3052
rect 14274 3000 14280 3052
rect 14332 3049 14338 3052
rect 14568 3049 14596 3080
rect 14642 3068 14648 3080
rect 14700 3068 14706 3120
rect 14332 3003 14344 3049
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 14332 3000 14338 3003
rect 8018 2932 8024 2984
rect 8076 2932 8082 2984
rect 14642 2932 14648 2984
rect 14700 2972 14706 2984
rect 15197 2975 15255 2981
rect 15197 2972 15209 2975
rect 14700 2944 15209 2972
rect 14700 2932 14706 2944
rect 15197 2941 15209 2944
rect 15243 2941 15255 2975
rect 15197 2935 15255 2941
rect 6638 2796 6644 2848
rect 6696 2836 6702 2848
rect 7837 2839 7895 2845
rect 7837 2836 7849 2839
rect 6696 2808 7849 2836
rect 6696 2796 6702 2808
rect 7837 2805 7849 2808
rect 7883 2805 7895 2839
rect 7837 2799 7895 2805
rect 13173 2839 13231 2845
rect 13173 2805 13185 2839
rect 13219 2836 13231 2839
rect 13906 2836 13912 2848
rect 13219 2808 13912 2836
rect 13219 2805 13231 2808
rect 13173 2799 13231 2805
rect 13906 2796 13912 2808
rect 13964 2796 13970 2848
rect 14550 2796 14556 2848
rect 14608 2836 14614 2848
rect 14645 2839 14703 2845
rect 14645 2836 14657 2839
rect 14608 2808 14657 2836
rect 14608 2796 14614 2808
rect 14645 2805 14657 2808
rect 14691 2805 14703 2839
rect 14645 2799 14703 2805
rect 1104 2746 17388 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 17388 2746
rect 1104 2672 17388 2694
rect 6089 2635 6147 2641
rect 6089 2601 6101 2635
rect 6135 2632 6147 2635
rect 6454 2632 6460 2644
rect 6135 2604 6460 2632
rect 6135 2601 6147 2604
rect 6089 2595 6147 2601
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 9122 2592 9128 2644
rect 9180 2592 9186 2644
rect 10226 2592 10232 2644
rect 10284 2632 10290 2644
rect 10413 2635 10471 2641
rect 10413 2632 10425 2635
rect 10284 2604 10425 2632
rect 10284 2592 10290 2604
rect 10413 2601 10425 2604
rect 10459 2601 10471 2635
rect 10413 2595 10471 2601
rect 14093 2635 14151 2641
rect 14093 2601 14105 2635
rect 14139 2632 14151 2635
rect 14274 2632 14280 2644
rect 14139 2604 14280 2632
rect 14139 2601 14151 2604
rect 14093 2595 14151 2601
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 14642 2496 14648 2508
rect 13924 2468 14648 2496
rect 13924 2440 13952 2468
rect 14642 2456 14648 2468
rect 14700 2456 14706 2508
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5868 2400 5917 2428
rect 5868 2388 5874 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 9088 2400 9321 2428
rect 9088 2388 9094 2400
rect 9309 2397 9321 2400
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10376 2400 10609 2428
rect 10376 2388 10382 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 13906 2388 13912 2440
rect 13964 2388 13970 2440
rect 14090 2388 14096 2440
rect 14148 2428 14154 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 14148 2400 14289 2428
rect 14148 2388 14154 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 14550 2388 14556 2440
rect 14608 2388 14614 2440
rect 14737 2431 14795 2437
rect 14737 2397 14749 2431
rect 14783 2428 14795 2431
rect 16022 2428 16028 2440
rect 14783 2400 16028 2428
rect 14783 2397 14795 2400
rect 14737 2391 14795 2397
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 13725 2295 13783 2301
rect 13725 2292 13737 2295
rect 13596 2264 13737 2292
rect 13596 2252 13602 2264
rect 13725 2261 13737 2264
rect 13771 2261 13783 2295
rect 13725 2255 13783 2261
rect 1104 2202 17388 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 17388 2202
rect 1104 2128 17388 2150
<< via1 >>
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 12900 17824 12952 17876
rect 13544 17824 13596 17876
rect 13268 17552 13320 17604
rect 14740 17552 14792 17604
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 14740 17323 14792 17332
rect 14740 17289 14749 17323
rect 14749 17289 14783 17323
rect 14783 17289 14792 17323
rect 14740 17280 14792 17289
rect 12532 17144 12584 17196
rect 15200 17212 15252 17264
rect 13636 17187 13688 17196
rect 13636 17153 13670 17187
rect 13670 17153 13688 17187
rect 13636 17144 13688 17153
rect 16764 17187 16816 17196
rect 16764 17153 16773 17187
rect 16773 17153 16807 17187
rect 16807 17153 16816 17187
rect 16764 17144 16816 17153
rect 13268 16983 13320 16992
rect 13268 16949 13277 16983
rect 13277 16949 13311 16983
rect 13311 16949 13320 16983
rect 13268 16940 13320 16949
rect 14004 16940 14056 16992
rect 15292 16940 15344 16992
rect 16488 16940 16540 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 12532 16779 12584 16788
rect 12532 16745 12541 16779
rect 12541 16745 12575 16779
rect 12575 16745 12584 16779
rect 12532 16736 12584 16745
rect 16764 16736 16816 16788
rect 13268 16600 13320 16652
rect 15200 16600 15252 16652
rect 12808 16507 12860 16516
rect 12808 16473 12817 16507
rect 12817 16473 12851 16507
rect 12851 16473 12860 16507
rect 12808 16464 12860 16473
rect 13084 16575 13136 16584
rect 13084 16541 13093 16575
rect 13093 16541 13127 16575
rect 13127 16541 13136 16575
rect 13084 16532 13136 16541
rect 14372 16532 14424 16584
rect 15292 16532 15344 16584
rect 15568 16575 15620 16584
rect 15568 16541 15577 16575
rect 15577 16541 15611 16575
rect 15611 16541 15620 16575
rect 15568 16532 15620 16541
rect 14096 16464 14148 16516
rect 13268 16396 13320 16448
rect 14188 16396 14240 16448
rect 14924 16439 14976 16448
rect 14924 16405 14933 16439
rect 14933 16405 14967 16439
rect 14967 16405 14976 16439
rect 14924 16396 14976 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 11980 16124 12032 16176
rect 8300 16056 8352 16108
rect 10232 16099 10284 16108
rect 10232 16065 10241 16099
rect 10241 16065 10275 16099
rect 10275 16065 10284 16099
rect 10232 16056 10284 16065
rect 10048 16031 10100 16040
rect 10048 15997 10057 16031
rect 10057 15997 10091 16031
rect 10091 15997 10100 16031
rect 10048 15988 10100 15997
rect 10968 16056 11020 16108
rect 13636 16235 13688 16244
rect 13636 16201 13645 16235
rect 13645 16201 13679 16235
rect 13679 16201 13688 16235
rect 13636 16192 13688 16201
rect 12440 16056 12492 16108
rect 11060 15920 11112 15972
rect 11888 15920 11940 15972
rect 13268 16099 13320 16108
rect 13268 16065 13277 16099
rect 13277 16065 13311 16099
rect 13311 16065 13320 16099
rect 13268 16056 13320 16065
rect 14004 16124 14056 16176
rect 14096 16099 14148 16108
rect 14096 16065 14105 16099
rect 14105 16065 14139 16099
rect 14139 16065 14148 16099
rect 14096 16056 14148 16065
rect 14188 16099 14240 16108
rect 14188 16065 14197 16099
rect 14197 16065 14231 16099
rect 14231 16065 14240 16099
rect 14188 16056 14240 16065
rect 14924 16192 14976 16244
rect 15568 16192 15620 16244
rect 15200 16124 15252 16176
rect 14004 15988 14056 16040
rect 14096 15920 14148 15972
rect 11612 15852 11664 15904
rect 12256 15895 12308 15904
rect 12256 15861 12265 15895
rect 12265 15861 12299 15895
rect 12299 15861 12308 15895
rect 12256 15852 12308 15861
rect 15476 15852 15528 15904
rect 16948 15895 17000 15904
rect 16948 15861 16957 15895
rect 16957 15861 16991 15895
rect 16991 15861 17000 15895
rect 16948 15852 17000 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 6184 15648 6236 15700
rect 7656 15648 7708 15700
rect 8300 15691 8352 15700
rect 8300 15657 8309 15691
rect 8309 15657 8343 15691
rect 8343 15657 8352 15691
rect 8300 15648 8352 15657
rect 9128 15691 9180 15700
rect 9128 15657 9137 15691
rect 9137 15657 9171 15691
rect 9171 15657 9180 15691
rect 9128 15648 9180 15657
rect 10232 15648 10284 15700
rect 7104 15580 7156 15632
rect 10968 15648 11020 15700
rect 11152 15648 11204 15700
rect 12256 15691 12308 15700
rect 12256 15657 12265 15691
rect 12265 15657 12299 15691
rect 12299 15657 12308 15691
rect 12256 15648 12308 15657
rect 12716 15648 12768 15700
rect 14188 15648 14240 15700
rect 15292 15648 15344 15700
rect 7932 15555 7984 15564
rect 7932 15521 7941 15555
rect 7941 15521 7975 15555
rect 7975 15521 7984 15555
rect 7932 15512 7984 15521
rect 5540 15376 5592 15428
rect 5908 15487 5960 15496
rect 5908 15453 5917 15487
rect 5917 15453 5951 15487
rect 5951 15453 5960 15487
rect 5908 15444 5960 15453
rect 8300 15444 8352 15496
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 9588 15444 9640 15496
rect 10232 15555 10284 15564
rect 10232 15521 10241 15555
rect 10241 15521 10275 15555
rect 10275 15521 10284 15555
rect 10232 15512 10284 15521
rect 11060 15580 11112 15632
rect 13268 15580 13320 15632
rect 15108 15580 15160 15632
rect 6828 15376 6880 15428
rect 10140 15419 10192 15428
rect 10140 15385 10149 15419
rect 10149 15385 10183 15419
rect 10183 15385 10192 15419
rect 10140 15376 10192 15385
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 11060 15376 11112 15428
rect 11704 15444 11756 15496
rect 15200 15512 15252 15564
rect 9680 15308 9732 15360
rect 14096 15376 14148 15428
rect 15752 15376 15804 15428
rect 12072 15308 12124 15360
rect 12808 15308 12860 15360
rect 15660 15308 15712 15360
rect 17040 15351 17092 15360
rect 17040 15317 17049 15351
rect 17049 15317 17083 15351
rect 17083 15317 17092 15351
rect 17040 15308 17092 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 7564 15104 7616 15156
rect 9128 15104 9180 15156
rect 6736 15036 6788 15088
rect 5724 14900 5776 14952
rect 6644 14943 6696 14952
rect 6644 14909 6653 14943
rect 6653 14909 6687 14943
rect 6687 14909 6696 14943
rect 6644 14900 6696 14909
rect 6828 15011 6880 15020
rect 6828 14977 6837 15011
rect 6837 14977 6871 15011
rect 6871 14977 6880 15011
rect 6828 14968 6880 14977
rect 7288 15036 7340 15088
rect 7288 14943 7340 14952
rect 7288 14909 7297 14943
rect 7297 14909 7331 14943
rect 7331 14909 7340 14943
rect 7288 14900 7340 14909
rect 5908 14832 5960 14884
rect 7564 14968 7616 15020
rect 7840 15011 7892 15020
rect 7840 14977 7849 15011
rect 7849 14977 7883 15011
rect 7883 14977 7892 15011
rect 7840 14968 7892 14977
rect 9128 14968 9180 15020
rect 9588 15011 9640 15020
rect 9588 14977 9597 15011
rect 9597 14977 9631 15011
rect 9631 14977 9640 15011
rect 9588 14968 9640 14977
rect 10416 15104 10468 15156
rect 11428 15036 11480 15088
rect 11152 15011 11204 15020
rect 11152 14977 11161 15011
rect 11161 14977 11195 15011
rect 11195 14977 11204 15011
rect 11152 14968 11204 14977
rect 12072 15011 12124 15020
rect 12072 14977 12081 15011
rect 12081 14977 12115 15011
rect 12115 14977 12124 15011
rect 12072 14968 12124 14977
rect 13544 14968 13596 15020
rect 6000 14807 6052 14816
rect 6000 14773 6009 14807
rect 6009 14773 6043 14807
rect 6043 14773 6052 14807
rect 6000 14764 6052 14773
rect 6368 14807 6420 14816
rect 6368 14773 6377 14807
rect 6377 14773 6411 14807
rect 6411 14773 6420 14807
rect 6368 14764 6420 14773
rect 6552 14807 6604 14816
rect 6552 14773 6561 14807
rect 6561 14773 6595 14807
rect 6595 14773 6604 14807
rect 7472 14832 7524 14884
rect 6552 14764 6604 14773
rect 7012 14764 7064 14816
rect 7840 14832 7892 14884
rect 8300 14900 8352 14952
rect 9956 14900 10008 14952
rect 12900 14900 12952 14952
rect 13360 14900 13412 14952
rect 14096 15011 14148 15020
rect 14096 14977 14105 15011
rect 14105 14977 14139 15011
rect 14139 14977 14148 15011
rect 14096 14968 14148 14977
rect 15752 15147 15804 15156
rect 15752 15113 15761 15147
rect 15761 15113 15795 15147
rect 15795 15113 15804 15147
rect 15752 15104 15804 15113
rect 16948 15147 17000 15156
rect 16948 15113 16957 15147
rect 16957 15113 16991 15147
rect 16991 15113 17000 15147
rect 16948 15104 17000 15113
rect 15384 15079 15436 15088
rect 15384 15045 15393 15079
rect 15393 15045 15427 15079
rect 15427 15045 15436 15079
rect 15384 15036 15436 15045
rect 15292 14968 15344 15020
rect 17040 14968 17092 15020
rect 14280 14943 14332 14952
rect 14280 14909 14289 14943
rect 14289 14909 14323 14943
rect 14323 14909 14332 14943
rect 14280 14900 14332 14909
rect 8116 14764 8168 14816
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 8208 14764 8260 14773
rect 8944 14764 8996 14816
rect 11152 14764 11204 14816
rect 11336 14807 11388 14816
rect 11336 14773 11345 14807
rect 11345 14773 11379 14807
rect 11379 14773 11388 14807
rect 11336 14764 11388 14773
rect 11980 14807 12032 14816
rect 11980 14773 11989 14807
rect 11989 14773 12023 14807
rect 12023 14773 12032 14807
rect 11980 14764 12032 14773
rect 13176 14807 13228 14816
rect 13176 14773 13185 14807
rect 13185 14773 13219 14807
rect 13219 14773 13228 14807
rect 13176 14764 13228 14773
rect 13360 14764 13412 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 6184 14560 6236 14612
rect 6828 14560 6880 14612
rect 8484 14603 8536 14612
rect 8484 14569 8493 14603
rect 8493 14569 8527 14603
rect 8527 14569 8536 14603
rect 8484 14560 8536 14569
rect 8760 14560 8812 14612
rect 9588 14560 9640 14612
rect 11428 14603 11480 14612
rect 6000 14492 6052 14544
rect 11428 14569 11437 14603
rect 11437 14569 11471 14603
rect 11471 14569 11480 14603
rect 11428 14560 11480 14569
rect 11244 14492 11296 14544
rect 9404 14424 9456 14476
rect 11336 14424 11388 14476
rect 3424 14356 3476 14408
rect 7196 14356 7248 14408
rect 8208 14399 8260 14408
rect 8208 14365 8217 14399
rect 8217 14365 8251 14399
rect 8251 14365 8260 14399
rect 8208 14356 8260 14365
rect 8300 14356 8352 14408
rect 6644 14288 6696 14340
rect 8392 14288 8444 14340
rect 9220 14356 9272 14408
rect 12072 14492 12124 14544
rect 13084 14492 13136 14544
rect 11796 14424 11848 14476
rect 15200 14424 15252 14476
rect 12992 14356 13044 14408
rect 13360 14356 13412 14408
rect 8944 14331 8996 14340
rect 8944 14297 8953 14331
rect 8953 14297 8987 14331
rect 8987 14297 8996 14331
rect 8944 14288 8996 14297
rect 4620 14220 4672 14272
rect 8300 14220 8352 14272
rect 12900 14288 12952 14340
rect 14188 14288 14240 14340
rect 15660 14288 15712 14340
rect 11060 14220 11112 14272
rect 12072 14220 12124 14272
rect 13820 14263 13872 14272
rect 13820 14229 13829 14263
rect 13829 14229 13863 14263
rect 13863 14229 13872 14263
rect 13820 14220 13872 14229
rect 16764 14220 16816 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 7012 14016 7064 14068
rect 3700 13948 3752 14000
rect 3148 13880 3200 13932
rect 3332 13923 3384 13932
rect 3332 13889 3341 13923
rect 3341 13889 3375 13923
rect 3375 13889 3384 13923
rect 3332 13880 3384 13889
rect 3424 13923 3476 13932
rect 3424 13889 3433 13923
rect 3433 13889 3467 13923
rect 3467 13889 3476 13923
rect 3424 13880 3476 13889
rect 3884 13880 3936 13932
rect 4160 13880 4212 13932
rect 5908 13880 5960 13932
rect 6828 13923 6880 13932
rect 6828 13889 6837 13923
rect 6837 13889 6871 13923
rect 6871 13889 6880 13923
rect 6828 13880 6880 13889
rect 7288 13948 7340 14000
rect 8208 14016 8260 14068
rect 8024 13948 8076 14000
rect 7196 13923 7248 13932
rect 7196 13889 7205 13923
rect 7205 13889 7239 13923
rect 7239 13889 7248 13923
rect 7196 13880 7248 13889
rect 8300 13880 8352 13932
rect 8392 13923 8444 13932
rect 8392 13889 8401 13923
rect 8401 13889 8435 13923
rect 8435 13889 8444 13923
rect 8392 13880 8444 13889
rect 10232 14016 10284 14068
rect 11060 14016 11112 14068
rect 13268 14016 13320 14068
rect 9404 13948 9456 14000
rect 5448 13744 5500 13796
rect 7840 13855 7892 13864
rect 7840 13821 7849 13855
rect 7849 13821 7883 13855
rect 7883 13821 7892 13855
rect 7840 13812 7892 13821
rect 9496 13880 9548 13932
rect 11612 13948 11664 14000
rect 15660 14059 15712 14068
rect 15660 14025 15669 14059
rect 15669 14025 15703 14059
rect 15703 14025 15712 14059
rect 15660 14016 15712 14025
rect 10140 13880 10192 13932
rect 6000 13676 6052 13728
rect 6828 13676 6880 13728
rect 7104 13676 7156 13728
rect 7564 13676 7616 13728
rect 8208 13744 8260 13796
rect 8760 13855 8812 13864
rect 8760 13821 8769 13855
rect 8769 13821 8803 13855
rect 8803 13821 8812 13855
rect 8760 13812 8812 13821
rect 9864 13855 9916 13864
rect 9864 13821 9873 13855
rect 9873 13821 9907 13855
rect 9907 13821 9916 13855
rect 9864 13812 9916 13821
rect 10508 13744 10560 13796
rect 11060 13880 11112 13932
rect 13912 13923 13964 13932
rect 13912 13889 13921 13923
rect 13921 13889 13955 13923
rect 13955 13889 13964 13923
rect 13912 13880 13964 13889
rect 11612 13855 11664 13864
rect 11612 13821 11621 13855
rect 11621 13821 11655 13855
rect 11655 13821 11664 13855
rect 11612 13812 11664 13821
rect 12440 13812 12492 13864
rect 12992 13744 13044 13796
rect 14740 13880 14792 13932
rect 16764 13923 16816 13932
rect 16764 13889 16773 13923
rect 16773 13889 16807 13923
rect 16807 13889 16816 13923
rect 16764 13880 16816 13889
rect 15752 13812 15804 13864
rect 15108 13744 15160 13796
rect 9220 13676 9272 13728
rect 9312 13719 9364 13728
rect 9312 13685 9321 13719
rect 9321 13685 9355 13719
rect 9355 13685 9364 13719
rect 9312 13676 9364 13685
rect 9588 13676 9640 13728
rect 9772 13676 9824 13728
rect 10876 13676 10928 13728
rect 11336 13676 11388 13728
rect 13820 13676 13872 13728
rect 15016 13676 15068 13728
rect 16948 13719 17000 13728
rect 16948 13685 16957 13719
rect 16957 13685 16991 13719
rect 16991 13685 17000 13719
rect 16948 13676 17000 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 4068 13404 4120 13456
rect 3148 13268 3200 13320
rect 3516 13336 3568 13388
rect 4712 13472 4764 13524
rect 4344 13404 4396 13456
rect 5448 13515 5500 13524
rect 5448 13481 5457 13515
rect 5457 13481 5491 13515
rect 5491 13481 5500 13515
rect 5448 13472 5500 13481
rect 3608 13268 3660 13320
rect 4068 13268 4120 13320
rect 5172 13336 5224 13388
rect 4344 13268 4396 13320
rect 4620 13311 4672 13320
rect 4620 13277 4629 13311
rect 4629 13277 4663 13311
rect 4663 13277 4672 13311
rect 4620 13268 4672 13277
rect 4712 13268 4764 13320
rect 5540 13404 5592 13456
rect 5816 13404 5868 13456
rect 6276 13404 6328 13456
rect 7012 13515 7064 13524
rect 7012 13481 7021 13515
rect 7021 13481 7055 13515
rect 7055 13481 7064 13515
rect 7012 13472 7064 13481
rect 7104 13472 7156 13524
rect 7840 13472 7892 13524
rect 8024 13515 8076 13524
rect 8024 13481 8033 13515
rect 8033 13481 8067 13515
rect 8067 13481 8076 13515
rect 8024 13472 8076 13481
rect 9772 13515 9824 13524
rect 6920 13404 6972 13456
rect 7288 13336 7340 13388
rect 3240 13243 3292 13252
rect 3240 13209 3249 13243
rect 3249 13209 3283 13243
rect 3283 13209 3292 13243
rect 3240 13200 3292 13209
rect 3792 13243 3844 13252
rect 3792 13209 3801 13243
rect 3801 13209 3835 13243
rect 3835 13209 3844 13243
rect 3792 13200 3844 13209
rect 3424 13132 3476 13184
rect 4160 13175 4212 13184
rect 4160 13141 4169 13175
rect 4169 13141 4203 13175
rect 4203 13141 4212 13175
rect 4160 13132 4212 13141
rect 4712 13132 4764 13184
rect 5356 13132 5408 13184
rect 6000 13311 6052 13320
rect 6000 13277 6009 13311
rect 6009 13277 6043 13311
rect 6043 13277 6052 13311
rect 6000 13268 6052 13277
rect 6460 13311 6512 13320
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 6092 13200 6144 13252
rect 6276 13243 6328 13252
rect 6276 13209 6285 13243
rect 6285 13209 6319 13243
rect 6319 13209 6328 13243
rect 6276 13200 6328 13209
rect 6736 13268 6788 13320
rect 7196 13268 7248 13320
rect 7564 13311 7616 13320
rect 7564 13277 7571 13311
rect 7571 13277 7616 13311
rect 7564 13268 7616 13277
rect 7748 13336 7800 13388
rect 6644 13200 6696 13252
rect 8024 13200 8076 13252
rect 6828 13175 6880 13184
rect 6828 13141 6837 13175
rect 6837 13141 6871 13175
rect 6871 13141 6880 13175
rect 6828 13132 6880 13141
rect 7012 13132 7064 13184
rect 9772 13481 9781 13515
rect 9781 13481 9815 13515
rect 9815 13481 9824 13515
rect 9772 13472 9824 13481
rect 10048 13472 10100 13524
rect 10508 13515 10560 13524
rect 10508 13481 10517 13515
rect 10517 13481 10551 13515
rect 10551 13481 10560 13515
rect 10508 13472 10560 13481
rect 12440 13472 12492 13524
rect 12992 13515 13044 13524
rect 12992 13481 13001 13515
rect 13001 13481 13035 13515
rect 13035 13481 13044 13515
rect 12992 13472 13044 13481
rect 13268 13472 13320 13524
rect 15200 13472 15252 13524
rect 9680 13336 9732 13388
rect 10048 13336 10100 13388
rect 10416 13336 10468 13388
rect 8208 13268 8260 13320
rect 9588 13311 9640 13320
rect 9588 13277 9597 13311
rect 9597 13277 9631 13311
rect 9631 13277 9640 13311
rect 9588 13268 9640 13277
rect 9772 13311 9824 13320
rect 9772 13277 9781 13311
rect 9781 13277 9815 13311
rect 9815 13277 9824 13311
rect 9772 13268 9824 13277
rect 10416 13243 10468 13252
rect 10416 13209 10425 13243
rect 10425 13209 10459 13243
rect 10459 13209 10468 13243
rect 10416 13200 10468 13209
rect 14004 13404 14056 13456
rect 12624 13379 12676 13388
rect 12624 13345 12633 13379
rect 12633 13345 12667 13379
rect 12667 13345 12676 13379
rect 12624 13336 12676 13345
rect 14280 13379 14332 13388
rect 14280 13345 14289 13379
rect 14289 13345 14323 13379
rect 14323 13345 14332 13379
rect 14280 13336 14332 13345
rect 15660 13379 15712 13388
rect 15660 13345 15669 13379
rect 15669 13345 15703 13379
rect 15703 13345 15712 13379
rect 15660 13336 15712 13345
rect 12532 13311 12584 13320
rect 12532 13277 12541 13311
rect 12541 13277 12575 13311
rect 12575 13277 12584 13311
rect 12532 13268 12584 13277
rect 12808 13311 12860 13320
rect 12808 13277 12817 13311
rect 12817 13277 12851 13311
rect 12851 13277 12860 13311
rect 12808 13268 12860 13277
rect 14464 13268 14516 13320
rect 15016 13311 15068 13320
rect 15016 13277 15025 13311
rect 15025 13277 15059 13311
rect 15059 13277 15068 13311
rect 15016 13268 15068 13277
rect 15384 13311 15436 13320
rect 15384 13277 15393 13311
rect 15393 13277 15427 13311
rect 15427 13277 15436 13311
rect 15384 13268 15436 13277
rect 9220 13132 9272 13184
rect 13268 13200 13320 13252
rect 14096 13243 14148 13252
rect 14096 13209 14105 13243
rect 14105 13209 14139 13243
rect 14139 13209 14148 13243
rect 14096 13200 14148 13209
rect 15200 13243 15252 13252
rect 15200 13209 15209 13243
rect 15209 13209 15243 13243
rect 15243 13209 15252 13243
rect 15200 13200 15252 13209
rect 15292 13243 15344 13252
rect 15292 13209 15301 13243
rect 15301 13209 15335 13243
rect 15335 13209 15344 13243
rect 15292 13200 15344 13209
rect 10692 13132 10744 13184
rect 12900 13132 12952 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 3792 12971 3844 12980
rect 3792 12937 3801 12971
rect 3801 12937 3835 12971
rect 3835 12937 3844 12971
rect 3792 12928 3844 12937
rect 4528 12928 4580 12980
rect 2872 12860 2924 12912
rect 5356 12860 5408 12912
rect 3056 12792 3108 12844
rect 3332 12792 3384 12844
rect 3608 12835 3660 12844
rect 3608 12801 3617 12835
rect 3617 12801 3651 12835
rect 3651 12801 3660 12835
rect 3608 12792 3660 12801
rect 4712 12835 4764 12844
rect 4712 12801 4721 12835
rect 4721 12801 4755 12835
rect 4755 12801 4764 12835
rect 4712 12792 4764 12801
rect 4620 12724 4672 12776
rect 5172 12792 5224 12844
rect 6092 12928 6144 12980
rect 6276 12860 6328 12912
rect 7012 12860 7064 12912
rect 7564 12928 7616 12980
rect 8208 12928 8260 12980
rect 10508 12928 10560 12980
rect 8760 12860 8812 12912
rect 10692 12860 10744 12912
rect 5632 12724 5684 12776
rect 5816 12835 5868 12844
rect 5816 12801 5825 12835
rect 5825 12801 5859 12835
rect 5859 12801 5868 12835
rect 5816 12792 5868 12801
rect 6092 12792 6144 12844
rect 6460 12792 6512 12844
rect 7104 12835 7156 12844
rect 7104 12801 7113 12835
rect 7113 12801 7147 12835
rect 7147 12801 7156 12835
rect 7104 12792 7156 12801
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 7380 12835 7432 12844
rect 7380 12801 7389 12835
rect 7389 12801 7423 12835
rect 7423 12801 7432 12835
rect 7380 12792 7432 12801
rect 7840 12792 7892 12844
rect 10508 12792 10560 12844
rect 10876 12792 10928 12844
rect 8024 12724 8076 12776
rect 8944 12724 8996 12776
rect 12440 12928 12492 12980
rect 12532 12928 12584 12980
rect 12348 12903 12400 12912
rect 12348 12869 12357 12903
rect 12357 12869 12391 12903
rect 12391 12869 12400 12903
rect 12348 12860 12400 12869
rect 14096 12928 14148 12980
rect 14372 12928 14424 12980
rect 15384 12928 15436 12980
rect 16948 12971 17000 12980
rect 16948 12937 16957 12971
rect 16957 12937 16991 12971
rect 16991 12937 17000 12971
rect 16948 12928 17000 12937
rect 12440 12792 12492 12844
rect 12808 12792 12860 12844
rect 12900 12835 12952 12844
rect 12900 12801 12909 12835
rect 12909 12801 12943 12835
rect 12943 12801 12952 12835
rect 12900 12792 12952 12801
rect 15568 12860 15620 12912
rect 15752 12860 15804 12912
rect 13084 12792 13136 12844
rect 14464 12835 14516 12844
rect 14464 12801 14473 12835
rect 14473 12801 14507 12835
rect 14507 12801 14516 12835
rect 14464 12792 14516 12801
rect 7564 12656 7616 12708
rect 7932 12656 7984 12708
rect 9220 12656 9272 12708
rect 11428 12656 11480 12708
rect 6000 12588 6052 12640
rect 6276 12588 6328 12640
rect 12164 12588 12216 12640
rect 13268 12699 13320 12708
rect 13268 12665 13277 12699
rect 13277 12665 13311 12699
rect 13311 12665 13320 12699
rect 13268 12656 13320 12665
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 5724 12384 5776 12436
rect 6276 12384 6328 12436
rect 2596 12155 2648 12164
rect 2596 12121 2605 12155
rect 2605 12121 2639 12155
rect 2639 12121 2648 12155
rect 2596 12112 2648 12121
rect 2780 12223 2832 12232
rect 2780 12189 2789 12223
rect 2789 12189 2823 12223
rect 2823 12189 2832 12223
rect 2780 12180 2832 12189
rect 3884 12248 3936 12300
rect 2872 12112 2924 12164
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 3608 12180 3660 12232
rect 4620 12223 4672 12232
rect 4620 12189 4629 12223
rect 4629 12189 4663 12223
rect 4663 12189 4672 12223
rect 4620 12180 4672 12189
rect 6368 12316 6420 12368
rect 6828 12248 6880 12300
rect 7656 12384 7708 12436
rect 7932 12427 7984 12436
rect 7932 12393 7941 12427
rect 7941 12393 7975 12427
rect 7975 12393 7984 12427
rect 7932 12384 7984 12393
rect 8484 12384 8536 12436
rect 9220 12427 9272 12436
rect 9220 12393 9229 12427
rect 9229 12393 9263 12427
rect 9263 12393 9272 12427
rect 9220 12384 9272 12393
rect 9404 12316 9456 12368
rect 3056 12044 3108 12096
rect 4344 12112 4396 12164
rect 4436 12155 4488 12164
rect 4436 12121 4445 12155
rect 4445 12121 4479 12155
rect 4479 12121 4488 12155
rect 4436 12112 4488 12121
rect 4712 12112 4764 12164
rect 5080 12155 5132 12164
rect 5080 12121 5089 12155
rect 5089 12121 5123 12155
rect 5123 12121 5132 12155
rect 5080 12112 5132 12121
rect 5172 12155 5224 12164
rect 5172 12121 5181 12155
rect 5181 12121 5215 12155
rect 5215 12121 5224 12155
rect 5172 12112 5224 12121
rect 6368 12112 6420 12164
rect 4528 12044 4580 12096
rect 5264 12044 5316 12096
rect 6000 12044 6052 12096
rect 6460 12044 6512 12096
rect 6920 12223 6972 12232
rect 6920 12189 6929 12223
rect 6929 12189 6963 12223
rect 6963 12189 6972 12223
rect 6920 12180 6972 12189
rect 7104 12180 7156 12232
rect 7288 12223 7340 12232
rect 7288 12189 7297 12223
rect 7297 12189 7331 12223
rect 7331 12189 7340 12223
rect 7288 12180 7340 12189
rect 7380 12223 7432 12232
rect 7380 12189 7390 12223
rect 7390 12189 7424 12223
rect 7424 12189 7432 12223
rect 7380 12180 7432 12189
rect 7196 12112 7248 12164
rect 7656 12155 7708 12164
rect 7656 12121 7665 12155
rect 7665 12121 7699 12155
rect 7699 12121 7708 12155
rect 7656 12112 7708 12121
rect 7012 12044 7064 12096
rect 7104 12044 7156 12096
rect 8484 12248 8536 12300
rect 9220 12248 9272 12300
rect 10692 12384 10744 12436
rect 10876 12384 10928 12436
rect 12532 12427 12584 12436
rect 12532 12393 12541 12427
rect 12541 12393 12575 12427
rect 12575 12393 12584 12427
rect 12532 12384 12584 12393
rect 10968 12316 11020 12368
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 8944 12180 8996 12232
rect 8484 12112 8536 12164
rect 9036 12155 9088 12164
rect 9036 12121 9045 12155
rect 9045 12121 9079 12155
rect 9079 12121 9088 12155
rect 9036 12112 9088 12121
rect 9588 12155 9640 12164
rect 9588 12121 9597 12155
rect 9597 12121 9631 12155
rect 9631 12121 9640 12155
rect 9588 12112 9640 12121
rect 9772 12180 9824 12232
rect 9772 12044 9824 12096
rect 10600 12223 10652 12232
rect 10600 12189 10609 12223
rect 10609 12189 10643 12223
rect 10643 12189 10652 12223
rect 10600 12180 10652 12189
rect 11060 12223 11112 12232
rect 11060 12189 11069 12223
rect 11069 12189 11103 12223
rect 11103 12189 11112 12223
rect 11060 12180 11112 12189
rect 11152 12223 11204 12232
rect 11152 12189 11161 12223
rect 11161 12189 11195 12223
rect 11195 12189 11204 12223
rect 11152 12180 11204 12189
rect 11520 12248 11572 12300
rect 12164 12248 12216 12300
rect 12440 12291 12492 12300
rect 12440 12257 12449 12291
rect 12449 12257 12483 12291
rect 12483 12257 12492 12291
rect 12440 12248 12492 12257
rect 13268 12248 13320 12300
rect 11428 12223 11480 12232
rect 11428 12189 11444 12223
rect 11444 12189 11478 12223
rect 11478 12189 11480 12223
rect 11428 12180 11480 12189
rect 12072 12180 12124 12232
rect 12532 12223 12584 12232
rect 12532 12189 12541 12223
rect 12541 12189 12575 12223
rect 12575 12189 12584 12223
rect 12532 12180 12584 12189
rect 15108 12180 15160 12232
rect 15568 12248 15620 12300
rect 15384 12223 15436 12232
rect 15384 12189 15393 12223
rect 15393 12189 15427 12223
rect 15427 12189 15436 12223
rect 15384 12180 15436 12189
rect 15660 12223 15712 12232
rect 15660 12189 15669 12223
rect 15669 12189 15703 12223
rect 15703 12189 15712 12223
rect 15660 12180 15712 12189
rect 15752 12180 15804 12232
rect 10692 12044 10744 12096
rect 11336 12087 11388 12096
rect 11336 12053 11345 12087
rect 11345 12053 11379 12087
rect 11379 12053 11388 12087
rect 11336 12044 11388 12053
rect 14648 12112 14700 12164
rect 12716 12087 12768 12096
rect 12716 12053 12725 12087
rect 12725 12053 12759 12087
rect 12759 12053 12768 12087
rect 12716 12044 12768 12053
rect 15476 12044 15528 12096
rect 16580 12044 16632 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 3240 11840 3292 11892
rect 3792 11883 3844 11892
rect 3792 11849 3801 11883
rect 3801 11849 3835 11883
rect 3835 11849 3844 11883
rect 3792 11840 3844 11849
rect 4620 11840 4672 11892
rect 3884 11772 3936 11824
rect 3332 11704 3384 11756
rect 3516 11747 3568 11756
rect 3516 11713 3525 11747
rect 3525 11713 3559 11747
rect 3559 11713 3568 11747
rect 3516 11704 3568 11713
rect 3608 11747 3660 11756
rect 3608 11713 3617 11747
rect 3617 11713 3651 11747
rect 3651 11713 3660 11747
rect 3608 11704 3660 11713
rect 4344 11704 4396 11756
rect 4620 11704 4672 11756
rect 5356 11840 5408 11892
rect 6276 11840 6328 11892
rect 6736 11840 6788 11892
rect 5448 11704 5500 11756
rect 7196 11840 7248 11892
rect 7288 11840 7340 11892
rect 12532 11840 12584 11892
rect 7380 11772 7432 11824
rect 8116 11772 8168 11824
rect 14372 11840 14424 11892
rect 15384 11840 15436 11892
rect 4804 11636 4856 11688
rect 5908 11636 5960 11688
rect 7104 11704 7156 11756
rect 8668 11747 8720 11756
rect 8668 11713 8677 11747
rect 8677 11713 8711 11747
rect 8711 11713 8720 11747
rect 8668 11704 8720 11713
rect 8944 11704 8996 11756
rect 9036 11747 9088 11756
rect 9036 11713 9045 11747
rect 9045 11713 9079 11747
rect 9079 11713 9088 11747
rect 9036 11704 9088 11713
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 4436 11568 4488 11620
rect 7288 11636 7340 11688
rect 7472 11611 7524 11620
rect 7472 11577 7481 11611
rect 7481 11577 7515 11611
rect 7515 11577 7524 11611
rect 7472 11568 7524 11577
rect 7656 11568 7708 11620
rect 8484 11636 8536 11688
rect 9680 11636 9732 11688
rect 10324 11636 10376 11688
rect 14464 11815 14516 11824
rect 14464 11781 14473 11815
rect 14473 11781 14507 11815
rect 14507 11781 14516 11815
rect 14464 11772 14516 11781
rect 12256 11704 12308 11756
rect 9036 11568 9088 11620
rect 2596 11500 2648 11552
rect 5908 11500 5960 11552
rect 6000 11500 6052 11552
rect 10140 11500 10192 11552
rect 10968 11636 11020 11688
rect 10692 11500 10744 11552
rect 11520 11568 11572 11620
rect 13728 11704 13780 11756
rect 14372 11704 14424 11756
rect 15016 11747 15068 11756
rect 15016 11713 15025 11747
rect 15025 11713 15059 11747
rect 15059 11713 15068 11747
rect 15016 11704 15068 11713
rect 16580 11704 16632 11756
rect 16764 11704 16816 11756
rect 13452 11636 13504 11688
rect 14464 11636 14516 11688
rect 15292 11636 15344 11688
rect 14096 11568 14148 11620
rect 11336 11500 11388 11552
rect 13728 11543 13780 11552
rect 13728 11509 13737 11543
rect 13737 11509 13771 11543
rect 13771 11509 13780 11543
rect 13728 11500 13780 11509
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 14004 11500 14056 11552
rect 14924 11543 14976 11552
rect 14924 11509 14933 11543
rect 14933 11509 14967 11543
rect 14967 11509 14976 11543
rect 14924 11500 14976 11509
rect 15016 11543 15068 11552
rect 15016 11509 15025 11543
rect 15025 11509 15059 11543
rect 15059 11509 15068 11543
rect 15016 11500 15068 11509
rect 15108 11500 15160 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 3608 11296 3660 11348
rect 7380 11296 7432 11348
rect 7656 11296 7708 11348
rect 8116 11296 8168 11348
rect 10324 11296 10376 11348
rect 10508 11296 10560 11348
rect 6184 11228 6236 11280
rect 6460 11228 6512 11280
rect 7288 11228 7340 11280
rect 3884 11160 3936 11212
rect 4528 11092 4580 11144
rect 5264 11092 5316 11144
rect 5540 11092 5592 11144
rect 6276 11092 6328 11144
rect 6736 11092 6788 11144
rect 6920 11092 6972 11144
rect 7564 11160 7616 11212
rect 7472 11135 7524 11144
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 8024 11228 8076 11280
rect 4620 11024 4672 11076
rect 5632 11067 5684 11076
rect 5632 11033 5641 11067
rect 5641 11033 5675 11067
rect 5675 11033 5684 11067
rect 5632 11024 5684 11033
rect 7840 11024 7892 11076
rect 5356 10999 5408 11008
rect 5356 10965 5365 10999
rect 5365 10965 5399 10999
rect 5399 10965 5408 10999
rect 5356 10956 5408 10965
rect 7104 10956 7156 11008
rect 9772 11160 9824 11212
rect 10508 11160 10560 11212
rect 12532 11296 12584 11348
rect 12808 11296 12860 11348
rect 12900 11296 12952 11348
rect 13820 11296 13872 11348
rect 14004 11296 14056 11348
rect 15016 11296 15068 11348
rect 12072 11228 12124 11280
rect 13176 11228 13228 11280
rect 15200 11160 15252 11212
rect 15660 11203 15712 11212
rect 15660 11169 15669 11203
rect 15669 11169 15703 11203
rect 15703 11169 15712 11203
rect 15660 11160 15712 11169
rect 12900 11092 12952 11144
rect 13084 11135 13136 11144
rect 13084 11101 13093 11135
rect 13093 11101 13127 11135
rect 13127 11101 13136 11135
rect 13084 11092 13136 11101
rect 13176 11135 13228 11144
rect 13176 11101 13185 11135
rect 13185 11101 13219 11135
rect 13219 11101 13228 11135
rect 13176 11092 13228 11101
rect 13728 11092 13780 11144
rect 8116 11067 8168 11076
rect 8116 11033 8125 11067
rect 8125 11033 8159 11067
rect 8159 11033 8168 11067
rect 8116 11024 8168 11033
rect 8852 11024 8904 11076
rect 8944 10956 8996 11008
rect 9404 11024 9456 11076
rect 10324 11024 10376 11076
rect 10600 11024 10652 11076
rect 12072 11067 12124 11076
rect 12072 11033 12081 11067
rect 12081 11033 12115 11067
rect 12115 11033 12124 11067
rect 12072 11024 12124 11033
rect 12256 11067 12308 11076
rect 12256 11033 12265 11067
rect 12265 11033 12299 11067
rect 12299 11033 12308 11067
rect 12256 11024 12308 11033
rect 13820 11024 13872 11076
rect 14924 11092 14976 11144
rect 15292 11135 15344 11144
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 15108 11024 15160 11076
rect 15292 10956 15344 11008
rect 16580 10956 16632 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 3884 10684 3936 10736
rect 4528 10752 4580 10804
rect 5080 10752 5132 10804
rect 5356 10684 5408 10736
rect 5540 10684 5592 10736
rect 7472 10752 7524 10804
rect 2872 10616 2924 10668
rect 3056 10659 3108 10668
rect 3056 10625 3065 10659
rect 3065 10625 3099 10659
rect 3099 10625 3108 10659
rect 3056 10616 3108 10625
rect 3424 10659 3476 10668
rect 3424 10625 3433 10659
rect 3433 10625 3467 10659
rect 3467 10625 3476 10659
rect 3424 10616 3476 10625
rect 3516 10616 3568 10668
rect 3976 10616 4028 10668
rect 4436 10659 4488 10668
rect 4436 10625 4445 10659
rect 4445 10625 4479 10659
rect 4479 10625 4488 10659
rect 4436 10616 4488 10625
rect 4712 10616 4764 10668
rect 5264 10659 5316 10668
rect 5264 10625 5273 10659
rect 5273 10625 5307 10659
rect 5307 10625 5316 10659
rect 5264 10616 5316 10625
rect 6920 10616 6972 10668
rect 7656 10727 7708 10736
rect 7656 10693 7665 10727
rect 7665 10693 7699 10727
rect 7699 10693 7708 10727
rect 7656 10684 7708 10693
rect 8116 10684 8168 10736
rect 8576 10727 8628 10736
rect 8576 10693 8585 10727
rect 8585 10693 8619 10727
rect 8619 10693 8628 10727
rect 8576 10684 8628 10693
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 7288 10616 7340 10668
rect 7380 10616 7432 10668
rect 7748 10659 7800 10668
rect 7748 10625 7757 10659
rect 7757 10625 7791 10659
rect 7791 10625 7800 10659
rect 7748 10616 7800 10625
rect 8024 10616 8076 10668
rect 10600 10752 10652 10804
rect 15384 10752 15436 10804
rect 17224 10752 17276 10804
rect 10140 10684 10192 10736
rect 9772 10616 9824 10668
rect 12716 10684 12768 10736
rect 4620 10480 4672 10532
rect 3516 10412 3568 10464
rect 7656 10548 7708 10600
rect 10324 10591 10376 10600
rect 10324 10557 10333 10591
rect 10333 10557 10367 10591
rect 10367 10557 10376 10591
rect 10324 10548 10376 10557
rect 10692 10616 10744 10668
rect 10968 10616 11020 10668
rect 8116 10480 8168 10532
rect 12072 10616 12124 10668
rect 13544 10659 13596 10668
rect 13544 10625 13553 10659
rect 13553 10625 13587 10659
rect 13587 10625 13596 10659
rect 13544 10616 13596 10625
rect 16580 10616 16632 10668
rect 16672 10616 16724 10668
rect 5080 10412 5132 10464
rect 5724 10412 5776 10464
rect 8668 10412 8720 10464
rect 9312 10412 9364 10464
rect 10600 10455 10652 10464
rect 10600 10421 10609 10455
rect 10609 10421 10643 10455
rect 10643 10421 10652 10455
rect 10600 10412 10652 10421
rect 10876 10412 10928 10464
rect 13176 10548 13228 10600
rect 13728 10548 13780 10600
rect 14280 10480 14332 10532
rect 12808 10412 12860 10464
rect 14556 10412 14608 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 3424 10208 3476 10260
rect 4068 10208 4120 10260
rect 2228 10004 2280 10056
rect 4712 10140 4764 10192
rect 4988 10183 5040 10192
rect 4988 10149 4997 10183
rect 4997 10149 5031 10183
rect 5031 10149 5040 10183
rect 4988 10140 5040 10149
rect 4160 10047 4212 10056
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 5448 10072 5500 10124
rect 2136 9979 2188 9988
rect 2136 9945 2145 9979
rect 2145 9945 2179 9979
rect 2179 9945 2188 9979
rect 2136 9936 2188 9945
rect 2320 9936 2372 9988
rect 3976 9979 4028 9988
rect 3976 9945 3985 9979
rect 3985 9945 4019 9979
rect 4019 9945 4028 9979
rect 3976 9936 4028 9945
rect 5540 10004 5592 10056
rect 5908 10140 5960 10192
rect 6644 10140 6696 10192
rect 7104 10208 7156 10260
rect 9496 10251 9548 10260
rect 9496 10217 9505 10251
rect 9505 10217 9539 10251
rect 9539 10217 9548 10251
rect 9496 10208 9548 10217
rect 10968 10208 11020 10260
rect 11060 10208 11112 10260
rect 12624 10208 12676 10260
rect 6276 10072 6328 10124
rect 8668 10140 8720 10192
rect 8760 10140 8812 10192
rect 13912 10208 13964 10260
rect 14280 10208 14332 10260
rect 16948 10251 17000 10260
rect 16948 10217 16957 10251
rect 16957 10217 16991 10251
rect 16991 10217 17000 10251
rect 16948 10208 17000 10217
rect 5908 10047 5960 10056
rect 5908 10013 5917 10047
rect 5917 10013 5951 10047
rect 5951 10013 5960 10047
rect 5908 10004 5960 10013
rect 2688 9868 2740 9920
rect 4344 9911 4396 9920
rect 4344 9877 4353 9911
rect 4353 9877 4387 9911
rect 4387 9877 4396 9911
rect 4344 9868 4396 9877
rect 4712 9979 4764 9988
rect 4712 9945 4721 9979
rect 4721 9945 4755 9979
rect 4755 9945 4764 9979
rect 4712 9936 4764 9945
rect 4804 9868 4856 9920
rect 5448 9936 5500 9988
rect 6184 10047 6236 10056
rect 6184 10013 6193 10047
rect 6193 10013 6227 10047
rect 6227 10013 6236 10047
rect 6184 10004 6236 10013
rect 9496 10072 9548 10124
rect 10692 10072 10744 10124
rect 5908 9868 5960 9920
rect 6460 10004 6512 10056
rect 6828 9979 6880 9988
rect 6828 9945 6837 9979
rect 6837 9945 6871 9979
rect 6871 9945 6880 9979
rect 6828 9936 6880 9945
rect 6460 9868 6512 9920
rect 6736 9911 6788 9920
rect 6736 9877 6745 9911
rect 6745 9877 6779 9911
rect 6779 9877 6788 9911
rect 6736 9868 6788 9877
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 7104 10004 7156 10056
rect 7380 10047 7432 10056
rect 7380 10013 7389 10047
rect 7389 10013 7423 10047
rect 7423 10013 7432 10047
rect 7380 10004 7432 10013
rect 7472 10004 7524 10056
rect 8300 10004 8352 10056
rect 8484 10004 8536 10056
rect 9220 10047 9272 10056
rect 9220 10013 9229 10047
rect 9229 10013 9263 10047
rect 9263 10013 9272 10047
rect 9220 10004 9272 10013
rect 9312 10004 9364 10056
rect 10968 10072 11020 10124
rect 12164 10072 12216 10124
rect 12716 10072 12768 10124
rect 14648 10115 14700 10124
rect 14648 10081 14657 10115
rect 14657 10081 14691 10115
rect 14691 10081 14700 10115
rect 14648 10072 14700 10081
rect 7196 9979 7248 9988
rect 7196 9945 7205 9979
rect 7205 9945 7239 9979
rect 7239 9945 7248 9979
rect 7196 9936 7248 9945
rect 8116 9936 8168 9988
rect 10968 9936 11020 9988
rect 8852 9868 8904 9920
rect 9680 9868 9732 9920
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 13452 10047 13504 10056
rect 13452 10013 13461 10047
rect 13461 10013 13495 10047
rect 13495 10013 13504 10047
rect 13452 10004 13504 10013
rect 13636 10004 13688 10056
rect 14556 10047 14608 10056
rect 14556 10013 14565 10047
rect 14565 10013 14599 10047
rect 14599 10013 14608 10047
rect 14556 10004 14608 10013
rect 16396 10047 16448 10056
rect 16396 10013 16405 10047
rect 16405 10013 16439 10047
rect 16439 10013 16448 10047
rect 16396 10004 16448 10013
rect 16580 10004 16632 10056
rect 11152 9936 11204 9988
rect 11520 9979 11572 9988
rect 11520 9945 11529 9979
rect 11529 9945 11563 9979
rect 11563 9945 11572 9979
rect 11520 9936 11572 9945
rect 11888 9979 11940 9988
rect 11888 9945 11897 9979
rect 11897 9945 11931 9979
rect 11931 9945 11940 9979
rect 11888 9936 11940 9945
rect 12992 9979 13044 9988
rect 12992 9945 13001 9979
rect 13001 9945 13035 9979
rect 13035 9945 13044 9979
rect 12992 9936 13044 9945
rect 13268 9979 13320 9988
rect 13268 9945 13277 9979
rect 13277 9945 13311 9979
rect 13311 9945 13320 9979
rect 13268 9936 13320 9945
rect 13084 9868 13136 9920
rect 14096 9868 14148 9920
rect 15016 9868 15068 9920
rect 16488 9868 16540 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 2136 9664 2188 9716
rect 3516 9664 3568 9716
rect 4344 9664 4396 9716
rect 2228 9596 2280 9648
rect 5724 9596 5776 9648
rect 6276 9596 6328 9648
rect 7104 9664 7156 9716
rect 7380 9664 7432 9716
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 2688 9528 2740 9580
rect 6644 9571 6696 9580
rect 6644 9537 6653 9571
rect 6653 9537 6687 9571
rect 6687 9537 6696 9571
rect 7564 9639 7616 9648
rect 7564 9605 7573 9639
rect 7573 9605 7607 9639
rect 7607 9605 7616 9639
rect 7564 9596 7616 9605
rect 7656 9639 7708 9648
rect 7656 9605 7665 9639
rect 7665 9605 7699 9639
rect 7699 9605 7708 9639
rect 7656 9596 7708 9605
rect 6644 9528 6696 9537
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 3976 9460 4028 9512
rect 5724 9503 5776 9512
rect 5724 9469 5733 9503
rect 5733 9469 5767 9503
rect 5767 9469 5776 9503
rect 5724 9460 5776 9469
rect 4620 9392 4672 9444
rect 6552 9460 6604 9512
rect 6920 9460 6972 9512
rect 7932 9528 7984 9580
rect 8300 9639 8352 9648
rect 8300 9605 8309 9639
rect 8309 9605 8343 9639
rect 8343 9605 8352 9639
rect 8300 9596 8352 9605
rect 8668 9664 8720 9716
rect 9220 9639 9272 9648
rect 9220 9605 9229 9639
rect 9229 9605 9263 9639
rect 9263 9605 9272 9639
rect 9220 9596 9272 9605
rect 10416 9596 10468 9648
rect 10968 9596 11020 9648
rect 12992 9664 13044 9716
rect 12808 9596 12860 9648
rect 13268 9596 13320 9648
rect 8392 9571 8444 9580
rect 8392 9537 8401 9571
rect 8401 9537 8435 9571
rect 8435 9537 8444 9571
rect 8392 9528 8444 9537
rect 7012 9392 7064 9444
rect 5356 9324 5408 9376
rect 6644 9367 6696 9376
rect 6644 9333 6653 9367
rect 6653 9333 6687 9367
rect 6687 9333 6696 9367
rect 6644 9324 6696 9333
rect 6736 9324 6788 9376
rect 8852 9528 8904 9580
rect 8944 9571 8996 9580
rect 8944 9537 8953 9571
rect 8953 9537 8987 9571
rect 8987 9537 8996 9571
rect 8944 9528 8996 9537
rect 9128 9528 9180 9580
rect 8576 9367 8628 9376
rect 8576 9333 8585 9367
rect 8585 9333 8619 9367
rect 8619 9333 8628 9367
rect 8576 9324 8628 9333
rect 8668 9367 8720 9376
rect 8668 9333 8677 9367
rect 8677 9333 8711 9367
rect 8711 9333 8720 9367
rect 8668 9324 8720 9333
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 9220 9460 9272 9512
rect 9956 9503 10008 9512
rect 9956 9469 9965 9503
rect 9965 9469 9999 9503
rect 9999 9469 10008 9503
rect 9956 9460 10008 9469
rect 9312 9392 9364 9444
rect 10232 9392 10284 9444
rect 13176 9528 13228 9580
rect 13912 9528 13964 9580
rect 15200 9528 15252 9580
rect 16120 9528 16172 9580
rect 10784 9460 10836 9512
rect 11152 9460 11204 9512
rect 14188 9460 14240 9512
rect 14648 9503 14700 9512
rect 14648 9469 14657 9503
rect 14657 9469 14691 9503
rect 14691 9469 14700 9503
rect 14648 9460 14700 9469
rect 11244 9435 11296 9444
rect 11244 9401 11253 9435
rect 11253 9401 11287 9435
rect 11287 9401 11296 9435
rect 11244 9392 11296 9401
rect 9772 9324 9824 9376
rect 10140 9324 10192 9376
rect 10876 9324 10928 9376
rect 11428 9324 11480 9376
rect 14740 9367 14792 9376
rect 14740 9333 14749 9367
rect 14749 9333 14783 9367
rect 14783 9333 14792 9367
rect 14740 9324 14792 9333
rect 14924 9367 14976 9376
rect 14924 9333 14933 9367
rect 14933 9333 14967 9367
rect 14967 9333 14976 9367
rect 14924 9324 14976 9333
rect 16488 9367 16540 9376
rect 16488 9333 16497 9367
rect 16497 9333 16531 9367
rect 16531 9333 16540 9367
rect 16488 9324 16540 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 6184 9120 6236 9172
rect 6368 9120 6420 9172
rect 6644 9120 6696 9172
rect 8760 9120 8812 9172
rect 9036 9120 9088 9172
rect 9220 9120 9272 9172
rect 2688 8984 2740 9036
rect 2228 8959 2280 8968
rect 2228 8925 2237 8959
rect 2237 8925 2271 8959
rect 2271 8925 2280 8959
rect 3976 9052 4028 9104
rect 3608 8984 3660 9036
rect 2228 8916 2280 8925
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 3332 8959 3384 8968
rect 3332 8925 3341 8959
rect 3341 8925 3375 8959
rect 3375 8925 3384 8959
rect 3332 8916 3384 8925
rect 3424 8916 3476 8968
rect 4804 8916 4856 8968
rect 5448 8984 5500 9036
rect 2136 8848 2188 8900
rect 2412 8891 2464 8900
rect 2412 8857 2421 8891
rect 2421 8857 2455 8891
rect 2455 8857 2464 8891
rect 2412 8848 2464 8857
rect 3056 8780 3108 8832
rect 3700 8848 3752 8900
rect 4620 8848 4672 8900
rect 5632 8916 5684 8968
rect 5816 8984 5868 9036
rect 8944 9052 8996 9104
rect 5908 8959 5960 8968
rect 5908 8925 5917 8959
rect 5917 8925 5951 8959
rect 5951 8925 5960 8959
rect 5908 8916 5960 8925
rect 3884 8780 3936 8832
rect 4160 8823 4212 8832
rect 4160 8789 4169 8823
rect 4169 8789 4203 8823
rect 4203 8789 4212 8823
rect 4160 8780 4212 8789
rect 5448 8848 5500 8900
rect 6276 8916 6328 8968
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 6644 8916 6696 8968
rect 7380 8916 7432 8968
rect 7564 8916 7616 8968
rect 8024 8984 8076 9036
rect 8300 9027 8352 9036
rect 8300 8993 8309 9027
rect 8309 8993 8343 9027
rect 8343 8993 8352 9027
rect 8300 8984 8352 8993
rect 8392 8984 8444 9036
rect 13176 9120 13228 9172
rect 13360 9163 13412 9172
rect 13360 9129 13369 9163
rect 13369 9129 13403 9163
rect 13403 9129 13412 9163
rect 13360 9120 13412 9129
rect 13912 9120 13964 9172
rect 14096 9163 14148 9172
rect 14096 9129 14105 9163
rect 14105 9129 14139 9163
rect 14139 9129 14148 9163
rect 14096 9120 14148 9129
rect 14648 9120 14700 9172
rect 16120 9163 16172 9172
rect 16120 9129 16129 9163
rect 16129 9129 16163 9163
rect 16163 9129 16172 9163
rect 16120 9120 16172 9129
rect 11244 9052 11296 9104
rect 11796 9052 11848 9104
rect 13268 9052 13320 9104
rect 13544 9052 13596 9104
rect 9772 8984 9824 9036
rect 10416 8984 10468 9036
rect 10692 8984 10744 9036
rect 14188 9027 14240 9036
rect 14188 8993 14197 9027
rect 14197 8993 14231 9027
rect 14231 8993 14240 9027
rect 14188 8984 14240 8993
rect 15752 8984 15804 9036
rect 8484 8959 8536 8968
rect 5908 8780 5960 8832
rect 6736 8891 6788 8900
rect 6736 8857 6745 8891
rect 6745 8857 6779 8891
rect 6779 8857 6788 8891
rect 6736 8848 6788 8857
rect 7288 8848 7340 8900
rect 7656 8891 7708 8900
rect 7656 8857 7665 8891
rect 7665 8857 7699 8891
rect 7699 8857 7708 8891
rect 7656 8848 7708 8857
rect 6184 8780 6236 8832
rect 8484 8925 8493 8959
rect 8493 8925 8527 8959
rect 8527 8925 8536 8959
rect 8484 8916 8536 8925
rect 8576 8916 8628 8968
rect 11520 8916 11572 8968
rect 12532 8916 12584 8968
rect 8852 8848 8904 8900
rect 9588 8848 9640 8900
rect 12992 8848 13044 8900
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 13636 8916 13688 8968
rect 14556 8916 14608 8968
rect 14924 8916 14976 8968
rect 16488 8984 16540 9036
rect 14188 8848 14240 8900
rect 15292 8848 15344 8900
rect 8300 8780 8352 8832
rect 8576 8780 8628 8832
rect 9772 8780 9824 8832
rect 10048 8780 10100 8832
rect 10968 8780 11020 8832
rect 11796 8780 11848 8832
rect 11888 8780 11940 8832
rect 14372 8780 14424 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 2412 8619 2464 8628
rect 2412 8585 2421 8619
rect 2421 8585 2455 8619
rect 2455 8585 2464 8619
rect 2412 8576 2464 8585
rect 2872 8576 2924 8628
rect 2964 8576 3016 8628
rect 6736 8576 6788 8628
rect 7840 8576 7892 8628
rect 8300 8576 8352 8628
rect 9036 8576 9088 8628
rect 9864 8576 9916 8628
rect 10692 8619 10744 8628
rect 10692 8585 10701 8619
rect 10701 8585 10735 8619
rect 10735 8585 10744 8619
rect 10692 8576 10744 8585
rect 11888 8619 11940 8628
rect 11888 8585 11897 8619
rect 11897 8585 11931 8619
rect 11931 8585 11940 8619
rect 11888 8576 11940 8585
rect 12992 8619 13044 8628
rect 12992 8585 13001 8619
rect 13001 8585 13035 8619
rect 13035 8585 13044 8619
rect 12992 8576 13044 8585
rect 13452 8619 13504 8628
rect 13452 8585 13461 8619
rect 13461 8585 13495 8619
rect 13495 8585 13504 8619
rect 13452 8576 13504 8585
rect 2228 8551 2280 8560
rect 2228 8517 2237 8551
rect 2237 8517 2271 8551
rect 2271 8517 2280 8551
rect 2228 8508 2280 8517
rect 2688 8508 2740 8560
rect 3516 8508 3568 8560
rect 5540 8508 5592 8560
rect 6644 8508 6696 8560
rect 3056 8440 3108 8492
rect 4988 8483 5040 8492
rect 4988 8449 4997 8483
rect 4997 8449 5031 8483
rect 5031 8449 5040 8483
rect 4988 8440 5040 8449
rect 7380 8508 7432 8560
rect 9588 8508 9640 8560
rect 9772 8551 9824 8560
rect 9772 8517 9781 8551
rect 9781 8517 9815 8551
rect 9815 8517 9824 8551
rect 9772 8508 9824 8517
rect 2136 8304 2188 8356
rect 5264 8372 5316 8424
rect 4068 8304 4120 8356
rect 5356 8347 5408 8356
rect 5356 8313 5365 8347
rect 5365 8313 5399 8347
rect 5399 8313 5408 8347
rect 5356 8304 5408 8313
rect 7564 8440 7616 8492
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 7840 8483 7892 8492
rect 7840 8449 7849 8483
rect 7849 8449 7883 8483
rect 7883 8449 7892 8483
rect 7840 8440 7892 8449
rect 8024 8440 8076 8492
rect 8300 8483 8352 8492
rect 8300 8449 8309 8483
rect 8309 8449 8343 8483
rect 8343 8449 8352 8483
rect 8300 8440 8352 8449
rect 9404 8440 9456 8492
rect 10600 8508 10652 8560
rect 11060 8508 11112 8560
rect 5816 8372 5868 8424
rect 10232 8440 10284 8492
rect 10416 8440 10468 8492
rect 10692 8440 10744 8492
rect 11520 8483 11572 8492
rect 11520 8449 11529 8483
rect 11529 8449 11563 8483
rect 11563 8449 11572 8483
rect 11520 8440 11572 8449
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 12900 8440 12952 8492
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 15292 8576 15344 8628
rect 15476 8576 15528 8628
rect 16948 8619 17000 8628
rect 16948 8585 16957 8619
rect 16957 8585 16991 8619
rect 16991 8585 17000 8619
rect 16948 8576 17000 8585
rect 9956 8415 10008 8424
rect 9956 8381 9965 8415
rect 9965 8381 9999 8415
rect 9999 8381 10008 8415
rect 9956 8372 10008 8381
rect 10968 8372 11020 8424
rect 11704 8372 11756 8424
rect 12624 8372 12676 8424
rect 6184 8304 6236 8356
rect 6920 8304 6972 8356
rect 7564 8304 7616 8356
rect 7932 8304 7984 8356
rect 11152 8304 11204 8356
rect 12992 8372 13044 8424
rect 13268 8372 13320 8424
rect 13452 8372 13504 8424
rect 14556 8440 14608 8492
rect 15200 8483 15252 8492
rect 15200 8449 15209 8483
rect 15209 8449 15243 8483
rect 15243 8449 15252 8483
rect 15200 8440 15252 8449
rect 15292 8440 15344 8492
rect 15752 8508 15804 8560
rect 16856 8440 16908 8492
rect 17040 8372 17092 8424
rect 3792 8236 3844 8288
rect 4160 8236 4212 8288
rect 5080 8236 5132 8288
rect 5908 8236 5960 8288
rect 8576 8236 8628 8288
rect 9312 8236 9364 8288
rect 9772 8279 9824 8288
rect 9772 8245 9781 8279
rect 9781 8245 9815 8279
rect 9815 8245 9824 8279
rect 9772 8236 9824 8245
rect 10140 8236 10192 8288
rect 10600 8236 10652 8288
rect 11336 8236 11388 8288
rect 11888 8236 11940 8288
rect 12624 8279 12676 8288
rect 12624 8245 12633 8279
rect 12633 8245 12667 8279
rect 12667 8245 12676 8279
rect 12624 8236 12676 8245
rect 12992 8236 13044 8288
rect 14004 8347 14056 8356
rect 14004 8313 14013 8347
rect 14013 8313 14047 8347
rect 14047 8313 14056 8347
rect 14004 8304 14056 8313
rect 13820 8236 13872 8288
rect 15752 8279 15804 8288
rect 15752 8245 15761 8279
rect 15761 8245 15795 8279
rect 15795 8245 15804 8279
rect 15752 8236 15804 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 2780 8032 2832 8084
rect 3608 8075 3660 8084
rect 3608 8041 3617 8075
rect 3617 8041 3651 8075
rect 3651 8041 3660 8075
rect 3608 8032 3660 8041
rect 2688 7964 2740 8016
rect 3700 7964 3752 8016
rect 2964 7896 3016 7948
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2044 7828 2096 7837
rect 2780 7803 2832 7812
rect 2780 7769 2789 7803
rect 2789 7769 2823 7803
rect 2823 7769 2832 7803
rect 2780 7760 2832 7769
rect 3148 7828 3200 7880
rect 3884 7871 3936 7880
rect 3884 7837 3893 7871
rect 3893 7837 3927 7871
rect 3927 7837 3936 7871
rect 3884 7828 3936 7837
rect 4068 7896 4120 7948
rect 5356 7964 5408 8016
rect 5540 7964 5592 8016
rect 5816 7964 5868 8016
rect 6092 8032 6144 8084
rect 9772 8032 9824 8084
rect 6276 7964 6328 8016
rect 6644 7964 6696 8016
rect 4804 7828 4856 7880
rect 5632 7896 5684 7948
rect 5080 7871 5132 7880
rect 5080 7837 5089 7871
rect 5089 7837 5123 7871
rect 5123 7837 5132 7871
rect 5080 7828 5132 7837
rect 5356 7871 5408 7880
rect 5356 7837 5365 7871
rect 5365 7837 5399 7871
rect 5399 7837 5408 7871
rect 5356 7828 5408 7837
rect 2964 7760 3016 7812
rect 4436 7803 4488 7812
rect 4436 7769 4445 7803
rect 4445 7769 4479 7803
rect 4479 7769 4488 7803
rect 4436 7760 4488 7769
rect 2688 7735 2740 7744
rect 2688 7701 2697 7735
rect 2697 7701 2731 7735
rect 2731 7701 2740 7735
rect 2688 7692 2740 7701
rect 2872 7692 2924 7744
rect 3976 7692 4028 7744
rect 5632 7760 5684 7812
rect 5356 7692 5408 7744
rect 5908 7828 5960 7880
rect 6184 7828 6236 7880
rect 7472 7896 7524 7948
rect 8392 7964 8444 8016
rect 11336 8032 11388 8084
rect 11428 8075 11480 8084
rect 11428 8041 11437 8075
rect 11437 8041 11471 8075
rect 11471 8041 11480 8075
rect 11428 8032 11480 8041
rect 11520 8032 11572 8084
rect 13820 8032 13872 8084
rect 14648 8032 14700 8084
rect 15016 8075 15068 8084
rect 15016 8041 15025 8075
rect 15025 8041 15059 8075
rect 15059 8041 15068 8075
rect 15016 8032 15068 8041
rect 15200 8032 15252 8084
rect 17040 8075 17092 8084
rect 17040 8041 17049 8075
rect 17049 8041 17083 8075
rect 17083 8041 17092 8075
rect 17040 8032 17092 8041
rect 7380 7871 7432 7880
rect 7380 7837 7387 7871
rect 7387 7837 7432 7871
rect 7380 7828 7432 7837
rect 7564 7871 7616 7880
rect 7564 7837 7573 7871
rect 7573 7837 7607 7871
rect 7607 7837 7616 7871
rect 7564 7828 7616 7837
rect 9772 7896 9824 7948
rect 7932 7871 7984 7880
rect 7932 7837 7941 7871
rect 7941 7837 7975 7871
rect 7975 7837 7984 7871
rect 7932 7828 7984 7837
rect 8024 7828 8076 7880
rect 8208 7871 8260 7880
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 8484 7828 8536 7880
rect 10508 7964 10560 8016
rect 9956 7896 10008 7948
rect 11520 7896 11572 7948
rect 10324 7828 10376 7880
rect 11060 7871 11112 7880
rect 11060 7837 11069 7871
rect 11069 7837 11103 7871
rect 11103 7837 11112 7871
rect 11060 7828 11112 7837
rect 11336 7871 11388 7880
rect 11336 7837 11345 7871
rect 11345 7837 11379 7871
rect 11379 7837 11388 7871
rect 11336 7828 11388 7837
rect 12900 7896 12952 7948
rect 6552 7692 6604 7744
rect 8668 7760 8720 7812
rect 8024 7692 8076 7744
rect 9220 7735 9272 7744
rect 9220 7701 9229 7735
rect 9229 7701 9263 7735
rect 9263 7701 9272 7735
rect 9220 7692 9272 7701
rect 10048 7760 10100 7812
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 13268 7803 13320 7812
rect 13268 7769 13277 7803
rect 13277 7769 13311 7803
rect 13311 7769 13320 7803
rect 13268 7760 13320 7769
rect 10140 7692 10192 7744
rect 10600 7692 10652 7744
rect 12808 7692 12860 7744
rect 15016 7871 15068 7880
rect 15016 7837 15025 7871
rect 15025 7837 15059 7871
rect 15059 7837 15068 7871
rect 15016 7828 15068 7837
rect 15660 7871 15712 7880
rect 15660 7837 15669 7871
rect 15669 7837 15703 7871
rect 15703 7837 15712 7871
rect 15660 7828 15712 7837
rect 15752 7828 15804 7880
rect 15568 7760 15620 7812
rect 14740 7692 14792 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 2596 7488 2648 7540
rect 2872 7488 2924 7540
rect 3516 7488 3568 7540
rect 3884 7531 3936 7540
rect 3884 7497 3893 7531
rect 3893 7497 3927 7531
rect 3927 7497 3936 7531
rect 3884 7488 3936 7497
rect 3976 7531 4028 7540
rect 3976 7497 3985 7531
rect 3985 7497 4019 7531
rect 4019 7497 4028 7531
rect 3976 7488 4028 7497
rect 4804 7488 4856 7540
rect 4988 7488 5040 7540
rect 2780 7420 2832 7472
rect 3148 7420 3200 7472
rect 3332 7420 3384 7472
rect 3424 7463 3476 7472
rect 3424 7429 3433 7463
rect 3433 7429 3467 7463
rect 3467 7429 3476 7463
rect 3424 7420 3476 7429
rect 3608 7463 3660 7472
rect 3608 7429 3617 7463
rect 3617 7429 3651 7463
rect 3651 7429 3660 7463
rect 3608 7420 3660 7429
rect 4068 7463 4120 7472
rect 4068 7429 4077 7463
rect 4077 7429 4111 7463
rect 4111 7429 4120 7463
rect 4068 7420 4120 7429
rect 5448 7488 5500 7540
rect 9128 7488 9180 7540
rect 9312 7531 9364 7540
rect 9312 7497 9321 7531
rect 9321 7497 9355 7531
rect 9355 7497 9364 7531
rect 9312 7488 9364 7497
rect 10048 7531 10100 7540
rect 10048 7497 10057 7531
rect 10057 7497 10091 7531
rect 10091 7497 10100 7531
rect 10048 7488 10100 7497
rect 11336 7488 11388 7540
rect 2044 7352 2096 7404
rect 2596 7352 2648 7404
rect 2688 7395 2740 7404
rect 2688 7361 2697 7395
rect 2697 7361 2731 7395
rect 2731 7361 2740 7395
rect 2688 7352 2740 7361
rect 2964 7352 3016 7404
rect 4436 7395 4488 7404
rect 4436 7361 4445 7395
rect 4445 7361 4479 7395
rect 4479 7361 4488 7395
rect 4436 7352 4488 7361
rect 4620 7395 4672 7404
rect 4620 7361 4629 7395
rect 4629 7361 4663 7395
rect 4663 7361 4672 7395
rect 4620 7352 4672 7361
rect 4068 7284 4120 7336
rect 3792 7216 3844 7268
rect 5080 7395 5132 7404
rect 5080 7361 5089 7395
rect 5089 7361 5123 7395
rect 5123 7361 5132 7395
rect 5080 7352 5132 7361
rect 6092 7420 6144 7472
rect 9772 7420 9824 7472
rect 10232 7420 10284 7472
rect 11244 7420 11296 7472
rect 15568 7488 15620 7540
rect 15936 7531 15988 7540
rect 15936 7497 15945 7531
rect 15945 7497 15979 7531
rect 15979 7497 15988 7531
rect 15936 7488 15988 7497
rect 16304 7531 16356 7540
rect 16304 7497 16313 7531
rect 16313 7497 16347 7531
rect 16347 7497 16356 7531
rect 16304 7488 16356 7497
rect 16948 7531 17000 7540
rect 16948 7497 16957 7531
rect 16957 7497 16991 7531
rect 16991 7497 17000 7531
rect 16948 7488 17000 7497
rect 5448 7395 5500 7404
rect 5448 7361 5457 7395
rect 5457 7361 5491 7395
rect 5491 7361 5500 7395
rect 5448 7352 5500 7361
rect 5632 7352 5684 7404
rect 8392 7352 8444 7404
rect 8852 7395 8904 7404
rect 8852 7361 8861 7395
rect 8861 7361 8895 7395
rect 8895 7361 8904 7395
rect 8852 7352 8904 7361
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 9312 7352 9364 7404
rect 9864 7395 9916 7404
rect 9864 7361 9873 7395
rect 9873 7361 9907 7395
rect 9907 7361 9916 7395
rect 9864 7352 9916 7361
rect 10140 7395 10192 7404
rect 10140 7361 10149 7395
rect 10149 7361 10183 7395
rect 10183 7361 10192 7395
rect 10140 7352 10192 7361
rect 11796 7395 11848 7404
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 11796 7352 11848 7361
rect 12072 7395 12124 7404
rect 12072 7361 12081 7395
rect 12081 7361 12115 7395
rect 12115 7361 12124 7395
rect 12072 7352 12124 7361
rect 5540 7284 5592 7336
rect 7472 7284 7524 7336
rect 8944 7327 8996 7336
rect 8944 7293 8953 7327
rect 8953 7293 8987 7327
rect 8987 7293 8996 7327
rect 8944 7284 8996 7293
rect 11428 7284 11480 7336
rect 12808 7463 12860 7472
rect 12808 7429 12817 7463
rect 12817 7429 12851 7463
rect 12851 7429 12860 7463
rect 12808 7420 12860 7429
rect 12348 7395 12400 7404
rect 12348 7361 12357 7395
rect 12357 7361 12391 7395
rect 12391 7361 12400 7395
rect 12348 7352 12400 7361
rect 16120 7395 16172 7404
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 16488 7395 16540 7404
rect 16488 7361 16497 7395
rect 16497 7361 16531 7395
rect 16531 7361 16540 7395
rect 16488 7352 16540 7361
rect 17040 7352 17092 7404
rect 9404 7216 9456 7268
rect 5356 7148 5408 7200
rect 8668 7148 8720 7200
rect 9312 7148 9364 7200
rect 14372 7284 14424 7336
rect 12532 7216 12584 7268
rect 13084 7216 13136 7268
rect 11060 7148 11112 7200
rect 11612 7191 11664 7200
rect 11612 7157 11621 7191
rect 11621 7157 11655 7191
rect 11655 7157 11664 7191
rect 11612 7148 11664 7157
rect 11888 7148 11940 7200
rect 12992 7191 13044 7200
rect 12992 7157 13001 7191
rect 13001 7157 13035 7191
rect 13035 7157 13044 7191
rect 12992 7148 13044 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 3332 6944 3384 6996
rect 6092 6944 6144 6996
rect 7564 6944 7616 6996
rect 7104 6876 7156 6928
rect 8760 6944 8812 6996
rect 9588 6944 9640 6996
rect 9956 6944 10008 6996
rect 11152 6987 11204 6996
rect 11152 6953 11161 6987
rect 11161 6953 11195 6987
rect 11195 6953 11204 6987
rect 11152 6944 11204 6953
rect 12072 6944 12124 6996
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 4068 6740 4120 6792
rect 4804 6783 4856 6792
rect 4804 6749 4813 6783
rect 4813 6749 4847 6783
rect 4847 6749 4856 6783
rect 4804 6740 4856 6749
rect 4988 6783 5040 6792
rect 4988 6749 4997 6783
rect 4997 6749 5031 6783
rect 5031 6749 5040 6783
rect 4988 6740 5040 6749
rect 5356 6740 5408 6792
rect 1676 6715 1728 6724
rect 1676 6681 1710 6715
rect 1710 6681 1728 6715
rect 1676 6672 1728 6681
rect 4712 6672 4764 6724
rect 5908 6783 5960 6792
rect 5908 6749 5917 6783
rect 5917 6749 5951 6783
rect 5951 6749 5960 6783
rect 5908 6740 5960 6749
rect 6368 6808 6420 6860
rect 7196 6808 7248 6860
rect 7288 6740 7340 6792
rect 6276 6672 6328 6724
rect 7196 6715 7248 6724
rect 7196 6681 7205 6715
rect 7205 6681 7239 6715
rect 7239 6681 7248 6715
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 8392 6876 8444 6928
rect 9404 6919 9456 6928
rect 9404 6885 9413 6919
rect 9413 6885 9447 6919
rect 9447 6885 9456 6919
rect 9404 6876 9456 6885
rect 7840 6740 7892 6792
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 7196 6672 7248 6681
rect 5632 6604 5684 6656
rect 7932 6672 7984 6724
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 8852 6740 8904 6792
rect 10140 6808 10192 6860
rect 10968 6808 11020 6860
rect 11244 6851 11296 6860
rect 11244 6817 11253 6851
rect 11253 6817 11287 6851
rect 11287 6817 11296 6851
rect 11244 6808 11296 6817
rect 12256 6808 12308 6860
rect 12900 6808 12952 6860
rect 13176 6851 13228 6860
rect 13176 6817 13185 6851
rect 13185 6817 13219 6851
rect 13219 6817 13228 6851
rect 13176 6808 13228 6817
rect 14096 6944 14148 6996
rect 15016 6944 15068 6996
rect 13912 6808 13964 6860
rect 11336 6740 11388 6792
rect 11428 6783 11480 6792
rect 11428 6749 11437 6783
rect 11437 6749 11471 6783
rect 11471 6749 11480 6783
rect 11428 6740 11480 6749
rect 8944 6715 8996 6724
rect 8944 6681 8953 6715
rect 8953 6681 8987 6715
rect 8987 6681 8996 6715
rect 8944 6672 8996 6681
rect 9588 6672 9640 6724
rect 9772 6672 9824 6724
rect 11152 6715 11204 6724
rect 11152 6681 11161 6715
rect 11161 6681 11195 6715
rect 11195 6681 11204 6715
rect 11152 6672 11204 6681
rect 12532 6672 12584 6724
rect 12624 6672 12676 6724
rect 9864 6604 9916 6656
rect 12164 6604 12216 6656
rect 13636 6672 13688 6724
rect 14372 6715 14424 6724
rect 14372 6681 14381 6715
rect 14381 6681 14415 6715
rect 14415 6681 14424 6715
rect 14372 6672 14424 6681
rect 13360 6647 13412 6656
rect 13360 6613 13369 6647
rect 13369 6613 13403 6647
rect 13403 6613 13412 6647
rect 13360 6604 13412 6613
rect 13820 6604 13872 6656
rect 14188 6604 14240 6656
rect 15660 6783 15712 6792
rect 15660 6749 15669 6783
rect 15669 6749 15703 6783
rect 15703 6749 15712 6783
rect 15660 6740 15712 6749
rect 15752 6672 15804 6724
rect 16488 6604 16540 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 1676 6400 1728 6452
rect 3792 6400 3844 6452
rect 6276 6400 6328 6452
rect 7748 6400 7800 6452
rect 8852 6400 8904 6452
rect 8944 6400 8996 6452
rect 9312 6400 9364 6452
rect 9588 6400 9640 6452
rect 11336 6400 11388 6452
rect 12624 6400 12676 6452
rect 12716 6400 12768 6452
rect 13636 6400 13688 6452
rect 13728 6443 13780 6452
rect 13728 6409 13737 6443
rect 13737 6409 13771 6443
rect 13771 6409 13780 6443
rect 13728 6400 13780 6409
rect 848 6264 900 6316
rect 1860 6307 1912 6316
rect 1860 6273 1869 6307
rect 1869 6273 1903 6307
rect 1903 6273 1912 6307
rect 1860 6264 1912 6273
rect 3700 6332 3752 6384
rect 3424 6264 3476 6316
rect 2872 6196 2924 6248
rect 3884 6264 3936 6316
rect 4804 6332 4856 6384
rect 7196 6332 7248 6384
rect 7564 6375 7616 6384
rect 7564 6341 7573 6375
rect 7573 6341 7607 6375
rect 7607 6341 7616 6375
rect 7564 6332 7616 6341
rect 7840 6332 7892 6384
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 4712 6264 4764 6316
rect 3608 6239 3660 6248
rect 3608 6205 3617 6239
rect 3617 6205 3651 6239
rect 3651 6205 3660 6239
rect 3608 6196 3660 6205
rect 3976 6196 4028 6248
rect 4804 6239 4856 6248
rect 4804 6205 4813 6239
rect 4813 6205 4847 6239
rect 4847 6205 4856 6239
rect 4804 6196 4856 6205
rect 5264 6307 5316 6316
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 5448 6307 5500 6316
rect 5448 6273 5462 6307
rect 5462 6273 5496 6307
rect 5496 6273 5500 6307
rect 5448 6264 5500 6273
rect 7104 6264 7156 6316
rect 6000 6196 6052 6248
rect 7288 6196 7340 6248
rect 7748 6307 7800 6316
rect 7748 6273 7757 6307
rect 7757 6273 7791 6307
rect 7791 6273 7800 6307
rect 7748 6264 7800 6273
rect 8760 6332 8812 6384
rect 12072 6332 12124 6384
rect 12992 6332 13044 6384
rect 15476 6400 15528 6452
rect 15752 6443 15804 6452
rect 15752 6409 15761 6443
rect 15761 6409 15795 6443
rect 15795 6409 15804 6443
rect 15752 6400 15804 6409
rect 3792 6128 3844 6180
rect 7196 6128 7248 6180
rect 7840 6196 7892 6248
rect 7564 6128 7616 6180
rect 8300 6307 8352 6316
rect 8300 6273 8309 6307
rect 8309 6273 8343 6307
rect 8343 6273 8352 6307
rect 8300 6264 8352 6273
rect 8484 6264 8536 6316
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 9864 6264 9916 6316
rect 10048 6264 10100 6316
rect 13360 6307 13412 6316
rect 13360 6273 13369 6307
rect 13369 6273 13403 6307
rect 13403 6273 13412 6307
rect 13360 6264 13412 6273
rect 13636 6307 13688 6316
rect 13636 6273 13645 6307
rect 13645 6273 13679 6307
rect 13679 6273 13688 6307
rect 13636 6264 13688 6273
rect 8852 6196 8904 6248
rect 10048 6128 10100 6180
rect 11428 6128 11480 6180
rect 12900 6128 12952 6180
rect 13728 6128 13780 6180
rect 15292 6264 15344 6316
rect 16488 6307 16540 6316
rect 16488 6273 16497 6307
rect 16497 6273 16531 6307
rect 16531 6273 16540 6307
rect 16488 6264 16540 6273
rect 16764 6307 16816 6316
rect 16764 6273 16773 6307
rect 16773 6273 16807 6307
rect 16807 6273 16816 6307
rect 16764 6264 16816 6273
rect 16948 6171 17000 6180
rect 16948 6137 16957 6171
rect 16957 6137 16991 6171
rect 16991 6137 17000 6171
rect 16948 6128 17000 6137
rect 1676 6103 1728 6112
rect 1676 6069 1685 6103
rect 1685 6069 1719 6103
rect 1719 6069 1728 6103
rect 1676 6060 1728 6069
rect 6368 6060 6420 6112
rect 7288 6060 7340 6112
rect 7472 6060 7524 6112
rect 8392 6060 8444 6112
rect 8668 6060 8720 6112
rect 11612 6060 11664 6112
rect 13636 6103 13688 6112
rect 13636 6069 13645 6103
rect 13645 6069 13679 6103
rect 13679 6069 13688 6103
rect 13636 6060 13688 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 2780 5899 2832 5908
rect 2780 5865 2789 5899
rect 2789 5865 2823 5899
rect 2823 5865 2832 5899
rect 2780 5856 2832 5865
rect 4712 5856 4764 5908
rect 3608 5788 3660 5840
rect 7380 5856 7432 5908
rect 8300 5856 8352 5908
rect 8484 5899 8536 5908
rect 8484 5865 8493 5899
rect 8493 5865 8527 5899
rect 8527 5865 8536 5899
rect 8484 5856 8536 5865
rect 9036 5856 9088 5908
rect 9588 5856 9640 5908
rect 10600 5899 10652 5908
rect 10600 5865 10609 5899
rect 10609 5865 10643 5899
rect 10643 5865 10652 5899
rect 10600 5856 10652 5865
rect 11612 5899 11664 5908
rect 11612 5865 11621 5899
rect 11621 5865 11655 5899
rect 11655 5865 11664 5899
rect 11612 5856 11664 5865
rect 12348 5856 12400 5908
rect 13728 5856 13780 5908
rect 14464 5856 14516 5908
rect 16856 5856 16908 5908
rect 3792 5720 3844 5772
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 1676 5695 1728 5704
rect 1676 5661 1710 5695
rect 1710 5661 1728 5695
rect 1676 5652 1728 5661
rect 3424 5652 3476 5704
rect 3976 5652 4028 5704
rect 5724 5788 5776 5840
rect 6644 5788 6696 5840
rect 5632 5652 5684 5704
rect 6460 5720 6512 5772
rect 6276 5695 6328 5704
rect 6276 5661 6278 5695
rect 6278 5661 6312 5695
rect 6312 5661 6328 5695
rect 6276 5652 6328 5661
rect 6368 5695 6420 5704
rect 6368 5661 6377 5695
rect 6377 5661 6411 5695
rect 6411 5661 6420 5695
rect 6368 5652 6420 5661
rect 6552 5695 6604 5704
rect 6552 5661 6561 5695
rect 6561 5661 6595 5695
rect 6595 5661 6604 5695
rect 6552 5652 6604 5661
rect 7564 5788 7616 5840
rect 7840 5788 7892 5840
rect 7380 5720 7432 5772
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 9404 5788 9456 5840
rect 15292 5788 15344 5840
rect 8208 5652 8260 5704
rect 8392 5652 8444 5704
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 3332 5584 3384 5636
rect 3884 5584 3936 5636
rect 5724 5627 5776 5636
rect 5724 5593 5733 5627
rect 5733 5593 5767 5627
rect 5767 5593 5776 5627
rect 5724 5584 5776 5593
rect 3700 5516 3752 5568
rect 4068 5516 4120 5568
rect 4620 5516 4672 5568
rect 6092 5516 6144 5568
rect 6736 5584 6788 5636
rect 7104 5627 7156 5636
rect 7104 5593 7113 5627
rect 7113 5593 7147 5627
rect 7147 5593 7156 5627
rect 7104 5584 7156 5593
rect 10416 5652 10468 5704
rect 10232 5627 10284 5636
rect 10232 5593 10241 5627
rect 10241 5593 10275 5627
rect 10275 5593 10284 5627
rect 10232 5584 10284 5593
rect 10508 5627 10560 5636
rect 10508 5593 10517 5627
rect 10517 5593 10551 5627
rect 10551 5593 10560 5627
rect 10508 5584 10560 5593
rect 10876 5652 10928 5704
rect 12348 5720 12400 5772
rect 14188 5763 14240 5772
rect 14188 5729 14197 5763
rect 14197 5729 14231 5763
rect 14231 5729 14240 5763
rect 14188 5720 14240 5729
rect 11060 5584 11112 5636
rect 11520 5652 11572 5704
rect 13544 5695 13596 5704
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 13636 5652 13688 5704
rect 15476 5720 15528 5772
rect 9036 5516 9088 5568
rect 10600 5516 10652 5568
rect 12624 5584 12676 5636
rect 13360 5584 13412 5636
rect 14096 5627 14148 5636
rect 14096 5593 14105 5627
rect 14105 5593 14139 5627
rect 14139 5593 14148 5627
rect 14096 5584 14148 5593
rect 15660 5695 15712 5704
rect 15660 5661 15669 5695
rect 15669 5661 15703 5695
rect 15703 5661 15712 5695
rect 15660 5652 15712 5661
rect 15292 5627 15344 5636
rect 15292 5593 15301 5627
rect 15301 5593 15335 5627
rect 15335 5593 15344 5627
rect 15292 5584 15344 5593
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 3056 5312 3108 5364
rect 1492 5176 1544 5228
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 3792 5244 3844 5296
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 3424 5108 3476 5160
rect 3700 5219 3752 5228
rect 3700 5185 3709 5219
rect 3709 5185 3743 5219
rect 3743 5185 3752 5219
rect 3700 5176 3752 5185
rect 3976 5219 4028 5228
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 4252 5176 4304 5228
rect 4804 5219 4856 5228
rect 4804 5185 4813 5219
rect 4813 5185 4847 5219
rect 4847 5185 4856 5219
rect 4804 5176 4856 5185
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 5172 5176 5224 5228
rect 5356 5176 5408 5228
rect 5632 5219 5684 5228
rect 5632 5185 5646 5219
rect 5646 5185 5680 5219
rect 5680 5185 5684 5219
rect 5632 5176 5684 5185
rect 5816 5176 5868 5228
rect 6000 5108 6052 5160
rect 3700 5040 3752 5092
rect 3884 5040 3936 5092
rect 4068 5040 4120 5092
rect 6368 5219 6420 5228
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 6552 5219 6604 5228
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 6552 5176 6604 5185
rect 7380 5287 7432 5296
rect 7380 5253 7389 5287
rect 7389 5253 7423 5287
rect 7423 5253 7432 5287
rect 7380 5244 7432 5253
rect 7932 5244 7984 5296
rect 6460 5108 6512 5160
rect 7104 5176 7156 5228
rect 7564 5219 7616 5228
rect 7564 5185 7573 5219
rect 7573 5185 7607 5219
rect 7607 5185 7616 5219
rect 7564 5176 7616 5185
rect 7656 5176 7708 5228
rect 7840 5219 7892 5228
rect 7840 5185 7849 5219
rect 7849 5185 7883 5219
rect 7883 5185 7892 5219
rect 7840 5176 7892 5185
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 8208 5219 8260 5228
rect 8208 5185 8217 5219
rect 8217 5185 8251 5219
rect 8251 5185 8260 5219
rect 8208 5176 8260 5185
rect 8484 5219 8536 5228
rect 8484 5185 8493 5219
rect 8493 5185 8527 5219
rect 8527 5185 8536 5219
rect 8484 5176 8536 5185
rect 8668 5355 8720 5364
rect 8668 5321 8677 5355
rect 8677 5321 8711 5355
rect 8711 5321 8720 5355
rect 8668 5312 8720 5321
rect 10508 5312 10560 5364
rect 11980 5312 12032 5364
rect 9036 5219 9088 5228
rect 9036 5185 9045 5219
rect 9045 5185 9079 5219
rect 9079 5185 9088 5219
rect 9036 5176 9088 5185
rect 9128 5176 9180 5228
rect 6092 4972 6144 5024
rect 8024 4972 8076 5024
rect 10324 5244 10376 5296
rect 12348 5312 12400 5364
rect 15292 5312 15344 5364
rect 16948 5355 17000 5364
rect 16948 5321 16957 5355
rect 16957 5321 16991 5355
rect 16991 5321 17000 5355
rect 16948 5312 17000 5321
rect 9680 5176 9732 5228
rect 9772 5219 9824 5228
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5176 9824 5185
rect 10140 5176 10192 5228
rect 12256 5287 12308 5296
rect 12256 5253 12265 5287
rect 12265 5253 12299 5287
rect 12299 5253 12308 5287
rect 12256 5244 12308 5253
rect 11796 5176 11848 5228
rect 12440 5219 12492 5228
rect 12440 5185 12449 5219
rect 12449 5185 12483 5219
rect 12483 5185 12492 5219
rect 12440 5176 12492 5185
rect 12716 5219 12768 5228
rect 12716 5185 12725 5219
rect 12725 5185 12759 5219
rect 12759 5185 12768 5219
rect 12716 5176 12768 5185
rect 15292 5176 15344 5228
rect 15752 5176 15804 5228
rect 13268 5108 13320 5160
rect 16856 5108 16908 5160
rect 15476 5040 15528 5092
rect 9680 5015 9732 5024
rect 9680 4981 9689 5015
rect 9689 4981 9723 5015
rect 9723 4981 9732 5015
rect 9680 4972 9732 4981
rect 10048 5015 10100 5024
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 13728 4972 13780 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 3240 4768 3292 4820
rect 3792 4768 3844 4820
rect 3976 4811 4028 4820
rect 3976 4777 3985 4811
rect 3985 4777 4019 4811
rect 4019 4777 4028 4811
rect 3976 4768 4028 4777
rect 4068 4768 4120 4820
rect 4896 4768 4948 4820
rect 5356 4768 5408 4820
rect 6552 4768 6604 4820
rect 5908 4700 5960 4752
rect 6736 4700 6788 4752
rect 7104 4700 7156 4752
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 3056 4564 3108 4616
rect 1676 4539 1728 4548
rect 1676 4505 1710 4539
rect 1710 4505 1728 4539
rect 1676 4496 1728 4505
rect 3700 4496 3752 4548
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4068 4564 4120 4573
rect 6460 4632 6512 4684
rect 6828 4632 6880 4684
rect 9772 4768 9824 4820
rect 9496 4700 9548 4752
rect 10692 4700 10744 4752
rect 8024 4632 8076 4684
rect 8576 4632 8628 4684
rect 16580 4768 16632 4820
rect 16764 4768 16816 4820
rect 7840 4607 7892 4616
rect 7840 4573 7849 4607
rect 7849 4573 7883 4607
rect 7883 4573 7892 4607
rect 7840 4564 7892 4573
rect 7656 4496 7708 4548
rect 8116 4564 8168 4616
rect 9956 4564 10008 4616
rect 10876 4564 10928 4616
rect 13452 4564 13504 4616
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 14004 4564 14056 4616
rect 15476 4632 15528 4684
rect 15384 4607 15436 4616
rect 15384 4573 15393 4607
rect 15393 4573 15427 4607
rect 15427 4573 15436 4607
rect 15384 4564 15436 4573
rect 15660 4607 15712 4616
rect 15660 4573 15669 4607
rect 15669 4573 15703 4607
rect 15703 4573 15712 4607
rect 15660 4564 15712 4573
rect 5632 4428 5684 4480
rect 6368 4428 6420 4480
rect 9680 4428 9732 4480
rect 10140 4428 10192 4480
rect 11152 4428 11204 4480
rect 13544 4428 13596 4480
rect 15200 4428 15252 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 1492 4224 1544 4276
rect 1676 4267 1728 4276
rect 1676 4233 1685 4267
rect 1685 4233 1719 4267
rect 1719 4233 1728 4267
rect 1676 4224 1728 4233
rect 6092 4224 6144 4276
rect 7656 4267 7708 4276
rect 7656 4233 7665 4267
rect 7665 4233 7699 4267
rect 7699 4233 7708 4267
rect 7656 4224 7708 4233
rect 9680 4224 9732 4276
rect 10968 4224 11020 4276
rect 7472 4156 7524 4208
rect 8208 4156 8260 4208
rect 10140 4199 10192 4208
rect 10140 4165 10149 4199
rect 10149 4165 10183 4199
rect 10183 4165 10192 4199
rect 10140 4156 10192 4165
rect 10876 4199 10928 4208
rect 10876 4165 10885 4199
rect 10885 4165 10919 4199
rect 10919 4165 10928 4199
rect 10876 4156 10928 4165
rect 1308 4088 1360 4140
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 6368 4131 6420 4140
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 6736 4088 6788 4140
rect 9128 4088 9180 4140
rect 9404 4131 9456 4140
rect 9404 4097 9413 4131
rect 9413 4097 9447 4131
rect 9447 4097 9456 4131
rect 9404 4088 9456 4097
rect 9496 4088 9548 4140
rect 10324 4088 10376 4140
rect 7196 4020 7248 4072
rect 7472 4063 7524 4072
rect 7472 4029 7481 4063
rect 7481 4029 7515 4063
rect 7515 4029 7524 4063
rect 7472 4020 7524 4029
rect 7840 4020 7892 4072
rect 10600 4088 10652 4140
rect 10692 4063 10744 4072
rect 10692 4029 10701 4063
rect 10701 4029 10735 4063
rect 10735 4029 10744 4063
rect 10692 4020 10744 4029
rect 10784 4020 10836 4072
rect 12072 4199 12124 4208
rect 12072 4165 12081 4199
rect 12081 4165 12115 4199
rect 12115 4165 12124 4199
rect 12072 4156 12124 4165
rect 13636 4156 13688 4208
rect 14096 4199 14148 4208
rect 14096 4165 14105 4199
rect 14105 4165 14139 4199
rect 14139 4165 14148 4199
rect 14096 4156 14148 4165
rect 13544 4131 13596 4140
rect 13544 4097 13553 4131
rect 13553 4097 13587 4131
rect 13587 4097 13596 4131
rect 13544 4088 13596 4097
rect 13820 4131 13872 4140
rect 13820 4097 13829 4131
rect 13829 4097 13863 4131
rect 13863 4097 13872 4131
rect 13820 4088 13872 4097
rect 14004 4131 14056 4140
rect 14004 4097 14013 4131
rect 14013 4097 14047 4131
rect 14047 4097 14056 4131
rect 14004 4088 14056 4097
rect 13360 4020 13412 4072
rect 15200 4224 15252 4276
rect 15384 4224 15436 4276
rect 14740 4131 14792 4140
rect 14740 4097 14749 4131
rect 14749 4097 14783 4131
rect 14783 4097 14792 4131
rect 14740 4088 14792 4097
rect 15752 4131 15804 4140
rect 15752 4097 15761 4131
rect 15761 4097 15795 4131
rect 15795 4097 15804 4131
rect 15752 4088 15804 4097
rect 16764 4088 16816 4140
rect 15292 4020 15344 4072
rect 7840 3927 7892 3936
rect 7840 3893 7849 3927
rect 7849 3893 7883 3927
rect 7883 3893 7892 3927
rect 7840 3884 7892 3893
rect 8944 3884 8996 3936
rect 9496 3884 9548 3936
rect 9864 3884 9916 3936
rect 9956 3927 10008 3936
rect 9956 3893 9965 3927
rect 9965 3893 9999 3927
rect 9999 3893 10008 3927
rect 9956 3884 10008 3893
rect 10324 3884 10376 3936
rect 14004 3884 14056 3936
rect 14556 3927 14608 3936
rect 14556 3893 14565 3927
rect 14565 3893 14599 3927
rect 14599 3893 14608 3927
rect 14556 3884 14608 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 6828 3680 6880 3732
rect 7472 3680 7524 3732
rect 7840 3680 7892 3732
rect 8116 3612 8168 3664
rect 8208 3612 8260 3664
rect 7472 3476 7524 3528
rect 8024 3476 8076 3528
rect 9128 3723 9180 3732
rect 9128 3689 9137 3723
rect 9137 3689 9171 3723
rect 9171 3689 9180 3723
rect 9128 3680 9180 3689
rect 10968 3723 11020 3732
rect 10968 3689 10977 3723
rect 10977 3689 11011 3723
rect 11011 3689 11020 3723
rect 10968 3680 11020 3689
rect 12348 3723 12400 3732
rect 12348 3689 12357 3723
rect 12357 3689 12391 3723
rect 12391 3689 12400 3723
rect 12348 3680 12400 3689
rect 12532 3723 12584 3732
rect 12532 3689 12541 3723
rect 12541 3689 12575 3723
rect 12575 3689 12584 3723
rect 12532 3680 12584 3689
rect 15752 3680 15804 3732
rect 16488 3680 16540 3732
rect 9956 3612 10008 3664
rect 12256 3587 12308 3596
rect 12256 3553 12265 3587
rect 12265 3553 12299 3587
rect 12299 3553 12308 3587
rect 12256 3544 12308 3553
rect 7196 3408 7248 3460
rect 8116 3408 8168 3460
rect 9404 3476 9456 3528
rect 9956 3408 10008 3460
rect 11152 3476 11204 3528
rect 12072 3519 12124 3528
rect 12072 3485 12081 3519
rect 12081 3485 12115 3519
rect 12115 3485 12124 3519
rect 12072 3476 12124 3485
rect 7288 3383 7340 3392
rect 7288 3349 7297 3383
rect 7297 3349 7331 3383
rect 7331 3349 7340 3383
rect 7288 3340 7340 3349
rect 7564 3340 7616 3392
rect 9312 3340 9364 3392
rect 9496 3340 9548 3392
rect 14648 3519 14700 3528
rect 14648 3485 14657 3519
rect 14657 3485 14691 3519
rect 14691 3485 14700 3519
rect 14648 3476 14700 3485
rect 15660 3476 15712 3528
rect 15936 3476 15988 3528
rect 14556 3408 14608 3460
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 7840 3136 7892 3188
rect 9956 3136 10008 3188
rect 11152 3136 11204 3188
rect 1400 3068 1452 3120
rect 6460 3000 6512 3052
rect 7840 3000 7892 3052
rect 8208 3043 8260 3052
rect 8208 3009 8217 3043
rect 8217 3009 8251 3043
rect 8251 3009 8260 3043
rect 8208 3000 8260 3009
rect 9220 3068 9272 3120
rect 9128 3000 9180 3052
rect 10232 3043 10284 3052
rect 10232 3009 10266 3043
rect 10266 3009 10284 3043
rect 10232 3000 10284 3009
rect 14280 3043 14332 3052
rect 14648 3068 14700 3120
rect 14280 3009 14298 3043
rect 14298 3009 14332 3043
rect 14280 3000 14332 3009
rect 8024 2975 8076 2984
rect 8024 2941 8033 2975
rect 8033 2941 8067 2975
rect 8067 2941 8076 2975
rect 8024 2932 8076 2941
rect 14648 2932 14700 2984
rect 6644 2796 6696 2848
rect 13912 2796 13964 2848
rect 14556 2796 14608 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 6460 2592 6512 2644
rect 9128 2635 9180 2644
rect 9128 2601 9137 2635
rect 9137 2601 9171 2635
rect 9171 2601 9180 2635
rect 9128 2592 9180 2601
rect 10232 2592 10284 2644
rect 14280 2592 14332 2644
rect 14648 2456 14700 2508
rect 5816 2388 5868 2440
rect 9036 2388 9088 2440
rect 10324 2388 10376 2440
rect 13912 2431 13964 2440
rect 13912 2397 13921 2431
rect 13921 2397 13955 2431
rect 13955 2397 13964 2431
rect 13912 2388 13964 2397
rect 14096 2388 14148 2440
rect 14556 2431 14608 2440
rect 14556 2397 14565 2431
rect 14565 2397 14599 2431
rect 14599 2397 14608 2431
rect 14556 2388 14608 2397
rect 16028 2388 16080 2440
rect 13544 2252 13596 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 12898 19858 12954 20658
rect 13542 19858 13598 20658
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 12912 17882 12940 19858
rect 13556 17882 13584 19858
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 13544 17876 13596 17882
rect 13544 17818 13596 17824
rect 13268 17604 13320 17610
rect 13268 17546 13320 17552
rect 14740 17604 14792 17610
rect 14740 17546 14792 17552
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 8574 17096 8630 17105
rect 8574 17031 8630 17040
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 8312 15706 8340 16050
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3436 13938 3464 14350
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 3700 14000 3752 14006
rect 3700 13942 3752 13948
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3160 13326 3188 13874
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2596 12164 2648 12170
rect 2596 12106 2648 12112
rect 2608 11558 2636 12106
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2792 10169 2820 12174
rect 2884 12170 2912 12854
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 3252 12832 3280 13194
rect 3344 13172 3372 13874
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3424 13184 3476 13190
rect 3344 13144 3424 13172
rect 3424 13126 3476 13132
rect 3332 12844 3384 12850
rect 3252 12804 3332 12832
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 2884 10674 2912 12106
rect 3068 12102 3096 12786
rect 3252 12238 3280 12804
rect 3332 12786 3384 12792
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 3068 10674 3096 12038
rect 3252 11898 3280 12174
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3252 11665 3280 11834
rect 3332 11756 3384 11762
rect 3436 11744 3464 13126
rect 3528 11762 3556 13330
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 3620 12850 3648 13262
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3620 12238 3648 12786
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3620 11762 3648 12174
rect 3384 11716 3464 11744
rect 3332 11698 3384 11704
rect 3238 11656 3294 11665
rect 3238 11591 3294 11600
rect 3436 10674 3464 11716
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3528 10674 3556 11698
rect 3620 11354 3648 11698
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3712 10724 3740 13942
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 3792 13252 3844 13258
rect 3792 13194 3844 13200
rect 3804 12986 3832 13194
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3896 12434 3924 13874
rect 4172 13818 4200 13874
rect 4080 13790 4200 13818
rect 4080 13462 4108 13790
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 4344 13456 4396 13462
rect 4632 13410 4660 14214
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5460 13530 5488 13738
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 4344 13398 4396 13404
rect 4080 13326 4108 13398
rect 4356 13326 4384 13398
rect 4540 13382 4660 13410
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4172 12889 4200 13126
rect 4540 12986 4568 13382
rect 4724 13326 4752 13466
rect 5552 13462 5580 15370
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5172 13388 5224 13394
rect 5224 13348 5304 13376
rect 5172 13330 5224 13336
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4158 12880 4214 12889
rect 4158 12815 4214 12824
rect 4632 12782 4660 13262
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4724 12850 4752 13126
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4712 12844 4764 12850
rect 5172 12844 5224 12850
rect 4764 12804 4844 12832
rect 4712 12786 4764 12792
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3896 12406 4016 12434
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 3804 11801 3832 11834
rect 3896 11830 3924 12242
rect 3884 11824 3936 11830
rect 3790 11792 3846 11801
rect 3884 11766 3936 11772
rect 3790 11727 3846 11736
rect 3896 11218 3924 11766
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3884 10736 3936 10742
rect 3712 10696 3884 10724
rect 3884 10678 3936 10684
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 2778 10160 2834 10169
rect 2778 10095 2834 10104
rect 2228 10056 2280 10062
rect 2228 9998 2280 10004
rect 2136 9988 2188 9994
rect 2136 9930 2188 9936
rect 2148 9722 2176 9930
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 2148 8906 2176 9658
rect 2240 9654 2268 9998
rect 2320 9988 2372 9994
rect 2320 9930 2372 9936
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2240 8974 2268 9590
rect 2332 9586 2360 9930
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2700 9586 2728 9862
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2332 8922 2360 9522
rect 2700 9042 2728 9522
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2136 8900 2188 8906
rect 2136 8842 2188 8848
rect 2148 8362 2176 8842
rect 2240 8566 2268 8910
rect 2332 8906 2452 8922
rect 2332 8900 2464 8906
rect 2332 8894 2412 8900
rect 2412 8842 2464 8848
rect 2424 8634 2452 8842
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2700 8566 2728 8978
rect 2884 8634 2912 10610
rect 3068 8838 3096 10610
rect 3436 10577 3464 10610
rect 3422 10568 3478 10577
rect 3422 10503 3478 10512
rect 3436 10266 3464 10503
rect 3528 10470 3556 10610
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3528 9722 3556 10406
rect 3896 9976 3924 10678
rect 3988 10674 4016 12406
rect 4632 12238 4660 12718
rect 4620 12232 4672 12238
rect 4526 12200 4582 12209
rect 4344 12164 4396 12170
rect 4344 12106 4396 12112
rect 4436 12164 4488 12170
rect 4620 12174 4672 12180
rect 4526 12135 4582 12144
rect 4436 12106 4488 12112
rect 4356 11762 4384 12106
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4448 11626 4476 12106
rect 4540 12102 4568 12135
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4632 11898 4660 12174
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4436 11620 4488 11626
rect 4436 11562 4488 11568
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4540 10810 4568 11086
rect 4632 11082 4660 11698
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4434 10704 4490 10713
rect 3976 10668 4028 10674
rect 4724 10674 4752 12106
rect 4816 11694 4844 12804
rect 5276 12832 5304 13348
rect 5630 13288 5686 13297
rect 5630 13223 5686 13232
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5368 12918 5396 13126
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5224 12804 5304 12832
rect 5172 12786 5224 12792
rect 5078 12744 5134 12753
rect 5078 12679 5134 12688
rect 5092 12170 5120 12679
rect 5184 12170 5212 12786
rect 5644 12782 5672 13223
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 5630 12608 5686 12617
rect 5630 12543 5686 12552
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 5172 12164 5224 12170
rect 5172 12106 5224 12112
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4434 10639 4436 10648
rect 3976 10610 4028 10616
rect 4488 10639 4490 10648
rect 4712 10668 4764 10674
rect 4436 10610 4488 10616
rect 4712 10610 4764 10616
rect 3988 10248 4016 10610
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4068 10260 4120 10266
rect 3988 10220 4068 10248
rect 4068 10202 4120 10208
rect 4080 10044 4108 10202
rect 4160 10056 4212 10062
rect 4080 10016 4160 10044
rect 4160 9998 4212 10004
rect 3976 9988 4028 9994
rect 3896 9948 3976 9976
rect 3976 9930 4028 9936
rect 3516 9716 3568 9722
rect 3516 9658 3568 9664
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2228 8560 2280 8566
rect 2228 8502 2280 8508
rect 2688 8560 2740 8566
rect 2740 8520 2820 8548
rect 2688 8502 2740 8508
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 2792 8090 2820 8520
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2688 8016 2740 8022
rect 2608 7964 2688 7970
rect 2740 7964 2820 7970
rect 2608 7942 2820 7964
rect 2976 7954 3004 8570
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2056 7410 2084 7822
rect 2608 7546 2636 7942
rect 2792 7818 2820 7942
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2780 7812 2832 7818
rect 2780 7754 2832 7760
rect 2964 7812 3016 7818
rect 2964 7754 3016 7760
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2608 7410 2636 7482
rect 2700 7410 2728 7686
rect 2884 7546 2912 7686
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2780 7472 2832 7478
rect 2780 7414 2832 7420
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 846 6352 902 6361
rect 846 6287 848 6296
rect 900 6287 902 6296
rect 848 6258 900 6264
rect 1412 5710 1440 6734
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 1688 6458 1716 6666
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1688 5710 1716 6054
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1412 5166 1440 5646
rect 1872 5545 1900 6258
rect 2792 5914 2820 7414
rect 2884 6254 2912 7482
rect 2976 7410 3004 7754
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 1858 5536 1914 5545
rect 1858 5471 1914 5480
rect 3068 5370 3096 8434
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3160 7478 3188 7822
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1306 4856 1362 4865
rect 1306 4791 1362 4800
rect 1320 4146 1348 4791
rect 1412 4622 1440 5102
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1308 4140 1360 4146
rect 1308 4082 1360 4088
rect 1412 3126 1440 4558
rect 1504 4282 1532 5170
rect 3068 4622 3096 5306
rect 3252 4826 3280 8910
rect 3344 7478 3372 8910
rect 3436 7478 3464 8910
rect 3528 8566 3556 9658
rect 3988 9518 4016 9930
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4356 9722 4384 9862
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 4632 9450 4660 10474
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 4724 9994 4752 10134
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4816 9926 4844 11630
rect 5276 11393 5304 12038
rect 5354 11928 5410 11937
rect 5354 11863 5356 11872
rect 5408 11863 5410 11872
rect 5356 11834 5408 11840
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5354 11520 5410 11529
rect 5354 11455 5410 11464
rect 5262 11384 5318 11393
rect 5262 11319 5318 11328
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5276 10985 5304 11086
rect 5368 11014 5396 11455
rect 5356 11008 5408 11014
rect 5262 10976 5318 10985
rect 5356 10950 5408 10956
rect 4874 10908 5182 10917
rect 5262 10911 5318 10920
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 5092 10470 5120 10746
rect 5356 10736 5408 10742
rect 5356 10678 5408 10684
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5276 10577 5304 10610
rect 5262 10568 5318 10577
rect 5262 10503 5318 10512
rect 5080 10464 5132 10470
rect 4986 10432 5042 10441
rect 5080 10406 5132 10412
rect 4986 10367 5042 10376
rect 5000 10198 5028 10367
rect 4988 10192 5040 10198
rect 4988 10134 5040 10140
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4620 9444 4672 9450
rect 4620 9386 4672 9392
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4816 9217 4844 9862
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4802 9208 4858 9217
rect 4802 9143 4858 9152
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3516 8560 3568 8566
rect 3516 8502 3568 8508
rect 3620 8412 3648 8978
rect 3700 8900 3752 8906
rect 3700 8842 3752 8848
rect 3528 8384 3648 8412
rect 3528 7546 3556 8384
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3620 7478 3648 8026
rect 3712 8022 3740 8842
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3700 8016 3752 8022
rect 3700 7958 3752 7964
rect 3332 7472 3384 7478
rect 3332 7414 3384 7420
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3608 7472 3660 7478
rect 3608 7414 3660 7420
rect 3344 7002 3372 7414
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 3436 6322 3464 7414
rect 3712 6390 3740 7958
rect 3804 7274 3832 8230
rect 3896 7886 3924 8774
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3896 7546 3924 7822
rect 3988 7750 4016 9046
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4080 7954 4108 8298
rect 4172 8294 4200 8774
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3988 7546 4016 7686
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 4080 7478 4108 7890
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 4448 7410 4476 7754
rect 4632 7410 4660 8842
rect 4816 7886 4844 8910
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4986 8528 5042 8537
rect 4986 8463 4988 8472
rect 5040 8463 5042 8472
rect 4988 8434 5040 8440
rect 5276 8430 5304 10503
rect 5368 9489 5396 10678
rect 5460 10588 5488 11698
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5552 10742 5580 11086
rect 5644 11082 5672 12543
rect 5736 12442 5764 14894
rect 5920 14890 5948 15438
rect 5908 14884 5960 14890
rect 5908 14826 5960 14832
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 6012 14550 6040 14758
rect 6196 14618 6224 15642
rect 7104 15632 7156 15638
rect 7104 15574 7156 15580
rect 7286 15600 7342 15609
rect 6828 15428 6880 15434
rect 6828 15370 6880 15376
rect 6736 15088 6788 15094
rect 6736 15030 6788 15036
rect 6644 14952 6696 14958
rect 6642 14920 6644 14929
rect 6696 14920 6698 14929
rect 6642 14855 6698 14864
rect 6368 14816 6420 14822
rect 6552 14816 6604 14822
rect 6368 14758 6420 14764
rect 6550 14784 6552 14793
rect 6604 14784 6606 14793
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 6000 14544 6052 14550
rect 6000 14486 6052 14492
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5828 12850 5856 13398
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5828 12753 5856 12786
rect 5814 12744 5870 12753
rect 5814 12679 5870 12688
rect 5724 12436 5776 12442
rect 5920 12434 5948 13874
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6012 13326 6040 13670
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 6012 12646 6040 13262
rect 6092 13252 6144 13258
rect 6092 13194 6144 13200
rect 6104 12986 6132 13194
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 6104 12481 6132 12786
rect 5724 12378 5776 12384
rect 5828 12406 5948 12434
rect 6090 12472 6146 12481
rect 6090 12407 6146 12416
rect 5736 12345 5764 12378
rect 5722 12336 5778 12345
rect 5722 12271 5778 12280
rect 5632 11076 5684 11082
rect 5684 11036 5764 11064
rect 5632 11018 5684 11024
rect 5630 10976 5686 10985
rect 5630 10911 5686 10920
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5460 10560 5580 10588
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5460 9994 5488 10066
rect 5552 10062 5580 10560
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 5354 9480 5410 9489
rect 5354 9415 5410 9424
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5368 8945 5396 9318
rect 5460 9042 5488 9930
rect 5644 9761 5672 10911
rect 5736 10577 5764 11036
rect 5722 10568 5778 10577
rect 5722 10503 5778 10512
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5630 9752 5686 9761
rect 5630 9687 5686 9696
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5644 8974 5672 9687
rect 5736 9654 5764 10406
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5632 8968 5684 8974
rect 5354 8936 5410 8945
rect 5632 8910 5684 8916
rect 5354 8871 5410 8880
rect 5448 8900 5500 8906
rect 5500 8860 5580 8888
rect 5448 8842 5500 8848
rect 5552 8566 5580 8860
rect 5540 8560 5592 8566
rect 5446 8528 5502 8537
rect 5540 8502 5592 8508
rect 5446 8463 5502 8472
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5354 8392 5410 8401
rect 5354 8327 5356 8336
rect 5408 8327 5410 8336
rect 5356 8298 5408 8304
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 7886 5120 8230
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 5368 7886 5396 7958
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 5080 7880 5132 7886
rect 5356 7880 5408 7886
rect 5132 7840 5304 7868
rect 5080 7822 5132 7828
rect 4816 7546 4844 7822
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 3792 7268 3844 7274
rect 3792 7210 3844 7216
rect 3804 6458 3832 7210
rect 4080 6798 4108 7278
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 5000 6798 5028 7482
rect 5080 7404 5132 7410
rect 5276 7392 5304 7840
rect 5356 7822 5408 7828
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5132 7364 5304 7392
rect 5080 7346 5132 7352
rect 5368 7206 5396 7686
rect 5460 7546 5488 8463
rect 5552 8022 5580 8502
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4988 6792 5040 6798
rect 5356 6792 5408 6798
rect 5040 6752 5304 6780
rect 4988 6734 5040 6740
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3700 6384 3752 6390
rect 3700 6326 3752 6332
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3436 5710 3464 6258
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3620 5846 3648 6190
rect 3608 5840 3660 5846
rect 3608 5782 3660 5788
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3344 5234 3372 5578
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3436 5166 3464 5646
rect 3712 5574 3740 6326
rect 3804 6186 3832 6394
rect 4724 6322 4752 6666
rect 4816 6390 4844 6734
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 5276 6322 5304 6752
rect 5460 6780 5488 7346
rect 5552 7342 5580 7958
rect 5644 7954 5672 8910
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5632 7812 5684 7818
rect 5632 7754 5684 7760
rect 5644 7410 5672 7754
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5408 6752 5488 6780
rect 5356 6734 5408 6740
rect 5460 6322 5488 6752
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 3792 6180 3844 6186
rect 3792 6122 3844 6128
rect 3804 5778 3832 6122
rect 3792 5772 3844 5778
rect 3792 5714 3844 5720
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3712 5234 3740 5510
rect 3804 5302 3832 5714
rect 3896 5642 3924 6258
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3988 5710 4016 6190
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 3792 5296 3844 5302
rect 3792 5238 3844 5244
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3712 5098 3740 5170
rect 3700 5092 3752 5098
rect 3700 5034 3752 5040
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 3712 4554 3740 5034
rect 3804 4826 3832 5238
rect 3896 5098 3924 5578
rect 3988 5234 4016 5646
rect 4632 5574 4660 6258
rect 4724 5914 4752 6258
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 3976 5228 4028 5234
rect 4080 5216 4108 5510
rect 4816 5234 4844 6190
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5170 5264 5226 5273
rect 4252 5228 4304 5234
rect 4080 5188 4252 5216
rect 3976 5170 4028 5176
rect 4252 5170 4304 5176
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4896 5228 4948 5234
rect 5170 5199 5172 5208
rect 4896 5170 4948 5176
rect 5224 5199 5226 5208
rect 5276 5216 5304 6258
rect 5356 5228 5408 5234
rect 5276 5188 5356 5216
rect 5172 5170 5224 5176
rect 5460 5216 5488 6258
rect 5552 5692 5580 7278
rect 5630 6760 5686 6769
rect 5630 6695 5686 6704
rect 5644 6662 5672 6695
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5736 5846 5764 9454
rect 5828 9042 5856 12406
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5908 11688 5960 11694
rect 5906 11656 5908 11665
rect 5960 11656 5962 11665
rect 5906 11591 5962 11600
rect 6012 11558 6040 12038
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 5920 10198 5948 11494
rect 5908 10192 5960 10198
rect 5908 10134 5960 10140
rect 5908 10056 5960 10062
rect 5960 10016 6040 10044
rect 5908 9998 5960 10004
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5828 8430 5856 8978
rect 5920 8974 5948 9862
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5920 8838 5948 8910
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5920 8294 5948 8774
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5816 8016 5868 8022
rect 5816 7958 5868 7964
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5632 5704 5684 5710
rect 5552 5664 5632 5692
rect 5632 5646 5684 5652
rect 5722 5672 5778 5681
rect 5722 5607 5724 5616
rect 5776 5607 5778 5616
rect 5724 5578 5776 5584
rect 5828 5409 5856 7958
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5920 6798 5948 7822
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5814 5400 5870 5409
rect 5814 5335 5870 5344
rect 5828 5234 5856 5335
rect 5632 5228 5684 5234
rect 5460 5188 5632 5216
rect 5356 5170 5408 5176
rect 5632 5170 5684 5176
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 3884 5092 3936 5098
rect 3884 5034 3936 5040
rect 3988 4826 4016 5170
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 4080 4826 4108 5034
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4908 4826 4936 5170
rect 5368 4826 5396 5170
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 4080 4622 4108 4762
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 1688 4282 1716 4490
rect 5644 4486 5672 5170
rect 5920 4758 5948 6734
rect 6012 6254 6040 10016
rect 6104 8090 6132 12407
rect 6196 11286 6224 14554
rect 6276 13456 6328 13462
rect 6274 13424 6276 13433
rect 6328 13424 6330 13433
rect 6274 13359 6330 13368
rect 6276 13252 6328 13258
rect 6276 13194 6328 13200
rect 6288 12918 6316 13194
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6288 12646 6316 12854
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6288 11898 6316 12378
rect 6380 12374 6408 14758
rect 6550 14719 6606 14728
rect 6644 14340 6696 14346
rect 6644 14282 6696 14288
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6472 12850 6500 13262
rect 6656 13258 6684 14282
rect 6748 13326 6776 15030
rect 6840 15026 6868 15370
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6840 14618 6868 14962
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 7024 14074 7052 14758
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 6840 13734 6868 13874
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 7024 13530 7052 14010
rect 7116 13818 7144 15574
rect 7286 15535 7342 15544
rect 7300 15094 7328 15535
rect 7564 15156 7616 15162
rect 7484 15116 7564 15144
rect 7288 15088 7340 15094
rect 7288 15030 7340 15036
rect 7300 14958 7328 15030
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7484 14890 7512 15116
rect 7564 15098 7616 15104
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7472 14884 7524 14890
rect 7472 14826 7524 14832
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7208 13938 7236 14350
rect 7288 14000 7340 14006
rect 7288 13942 7340 13948
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 7116 13790 7236 13818
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7116 13530 7144 13670
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6748 13138 6776 13262
rect 6564 13110 6776 13138
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6368 12368 6420 12374
rect 6368 12310 6420 12316
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6274 11656 6330 11665
rect 6274 11591 6330 11600
rect 6184 11280 6236 11286
rect 6184 11222 6236 11228
rect 6288 11150 6316 11591
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6274 10160 6330 10169
rect 6274 10095 6276 10104
rect 6328 10095 6330 10104
rect 6276 10066 6328 10072
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6274 10024 6330 10033
rect 6196 9353 6224 9998
rect 6274 9959 6330 9968
rect 6288 9654 6316 9959
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6182 9344 6238 9353
rect 6182 9279 6238 9288
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6196 8838 6224 9114
rect 6288 8974 6316 9590
rect 6380 9330 6408 12106
rect 6460 12096 6512 12102
rect 6458 12064 6460 12073
rect 6512 12064 6514 12073
rect 6458 11999 6514 12008
rect 6460 11280 6512 11286
rect 6460 11222 6512 11228
rect 6472 10062 6500 11222
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6472 9625 6500 9862
rect 6458 9616 6514 9625
rect 6458 9551 6514 9560
rect 6564 9518 6592 13110
rect 6840 12306 6868 13126
rect 6932 12617 6960 13398
rect 7208 13326 7236 13790
rect 7300 13394 7328 13942
rect 7576 13734 7604 14962
rect 7564 13728 7616 13734
rect 7564 13670 7616 13676
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7196 13320 7248 13326
rect 7194 13288 7196 13297
rect 7248 13288 7250 13297
rect 7194 13223 7250 13232
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 7024 12918 7052 13126
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 7300 12850 7328 13330
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7576 12986 7604 13262
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 6918 12608 6974 12617
rect 6918 12543 6974 12552
rect 7116 12424 7144 12786
rect 7300 12617 7328 12786
rect 7392 12753 7420 12786
rect 7378 12744 7434 12753
rect 7576 12714 7604 12922
rect 7378 12679 7434 12688
rect 7564 12708 7616 12714
rect 7286 12608 7342 12617
rect 7286 12543 7342 12552
rect 6932 12396 7144 12424
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6932 12238 6960 12396
rect 7392 12322 7420 12679
rect 7564 12650 7616 12656
rect 7562 12608 7618 12617
rect 7562 12543 7618 12552
rect 7024 12294 7420 12322
rect 6920 12232 6972 12238
rect 6734 12200 6790 12209
rect 6734 12135 6790 12144
rect 6840 12180 6920 12186
rect 6840 12174 6972 12180
rect 6840 12158 6960 12174
rect 6748 11898 6776 12135
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6748 10452 6776 11086
rect 6840 10656 6868 12158
rect 7024 12102 7052 12294
rect 7104 12232 7156 12238
rect 7102 12200 7104 12209
rect 7288 12232 7340 12238
rect 7156 12200 7158 12209
rect 7288 12174 7340 12180
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7102 12135 7158 12144
rect 7196 12164 7248 12170
rect 7116 12102 7144 12135
rect 7196 12106 7248 12112
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 6918 11248 6974 11257
rect 6918 11183 6974 11192
rect 6932 11150 6960 11183
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 7024 10996 7052 12038
rect 7208 11898 7236 12106
rect 7300 11898 7328 12174
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7116 11121 7144 11698
rect 7102 11112 7158 11121
rect 7102 11047 7158 11056
rect 7104 11008 7156 11014
rect 7024 10968 7104 10996
rect 7104 10950 7156 10956
rect 7116 10674 7144 10950
rect 6920 10668 6972 10674
rect 6840 10628 6920 10656
rect 7104 10668 7156 10674
rect 6972 10628 7052 10656
rect 6920 10610 6972 10616
rect 6748 10424 6960 10452
rect 6642 10296 6698 10305
rect 6642 10231 6698 10240
rect 6656 10198 6684 10231
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6552 9512 6604 9518
rect 6656 9489 6684 9522
rect 6552 9454 6604 9460
rect 6642 9480 6698 9489
rect 6642 9415 6698 9424
rect 6748 9382 6776 9862
rect 6644 9376 6696 9382
rect 6380 9302 6500 9330
rect 6644 9318 6696 9324
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6196 7970 6224 8298
rect 6288 8022 6316 8910
rect 6104 7942 6224 7970
rect 6276 8016 6328 8022
rect 6276 7958 6328 7964
rect 6104 7478 6132 7942
rect 6184 7880 6236 7886
rect 6288 7868 6316 7958
rect 6236 7840 6316 7868
rect 6184 7822 6236 7828
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 6092 6996 6144 7002
rect 6092 6938 6144 6944
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 6104 5574 6132 6938
rect 6196 5681 6224 7822
rect 6380 6866 6408 9114
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 6288 6458 6316 6666
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6472 6361 6500 9302
rect 6656 9178 6684 9318
rect 6748 9217 6776 9318
rect 6734 9208 6790 9217
rect 6644 9172 6696 9178
rect 6734 9143 6790 9152
rect 6644 9114 6696 9120
rect 6550 9072 6606 9081
rect 6550 9007 6606 9016
rect 6564 8974 6592 9007
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6564 7750 6592 8910
rect 6656 8566 6684 8910
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6748 8634 6776 8842
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 6656 8022 6684 8502
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6458 6352 6514 6361
rect 6458 6287 6514 6296
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6380 5710 6408 6054
rect 6472 5778 6500 6287
rect 6644 5840 6696 5846
rect 6644 5782 6696 5788
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6276 5704 6328 5710
rect 6182 5672 6238 5681
rect 6276 5646 6328 5652
rect 6368 5704 6420 5710
rect 6552 5704 6604 5710
rect 6368 5646 6420 5652
rect 6458 5672 6514 5681
rect 6182 5607 6238 5616
rect 6092 5568 6144 5574
rect 6288 5545 6316 5646
rect 6552 5646 6604 5652
rect 6458 5607 6514 5616
rect 6092 5510 6144 5516
rect 6274 5536 6330 5545
rect 6274 5471 6330 5480
rect 6000 5160 6052 5166
rect 6288 5148 6316 5471
rect 6366 5400 6422 5409
rect 6366 5335 6422 5344
rect 6380 5234 6408 5335
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6472 5166 6500 5607
rect 6564 5545 6592 5646
rect 6550 5536 6606 5545
rect 6550 5471 6606 5480
rect 6550 5400 6606 5409
rect 6550 5335 6606 5344
rect 6564 5234 6592 5335
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6052 5120 6316 5148
rect 6460 5160 6512 5166
rect 6000 5102 6052 5108
rect 6460 5102 6512 5108
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 6104 4282 6132 4966
rect 6472 4690 6500 5102
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 1492 4276 1544 4282
rect 1492 4218 1544 4224
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 1858 4176 1914 4185
rect 6380 4146 6408 4422
rect 6564 4146 6592 4762
rect 1858 4111 1860 4120
rect 1912 4111 1914 4120
rect 6368 4140 6420 4146
rect 1860 4082 1912 4088
rect 6368 4082 6420 4088
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 1400 3120 1452 3126
rect 1400 3062 1452 3068
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 6472 2650 6500 2994
rect 6656 2854 6684 5782
rect 6734 5672 6790 5681
rect 6734 5607 6736 5616
rect 6788 5607 6790 5616
rect 6736 5578 6788 5584
rect 6736 4752 6788 4758
rect 6736 4694 6788 4700
rect 6748 4146 6776 4694
rect 6840 4690 6868 9930
rect 6932 9518 6960 10424
rect 7024 10169 7052 10628
rect 7104 10610 7156 10616
rect 7116 10266 7144 10610
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7010 10160 7066 10169
rect 7010 10095 7066 10104
rect 7024 10062 7052 10095
rect 7116 10062 7144 10202
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7208 9994 7236 11834
rect 7300 11801 7328 11834
rect 7392 11830 7420 12174
rect 7380 11824 7432 11830
rect 7286 11792 7342 11801
rect 7380 11766 7432 11772
rect 7286 11727 7342 11736
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7300 11529 7328 11630
rect 7286 11520 7342 11529
rect 7286 11455 7342 11464
rect 7392 11354 7420 11766
rect 7472 11620 7524 11626
rect 7472 11562 7524 11568
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7288 11280 7340 11286
rect 7288 11222 7340 11228
rect 7300 10674 7328 11222
rect 7392 10674 7420 11290
rect 7484 11150 7512 11562
rect 7576 11529 7604 12543
rect 7668 12442 7696 15642
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 7852 14890 7880 14962
rect 7840 14884 7892 14890
rect 7840 14826 7892 14832
rect 7840 13864 7892 13870
rect 7838 13832 7840 13841
rect 7892 13832 7894 13841
rect 7838 13767 7894 13776
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7668 11626 7696 12106
rect 7760 11665 7788 13330
rect 7852 12850 7880 13466
rect 7944 13376 7972 15506
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8312 14958 8340 15438
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8024 14000 8076 14006
rect 8128 13977 8156 14758
rect 8220 14414 8248 14758
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8220 14074 8248 14350
rect 8312 14278 8340 14350
rect 8392 14340 8444 14346
rect 8392 14282 8444 14288
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8024 13942 8076 13948
rect 8114 13968 8170 13977
rect 8036 13530 8064 13942
rect 8312 13938 8340 14214
rect 8404 13938 8432 14282
rect 8114 13903 8170 13912
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 7944 13348 8156 13376
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 8036 13161 8064 13194
rect 8022 13152 8078 13161
rect 8022 13087 8078 13096
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7746 11656 7802 11665
rect 7656 11620 7708 11626
rect 7746 11591 7802 11600
rect 7656 11562 7708 11568
rect 7562 11520 7618 11529
rect 7562 11455 7618 11464
rect 7576 11218 7604 11455
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7668 10849 7696 11290
rect 7852 11082 7880 12786
rect 8036 12782 8064 13087
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 7944 12442 7972 12650
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 8128 12050 8156 13348
rect 8220 13326 8248 13738
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 8036 12022 8156 12050
rect 7930 11520 7986 11529
rect 7930 11455 7986 11464
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7654 10840 7710 10849
rect 7484 10810 7654 10826
rect 7472 10804 7654 10810
rect 7524 10798 7654 10804
rect 7654 10775 7710 10784
rect 7472 10746 7524 10752
rect 7656 10736 7708 10742
rect 7470 10704 7526 10713
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7380 10668 7432 10674
rect 7656 10678 7708 10684
rect 7470 10639 7526 10648
rect 7380 10610 7432 10616
rect 7300 10554 7328 10610
rect 7484 10554 7512 10639
rect 7668 10606 7696 10678
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7300 10526 7512 10554
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6932 8362 6960 9454
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 7024 9217 7052 9386
rect 7010 9208 7066 9217
rect 7010 9143 7066 9152
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 7116 6934 7144 9658
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 7116 6322 7144 6870
rect 7208 6866 7236 9930
rect 7300 9602 7328 10526
rect 7378 10432 7434 10441
rect 7378 10367 7434 10376
rect 7562 10432 7618 10441
rect 7562 10367 7618 10376
rect 7392 10062 7420 10367
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7392 9722 7420 9998
rect 7484 9761 7512 9998
rect 7470 9752 7526 9761
rect 7380 9716 7432 9722
rect 7470 9687 7526 9696
rect 7380 9658 7432 9664
rect 7576 9654 7604 10367
rect 7668 9654 7696 10542
rect 7564 9648 7616 9654
rect 7484 9608 7564 9636
rect 7300 9586 7420 9602
rect 7300 9580 7432 9586
rect 7300 9574 7380 9580
rect 7380 9522 7432 9528
rect 7286 9344 7342 9353
rect 7286 9279 7342 9288
rect 7300 8906 7328 9279
rect 7392 8974 7420 9522
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7300 6798 7328 8842
rect 7392 8566 7420 8910
rect 7380 8560 7432 8566
rect 7484 8537 7512 9608
rect 7564 9590 7616 9596
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7668 9160 7696 9590
rect 7576 9132 7696 9160
rect 7576 8974 7604 9132
rect 7760 9081 7788 10610
rect 7852 9761 7880 11018
rect 7838 9752 7894 9761
rect 7838 9687 7894 9696
rect 7746 9072 7802 9081
rect 7746 9007 7802 9016
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7380 8502 7432 8508
rect 7470 8528 7526 8537
rect 7576 8498 7604 8910
rect 7656 8900 7708 8906
rect 7656 8842 7708 8848
rect 7668 8498 7696 8842
rect 7852 8634 7880 9687
rect 7944 9586 7972 11455
rect 8036 11370 8064 12022
rect 8114 11928 8170 11937
rect 8114 11863 8170 11872
rect 8128 11830 8156 11863
rect 8116 11824 8168 11830
rect 8116 11766 8168 11772
rect 8036 11354 8156 11370
rect 8036 11348 8168 11354
rect 8036 11342 8116 11348
rect 8116 11290 8168 11296
rect 8024 11280 8076 11286
rect 8024 11222 8076 11228
rect 8036 10713 8064 11222
rect 8220 11132 8248 12922
rect 8390 12472 8446 12481
rect 8496 12442 8524 14554
rect 8390 12407 8446 12416
rect 8484 12436 8536 12442
rect 8404 12238 8432 12407
rect 8484 12378 8536 12384
rect 8496 12306 8524 12378
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8496 11694 8524 12106
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8220 11104 8340 11132
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 8128 10742 8156 11018
rect 8116 10736 8168 10742
rect 8022 10704 8078 10713
rect 8312 10724 8340 11104
rect 8312 10696 8432 10724
rect 8116 10678 8168 10684
rect 8022 10639 8024 10648
rect 8076 10639 8078 10648
rect 8024 10610 8076 10616
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 8128 10305 8156 10474
rect 8114 10296 8170 10305
rect 8114 10231 8170 10240
rect 8404 10146 8432 10696
rect 8496 10554 8524 11630
rect 8588 10742 8616 17031
rect 12544 16794 12572 17138
rect 13280 16998 13308 17546
rect 14752 17338 14780 17546
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 15200 17264 15252 17270
rect 15200 17206 15252 17212
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 13280 16658 13308 16934
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 11980 16176 12032 16182
rect 11980 16118 12032 16124
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9140 15609 9168 15642
rect 9126 15600 9182 15609
rect 9126 15535 9182 15544
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9140 15162 9168 15438
rect 9128 15156 9180 15162
rect 9048 15116 9128 15144
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8772 13870 8800 14554
rect 8956 14346 8984 14758
rect 8944 14340 8996 14346
rect 8944 14282 8996 14288
rect 8956 14249 8984 14282
rect 8942 14240 8998 14249
rect 8942 14175 8998 14184
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8772 12918 8800 13806
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8942 12880 8998 12889
rect 8942 12815 8998 12824
rect 8956 12782 8984 12815
rect 8944 12776 8996 12782
rect 9048 12753 9076 15116
rect 9128 15098 9180 15104
rect 9600 15026 9628 15438
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 8944 12718 8996 12724
rect 9034 12744 9090 12753
rect 8956 12238 8984 12718
rect 9034 12679 9090 12688
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 9048 11762 9076 12106
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8496 10526 8616 10554
rect 8220 10118 8432 10146
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8022 9616 8078 9625
rect 7932 9580 7984 9586
rect 8022 9551 8078 9560
rect 7932 9522 7984 9528
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7470 8463 7526 8472
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7208 6390 7236 6666
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7208 6186 7236 6326
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 7300 6118 7328 6190
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7392 5914 7420 7822
rect 7484 7342 7512 7890
rect 7576 7886 7604 8298
rect 7654 8120 7710 8129
rect 7654 8055 7710 8064
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7576 7002 7604 7822
rect 7564 6996 7616 7002
rect 7484 6956 7564 6984
rect 7484 6497 7512 6956
rect 7564 6938 7616 6944
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7470 6488 7526 6497
rect 7470 6423 7526 6432
rect 7576 6390 7604 6734
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 7576 6186 7604 6326
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7104 5636 7156 5642
rect 7104 5578 7156 5584
rect 7116 5234 7144 5578
rect 7392 5302 7420 5714
rect 7380 5296 7432 5302
rect 7286 5264 7342 5273
rect 7104 5228 7156 5234
rect 7380 5238 7432 5244
rect 7286 5199 7342 5208
rect 7104 5170 7156 5176
rect 7116 4758 7144 5170
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6840 3738 6868 4626
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 7208 3466 7236 4014
rect 7196 3460 7248 3466
rect 7196 3402 7248 3408
rect 7300 3398 7328 5199
rect 7484 4298 7512 6054
rect 7576 5846 7604 6122
rect 7564 5840 7616 5846
rect 7564 5782 7616 5788
rect 7668 5710 7696 8055
rect 7852 6798 7880 8434
rect 7944 8362 7972 9522
rect 8036 9042 8064 9551
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8036 8498 8064 8978
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 8022 8120 8078 8129
rect 8022 8055 8078 8064
rect 8036 7886 8064 8055
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7840 6792 7892 6798
rect 7760 6752 7840 6780
rect 7760 6458 7788 6752
rect 7840 6734 7892 6740
rect 7944 6730 7972 7822
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 8036 6798 8064 7686
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 7932 6724 7984 6730
rect 7932 6666 7984 6672
rect 7838 6488 7894 6497
rect 7748 6452 7800 6458
rect 7838 6423 7894 6432
rect 7748 6394 7800 6400
rect 7760 6322 7788 6394
rect 7852 6390 7880 6423
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7852 5846 7880 6190
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7668 5409 7696 5646
rect 7654 5400 7710 5409
rect 7852 5352 7880 5782
rect 7654 5335 7710 5344
rect 7668 5234 7696 5335
rect 7760 5324 7880 5352
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7576 5114 7604 5170
rect 7760 5114 7788 5324
rect 7944 5302 7972 6666
rect 8036 5817 8064 6734
rect 8022 5808 8078 5817
rect 8022 5743 8078 5752
rect 8036 5409 8064 5743
rect 8022 5400 8078 5409
rect 8022 5335 8078 5344
rect 7932 5296 7984 5302
rect 7932 5238 7984 5244
rect 8036 5234 8064 5335
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7576 5086 7788 5114
rect 7852 4622 7880 5170
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 8036 4690 8064 4966
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 8128 4622 8156 9930
rect 8220 8129 8248 10118
rect 8300 10056 8352 10062
rect 8484 10056 8536 10062
rect 8352 10016 8432 10044
rect 8300 9998 8352 10004
rect 8298 9752 8354 9761
rect 8298 9687 8354 9696
rect 8312 9654 8340 9687
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8404 9586 8432 10016
rect 8482 10024 8484 10033
rect 8536 10024 8538 10033
rect 8482 9959 8538 9968
rect 8588 9908 8616 10526
rect 8680 10470 8708 11698
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 8760 10192 8812 10198
rect 8864 10169 8892 11018
rect 8956 11014 8984 11698
rect 9036 11620 9088 11626
rect 9036 11562 9088 11568
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8760 10134 8812 10140
rect 8850 10160 8906 10169
rect 8496 9880 8616 9908
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8390 9208 8446 9217
rect 8390 9143 8446 9152
rect 8404 9042 8432 9143
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8312 8945 8340 8978
rect 8496 8974 8524 9880
rect 8680 9722 8708 10134
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8680 9382 8708 9658
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8588 8974 8616 9318
rect 8772 9178 8800 10134
rect 8850 10095 8906 10104
rect 8864 9926 8892 10095
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8484 8968 8536 8974
rect 8298 8936 8354 8945
rect 8484 8910 8536 8916
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8298 8871 8354 8880
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8576 8832 8628 8838
rect 8628 8792 8708 8820
rect 8576 8774 8628 8780
rect 8312 8634 8340 8774
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8206 8120 8262 8129
rect 8206 8055 8262 8064
rect 8206 7984 8262 7993
rect 8206 7919 8262 7928
rect 8220 7886 8248 7919
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8220 5710 8248 7822
rect 8312 6322 8340 8434
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8392 8016 8444 8022
rect 8444 7976 8524 8004
rect 8392 7958 8444 7964
rect 8496 7886 8524 7976
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8404 7041 8432 7346
rect 8390 7032 8446 7041
rect 8390 6967 8446 6976
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 8404 6798 8432 6870
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8312 5914 8340 6258
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8404 5710 8432 6054
rect 8496 5914 8524 6258
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8220 5234 8248 5646
rect 8482 5264 8538 5273
rect 8208 5228 8260 5234
rect 8482 5199 8484 5208
rect 8208 5170 8260 5176
rect 8536 5199 8538 5208
rect 8484 5170 8536 5176
rect 8588 4690 8616 8230
rect 8680 7818 8708 8792
rect 8668 7812 8720 7818
rect 8668 7754 8720 7760
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8680 6372 8708 7142
rect 8772 7002 8800 9114
rect 8864 8906 8892 9522
rect 8956 9110 8984 9522
rect 9048 9466 9076 11562
rect 9140 9586 9168 14962
rect 9600 14618 9628 14962
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 9232 13734 9260 14350
rect 9416 14006 9444 14418
rect 9404 14000 9456 14006
rect 9404 13942 9456 13948
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9232 12714 9260 13126
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9232 12442 9260 12650
rect 9220 12436 9272 12442
rect 9324 12434 9352 13670
rect 9324 12406 9444 12434
rect 9220 12378 9272 12384
rect 9416 12374 9444 12406
rect 9404 12368 9456 12374
rect 9218 12336 9274 12345
rect 9404 12310 9456 12316
rect 9218 12271 9220 12280
rect 9272 12271 9274 12280
rect 9220 12242 9272 12248
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9324 10062 9352 10406
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9232 9654 9260 9998
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9220 9512 9272 9518
rect 9048 9438 9168 9466
rect 9220 9454 9272 9460
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8864 6798 8892 7346
rect 8956 7342 8984 9046
rect 9048 8634 9076 9114
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 8942 6760 8998 6769
rect 8864 6458 8892 6734
rect 8942 6695 8944 6704
rect 8996 6695 8998 6704
rect 8944 6666 8996 6672
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8760 6384 8812 6390
rect 8680 6344 8760 6372
rect 8680 6118 8708 6344
rect 8760 6326 8812 6332
rect 8864 6254 8892 6394
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8666 5400 8722 5409
rect 8666 5335 8668 5344
rect 8720 5335 8722 5344
rect 8668 5306 8720 5312
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 7484 4270 7604 4298
rect 7668 4282 7696 4490
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7484 4078 7512 4150
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7484 3738 7512 4014
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7484 3534 7512 3674
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7576 3398 7604 4270
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7852 3942 7880 4014
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7852 3738 7880 3878
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7852 3194 7880 3674
rect 8128 3670 8156 4558
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8220 3670 8248 4150
rect 8956 3942 8984 6394
rect 9048 5914 9076 8570
rect 9140 7546 9168 9438
rect 9232 9178 9260 9454
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9324 8294 9352 9386
rect 9416 8498 9444 11018
rect 9508 10266 9536 13874
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9600 13326 9628 13670
rect 9692 13394 9720 15302
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9784 13530 9812 13670
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9784 12345 9812 13262
rect 9770 12336 9826 12345
rect 9770 12271 9826 12280
rect 9772 12232 9824 12238
rect 9692 12192 9772 12220
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9048 5234 9076 5510
rect 9140 5234 9168 7346
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 9140 3738 9168 4082
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8024 3528 8076 3534
rect 8220 3482 8248 3606
rect 8024 3470 8076 3476
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7852 3058 7880 3130
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 8036 2990 8064 3470
rect 8128 3466 8248 3482
rect 8116 3460 8248 3466
rect 8168 3454 8248 3460
rect 8116 3402 8168 3408
rect 8220 3058 8248 3454
rect 9232 3126 9260 7686
rect 9310 7576 9366 7585
rect 9310 7511 9312 7520
rect 9364 7511 9366 7520
rect 9312 7482 9364 7488
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9324 7206 9352 7346
rect 9416 7274 9444 8434
rect 9404 7268 9456 7274
rect 9404 7210 9456 7216
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 9324 6458 9352 7142
rect 9404 6928 9456 6934
rect 9404 6870 9456 6876
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9310 6352 9366 6361
rect 9310 6287 9312 6296
rect 9364 6287 9366 6296
rect 9312 6258 9364 6264
rect 9416 5846 9444 6870
rect 9404 5840 9456 5846
rect 9310 5808 9366 5817
rect 9404 5782 9456 5788
rect 9310 5743 9366 5752
rect 9324 5710 9352 5743
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9324 3398 9352 5646
rect 9508 4758 9536 10066
rect 9600 8906 9628 12106
rect 9692 11694 9720 12192
rect 9772 12174 9824 12180
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9784 11218 9812 12038
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9586 8800 9642 8809
rect 9586 8735 9642 8744
rect 9600 8566 9628 8735
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9600 7002 9628 8502
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9600 6458 9628 6666
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9692 6202 9720 9862
rect 9784 9382 9812 10610
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9784 9042 9812 9318
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9784 8566 9812 8774
rect 9876 8634 9904 13806
rect 9968 9518 9996 14894
rect 10060 13530 10088 15982
rect 10244 15706 10272 16050
rect 10980 15706 11008 16050
rect 11060 15972 11112 15978
rect 11060 15914 11112 15920
rect 11888 15972 11940 15978
rect 11888 15914 11940 15920
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 11072 15638 11100 15914
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10140 15428 10192 15434
rect 10140 15370 10192 15376
rect 10152 15337 10180 15370
rect 10138 15328 10194 15337
rect 10138 15263 10194 15272
rect 10244 14074 10272 15506
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 15162 10456 15438
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9772 8560 9824 8566
rect 9968 8514 9996 9454
rect 10060 8838 10088 13330
rect 10152 12322 10180 13874
rect 10428 13394 10456 15098
rect 11072 14278 11100 15370
rect 11164 15026 11192 15642
rect 11428 15088 11480 15094
rect 11428 15030 11480 15036
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11164 14822 11192 14962
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11244 14544 11296 14550
rect 11244 14486 11296 14492
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11072 14074 11100 14214
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10508 13796 10560 13802
rect 10508 13738 10560 13744
rect 10520 13530 10548 13738
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10416 13388 10468 13394
rect 10468 13348 10548 13376
rect 10416 13330 10468 13336
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10152 12294 10272 12322
rect 10138 12200 10194 12209
rect 10138 12135 10194 12144
rect 10152 11558 10180 12135
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10152 10742 10180 11494
rect 10244 10985 10272 12294
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10336 11354 10364 11630
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10230 10976 10286 10985
rect 10230 10911 10286 10920
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 10336 10606 10364 11018
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10152 9382 10180 9522
rect 10230 9480 10286 9489
rect 10230 9415 10232 9424
rect 10284 9415 10286 9424
rect 10232 9386 10284 9392
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 9772 8502 9824 8508
rect 9876 8486 9996 8514
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9784 8090 9812 8230
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9784 7478 9812 7890
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 9876 7410 9904 8486
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9968 7954 9996 8366
rect 10152 8294 10180 9318
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 10060 7546 10088 7754
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10152 7410 10180 7686
rect 10244 7478 10272 8434
rect 10336 7886 10364 10542
rect 10428 9654 10456 13194
rect 10520 12986 10548 13348
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10704 12918 10732 13126
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10888 12850 10916 13670
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10520 12434 10548 12786
rect 10888 12442 10916 12786
rect 10966 12608 11022 12617
rect 10966 12543 11022 12552
rect 10692 12436 10744 12442
rect 10520 12406 10640 12434
rect 10612 12322 10640 12406
rect 10876 12436 10928 12442
rect 10744 12396 10824 12424
rect 10692 12378 10744 12384
rect 10612 12294 10732 12322
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10520 11354 10548 11698
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10428 8498 10456 8978
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10414 8392 10470 8401
rect 10414 8327 10470 8336
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 9770 7032 9826 7041
rect 9770 6967 9826 6976
rect 9784 6730 9812 6967
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9876 6662 9904 7346
rect 10152 7313 10180 7346
rect 10138 7304 10194 7313
rect 10138 7239 10194 7248
rect 10322 7304 10378 7313
rect 10322 7239 10378 7248
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9876 6322 9904 6598
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9692 6174 9904 6202
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9600 5216 9628 5850
rect 9680 5228 9732 5234
rect 9600 5188 9680 5216
rect 9680 5170 9732 5176
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9508 4146 9536 4694
rect 9692 4486 9720 4966
rect 9784 4826 9812 5170
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9692 4282 9720 4422
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9416 3534 9444 4082
rect 9876 3942 9904 6174
rect 9968 4622 9996 6938
rect 10230 6896 10286 6905
rect 10140 6860 10192 6866
rect 10230 6831 10286 6840
rect 10140 6802 10192 6808
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10060 6186 10088 6258
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 10060 5030 10088 6122
rect 10152 5234 10180 6802
rect 10244 5642 10272 6831
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10336 5302 10364 7239
rect 10428 5817 10456 8327
rect 10520 8022 10548 11154
rect 10612 11082 10640 12174
rect 10704 12102 10732 12294
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11558 10732 12038
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10612 10810 10640 11018
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10612 8566 10640 10406
rect 10704 10130 10732 10610
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10796 9518 10824 12396
rect 10876 12378 10928 12384
rect 10980 12374 11008 12543
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 11072 12238 11100 13874
rect 11060 12232 11112 12238
rect 11152 12232 11204 12238
rect 11060 12174 11112 12180
rect 11150 12200 11152 12209
rect 11204 12200 11206 12209
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10980 10674 11008 11630
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10704 8634 10732 8978
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10600 8288 10652 8294
rect 10600 8230 10652 8236
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 10612 7750 10640 8230
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10414 5808 10470 5817
rect 10414 5743 10470 5752
rect 10428 5710 10456 5743
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 10520 5370 10548 5578
rect 10612 5574 10640 5850
rect 10600 5568 10652 5574
rect 10600 5510 10652 5516
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10324 5296 10376 5302
rect 10324 5238 10376 5244
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10152 4214 10180 4422
rect 10140 4208 10192 4214
rect 10140 4150 10192 4156
rect 10612 4146 10640 5510
rect 10704 4758 10732 8434
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10336 3942 10364 4082
rect 10796 4078 10824 9454
rect 10888 9382 10916 10406
rect 11072 10266 11100 12174
rect 11150 12135 11206 12144
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10980 10130 11008 10202
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 10980 9761 11008 9930
rect 10966 9752 11022 9761
rect 10966 9687 11022 9696
rect 10980 9654 11008 9687
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 11164 9518 11192 9930
rect 11152 9512 11204 9518
rect 11150 9480 11152 9489
rect 11204 9480 11206 9489
rect 11256 9450 11284 14486
rect 11348 14482 11376 14758
rect 11440 14618 11468 15030
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 11348 13734 11376 14418
rect 11624 14006 11652 15846
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11612 14000 11664 14006
rect 11612 13942 11664 13948
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11428 12708 11480 12714
rect 11428 12650 11480 12656
rect 11440 12238 11468 12650
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11348 11937 11376 12038
rect 11334 11928 11390 11937
rect 11334 11863 11390 11872
rect 11532 11626 11560 12242
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11150 9415 11206 9424
rect 11244 9444 11296 9450
rect 11244 9386 11296 9392
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 11244 9104 11296 9110
rect 11244 9046 11296 9052
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10980 8430 11008 8774
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 10968 8424 11020 8430
rect 10966 8392 10968 8401
rect 11020 8392 11022 8401
rect 10966 8327 11022 8336
rect 11072 7886 11100 8502
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 11072 7290 11100 7822
rect 10980 7262 11100 7290
rect 10980 6866 11008 7262
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10874 6488 10930 6497
rect 10874 6423 10930 6432
rect 10888 5710 10916 6423
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 11072 5642 11100 7142
rect 11164 7002 11192 8298
rect 11256 8106 11284 9046
rect 11348 8294 11376 11494
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11256 8090 11376 8106
rect 11440 8090 11468 9318
rect 11532 8974 11560 9930
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11532 8090 11560 8434
rect 11256 8084 11388 8090
rect 11256 8078 11336 8084
rect 11336 8026 11388 8032
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11242 7712 11298 7721
rect 11242 7647 11298 7656
rect 11256 7478 11284 7647
rect 11348 7546 11376 7822
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11440 7342 11468 8026
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11242 6896 11298 6905
rect 11242 6831 11244 6840
rect 11296 6831 11298 6840
rect 11244 6802 11296 6808
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11164 6633 11192 6666
rect 11150 6624 11206 6633
rect 11150 6559 11206 6568
rect 11348 6458 11376 6734
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11440 6186 11468 6734
rect 11428 6180 11480 6186
rect 11428 6122 11480 6128
rect 11532 5710 11560 7890
rect 11624 7206 11652 13806
rect 11716 8430 11744 15438
rect 11796 14476 11848 14482
rect 11796 14418 11848 14424
rect 11808 9110 11836 14418
rect 11900 9994 11928 15914
rect 11992 14822 12020 16118
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12268 15706 12296 15846
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 12084 15026 12112 15302
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11900 9897 11928 9930
rect 11886 9888 11942 9897
rect 11886 9823 11942 9832
rect 11796 9104 11848 9110
rect 11796 9046 11848 9052
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11808 7410 11836 8774
rect 11900 8634 11928 8774
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11624 5914 11652 6054
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 11808 5234 11836 7346
rect 11900 7206 11928 8230
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11992 5370 12020 14758
rect 12084 14550 12112 14962
rect 12072 14544 12124 14550
rect 12072 14486 12124 14492
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 12084 12238 12112 14214
rect 12452 13988 12480 16050
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12452 13960 12572 13988
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12452 13530 12480 13806
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12544 13326 12572 13960
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12348 12912 12400 12918
rect 12346 12880 12348 12889
rect 12400 12880 12402 12889
rect 12452 12850 12480 12922
rect 12346 12815 12402 12824
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12346 12744 12402 12753
rect 12346 12679 12402 12688
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12176 12306 12204 12582
rect 12360 12424 12388 12679
rect 12544 12481 12572 12922
rect 12530 12472 12586 12481
rect 12360 12396 12480 12424
rect 12530 12407 12532 12416
rect 12452 12306 12480 12396
rect 12584 12407 12586 12416
rect 12532 12378 12584 12384
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12544 11898 12572 12174
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12070 11384 12126 11393
rect 12070 11319 12126 11328
rect 12084 11286 12112 11319
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 12268 11082 12296 11698
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 12084 10674 12112 11018
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12084 7002 12112 7346
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12176 6662 12204 10066
rect 12544 8974 12572 11290
rect 12636 10305 12664 13330
rect 12728 12434 12756 15642
rect 12820 15366 12848 16458
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12912 14346 12940 14894
rect 13096 14550 13124 16526
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13280 16114 13308 16390
rect 13648 16250 13676 17138
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 13636 16244 13688 16250
rect 13636 16186 13688 16192
rect 14016 16182 14044 16934
rect 15212 16658 15240 17206
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14096 16516 14148 16522
rect 14096 16458 14148 16464
rect 14004 16176 14056 16182
rect 14004 16118 14056 16124
rect 14108 16114 14136 16458
rect 14188 16448 14240 16454
rect 14188 16390 14240 16396
rect 14200 16114 14228 16390
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 14096 16108 14148 16114
rect 14096 16050 14148 16056
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 13280 15638 13308 16050
rect 14004 16040 14056 16046
rect 14200 15994 14228 16050
rect 14004 15982 14056 15988
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13360 14952 13412 14958
rect 13280 14912 13360 14940
rect 13176 14816 13228 14822
rect 13280 14804 13308 14912
rect 13360 14894 13412 14900
rect 13228 14776 13308 14804
rect 13360 14816 13412 14822
rect 13176 14758 13228 14764
rect 13360 14758 13412 14764
rect 13084 14544 13136 14550
rect 13084 14486 13136 14492
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 13004 13802 13032 14350
rect 12992 13796 13044 13802
rect 12992 13738 13044 13744
rect 13004 13530 13032 13738
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12820 12850 12848 13262
rect 12900 13184 12952 13190
rect 12952 13132 13032 13138
rect 12900 13126 13032 13132
rect 12912 13110 13032 13126
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12728 12406 12848 12434
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12728 10742 12756 12038
rect 12820 11354 12848 12406
rect 12912 11354 12940 12786
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12912 11150 12940 11290
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12806 10840 12862 10849
rect 12806 10775 12862 10784
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12820 10470 12848 10775
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12622 10296 12678 10305
rect 12622 10231 12624 10240
rect 12676 10231 12678 10240
rect 12624 10202 12676 10208
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12544 8498 12572 8910
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12636 8294 12664 8366
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10888 4214 10916 4558
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10692 4072 10744 4078
rect 10690 4040 10692 4049
rect 10784 4072 10836 4078
rect 10744 4040 10746 4049
rect 10784 4014 10836 4020
rect 10690 3975 10746 3984
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9508 3398 9536 3878
rect 9968 3670 9996 3878
rect 10980 3738 11008 4218
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9968 3466 9996 3606
rect 11164 3534 11192 4422
rect 12084 4214 12112 6326
rect 12268 5302 12296 6802
rect 12360 5914 12388 7346
rect 12530 7304 12586 7313
rect 12530 7239 12532 7248
rect 12584 7239 12586 7248
rect 12532 7210 12584 7216
rect 12544 6730 12572 7210
rect 12636 6730 12664 8230
rect 12532 6724 12584 6730
rect 12532 6666 12584 6672
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12360 5370 12388 5714
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 12072 4208 12124 4214
rect 12072 4150 12124 4156
rect 12084 3534 12112 4150
rect 12268 3602 12296 5238
rect 12360 3738 12388 5306
rect 12440 5228 12492 5234
rect 12544 5216 12572 6666
rect 12636 6458 12664 6666
rect 12728 6458 12756 10066
rect 12820 10062 12848 10406
rect 13004 10112 13032 13110
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 13096 12617 13124 12786
rect 13082 12608 13138 12617
rect 13082 12543 13138 12552
rect 13188 11286 13216 14758
rect 13372 14414 13400 14758
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13280 13530 13308 14010
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13280 12714 13308 13194
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13176 11280 13228 11286
rect 13176 11222 13228 11228
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 12912 10084 13032 10112
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12820 7834 12848 9590
rect 12912 8498 12940 10084
rect 12992 9988 13044 9994
rect 12992 9930 13044 9936
rect 13004 9722 13032 9930
rect 13096 9926 13124 11086
rect 13188 10606 13216 11086
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 13174 10160 13230 10169
rect 13174 10095 13230 10104
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13188 9738 13216 10095
rect 13280 9994 13308 12242
rect 13268 9988 13320 9994
rect 13268 9930 13320 9936
rect 12992 9716 13044 9722
rect 13188 9710 13308 9738
rect 12992 9658 13044 9664
rect 13280 9654 13308 9710
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13188 9178 13216 9522
rect 13372 9178 13400 14350
rect 13556 12434 13584 14962
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13832 13734 13860 14214
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13556 12406 13676 12434
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13464 10062 13492 11630
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 12992 8900 13044 8906
rect 12992 8842 13044 8848
rect 13004 8634 13032 8842
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 12912 7954 12940 8434
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 13004 8294 13032 8366
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12820 7806 12940 7834
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12820 7478 12848 7686
rect 12808 7472 12860 7478
rect 12808 7414 12860 7420
rect 12912 6866 12940 7806
rect 13096 7274 13124 8434
rect 13084 7268 13136 7274
rect 13084 7210 13136 7216
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12728 5794 12756 6394
rect 12912 6186 12940 6802
rect 13004 6390 13032 7142
rect 13188 6866 13216 9114
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13280 8430 13308 9046
rect 13464 8634 13492 9998
rect 13556 9110 13584 10610
rect 13648 10169 13676 12406
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13740 11558 13768 11698
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13740 11150 13768 11494
rect 13832 11354 13860 11494
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13634 10160 13690 10169
rect 13634 10095 13690 10104
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13648 9761 13676 9998
rect 13634 9752 13690 9761
rect 13634 9687 13690 9696
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13648 8974 13676 9687
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13556 8650 13584 8910
rect 13452 8628 13504 8634
rect 13556 8622 13676 8650
rect 13452 8570 13504 8576
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13452 8424 13504 8430
rect 13556 8401 13584 8434
rect 13452 8366 13504 8372
rect 13542 8392 13598 8401
rect 13464 8242 13492 8366
rect 13542 8327 13598 8336
rect 13464 8214 13584 8242
rect 13556 7886 13584 8214
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 12636 5766 12756 5794
rect 12636 5642 12664 5766
rect 12714 5672 12770 5681
rect 12624 5636 12676 5642
rect 12714 5607 12770 5616
rect 12624 5578 12676 5584
rect 12728 5234 12756 5607
rect 12492 5188 12572 5216
rect 12716 5228 12768 5234
rect 12440 5170 12492 5176
rect 12716 5170 12768 5176
rect 13280 5166 13308 7754
rect 13648 6730 13676 8622
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 13360 6656 13412 6662
rect 13412 6616 13492 6644
rect 13648 6633 13676 6666
rect 13360 6598 13412 6604
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13372 5642 13400 6258
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 13268 5160 13320 5166
rect 13268 5102 13320 5108
rect 13464 4622 13492 6616
rect 13634 6624 13690 6633
rect 13634 6559 13690 6568
rect 13740 6458 13768 10542
rect 13832 8294 13860 11018
rect 13924 10266 13952 13874
rect 14016 13462 14044 15982
rect 14108 15978 14228 15994
rect 14096 15972 14228 15978
rect 14148 15966 14228 15972
rect 14096 15914 14148 15920
rect 14200 15706 14228 15966
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14096 15428 14148 15434
rect 14096 15370 14148 15376
rect 14108 15026 14136 15370
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14108 14929 14136 14962
rect 14280 14952 14332 14958
rect 14094 14920 14150 14929
rect 14280 14894 14332 14900
rect 14094 14855 14150 14864
rect 14188 14340 14240 14346
rect 14188 14282 14240 14288
rect 14004 13456 14056 13462
rect 14004 13398 14056 13404
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 14108 12986 14136 13194
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14200 12866 14228 14282
rect 14292 13394 14320 14894
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14016 12838 14228 12866
rect 14016 11558 14044 12838
rect 14096 11620 14148 11626
rect 14096 11562 14148 11568
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 13924 9178 13952 9522
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 14016 8514 14044 11290
rect 14108 9926 14136 11562
rect 14292 10538 14320 13330
rect 14384 12986 14412 16526
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14936 16250 14964 16390
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 15212 16182 15240 16594
rect 15304 16590 15332 16934
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15580 16250 15608 16526
rect 16500 16425 16528 16934
rect 16776 16794 16804 17138
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16486 16416 16542 16425
rect 16486 16351 16542 16360
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 15108 15632 15160 15638
rect 15108 15574 15160 15580
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14476 12850 14504 13262
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14476 12434 14504 12786
rect 14384 12406 14504 12434
rect 14384 11898 14412 12406
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 14462 11928 14518 11937
rect 14372 11892 14424 11898
rect 14462 11863 14518 11872
rect 14372 11834 14424 11840
rect 14476 11830 14504 11863
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14280 10532 14332 10538
rect 14280 10474 14332 10480
rect 14278 10296 14334 10305
rect 14278 10231 14280 10240
rect 14332 10231 14334 10240
rect 14280 10202 14332 10208
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14108 9178 14136 9862
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14200 9042 14228 9454
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14188 8900 14240 8906
rect 14188 8842 14240 8848
rect 13924 8486 14044 8514
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13832 8090 13860 8230
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13924 6866 13952 8486
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13648 6322 13676 6394
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13648 6202 13676 6258
rect 13648 6186 13768 6202
rect 13648 6180 13780 6186
rect 13648 6174 13728 6180
rect 13728 6122 13780 6128
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13542 5808 13598 5817
rect 13542 5743 13598 5752
rect 13556 5710 13584 5743
rect 13648 5710 13676 6054
rect 13740 5914 13768 6122
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13740 4622 13768 4966
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13464 4162 13492 4558
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13372 4134 13492 4162
rect 13556 4146 13584 4422
rect 13636 4208 13688 4214
rect 13740 4196 13768 4558
rect 13688 4168 13768 4196
rect 13636 4150 13688 4156
rect 13832 4146 13860 6598
rect 14016 4622 14044 8298
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14108 5642 14136 6938
rect 14200 6662 14228 8842
rect 14384 8838 14412 11698
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14384 6730 14412 7278
rect 14372 6724 14424 6730
rect 14372 6666 14424 6672
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14476 5914 14504 11630
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14568 10062 14596 10406
rect 14660 10130 14688 12106
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14660 9602 14688 10066
rect 14568 9574 14688 9602
rect 14568 8974 14596 9574
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14660 9178 14688 9454
rect 14752 9382 14780 13874
rect 15120 13802 15148 15574
rect 15212 15570 15240 16118
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 15212 14482 15240 15506
rect 15304 15026 15332 15642
rect 15384 15088 15436 15094
rect 15488 15042 15516 15846
rect 16960 15745 16988 15846
rect 16946 15736 17002 15745
rect 16946 15671 17002 15680
rect 15752 15428 15804 15434
rect 15752 15370 15804 15376
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15436 15036 15516 15042
rect 15384 15030 15516 15036
rect 15292 15020 15344 15026
rect 15396 15014 15516 15030
rect 15292 14962 15344 14968
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15028 13326 15056 13670
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 15120 13240 15148 13738
rect 15212 13530 15240 14418
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15304 13258 15332 14962
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15200 13252 15252 13258
rect 15120 13212 15200 13240
rect 15200 13194 15252 13200
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 15108 12232 15160 12238
rect 15014 12200 15070 12209
rect 15108 12174 15160 12180
rect 15014 12135 15070 12144
rect 15028 11762 15056 12135
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 15120 11558 15148 12174
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 14936 11150 14964 11494
rect 15028 11354 15056 11494
rect 15212 11370 15240 13194
rect 15304 11694 15332 13194
rect 15396 12986 15424 13262
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15396 11898 15424 12174
rect 15488 12102 15516 15014
rect 15672 14498 15700 15302
rect 15764 15162 15792 15370
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 16960 15065 16988 15098
rect 16946 15056 17002 15065
rect 17052 15026 17080 15302
rect 16946 14991 17002 15000
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 15672 14470 15792 14498
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15672 14074 15700 14282
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15764 13870 15792 14470
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16776 13938 16804 14214
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15580 12306 15608 12854
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15672 12238 15700 13330
rect 15764 12918 15792 13806
rect 16948 13728 17000 13734
rect 16946 13696 16948 13705
rect 17000 13696 17002 13705
rect 16946 13631 17002 13640
rect 16946 13016 17002 13025
rect 16946 12951 16948 12960
rect 17000 12951 17002 12960
rect 16948 12922 17000 12928
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15476 12096 15528 12102
rect 15528 12044 15608 12050
rect 15476 12038 15608 12044
rect 15488 12022 15608 12038
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15120 11342 15240 11370
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 15120 11082 15148 11342
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14568 8498 14596 8910
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14660 8090 14688 9114
rect 14936 8974 14964 9318
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 15028 8090 15056 9862
rect 15212 9586 15240 11154
rect 15304 11150 15332 11630
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15304 8906 15332 10950
rect 15396 10810 15424 11086
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15580 10690 15608 12022
rect 15672 11218 15700 12174
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15396 10662 15608 10690
rect 15292 8900 15344 8906
rect 15292 8842 15344 8848
rect 15304 8634 15332 8842
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15212 8090 15240 8434
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14186 5808 14242 5817
rect 14186 5743 14188 5752
rect 14240 5743 14242 5752
rect 14188 5714 14240 5720
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 14200 4434 14228 5714
rect 14016 4406 14228 4434
rect 14016 4146 14044 4406
rect 14096 4208 14148 4214
rect 14096 4150 14148 4156
rect 13544 4140 13596 4146
rect 13372 4078 13400 4134
rect 13544 4082 13596 4088
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 14016 3942 14044 4082
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 12530 3768 12586 3777
rect 12348 3732 12400 3738
rect 12530 3703 12532 3712
rect 12348 3674 12400 3680
rect 12584 3703 12586 3712
rect 12532 3674 12584 3680
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 9956 3460 10008 3466
rect 9956 3402 10008 3408
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9968 3194 9996 3402
rect 11164 3194 11192 3470
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 9140 2650 9168 2994
rect 10244 2650 10272 2994
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 13924 2446 13952 2790
rect 14108 2446 14136 4150
rect 14752 4146 14780 7686
rect 15028 7002 15056 7822
rect 15016 6996 15068 7002
rect 15016 6938 15068 6944
rect 15304 6322 15332 8434
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 15304 5846 15332 6258
rect 15292 5840 15344 5846
rect 15212 5788 15292 5794
rect 15212 5782 15344 5788
rect 15212 5766 15332 5782
rect 15212 4486 15240 5766
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15304 5370 15332 5578
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15292 5228 15344 5234
rect 15396 5216 15424 10662
rect 15764 9042 15792 12174
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16592 11762 16620 12038
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16592 11098 16620 11698
rect 16592 11070 16712 11098
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16592 10674 16620 10950
rect 16684 10674 16712 11070
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16592 10062 16620 10610
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16132 9178 16160 9522
rect 16408 9466 16436 9998
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16500 9625 16528 9862
rect 16486 9616 16542 9625
rect 16486 9551 16542 9560
rect 16408 9438 16528 9466
rect 16500 9382 16528 9438
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 16500 9042 16528 9318
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15488 6458 15516 8570
rect 15764 8566 15792 8978
rect 15752 8560 15804 8566
rect 15752 8502 15804 8508
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 15764 7886 15792 8230
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15580 7546 15608 7754
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15672 6798 15700 7822
rect 16302 7576 16358 7585
rect 15936 7540 15988 7546
rect 16302 7511 16304 7520
rect 15936 7482 15988 7488
rect 16356 7511 16358 7520
rect 16304 7482 16356 7488
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15488 5778 15516 6394
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15344 5188 15424 5216
rect 15292 5170 15344 5176
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15212 4282 15240 4422
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 15304 4078 15332 5170
rect 15488 5098 15516 5714
rect 15672 5710 15700 6734
rect 15752 6724 15804 6730
rect 15752 6666 15804 6672
rect 15764 6458 15792 6666
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15476 5092 15528 5098
rect 15476 5034 15528 5040
rect 15488 4690 15516 5034
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 15672 4622 15700 5646
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 15396 4282 15424 4558
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14568 3466 14596 3878
rect 15672 3534 15700 4558
rect 15764 4146 15792 5170
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15764 3738 15792 4082
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15948 3534 15976 7482
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16132 6905 16160 7346
rect 16118 6896 16174 6905
rect 16118 6831 16174 6840
rect 16500 6662 16528 7346
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16500 6322 16528 6598
rect 16776 6474 16804 11698
rect 17222 11656 17278 11665
rect 17222 11591 17278 11600
rect 16946 10976 17002 10985
rect 16946 10911 17002 10920
rect 16960 10266 16988 10911
rect 17236 10810 17264 11591
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 16946 8936 17002 8945
rect 16946 8871 17002 8880
rect 16960 8634 16988 8871
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16592 6446 16804 6474
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16592 4826 16620 6446
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 16776 4826 16804 6258
rect 16868 5914 16896 8434
rect 17040 8424 17092 8430
rect 17040 8366 17092 8372
rect 16946 8256 17002 8265
rect 16946 8191 17002 8200
rect 16960 7546 16988 8191
rect 17052 8090 17080 8366
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17052 7410 17080 8026
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16946 6216 17002 6225
rect 16946 6151 16948 6160
rect 17000 6151 17002 6160
rect 16948 6122 17000 6128
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16868 5166 16896 5850
rect 16946 5536 17002 5545
rect 16946 5471 17002 5480
rect 16960 5370 16988 5471
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 16592 4162 16620 4762
rect 16500 4134 16620 4162
rect 16776 4146 16804 4762
rect 16764 4140 16816 4146
rect 16500 3738 16528 4134
rect 16764 4082 16816 4088
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15936 3528 15988 3534
rect 15988 3488 16068 3516
rect 15936 3470 15988 3476
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 14660 3126 14688 3470
rect 14648 3120 14700 3126
rect 14648 3062 14700 3068
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14292 2650 14320 2994
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14568 2446 14596 2790
rect 14660 2514 14688 2926
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 16040 2446 16068 3488
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5828 800 5856 2382
rect 9048 800 9076 2382
rect 10336 800 10364 2382
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13556 800 13584 2246
rect 5814 0 5870 800
rect 9034 0 9090 800
rect 10322 0 10378 800
rect 13542 0 13598 800
<< via2 >>
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 8574 17040 8630 17096
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 3238 11600 3294 11656
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4158 12824 4214 12880
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 3790 11736 3846 11792
rect 2778 10104 2834 10160
rect 3422 10512 3478 10568
rect 4526 12144 4582 12200
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4434 10668 4490 10704
rect 5630 13232 5686 13288
rect 5078 12688 5134 12744
rect 5630 12552 5686 12608
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4434 10648 4436 10668
rect 4436 10648 4488 10668
rect 4488 10648 4490 10668
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 846 6316 902 6352
rect 846 6296 848 6316
rect 848 6296 900 6316
rect 900 6296 902 6316
rect 1858 5480 1914 5536
rect 1306 4800 1362 4856
rect 5354 11892 5410 11928
rect 5354 11872 5356 11892
rect 5356 11872 5408 11892
rect 5408 11872 5410 11892
rect 5354 11464 5410 11520
rect 5262 11328 5318 11384
rect 5262 10920 5318 10976
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 5262 10512 5318 10568
rect 4986 10376 5042 10432
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4802 9152 4858 9208
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4986 8492 5042 8528
rect 4986 8472 4988 8492
rect 4988 8472 5040 8492
rect 5040 8472 5042 8492
rect 6642 14900 6644 14920
rect 6644 14900 6696 14920
rect 6696 14900 6698 14920
rect 6642 14864 6698 14900
rect 6550 14764 6552 14784
rect 6552 14764 6604 14784
rect 6604 14764 6606 14784
rect 5814 12688 5870 12744
rect 6090 12416 6146 12472
rect 5722 12280 5778 12336
rect 5630 10920 5686 10976
rect 5354 9424 5410 9480
rect 5722 10512 5778 10568
rect 5630 9696 5686 9752
rect 5354 8880 5410 8936
rect 5446 8472 5502 8528
rect 5354 8356 5410 8392
rect 5354 8336 5356 8356
rect 5356 8336 5408 8356
rect 5408 8336 5410 8356
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 5170 5228 5226 5264
rect 5170 5208 5172 5228
rect 5172 5208 5224 5228
rect 5224 5208 5226 5228
rect 5630 6704 5686 6760
rect 5906 11636 5908 11656
rect 5908 11636 5960 11656
rect 5960 11636 5962 11656
rect 5906 11600 5962 11636
rect 5722 5636 5778 5672
rect 5722 5616 5724 5636
rect 5724 5616 5776 5636
rect 5776 5616 5778 5636
rect 5814 5344 5870 5400
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 6274 13404 6276 13424
rect 6276 13404 6328 13424
rect 6328 13404 6330 13424
rect 6274 13368 6330 13404
rect 6550 14728 6606 14764
rect 7286 15544 7342 15600
rect 6274 11600 6330 11656
rect 6274 10124 6330 10160
rect 6274 10104 6276 10124
rect 6276 10104 6328 10124
rect 6328 10104 6330 10124
rect 6274 9968 6330 10024
rect 6182 9288 6238 9344
rect 6458 12044 6460 12064
rect 6460 12044 6512 12064
rect 6512 12044 6514 12064
rect 6458 12008 6514 12044
rect 6458 9560 6514 9616
rect 7194 13268 7196 13288
rect 7196 13268 7248 13288
rect 7248 13268 7250 13288
rect 7194 13232 7250 13268
rect 6918 12552 6974 12608
rect 7378 12688 7434 12744
rect 7286 12552 7342 12608
rect 7562 12552 7618 12608
rect 6734 12144 6790 12200
rect 7102 12180 7104 12200
rect 7104 12180 7156 12200
rect 7156 12180 7158 12200
rect 7102 12144 7158 12180
rect 6918 11192 6974 11248
rect 7102 11056 7158 11112
rect 6642 10240 6698 10296
rect 6642 9424 6698 9480
rect 6734 9152 6790 9208
rect 6550 9016 6606 9072
rect 6458 6296 6514 6352
rect 6182 5616 6238 5672
rect 6458 5616 6514 5672
rect 6274 5480 6330 5536
rect 6366 5344 6422 5400
rect 6550 5480 6606 5536
rect 6550 5344 6606 5400
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 1858 4140 1914 4176
rect 1858 4120 1860 4140
rect 1860 4120 1912 4140
rect 1912 4120 1914 4140
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 6734 5636 6790 5672
rect 6734 5616 6736 5636
rect 6736 5616 6788 5636
rect 6788 5616 6790 5636
rect 7010 10104 7066 10160
rect 7286 11736 7342 11792
rect 7286 11464 7342 11520
rect 7838 13812 7840 13832
rect 7840 13812 7892 13832
rect 7892 13812 7894 13832
rect 7838 13776 7894 13812
rect 8114 13912 8170 13968
rect 8022 13096 8078 13152
rect 7746 11600 7802 11656
rect 7562 11464 7618 11520
rect 7930 11464 7986 11520
rect 7654 10784 7710 10840
rect 7470 10648 7526 10704
rect 7010 9152 7066 9208
rect 7378 10376 7434 10432
rect 7562 10376 7618 10432
rect 7470 9696 7526 9752
rect 7286 9288 7342 9344
rect 7838 9696 7894 9752
rect 7746 9016 7802 9072
rect 7470 8472 7526 8528
rect 8114 11872 8170 11928
rect 8390 12416 8446 12472
rect 8022 10668 8078 10704
rect 8022 10648 8024 10668
rect 8024 10648 8076 10668
rect 8076 10648 8078 10668
rect 8114 10240 8170 10296
rect 9126 15544 9182 15600
rect 8942 14184 8998 14240
rect 8942 12824 8998 12880
rect 9034 12688 9090 12744
rect 8022 9560 8078 9616
rect 7654 8064 7710 8120
rect 7470 6432 7526 6488
rect 7286 5208 7342 5264
rect 8022 8064 8078 8120
rect 7838 6432 7894 6488
rect 7654 5344 7710 5400
rect 8022 5752 8078 5808
rect 8022 5344 8078 5400
rect 8298 9696 8354 9752
rect 8482 10004 8484 10024
rect 8484 10004 8536 10024
rect 8536 10004 8538 10024
rect 8482 9968 8538 10004
rect 8390 9152 8446 9208
rect 8850 10104 8906 10160
rect 8298 8880 8354 8936
rect 8206 8064 8262 8120
rect 8206 7928 8262 7984
rect 8390 6976 8446 7032
rect 8482 5228 8538 5264
rect 8482 5208 8484 5228
rect 8484 5208 8536 5228
rect 8536 5208 8538 5228
rect 9218 12300 9274 12336
rect 9218 12280 9220 12300
rect 9220 12280 9272 12300
rect 9272 12280 9274 12300
rect 8942 6724 8998 6760
rect 8942 6704 8944 6724
rect 8944 6704 8996 6724
rect 8996 6704 8998 6724
rect 8666 5364 8722 5400
rect 8666 5344 8668 5364
rect 8668 5344 8720 5364
rect 8720 5344 8722 5364
rect 9770 12280 9826 12336
rect 9310 7540 9366 7576
rect 9310 7520 9312 7540
rect 9312 7520 9364 7540
rect 9364 7520 9366 7540
rect 9310 6316 9366 6352
rect 9310 6296 9312 6316
rect 9312 6296 9364 6316
rect 9364 6296 9366 6316
rect 9310 5752 9366 5808
rect 9586 8744 9642 8800
rect 10138 15272 10194 15328
rect 10138 12144 10194 12200
rect 10230 10920 10286 10976
rect 10230 9444 10286 9480
rect 10230 9424 10232 9444
rect 10232 9424 10284 9444
rect 10284 9424 10286 9444
rect 10966 12552 11022 12608
rect 10414 8336 10470 8392
rect 9770 6976 9826 7032
rect 10138 7248 10194 7304
rect 10322 7248 10378 7304
rect 10230 6840 10286 6896
rect 11150 12180 11152 12200
rect 11152 12180 11204 12200
rect 11204 12180 11206 12200
rect 10414 5752 10470 5808
rect 11150 12144 11206 12180
rect 10966 9696 11022 9752
rect 11150 9460 11152 9480
rect 11152 9460 11204 9480
rect 11204 9460 11206 9480
rect 11150 9424 11206 9460
rect 11334 11872 11390 11928
rect 10966 8372 10968 8392
rect 10968 8372 11020 8392
rect 11020 8372 11022 8392
rect 10966 8336 11022 8372
rect 10874 6432 10930 6488
rect 11242 7656 11298 7712
rect 11242 6860 11298 6896
rect 11242 6840 11244 6860
rect 11244 6840 11296 6860
rect 11296 6840 11298 6860
rect 11150 6568 11206 6624
rect 11886 9832 11942 9888
rect 12346 12860 12348 12880
rect 12348 12860 12400 12880
rect 12400 12860 12402 12880
rect 12346 12824 12402 12860
rect 12346 12688 12402 12744
rect 12530 12436 12586 12472
rect 12530 12416 12532 12436
rect 12532 12416 12584 12436
rect 12584 12416 12586 12436
rect 12070 11328 12126 11384
rect 12806 10784 12862 10840
rect 12622 10260 12678 10296
rect 12622 10240 12624 10260
rect 12624 10240 12676 10260
rect 12676 10240 12678 10260
rect 10690 4020 10692 4040
rect 10692 4020 10744 4040
rect 10744 4020 10746 4040
rect 10690 3984 10746 4020
rect 12530 7268 12586 7304
rect 12530 7248 12532 7268
rect 12532 7248 12584 7268
rect 12584 7248 12586 7268
rect 13082 12552 13138 12608
rect 13174 10104 13230 10160
rect 13634 10104 13690 10160
rect 13634 9696 13690 9752
rect 13542 8336 13598 8392
rect 12714 5616 12770 5672
rect 13634 6568 13690 6624
rect 14094 14864 14150 14920
rect 16486 16360 16542 16416
rect 14462 11872 14518 11928
rect 14278 10260 14334 10296
rect 14278 10240 14280 10260
rect 14280 10240 14332 10260
rect 14332 10240 14334 10260
rect 13542 5752 13598 5808
rect 16946 15680 17002 15736
rect 15014 12144 15070 12200
rect 16946 15000 17002 15056
rect 16946 13676 16948 13696
rect 16948 13676 17000 13696
rect 17000 13676 17002 13696
rect 16946 13640 17002 13676
rect 16946 12980 17002 13016
rect 16946 12960 16948 12980
rect 16948 12960 17000 12980
rect 17000 12960 17002 12980
rect 14186 5772 14242 5808
rect 14186 5752 14188 5772
rect 14188 5752 14240 5772
rect 14240 5752 14242 5772
rect 12530 3732 12586 3768
rect 12530 3712 12532 3732
rect 12532 3712 12584 3732
rect 12584 3712 12586 3732
rect 16486 9560 16542 9616
rect 16302 7540 16358 7576
rect 16302 7520 16304 7540
rect 16304 7520 16356 7540
rect 16356 7520 16358 7540
rect 16118 6840 16174 6896
rect 17222 11600 17278 11656
rect 16946 10920 17002 10976
rect 16946 8880 17002 8936
rect 16946 8200 17002 8256
rect 16946 6180 17002 6216
rect 16946 6160 16948 6180
rect 16948 6160 17000 6180
rect 17000 6160 17002 6180
rect 16946 5480 17002 5536
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 0 17098 800 17128
rect 8569 17098 8635 17101
rect 0 17096 8635 17098
rect 0 17040 8574 17096
rect 8630 17040 8635 17096
rect 0 17038 8635 17040
rect 0 17008 800 17038
rect 8569 17035 8635 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 16481 16418 16547 16421
rect 17714 16418 18514 16448
rect 16481 16416 18514 16418
rect 16481 16360 16486 16416
rect 16542 16360 18514 16416
rect 16481 16358 18514 16360
rect 16481 16355 16547 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 17714 16328 18514 16358
rect 4870 16287 5186 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 16941 15738 17007 15741
rect 17714 15738 18514 15768
rect 16941 15736 18514 15738
rect 16941 15680 16946 15736
rect 17002 15680 18514 15736
rect 16941 15678 18514 15680
rect 16941 15675 17007 15678
rect 17714 15648 18514 15678
rect 7281 15602 7347 15605
rect 9121 15602 9187 15605
rect 7281 15600 9187 15602
rect 7281 15544 7286 15600
rect 7342 15544 9126 15600
rect 9182 15544 9187 15600
rect 7281 15542 9187 15544
rect 7281 15539 7347 15542
rect 9121 15539 9187 15542
rect 9622 15268 9628 15332
rect 9692 15330 9698 15332
rect 10133 15330 10199 15333
rect 9692 15328 10199 15330
rect 9692 15272 10138 15328
rect 10194 15272 10199 15328
rect 9692 15270 10199 15272
rect 9692 15268 9698 15270
rect 10133 15267 10199 15270
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 16941 15058 17007 15061
rect 17714 15058 18514 15088
rect 16941 15056 18514 15058
rect 16941 15000 16946 15056
rect 17002 15000 18514 15056
rect 16941 14998 18514 15000
rect 16941 14995 17007 14998
rect 17714 14968 18514 14998
rect 6637 14924 6703 14925
rect 6637 14922 6684 14924
rect 6592 14920 6684 14922
rect 6592 14864 6642 14920
rect 6592 14862 6684 14864
rect 6637 14860 6684 14862
rect 6748 14860 6754 14924
rect 14089 14922 14155 14925
rect 14222 14922 14228 14924
rect 14089 14920 14228 14922
rect 14089 14864 14094 14920
rect 14150 14864 14228 14920
rect 14089 14862 14228 14864
rect 6637 14859 6703 14860
rect 14089 14859 14155 14862
rect 14222 14860 14228 14862
rect 14292 14860 14298 14924
rect 6310 14724 6316 14788
rect 6380 14786 6386 14788
rect 6545 14786 6611 14789
rect 6380 14784 6611 14786
rect 6380 14728 6550 14784
rect 6606 14728 6611 14784
rect 6380 14726 6611 14728
rect 6380 14724 6386 14726
rect 6545 14723 6611 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 8937 14244 9003 14245
rect 8886 14180 8892 14244
rect 8956 14242 9003 14244
rect 8956 14240 9048 14242
rect 8998 14184 9048 14240
rect 8956 14182 9048 14184
rect 8956 14180 9003 14182
rect 8937 14179 9003 14180
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 8109 13970 8175 13973
rect 9070 13970 9076 13972
rect 8109 13968 9076 13970
rect 8109 13912 8114 13968
rect 8170 13912 9076 13968
rect 8109 13910 9076 13912
rect 8109 13907 8175 13910
rect 9070 13908 9076 13910
rect 9140 13908 9146 13972
rect 7833 13834 7899 13837
rect 9254 13834 9260 13836
rect 7833 13832 9260 13834
rect 7833 13776 7838 13832
rect 7894 13776 9260 13832
rect 7833 13774 9260 13776
rect 7833 13771 7899 13774
rect 9254 13772 9260 13774
rect 9324 13772 9330 13836
rect 16941 13698 17007 13701
rect 17714 13698 18514 13728
rect 16941 13696 18514 13698
rect 16941 13640 16946 13696
rect 17002 13640 18514 13696
rect 16941 13638 18514 13640
rect 16941 13635 17007 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 17714 13608 18514 13638
rect 4210 13567 4526 13568
rect 6269 13426 6335 13429
rect 6494 13426 6500 13428
rect 6269 13424 6500 13426
rect 6269 13368 6274 13424
rect 6330 13368 6500 13424
rect 6269 13366 6500 13368
rect 6269 13363 6335 13366
rect 6494 13364 6500 13366
rect 6564 13364 6570 13428
rect 5625 13290 5691 13293
rect 7189 13290 7255 13293
rect 5625 13288 7255 13290
rect 5625 13232 5630 13288
rect 5686 13232 7194 13288
rect 7250 13232 7255 13288
rect 5625 13230 7255 13232
rect 5625 13227 5691 13230
rect 7189 13227 7255 13230
rect 8017 13154 8083 13157
rect 8150 13154 8156 13156
rect 8017 13152 8156 13154
rect 8017 13096 8022 13152
rect 8078 13096 8156 13152
rect 8017 13094 8156 13096
rect 8017 13091 8083 13094
rect 8150 13092 8156 13094
rect 8220 13092 8226 13156
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 16941 13018 17007 13021
rect 17714 13018 18514 13048
rect 16941 13016 18514 13018
rect 16941 12960 16946 13016
rect 17002 12960 18514 13016
rect 16941 12958 18514 12960
rect 16941 12955 17007 12958
rect 17714 12928 18514 12958
rect 4153 12882 4219 12885
rect 8937 12882 9003 12885
rect 4153 12880 9003 12882
rect 4153 12824 4158 12880
rect 4214 12824 8942 12880
rect 8998 12824 9003 12880
rect 4153 12822 9003 12824
rect 4153 12819 4219 12822
rect 8937 12819 9003 12822
rect 12198 12820 12204 12884
rect 12268 12882 12274 12884
rect 12341 12882 12407 12885
rect 12268 12880 12407 12882
rect 12268 12824 12346 12880
rect 12402 12824 12407 12880
rect 12268 12822 12407 12824
rect 12268 12820 12274 12822
rect 12341 12819 12407 12822
rect 5073 12746 5139 12749
rect 5809 12746 5875 12749
rect 7373 12746 7439 12749
rect 5073 12744 7439 12746
rect 5073 12688 5078 12744
rect 5134 12688 5814 12744
rect 5870 12688 7378 12744
rect 7434 12688 7439 12744
rect 5073 12686 7439 12688
rect 5073 12683 5139 12686
rect 5809 12683 5875 12686
rect 7373 12683 7439 12686
rect 9029 12746 9095 12749
rect 12341 12746 12407 12749
rect 9029 12744 12407 12746
rect 9029 12688 9034 12744
rect 9090 12688 12346 12744
rect 12402 12688 12407 12744
rect 9029 12686 12407 12688
rect 9029 12683 9095 12686
rect 12341 12683 12407 12686
rect 5625 12610 5691 12613
rect 6913 12610 6979 12613
rect 5625 12608 6979 12610
rect 5625 12552 5630 12608
rect 5686 12552 6918 12608
rect 6974 12552 6979 12608
rect 5625 12550 6979 12552
rect 5625 12547 5691 12550
rect 6913 12547 6979 12550
rect 7281 12610 7347 12613
rect 7557 12610 7623 12613
rect 7281 12608 7623 12610
rect 7281 12552 7286 12608
rect 7342 12552 7562 12608
rect 7618 12552 7623 12608
rect 7281 12550 7623 12552
rect 7281 12547 7347 12550
rect 7557 12547 7623 12550
rect 10961 12610 11027 12613
rect 13077 12610 13143 12613
rect 10961 12608 13143 12610
rect 10961 12552 10966 12608
rect 11022 12552 13082 12608
rect 13138 12552 13143 12608
rect 10961 12550 13143 12552
rect 10961 12547 11027 12550
rect 13077 12547 13143 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 6085 12474 6151 12477
rect 8385 12474 8451 12477
rect 12525 12474 12591 12477
rect 6085 12472 12591 12474
rect 6085 12416 6090 12472
rect 6146 12416 8390 12472
rect 8446 12416 12530 12472
rect 12586 12416 12591 12472
rect 6085 12414 12591 12416
rect 6085 12411 6151 12414
rect 8385 12411 8451 12414
rect 12525 12411 12591 12414
rect 5717 12338 5783 12341
rect 9213 12338 9279 12341
rect 5717 12336 9279 12338
rect 5717 12280 5722 12336
rect 5778 12280 9218 12336
rect 9274 12280 9279 12336
rect 5717 12278 9279 12280
rect 5717 12275 5783 12278
rect 9213 12275 9279 12278
rect 9765 12338 9831 12341
rect 9765 12336 9874 12338
rect 9765 12280 9770 12336
rect 9826 12280 9874 12336
rect 9765 12275 9874 12280
rect 4521 12202 4587 12205
rect 6494 12202 6500 12204
rect 4521 12200 6500 12202
rect 4521 12144 4526 12200
rect 4582 12144 6500 12200
rect 4521 12142 6500 12144
rect 4521 12139 4587 12142
rect 6494 12140 6500 12142
rect 6564 12140 6570 12204
rect 6729 12202 6795 12205
rect 7097 12202 7163 12205
rect 7230 12202 7236 12204
rect 6729 12200 7236 12202
rect 6729 12144 6734 12200
rect 6790 12144 7102 12200
rect 7158 12144 7236 12200
rect 6729 12142 7236 12144
rect 6729 12139 6795 12142
rect 7097 12139 7163 12142
rect 7230 12140 7236 12142
rect 7300 12140 7306 12204
rect 9814 12202 9874 12275
rect 10133 12202 10199 12205
rect 11145 12202 11211 12205
rect 15009 12202 15075 12205
rect 9814 12200 11211 12202
rect 9814 12144 10138 12200
rect 10194 12144 11150 12200
rect 11206 12144 11211 12200
rect 9814 12142 11211 12144
rect 10133 12139 10199 12142
rect 11145 12139 11211 12142
rect 12390 12200 15075 12202
rect 12390 12144 15014 12200
rect 15070 12144 15075 12200
rect 12390 12142 15075 12144
rect 6453 12066 6519 12069
rect 12390 12066 12450 12142
rect 15009 12139 15075 12142
rect 6453 12064 12450 12066
rect 6453 12008 6458 12064
rect 6514 12008 12450 12064
rect 6453 12006 12450 12008
rect 6453 12003 6519 12006
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 5349 11930 5415 11933
rect 8109 11930 8175 11933
rect 5349 11928 8175 11930
rect 5349 11872 5354 11928
rect 5410 11872 8114 11928
rect 8170 11872 8175 11928
rect 5349 11870 8175 11872
rect 5349 11867 5415 11870
rect 8109 11867 8175 11870
rect 11329 11930 11395 11933
rect 14457 11930 14523 11933
rect 11329 11928 14523 11930
rect 11329 11872 11334 11928
rect 11390 11872 14462 11928
rect 14518 11872 14523 11928
rect 11329 11870 14523 11872
rect 11329 11867 11395 11870
rect 14457 11867 14523 11870
rect 3785 11794 3851 11797
rect 7281 11794 7347 11797
rect 3785 11792 7347 11794
rect 3785 11736 3790 11792
rect 3846 11736 7286 11792
rect 7342 11736 7347 11792
rect 3785 11734 7347 11736
rect 3785 11731 3851 11734
rect 7281 11731 7347 11734
rect 3233 11658 3299 11661
rect 5901 11658 5967 11661
rect 3233 11656 5967 11658
rect 3233 11600 3238 11656
rect 3294 11600 5906 11656
rect 5962 11600 5967 11656
rect 3233 11598 5967 11600
rect 3233 11595 3299 11598
rect 5901 11595 5967 11598
rect 6269 11658 6335 11661
rect 7741 11658 7807 11661
rect 6269 11656 7807 11658
rect 6269 11600 6274 11656
rect 6330 11600 7746 11656
rect 7802 11600 7807 11656
rect 6269 11598 7807 11600
rect 6269 11595 6335 11598
rect 7741 11595 7807 11598
rect 17217 11658 17283 11661
rect 17714 11658 18514 11688
rect 17217 11656 18514 11658
rect 17217 11600 17222 11656
rect 17278 11600 18514 11656
rect 17217 11598 18514 11600
rect 17217 11595 17283 11598
rect 17714 11568 18514 11598
rect 5349 11522 5415 11525
rect 7281 11522 7347 11525
rect 5349 11520 7347 11522
rect 5349 11464 5354 11520
rect 5410 11464 7286 11520
rect 7342 11464 7347 11520
rect 5349 11462 7347 11464
rect 5349 11459 5415 11462
rect 7281 11459 7347 11462
rect 7557 11522 7623 11525
rect 7925 11522 7991 11525
rect 7557 11520 7991 11522
rect 7557 11464 7562 11520
rect 7618 11464 7930 11520
rect 7986 11464 7991 11520
rect 7557 11462 7991 11464
rect 7557 11459 7623 11462
rect 7925 11459 7991 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 5257 11386 5323 11389
rect 10910 11386 10916 11388
rect 5257 11384 10916 11386
rect 5257 11328 5262 11384
rect 5318 11328 10916 11384
rect 5257 11326 10916 11328
rect 5257 11323 5323 11326
rect 10910 11324 10916 11326
rect 10980 11386 10986 11388
rect 12065 11386 12131 11389
rect 10980 11384 12131 11386
rect 10980 11328 12070 11384
rect 12126 11328 12131 11384
rect 10980 11326 12131 11328
rect 10980 11324 10986 11326
rect 12065 11323 12131 11326
rect 6913 11250 6979 11253
rect 6913 11248 7850 11250
rect 6913 11192 6918 11248
rect 6974 11192 7850 11248
rect 6913 11190 7850 11192
rect 6913 11187 6979 11190
rect 6862 11052 6868 11116
rect 6932 11114 6938 11116
rect 7097 11114 7163 11117
rect 6932 11112 7163 11114
rect 6932 11056 7102 11112
rect 7158 11056 7163 11112
rect 6932 11054 7163 11056
rect 7790 11114 7850 11190
rect 9070 11114 9076 11116
rect 7790 11054 9076 11114
rect 6932 11052 6938 11054
rect 7097 11051 7163 11054
rect 9070 11052 9076 11054
rect 9140 11052 9146 11116
rect 5257 10978 5323 10981
rect 5625 10978 5691 10981
rect 10225 10978 10291 10981
rect 10358 10978 10364 10980
rect 5257 10976 5691 10978
rect 5257 10920 5262 10976
rect 5318 10920 5630 10976
rect 5686 10920 5691 10976
rect 5257 10918 5691 10920
rect 5257 10915 5323 10918
rect 5625 10915 5691 10918
rect 7238 10976 10364 10978
rect 7238 10920 10230 10976
rect 10286 10920 10364 10976
rect 7238 10918 10364 10920
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 4429 10706 4495 10709
rect 7238 10706 7298 10918
rect 10225 10915 10291 10918
rect 10358 10916 10364 10918
rect 10428 10916 10434 10980
rect 16941 10978 17007 10981
rect 17714 10978 18514 11008
rect 16941 10976 18514 10978
rect 16941 10920 16946 10976
rect 17002 10920 18514 10976
rect 16941 10918 18514 10920
rect 16941 10915 17007 10918
rect 17714 10888 18514 10918
rect 7649 10842 7715 10845
rect 12801 10842 12867 10845
rect 7649 10840 12867 10842
rect 7649 10784 7654 10840
rect 7710 10784 12806 10840
rect 12862 10784 12867 10840
rect 7649 10782 12867 10784
rect 7649 10779 7715 10782
rect 12801 10779 12867 10782
rect 4429 10704 7298 10706
rect 4429 10648 4434 10704
rect 4490 10648 7298 10704
rect 4429 10646 7298 10648
rect 7465 10706 7531 10709
rect 8017 10706 8083 10709
rect 7465 10704 8083 10706
rect 7465 10648 7470 10704
rect 7526 10648 8022 10704
rect 8078 10648 8083 10704
rect 7465 10646 8083 10648
rect 4429 10643 4495 10646
rect 7465 10643 7531 10646
rect 8017 10643 8083 10646
rect 3417 10570 3483 10573
rect 5257 10570 5323 10573
rect 3417 10568 5323 10570
rect 3417 10512 3422 10568
rect 3478 10512 5262 10568
rect 5318 10512 5323 10568
rect 3417 10510 5323 10512
rect 3417 10507 3483 10510
rect 5257 10507 5323 10510
rect 5717 10570 5783 10573
rect 5717 10568 7620 10570
rect 5717 10512 5722 10568
rect 5778 10512 7620 10568
rect 5717 10510 7620 10512
rect 5717 10507 5783 10510
rect 7560 10437 7620 10510
rect 4981 10434 5047 10437
rect 4981 10432 6884 10434
rect 4981 10376 4986 10432
rect 5042 10376 6884 10432
rect 4981 10374 6884 10376
rect 4981 10371 5047 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 6310 10236 6316 10300
rect 6380 10298 6386 10300
rect 6637 10298 6703 10301
rect 6380 10296 6703 10298
rect 6380 10240 6642 10296
rect 6698 10240 6703 10296
rect 6380 10238 6703 10240
rect 6824 10298 6884 10374
rect 7230 10372 7236 10436
rect 7300 10434 7306 10436
rect 7373 10434 7439 10437
rect 7300 10432 7439 10434
rect 7300 10376 7378 10432
rect 7434 10376 7439 10432
rect 7300 10374 7439 10376
rect 7300 10372 7306 10374
rect 7373 10371 7439 10374
rect 7557 10432 7623 10437
rect 7557 10376 7562 10432
rect 7618 10376 7623 10432
rect 7557 10371 7623 10376
rect 8109 10298 8175 10301
rect 6824 10296 8175 10298
rect 6824 10240 8114 10296
rect 8170 10240 8175 10296
rect 6824 10238 8175 10240
rect 6380 10236 6386 10238
rect 6637 10235 6703 10238
rect 8109 10235 8175 10238
rect 12617 10298 12683 10301
rect 14273 10298 14339 10301
rect 12617 10296 14339 10298
rect 12617 10240 12622 10296
rect 12678 10240 14278 10296
rect 14334 10240 14339 10296
rect 12617 10238 14339 10240
rect 12617 10235 12683 10238
rect 14273 10235 14339 10238
rect 2773 10162 2839 10165
rect 6269 10162 6335 10165
rect 2773 10160 6335 10162
rect 2773 10104 2778 10160
rect 2834 10104 6274 10160
rect 6330 10104 6335 10160
rect 2773 10102 6335 10104
rect 2773 10099 2839 10102
rect 6269 10099 6335 10102
rect 7005 10162 7071 10165
rect 8845 10162 8911 10165
rect 7005 10160 8911 10162
rect 7005 10104 7010 10160
rect 7066 10104 8850 10160
rect 8906 10104 8911 10160
rect 7005 10102 8911 10104
rect 7005 10099 7071 10102
rect 8845 10099 8911 10102
rect 13169 10162 13235 10165
rect 13629 10162 13695 10165
rect 13169 10160 13695 10162
rect 13169 10104 13174 10160
rect 13230 10104 13634 10160
rect 13690 10104 13695 10160
rect 13169 10102 13695 10104
rect 13169 10099 13235 10102
rect 13629 10099 13695 10102
rect 6269 10026 6335 10029
rect 8477 10026 8543 10029
rect 6269 10024 8543 10026
rect 6269 9968 6274 10024
rect 6330 9968 8482 10024
rect 8538 9968 8543 10024
rect 6269 9966 8543 9968
rect 6269 9963 6335 9966
rect 8477 9963 8543 9966
rect 11881 9892 11947 9893
rect 11830 9828 11836 9892
rect 11900 9890 11947 9892
rect 11900 9888 11992 9890
rect 11942 9832 11992 9888
rect 11900 9830 11992 9832
rect 11900 9828 11947 9830
rect 11881 9827 11947 9828
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 5625 9754 5691 9757
rect 7465 9754 7531 9757
rect 5625 9752 7531 9754
rect 5625 9696 5630 9752
rect 5686 9696 7470 9752
rect 7526 9696 7531 9752
rect 5625 9694 7531 9696
rect 5625 9691 5691 9694
rect 7465 9691 7531 9694
rect 7833 9754 7899 9757
rect 8293 9754 8359 9757
rect 7833 9752 8359 9754
rect 7833 9696 7838 9752
rect 7894 9696 8298 9752
rect 8354 9696 8359 9752
rect 7833 9694 8359 9696
rect 7833 9691 7899 9694
rect 8293 9691 8359 9694
rect 10961 9754 11027 9757
rect 13629 9754 13695 9757
rect 10961 9752 13695 9754
rect 10961 9696 10966 9752
rect 11022 9696 13634 9752
rect 13690 9696 13695 9752
rect 10961 9694 13695 9696
rect 10961 9691 11027 9694
rect 13629 9691 13695 9694
rect 6453 9618 6519 9621
rect 8017 9618 8083 9621
rect 6453 9616 8083 9618
rect 6453 9560 6458 9616
rect 6514 9560 8022 9616
rect 8078 9560 8083 9616
rect 6453 9558 8083 9560
rect 6453 9555 6519 9558
rect 8017 9555 8083 9558
rect 16481 9618 16547 9621
rect 17714 9618 18514 9648
rect 16481 9616 18514 9618
rect 16481 9560 16486 9616
rect 16542 9560 18514 9616
rect 16481 9558 18514 9560
rect 16481 9555 16547 9558
rect 17714 9528 18514 9558
rect 5349 9482 5415 9485
rect 6637 9482 6703 9485
rect 5349 9480 6703 9482
rect 5349 9424 5354 9480
rect 5410 9424 6642 9480
rect 6698 9424 6703 9480
rect 5349 9422 6703 9424
rect 5349 9419 5415 9422
rect 6637 9419 6703 9422
rect 10225 9482 10291 9485
rect 11145 9482 11211 9485
rect 10225 9480 11211 9482
rect 10225 9424 10230 9480
rect 10286 9424 11150 9480
rect 11206 9424 11211 9480
rect 10225 9422 11211 9424
rect 10225 9419 10291 9422
rect 11145 9419 11211 9422
rect 6177 9346 6243 9349
rect 7281 9346 7347 9349
rect 6177 9344 7347 9346
rect 6177 9288 6182 9344
rect 6238 9288 7286 9344
rect 7342 9288 7347 9344
rect 6177 9286 7347 9288
rect 6177 9283 6243 9286
rect 7281 9283 7347 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4797 9210 4863 9213
rect 6729 9210 6795 9213
rect 4797 9208 6795 9210
rect 4797 9152 4802 9208
rect 4858 9152 6734 9208
rect 6790 9152 6795 9208
rect 4797 9150 6795 9152
rect 4797 9147 4863 9150
rect 6729 9147 6795 9150
rect 7005 9210 7071 9213
rect 8385 9210 8451 9213
rect 7005 9208 8451 9210
rect 7005 9152 7010 9208
rect 7066 9152 8390 9208
rect 8446 9152 8451 9208
rect 7005 9150 8451 9152
rect 7005 9147 7071 9150
rect 8385 9147 8451 9150
rect 6545 9074 6611 9077
rect 7741 9074 7807 9077
rect 6545 9072 7807 9074
rect 6545 9016 6550 9072
rect 6606 9016 7746 9072
rect 7802 9016 7807 9072
rect 6545 9014 7807 9016
rect 6545 9011 6611 9014
rect 7741 9011 7807 9014
rect 5349 8938 5415 8941
rect 8293 8938 8359 8941
rect 5349 8936 8359 8938
rect 5349 8880 5354 8936
rect 5410 8880 8298 8936
rect 8354 8880 8359 8936
rect 5349 8878 8359 8880
rect 5349 8875 5415 8878
rect 8293 8875 8359 8878
rect 16941 8938 17007 8941
rect 17714 8938 18514 8968
rect 16941 8936 18514 8938
rect 16941 8880 16946 8936
rect 17002 8880 18514 8936
rect 16941 8878 18514 8880
rect 16941 8875 17007 8878
rect 17714 8848 18514 8878
rect 6494 8740 6500 8804
rect 6564 8802 6570 8804
rect 9581 8802 9647 8805
rect 6564 8800 9647 8802
rect 6564 8744 9586 8800
rect 9642 8744 9647 8800
rect 6564 8742 9647 8744
rect 6564 8740 6570 8742
rect 9581 8739 9647 8742
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 4981 8530 5047 8533
rect 5441 8530 5507 8533
rect 7465 8530 7531 8533
rect 4981 8528 7531 8530
rect 4981 8472 4986 8528
rect 5042 8472 5446 8528
rect 5502 8472 7470 8528
rect 7526 8472 7531 8528
rect 4981 8470 7531 8472
rect 4981 8467 5047 8470
rect 5441 8467 5507 8470
rect 7465 8467 7531 8470
rect 10550 8470 12450 8530
rect 5349 8394 5415 8397
rect 10409 8394 10475 8397
rect 10550 8394 10610 8470
rect 5349 8392 10610 8394
rect 5349 8336 5354 8392
rect 5410 8336 10414 8392
rect 10470 8336 10610 8392
rect 5349 8334 10610 8336
rect 5349 8331 5415 8334
rect 10409 8331 10475 8334
rect 10726 8332 10732 8396
rect 10796 8394 10802 8396
rect 10961 8394 11027 8397
rect 10796 8392 11027 8394
rect 10796 8336 10966 8392
rect 11022 8336 11027 8392
rect 10796 8334 11027 8336
rect 12390 8394 12450 8470
rect 13537 8394 13603 8397
rect 12390 8392 13603 8394
rect 12390 8336 13542 8392
rect 13598 8336 13603 8392
rect 12390 8334 13603 8336
rect 10796 8332 10802 8334
rect 10961 8331 11027 8334
rect 13537 8331 13603 8334
rect 16941 8258 17007 8261
rect 17714 8258 18514 8288
rect 16941 8256 18514 8258
rect 16941 8200 16946 8256
rect 17002 8200 18514 8256
rect 16941 8198 18514 8200
rect 16941 8195 17007 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 17714 8168 18514 8198
rect 4210 8127 4526 8128
rect 7649 8122 7715 8125
rect 8017 8122 8083 8125
rect 8201 8122 8267 8125
rect 7649 8120 8267 8122
rect 7649 8064 7654 8120
rect 7710 8064 8022 8120
rect 8078 8064 8206 8120
rect 8262 8064 8267 8120
rect 7649 8062 8267 8064
rect 7649 8059 7715 8062
rect 8017 8059 8083 8062
rect 8201 8059 8267 8062
rect 8201 7988 8267 7989
rect 8150 7924 8156 7988
rect 8220 7986 8267 7988
rect 8220 7984 8312 7986
rect 8262 7928 8312 7984
rect 8220 7926 8312 7928
rect 8220 7924 8267 7926
rect 8201 7923 8267 7924
rect 9254 7652 9260 7716
rect 9324 7714 9330 7716
rect 11237 7714 11303 7717
rect 9324 7712 11303 7714
rect 9324 7656 11242 7712
rect 11298 7656 11303 7712
rect 9324 7654 11303 7656
rect 9324 7652 9330 7654
rect 11237 7651 11303 7654
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 9305 7578 9371 7581
rect 9622 7578 9628 7580
rect 9305 7576 9628 7578
rect 9305 7520 9310 7576
rect 9366 7520 9628 7576
rect 9305 7518 9628 7520
rect 9305 7515 9371 7518
rect 9622 7516 9628 7518
rect 9692 7516 9698 7580
rect 16297 7578 16363 7581
rect 17714 7578 18514 7608
rect 16297 7576 18514 7578
rect 16297 7520 16302 7576
rect 16358 7520 18514 7576
rect 16297 7518 18514 7520
rect 16297 7515 16363 7518
rect 17714 7488 18514 7518
rect 10133 7306 10199 7309
rect 10317 7306 10383 7309
rect 12525 7306 12591 7309
rect 10133 7304 12591 7306
rect 10133 7248 10138 7304
rect 10194 7248 10322 7304
rect 10378 7248 12530 7304
rect 12586 7248 12591 7304
rect 10133 7246 12591 7248
rect 10133 7243 10199 7246
rect 10317 7243 10383 7246
rect 12525 7243 12591 7246
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 8385 7034 8451 7037
rect 8702 7034 8708 7036
rect 8385 7032 8708 7034
rect 8385 6976 8390 7032
rect 8446 6976 8708 7032
rect 8385 6974 8708 6976
rect 8385 6971 8451 6974
rect 8702 6972 8708 6974
rect 8772 7034 8778 7036
rect 9765 7034 9831 7037
rect 8772 7032 9831 7034
rect 8772 6976 9770 7032
rect 9826 6976 9831 7032
rect 8772 6974 9831 6976
rect 8772 6972 8778 6974
rect 9765 6971 9831 6974
rect 10225 6898 10291 6901
rect 10910 6898 10916 6900
rect 10225 6896 10916 6898
rect 10225 6840 10230 6896
rect 10286 6840 10916 6896
rect 10225 6838 10916 6840
rect 10225 6835 10291 6838
rect 10910 6836 10916 6838
rect 10980 6898 10986 6900
rect 11237 6898 11303 6901
rect 10980 6896 11303 6898
rect 10980 6840 11242 6896
rect 11298 6840 11303 6896
rect 10980 6838 11303 6840
rect 10980 6836 10986 6838
rect 11237 6835 11303 6838
rect 16113 6898 16179 6901
rect 17714 6898 18514 6928
rect 16113 6896 18514 6898
rect 16113 6840 16118 6896
rect 16174 6840 18514 6896
rect 16113 6838 18514 6840
rect 16113 6835 16179 6838
rect 17714 6808 18514 6838
rect 5625 6762 5691 6765
rect 8937 6764 9003 6765
rect 6678 6762 6684 6764
rect 5625 6760 6684 6762
rect 5625 6704 5630 6760
rect 5686 6704 6684 6760
rect 5625 6702 6684 6704
rect 5625 6699 5691 6702
rect 6678 6700 6684 6702
rect 6748 6700 6754 6764
rect 8886 6700 8892 6764
rect 8956 6762 9003 6764
rect 8956 6760 12450 6762
rect 8998 6704 12450 6760
rect 8956 6702 12450 6704
rect 8956 6700 9003 6702
rect 6686 6626 6746 6700
rect 8937 6699 9003 6700
rect 11145 6626 11211 6629
rect 6686 6624 11211 6626
rect 6686 6568 11150 6624
rect 11206 6568 11211 6624
rect 6686 6566 11211 6568
rect 12390 6626 12450 6702
rect 13629 6626 13695 6629
rect 12390 6624 13695 6626
rect 12390 6568 13634 6624
rect 13690 6568 13695 6624
rect 12390 6566 13695 6568
rect 11145 6563 11211 6566
rect 13629 6563 13695 6566
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 7465 6490 7531 6493
rect 7833 6490 7899 6493
rect 7465 6488 7899 6490
rect 7465 6432 7470 6488
rect 7526 6432 7838 6488
rect 7894 6432 7899 6488
rect 7465 6430 7899 6432
rect 7465 6427 7531 6430
rect 7833 6427 7899 6430
rect 10358 6428 10364 6492
rect 10428 6490 10434 6492
rect 10869 6490 10935 6493
rect 10428 6488 10935 6490
rect 10428 6432 10874 6488
rect 10930 6432 10935 6488
rect 10428 6430 10935 6432
rect 10428 6428 10434 6430
rect 10869 6427 10935 6430
rect 841 6354 907 6357
rect 798 6352 907 6354
rect 798 6296 846 6352
rect 902 6296 907 6352
rect 798 6291 907 6296
rect 6453 6354 6519 6357
rect 9305 6354 9371 6357
rect 6453 6352 9371 6354
rect 6453 6296 6458 6352
rect 6514 6296 9310 6352
rect 9366 6296 9371 6352
rect 6453 6294 9371 6296
rect 6453 6291 6519 6294
rect 9305 6291 9371 6294
rect 798 6248 858 6291
rect 0 6158 858 6248
rect 16941 6218 17007 6221
rect 17714 6218 18514 6248
rect 16941 6216 18514 6218
rect 16941 6160 16946 6216
rect 17002 6160 18514 6216
rect 16941 6158 18514 6160
rect 0 6128 800 6158
rect 16941 6155 17007 6158
rect 17714 6128 18514 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 8017 5810 8083 5813
rect 5950 5808 8083 5810
rect 5950 5752 8022 5808
rect 8078 5752 8083 5808
rect 5950 5750 8083 5752
rect 5717 5674 5783 5677
rect 5950 5674 6010 5750
rect 8017 5747 8083 5750
rect 9070 5748 9076 5812
rect 9140 5810 9146 5812
rect 9305 5810 9371 5813
rect 9140 5808 9371 5810
rect 9140 5752 9310 5808
rect 9366 5752 9371 5808
rect 9140 5750 9371 5752
rect 9140 5748 9146 5750
rect 9305 5747 9371 5750
rect 10409 5810 10475 5813
rect 13537 5810 13603 5813
rect 14181 5812 14247 5813
rect 14181 5810 14228 5812
rect 10409 5808 13603 5810
rect 10409 5752 10414 5808
rect 10470 5752 13542 5808
rect 13598 5752 13603 5808
rect 10409 5750 13603 5752
rect 14136 5808 14228 5810
rect 14136 5752 14186 5808
rect 14136 5750 14228 5752
rect 10409 5747 10475 5750
rect 13537 5747 13603 5750
rect 14181 5748 14228 5750
rect 14292 5748 14298 5812
rect 14181 5747 14247 5748
rect 5717 5672 6010 5674
rect 5717 5616 5722 5672
rect 5778 5616 6010 5672
rect 5717 5614 6010 5616
rect 6177 5674 6243 5677
rect 6453 5674 6519 5677
rect 6177 5672 6519 5674
rect 6177 5616 6182 5672
rect 6238 5616 6458 5672
rect 6514 5616 6519 5672
rect 6177 5614 6519 5616
rect 5717 5611 5783 5614
rect 6177 5611 6243 5614
rect 6453 5611 6519 5614
rect 6729 5674 6795 5677
rect 11830 5674 11836 5676
rect 6729 5672 11836 5674
rect 6729 5616 6734 5672
rect 6790 5616 11836 5672
rect 6729 5614 11836 5616
rect 6729 5611 6795 5614
rect 11830 5612 11836 5614
rect 11900 5674 11906 5676
rect 12709 5674 12775 5677
rect 11900 5672 12775 5674
rect 11900 5616 12714 5672
rect 12770 5616 12775 5672
rect 11900 5614 12775 5616
rect 11900 5612 11906 5614
rect 12709 5611 12775 5614
rect 0 5538 800 5568
rect 1853 5538 1919 5541
rect 0 5536 1919 5538
rect 0 5480 1858 5536
rect 1914 5480 1919 5536
rect 0 5478 1919 5480
rect 0 5448 800 5478
rect 1853 5475 1919 5478
rect 6269 5538 6335 5541
rect 6545 5538 6611 5541
rect 6269 5536 6611 5538
rect 6269 5480 6274 5536
rect 6330 5480 6550 5536
rect 6606 5480 6611 5536
rect 6269 5478 6611 5480
rect 6269 5475 6335 5478
rect 6545 5475 6611 5478
rect 16941 5538 17007 5541
rect 17714 5538 18514 5568
rect 16941 5536 18514 5538
rect 16941 5480 16946 5536
rect 17002 5480 18514 5536
rect 16941 5478 18514 5480
rect 16941 5475 17007 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 17714 5448 18514 5478
rect 4870 5407 5186 5408
rect 5809 5402 5875 5405
rect 6361 5402 6427 5405
rect 6545 5402 6611 5405
rect 7649 5402 7715 5405
rect 5809 5400 6427 5402
rect 5809 5344 5814 5400
rect 5870 5344 6366 5400
rect 6422 5344 6427 5400
rect 5809 5342 6427 5344
rect 5809 5339 5875 5342
rect 6361 5339 6427 5342
rect 6502 5400 7715 5402
rect 6502 5344 6550 5400
rect 6606 5344 7654 5400
rect 7710 5344 7715 5400
rect 6502 5342 7715 5344
rect 6502 5339 6611 5342
rect 7649 5339 7715 5342
rect 8017 5402 8083 5405
rect 8661 5402 8727 5405
rect 8017 5400 8727 5402
rect 8017 5344 8022 5400
rect 8078 5344 8666 5400
rect 8722 5344 8727 5400
rect 8017 5342 8727 5344
rect 8017 5339 8083 5342
rect 8661 5339 8727 5342
rect 5165 5266 5231 5269
rect 6502 5266 6562 5339
rect 5165 5264 6562 5266
rect 5165 5208 5170 5264
rect 5226 5208 6562 5264
rect 5165 5206 6562 5208
rect 5165 5203 5231 5206
rect 6862 5204 6868 5268
rect 6932 5266 6938 5268
rect 7281 5266 7347 5269
rect 8477 5266 8543 5269
rect 6932 5264 8543 5266
rect 6932 5208 7286 5264
rect 7342 5208 8482 5264
rect 8538 5208 8543 5264
rect 6932 5206 8543 5208
rect 6932 5204 6938 5206
rect 7281 5203 7347 5206
rect 8477 5203 8543 5206
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 0 4178 800 4208
rect 1853 4178 1919 4181
rect 0 4176 1919 4178
rect 0 4120 1858 4176
rect 1914 4120 1919 4176
rect 0 4118 1919 4120
rect 0 4088 800 4118
rect 1853 4115 1919 4118
rect 10685 4044 10751 4045
rect 10685 4042 10732 4044
rect 10640 4040 10732 4042
rect 10640 3984 10690 4040
rect 10640 3982 10732 3984
rect 10685 3980 10732 3982
rect 10796 3980 10802 4044
rect 10685 3979 10751 3980
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 12198 3708 12204 3772
rect 12268 3770 12274 3772
rect 12525 3770 12591 3773
rect 12268 3768 12591 3770
rect 12268 3712 12530 3768
rect 12586 3712 12591 3768
rect 12268 3710 12591 3712
rect 12268 3708 12274 3710
rect 12525 3707 12591 3710
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 9628 15268 9692 15332
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 6684 14920 6748 14924
rect 6684 14864 6698 14920
rect 6698 14864 6748 14920
rect 6684 14860 6748 14864
rect 14228 14860 14292 14924
rect 6316 14724 6380 14788
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 8892 14240 8956 14244
rect 8892 14184 8942 14240
rect 8942 14184 8956 14240
rect 8892 14180 8956 14184
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 9076 13908 9140 13972
rect 9260 13772 9324 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 6500 13364 6564 13428
rect 8156 13092 8220 13156
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 12204 12820 12268 12884
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 6500 12140 6564 12204
rect 7236 12140 7300 12204
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 10916 11324 10980 11388
rect 6868 11052 6932 11116
rect 9076 11052 9140 11116
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 10364 10916 10428 10980
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 6316 10236 6380 10300
rect 7236 10372 7300 10436
rect 11836 9888 11900 9892
rect 11836 9832 11886 9888
rect 11886 9832 11900 9888
rect 11836 9828 11900 9832
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 6500 8740 6564 8804
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 10732 8332 10796 8396
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 8156 7984 8220 7988
rect 8156 7928 8206 7984
rect 8206 7928 8220 7984
rect 8156 7924 8220 7928
rect 9260 7652 9324 7716
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 9628 7516 9692 7580
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 8708 6972 8772 7036
rect 10916 6836 10980 6900
rect 6684 6700 6748 6764
rect 8892 6760 8956 6764
rect 8892 6704 8942 6760
rect 8942 6704 8956 6760
rect 8892 6700 8956 6704
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 10364 6428 10428 6492
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 9076 5748 9140 5812
rect 14228 5808 14292 5812
rect 14228 5752 14242 5808
rect 14242 5752 14292 5808
rect 14228 5748 14292 5752
rect 11836 5612 11900 5676
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 6868 5204 6932 5268
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 10732 4040 10796 4044
rect 10732 3984 10746 4040
rect 10746 3984 10796 4040
rect 10732 3980 10796 3984
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 12204 3708 12268 3772
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 17984 4528 18000
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 17440 5188 18000
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 9627 15332 9693 15333
rect 9627 15268 9628 15332
rect 9692 15268 9693 15332
rect 9627 15267 9693 15268
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 6683 14924 6749 14925
rect 6683 14860 6684 14924
rect 6748 14860 6749 14924
rect 6683 14859 6749 14860
rect 6315 14788 6381 14789
rect 6315 14724 6316 14788
rect 6380 14724 6381 14788
rect 6315 14723 6381 14724
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 6318 10301 6378 14723
rect 6499 13428 6565 13429
rect 6499 13364 6500 13428
rect 6564 13364 6565 13428
rect 6499 13363 6565 13364
rect 6502 12205 6562 13363
rect 6499 12204 6565 12205
rect 6499 12140 6500 12204
rect 6564 12140 6565 12204
rect 6499 12139 6565 12140
rect 6315 10300 6381 10301
rect 6315 10236 6316 10300
rect 6380 10236 6381 10300
rect 6315 10235 6381 10236
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 6502 8805 6562 12139
rect 6499 8804 6565 8805
rect 6499 8740 6500 8804
rect 6564 8740 6565 8804
rect 6499 8739 6565 8740
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 6686 6765 6746 14859
rect 8891 14244 8957 14245
rect 8891 14180 8892 14244
rect 8956 14180 8957 14244
rect 8891 14179 8957 14180
rect 8155 13156 8221 13157
rect 8155 13092 8156 13156
rect 8220 13092 8221 13156
rect 8155 13091 8221 13092
rect 7235 12204 7301 12205
rect 7235 12140 7236 12204
rect 7300 12140 7301 12204
rect 7235 12139 7301 12140
rect 6867 11116 6933 11117
rect 6867 11052 6868 11116
rect 6932 11052 6933 11116
rect 6867 11051 6933 11052
rect 6683 6764 6749 6765
rect 6683 6700 6684 6764
rect 6748 6700 6749 6764
rect 6683 6699 6749 6700
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 6870 5269 6930 11051
rect 7238 10437 7298 12139
rect 7235 10436 7301 10437
rect 7235 10372 7236 10436
rect 7300 10372 7301 10436
rect 7235 10371 7301 10372
rect 8158 7989 8218 13091
rect 8894 12450 8954 14179
rect 9075 13972 9141 13973
rect 9075 13908 9076 13972
rect 9140 13908 9141 13972
rect 9075 13907 9141 13908
rect 8710 12390 8954 12450
rect 8155 7988 8221 7989
rect 8155 7924 8156 7988
rect 8220 7924 8221 7988
rect 8155 7923 8221 7924
rect 8710 7037 8770 12390
rect 9078 11250 9138 13907
rect 9259 13836 9325 13837
rect 9259 13772 9260 13836
rect 9324 13772 9325 13836
rect 9259 13771 9325 13772
rect 8894 11190 9138 11250
rect 8707 7036 8773 7037
rect 8707 6972 8708 7036
rect 8772 6972 8773 7036
rect 8707 6971 8773 6972
rect 8894 6765 8954 11190
rect 9075 11116 9141 11117
rect 9075 11052 9076 11116
rect 9140 11052 9141 11116
rect 9075 11051 9141 11052
rect 8891 6764 8957 6765
rect 8891 6700 8892 6764
rect 8956 6700 8957 6764
rect 8891 6699 8957 6700
rect 9078 5813 9138 11051
rect 9262 7717 9322 13771
rect 9259 7716 9325 7717
rect 9259 7652 9260 7716
rect 9324 7652 9325 7716
rect 9259 7651 9325 7652
rect 9630 7581 9690 15267
rect 14227 14924 14293 14925
rect 14227 14860 14228 14924
rect 14292 14860 14293 14924
rect 14227 14859 14293 14860
rect 12203 12884 12269 12885
rect 12203 12820 12204 12884
rect 12268 12820 12269 12884
rect 12203 12819 12269 12820
rect 10915 11388 10981 11389
rect 10915 11324 10916 11388
rect 10980 11324 10981 11388
rect 10915 11323 10981 11324
rect 10363 10980 10429 10981
rect 10363 10916 10364 10980
rect 10428 10916 10429 10980
rect 10363 10915 10429 10916
rect 9627 7580 9693 7581
rect 9627 7516 9628 7580
rect 9692 7516 9693 7580
rect 9627 7515 9693 7516
rect 10366 6493 10426 10915
rect 10731 8396 10797 8397
rect 10731 8332 10732 8396
rect 10796 8332 10797 8396
rect 10731 8331 10797 8332
rect 10363 6492 10429 6493
rect 10363 6428 10364 6492
rect 10428 6428 10429 6492
rect 10363 6427 10429 6428
rect 9075 5812 9141 5813
rect 9075 5748 9076 5812
rect 9140 5748 9141 5812
rect 9075 5747 9141 5748
rect 6867 5268 6933 5269
rect 6867 5204 6868 5268
rect 6932 5204 6933 5268
rect 6867 5203 6933 5204
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 10734 4045 10794 8331
rect 10918 6901 10978 11323
rect 11835 9892 11901 9893
rect 11835 9828 11836 9892
rect 11900 9828 11901 9892
rect 11835 9827 11901 9828
rect 10915 6900 10981 6901
rect 10915 6836 10916 6900
rect 10980 6836 10981 6900
rect 10915 6835 10981 6836
rect 11838 5677 11898 9827
rect 11835 5676 11901 5677
rect 11835 5612 11836 5676
rect 11900 5612 11901 5676
rect 11835 5611 11901 5612
rect 10731 4044 10797 4045
rect 10731 3980 10732 4044
rect 10796 3980 10797 4044
rect 10731 3979 10797 3980
rect 12206 3773 12266 12819
rect 14230 5813 14290 14859
rect 14227 5812 14293 5813
rect 14227 5748 14228 5812
rect 14292 5748 14293 5812
rect 14227 5747 14293 5748
rect 12203 3772 12269 3773
rect 12203 3708 12204 3772
rect 12268 3708 12269 3772
rect 12203 3707 12269 3708
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1
transform 1 0 16100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _242_
timestamp 1
transform -1 0 8096 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_2  _243_
timestamp 1
transform -1 0 3036 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _244_
timestamp 1
transform 1 0 9200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_1  _245_
timestamp 1
transform 1 0 7084 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_2  _246_
timestamp 1
transform -1 0 3036 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _247_
timestamp 1
transform 1 0 4876 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _248_
timestamp 1
transform -1 0 4692 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_2  _249_
timestamp 1
transform 1 0 3588 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _250_
timestamp 1
transform 1 0 5520 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _251_
timestamp 1
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _252_
timestamp 1
transform -1 0 6808 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_2  _253_
timestamp 1
transform 1 0 2116 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_2  _254_
timestamp 1
transform -1 0 3128 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _255_
timestamp 1
transform 1 0 4876 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _256_
timestamp 1
transform 1 0 10396 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _257_
timestamp 1
transform 1 0 4876 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_2  _258_
timestamp 1
transform 1 0 2852 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__and4bb_2  _259_
timestamp 1
transform -1 0 4876 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _260_
timestamp 1
transform 1 0 5612 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _261_
timestamp 1
transform 1 0 8372 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _262_
timestamp 1
transform -1 0 9568 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_2  _263_
timestamp 1
transform 1 0 3404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__and3b_1  _264_
timestamp 1
transform 1 0 6716 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _265_
timestamp 1
transform 1 0 4508 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _266_
timestamp 1
transform 1 0 7820 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _267_
timestamp 1
transform -1 0 3404 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _268_
timestamp 1
transform -1 0 9476 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _269_
timestamp 1
transform 1 0 13248 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _270_
timestamp 1
transform 1 0 4692 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _271_
timestamp 1
transform 1 0 4784 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _272_
timestamp 1
transform 1 0 9476 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_1  _273_
timestamp 1
transform 1 0 5520 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_2  _274_
timestamp 1
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_2  _275_
timestamp 1
transform 1 0 2024 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _276_
timestamp 1
transform 1 0 6532 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _277_
timestamp 1
transform 1 0 7176 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _278_
timestamp 1
transform 1 0 3036 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _279_
timestamp 1
transform 1 0 4416 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _280_
timestamp 1
transform 1 0 9292 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_2  _281_
timestamp 1
transform 1 0 3772 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor4b_2  _282_
timestamp 1
transform 1 0 2024 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _283_
timestamp 1
transform 1 0 8004 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _284_
timestamp 1
transform 1 0 7912 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _285_
timestamp 1
transform 1 0 9660 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _286_
timestamp 1
transform 1 0 10764 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _287_
timestamp 1
transform 1 0 3036 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _288_
timestamp 1
transform 1 0 3220 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _289_
timestamp 1
transform 1 0 3772 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _290_
timestamp 1
transform 1 0 3220 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _291_
timestamp 1
transform 1 0 7268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _292_
timestamp 1
transform 1 0 4876 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _293_
timestamp 1
transform -1 0 6072 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _294_
timestamp 1
transform 1 0 8372 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _295_
timestamp 1
transform 1 0 7268 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _296_
timestamp 1
transform 1 0 7452 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _297_
timestamp 1
transform 1 0 8648 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _298_
timestamp 1
transform 1 0 9016 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _299_
timestamp 1
transform 1 0 7912 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _300_
timestamp 1
transform 1 0 5520 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _301_
timestamp 1
transform -1 0 11040 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _302_
timestamp 1
transform 1 0 7084 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _303_
timestamp 1
transform 1 0 6624 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _304_
timestamp 1
transform 1 0 11408 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _305_
timestamp 1
transform 1 0 6992 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _306_
timestamp 1
transform 1 0 6808 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _307_
timestamp 1
transform 1 0 12788 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _308_
timestamp 1
transform 1 0 6348 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _309_
timestamp 1
transform -1 0 10212 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _310_
timestamp 1
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _311_
timestamp 1
transform -1 0 14996 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_1  _312_
timestamp 1
transform 1 0 8004 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _313_
timestamp 1
transform 1 0 7820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _314_
timestamp 1
transform 1 0 8004 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _315_
timestamp 1
transform 1 0 7452 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _316_
timestamp 1
transform 1 0 7360 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _317_
timestamp 1
transform 1 0 7636 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _318_
timestamp 1
transform -1 0 14168 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _319_
timestamp 1
transform -1 0 13708 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _320_
timestamp 1
transform 1 0 2760 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _321_
timestamp 1
transform -1 0 6164 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _322_
timestamp 1
transform 1 0 3404 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _323_
timestamp 1
transform 1 0 3772 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _324_
timestamp 1
transform 1 0 4048 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _325_
timestamp 1
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _326_
timestamp 1
transform 1 0 13616 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _327_
timestamp 1
transform 1 0 7360 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _328_
timestamp 1
transform 1 0 7452 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _329_
timestamp 1
transform 1 0 10580 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _330_
timestamp 1
transform 1 0 7176 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _331_
timestamp 1
transform -1 0 12512 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _332_
timestamp 1
transform 1 0 13064 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _333_
timestamp 1
transform 1 0 12420 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _334_
timestamp 1
transform 1 0 6808 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _335_
timestamp 1
transform 1 0 3036 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _336_
timestamp 1
transform 1 0 7820 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _337_
timestamp 1
transform 1 0 2392 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _338_
timestamp 1
transform 1 0 5980 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _339_
timestamp 1
transform 1 0 7176 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _340_
timestamp 1
transform -1 0 13524 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _341_
timestamp 1
transform 1 0 7360 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _342_
timestamp 1
transform -1 0 6716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _343_
timestamp 1
transform 1 0 8004 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _344_
timestamp 1
transform 1 0 7360 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _345_
timestamp 1
transform 1 0 11040 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_1  _346_
timestamp 1
transform 1 0 5244 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _347_
timestamp 1
transform 1 0 5060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _348_
timestamp 1
transform 1 0 6348 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _349_
timestamp 1
transform -1 0 12788 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _350_
timestamp 1
transform 1 0 4232 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _351_
timestamp 1
transform 1 0 4784 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _352_
timestamp 1
transform 1 0 10028 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _353_
timestamp 1
transform 1 0 7544 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _354_
timestamp 1
transform 1 0 5060 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _355_
timestamp 1
transform -1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _356_
timestamp 1
transform 1 0 11868 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _357_
timestamp 1
transform 1 0 4508 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _358_
timestamp 1
transform 1 0 4416 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _359_
timestamp 1
transform 1 0 12052 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _360_
timestamp 1
transform 1 0 13800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _361_
timestamp 1
transform 1 0 4784 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _362_
timestamp 1
transform 1 0 5428 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _363_
timestamp 1
transform 1 0 4232 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _364_
timestamp 1
transform 1 0 4508 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _365_
timestamp 1
transform 1 0 11776 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _366_
timestamp 1
transform 1 0 5612 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a2111oi_1  _367_
timestamp 1
transform -1 0 10948 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a41oi_1  _368_
timestamp 1
transform -1 0 13800 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _369_
timestamp 1
transform 1 0 14076 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _370_
timestamp 1
transform -1 0 6348 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _371_
timestamp 1
transform 1 0 9292 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _372_
timestamp 1
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _373_
timestamp 1
transform 1 0 10396 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _374_
timestamp 1
transform 1 0 9292 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _375_
timestamp 1
transform 1 0 9752 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _376_
timestamp 1
transform 1 0 10488 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _377_
timestamp 1
transform 1 0 11316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _378_
timestamp 1
transform 1 0 14996 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _379_
timestamp 1
transform 1 0 11868 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _380_
timestamp 1
transform 1 0 9108 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _381_
timestamp 1
transform 1 0 12880 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _382_
timestamp 1
transform 1 0 12512 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _383_
timestamp 1
transform 1 0 10948 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _384_
timestamp 1
transform 1 0 5612 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _385_
timestamp 1
transform 1 0 9200 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _386_
timestamp 1
transform -1 0 11408 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _387_
timestamp 1
transform -1 0 11960 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _388_
timestamp 1
transform 1 0 8924 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _389_
timestamp 1
transform 1 0 11408 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _390_
timestamp 1
transform 1 0 9844 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _391_
timestamp 1
transform 1 0 10856 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _392_
timestamp 1
transform 1 0 12236 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _393_
timestamp 1
transform -1 0 13156 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _394_
timestamp 1
transform 1 0 10580 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _395_
timestamp 1
transform 1 0 10120 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _396_
timestamp 1
transform 1 0 11316 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _397_
timestamp 1
transform 1 0 11500 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _398_
timestamp 1
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _399_
timestamp 1
transform 1 0 13524 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _400_
timestamp 1
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _401_
timestamp 1
transform -1 0 11592 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _402_
timestamp 1
transform -1 0 7084 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _403_
timestamp 1
transform 1 0 10856 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _404_
timestamp 1
transform 1 0 14444 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _405_
timestamp 1
transform 1 0 14996 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _406_
timestamp 1
transform -1 0 14168 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _407_
timestamp 1
transform 1 0 13432 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _408_
timestamp 1
transform 1 0 10396 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _409_
timestamp 1
transform 1 0 13248 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _410_
timestamp 1
transform 1 0 13892 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _411_
timestamp 1
transform 1 0 15088 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _412_
timestamp 1
transform 1 0 11316 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _413_
timestamp 1
transform -1 0 12696 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _414_
timestamp 1
transform 1 0 9108 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _415_
timestamp 1
transform 1 0 4324 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _416_
timestamp 1
transform 1 0 10304 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _417_
timestamp 1
transform -1 0 9936 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _418_
timestamp 1
transform 1 0 9660 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _419_
timestamp 1
transform 1 0 8832 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _420_
timestamp 1
transform 1 0 10120 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _421_
timestamp 1
transform 1 0 12052 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _422_
timestamp 1
transform 1 0 13064 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _423_
timestamp 1
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _424_
timestamp 1
transform 1 0 13064 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _425_
timestamp 1
transform 1 0 13340 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _426_
timestamp 1
transform 1 0 13800 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _427_
timestamp 1
transform 1 0 7360 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _428_
timestamp 1
transform 1 0 8832 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _429_
timestamp 1
transform 1 0 9568 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _430_
timestamp 1
transform 1 0 10304 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _431_
timestamp 1
transform 1 0 14260 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _432_
timestamp 1
transform 1 0 14260 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _433_
timestamp 1
transform 1 0 14076 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _434_
timestamp 1
transform -1 0 6900 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _435_
timestamp 1
transform 1 0 6256 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _436_
timestamp 1
transform -1 0 7360 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _437_
timestamp 1
transform -1 0 6624 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _438_
timestamp 1
transform 1 0 14996 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _439_
timestamp 1
transform 1 0 14996 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _440_
timestamp 1
transform 1 0 7452 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _441_
timestamp 1
transform 1 0 12236 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _442_
timestamp 1
transform 1 0 13248 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _443_
timestamp 1
transform 1 0 14536 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _444_
timestamp 1
transform 1 0 14352 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _445_
timestamp 1
transform 1 0 14996 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _446_
timestamp 1
transform 1 0 15180 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _447_
timestamp 1
transform 1 0 11500 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _448_
timestamp 1
transform 1 0 11500 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _449_
timestamp 1
transform 1 0 12052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _450_
timestamp 1
transform 1 0 12328 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _451_
timestamp 1
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _452_
timestamp 1
transform 1 0 13892 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _453_
timestamp 1
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _454_
timestamp 1
transform 1 0 9752 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _455_
timestamp 1
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _456_
timestamp 1
transform 1 0 11132 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _457_
timestamp 1
transform 1 0 12052 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _458_
timestamp 1
transform 1 0 12604 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _459_
timestamp 1
transform 1 0 15180 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _460_
timestamp 1
transform 1 0 8648 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _461_
timestamp 1
transform 1 0 9292 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _462_
timestamp 1
transform 1 0 11868 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _463_
timestamp 1
transform 1 0 13156 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _464_
timestamp 1
transform 1 0 14168 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _465_
timestamp 1
transform 1 0 15180 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _466_
timestamp 1
transform -1 0 10948 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _467_
timestamp 1
transform 1 0 9568 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _468_
timestamp 1
transform 1 0 7820 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _469_
timestamp 1
transform 1 0 9936 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _470_
timestamp 1
transform 1 0 14444 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _471_
timestamp 1
transform 1 0 14996 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _472_
timestamp 1
transform 1 0 12512 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _473_
timestamp 1
transform 1 0 13248 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _474_
timestamp 1
transform 1 0 14536 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _475_
timestamp 1
transform 1 0 15548 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _476_
timestamp 1
transform 1 0 13524 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _477_
timestamp 1
transform 1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _478_
timestamp 1
transform -1 0 13984 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _479_
timestamp 1
transform 1 0 14996 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _480_
timestamp 1
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _481_
timestamp 1
transform 1 0 14536 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _482_
timestamp 1
transform 1 0 1380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _483_
timestamp 1
transform 1 0 1380 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _484_
timestamp 1
transform 1 0 1380 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _485_
timestamp 1
transform 1 0 1380 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _486_
timestamp 1
transform 1 0 9936 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _487_
timestamp 1
transform 1 0 6348 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _488_
timestamp 1
transform 1 0 8464 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _489_
timestamp 1
transform 1 0 15640 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _490_
timestamp 1
transform 1 0 11868 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _491_
timestamp 1
transform 1 0 15640 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _492_
timestamp 1
transform 1 0 15272 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _493_
timestamp 1
transform 1 0 13340 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _494_
timestamp 1
transform 1 0 15640 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _495_
timestamp 1
transform 1 0 15640 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _496_
timestamp 1
transform 1 0 15640 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _497_
timestamp 1
transform 1 0 14536 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _498_
timestamp 1
transform 1 0 15640 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _499_
timestamp 1
transform 1 0 15640 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _500_
timestamp 1
transform 1 0 15640 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _501_
timestamp 1
transform 1 0 15088 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _502_
timestamp 1
transform 1 0 15640 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _503_
timestamp 1
transform -1 0 14628 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _504_
timestamp 1
transform 1 0 14628 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk0
timestamp 1
transform 1 0 8556 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk0
timestamp 1
transform -1 0 10764 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk0
timestamp 1
transform 1 0 10212 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinv_2  clkload0
timestamp 1
transform -1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 1
transform 1 0 15456 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1
transform 1 0 7176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout28
timestamp 1
transform -1 0 6992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout30
timestamp 1
transform -1 0 8004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1
transform 1 0 7268 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout32
timestamp 1
transform -1 0 5796 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 1
transform 1 0 8280 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout34
timestamp 1
transform -1 0 5980 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 1
transform 1 0 8464 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout38
timestamp 1
transform -1 0 7820 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp 1
transform 1 0 9292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout41
timestamp 1
transform -1 0 7268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout43
timestamp 1
transform 1 0 8004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout44
timestamp 1
transform -1 0 6256 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 1
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout46
timestamp 1
transform -1 0 6992 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout47
timestamp 1
transform -1 0 11592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout48
timestamp 1
transform -1 0 2024 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout49
timestamp 1
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout50
timestamp 1
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout51
timestamp 1
transform 1 0 3312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout52
timestamp 1
transform 1 0 3128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout53
timestamp 1
transform 1 0 3312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout54
timestamp 1
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout55
timestamp 1
transform -1 0 3312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout56
timestamp 1
transform -1 0 14996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout57
timestamp 1
transform -1 0 17020 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_41
timestamp 1
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_49
timestamp 1
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_90
timestamp 1
transform 1 0 9384 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_98
timestamp 1
transform 1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_104
timestamp 1
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_125
timestamp 1
transform 1 0 12604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_133
timestamp 1
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_149
timestamp 1636968456
transform 1 0 14812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_161
timestamp 1
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_169
timestamp 1
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_173
timestamp 1
transform 1 0 17020 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_79
timestamp 1
transform 1 0 8372 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_125
timestamp 1
transform 1 0 12604 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_155
timestamp 1636968456
transform 1 0 15364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_169
timestamp 1
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_173
timestamp 1
transform 1 0 17020 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_53
timestamp 1
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_81
timestamp 1
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_92
timestamp 1
transform 1 0 9568 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_100
timestamp 1
transform 1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_114
timestamp 1
transform 1 0 11592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_118
timestamp 1
transform 1 0 11960 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_125
timestamp 1636968456
transform 1 0 12604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_137
timestamp 1
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_141
timestamp 1
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_166
timestamp 1
transform 1 0 16376 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_9
timestamp 1636968456
transform 1 0 1932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_21
timestamp 1636968456
transform 1 0 3036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_33
timestamp 1636968456
transform 1 0 4140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_45
timestamp 1
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_53
timestamp 1
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_76
timestamp 1636968456
transform 1 0 8096 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_91
timestamp 1
transform 1 0 9476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_113
timestamp 1
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_122
timestamp 1
transform 1 0 12328 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_130
timestamp 1
transform 1 0 13064 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_169
timestamp 1
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_173
timestamp 1
transform 1 0 17020 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_19
timestamp 1
transform 1 0 2852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_23
timestamp 1
transform 1 0 3220 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_53
timestamp 1
transform 1 0 5980 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_59
timestamp 1
transform 1 0 6532 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_64
timestamp 1
transform 1 0 6992 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_81
timestamp 1
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_85
timestamp 1
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_98
timestamp 1
transform 1 0 10120 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_106
timestamp 1
transform 1 0 10856 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_111
timestamp 1636968456
transform 1 0 11316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_123
timestamp 1636968456
transform 1 0 12420 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_135
timestamp 1
transform 1 0 13524 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_141
timestamp 1
transform 1 0 14076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_19
timestamp 1
transform 1 0 2852 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_51
timestamp 1
transform 1 0 5796 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_64
timestamp 1
transform 1 0 6992 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_84
timestamp 1
transform 1 0 8832 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_100
timestamp 1636968456
transform 1 0 10304 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_113
timestamp 1
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_127
timestamp 1636968456
transform 1 0 12788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_139
timestamp 1636968456
transform 1 0 13892 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_151
timestamp 1
transform 1 0 14996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_155
timestamp 1
transform 1 0 15364 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_169
timestamp 1
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_19
timestamp 1
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_38
timestamp 1
transform 1 0 4600 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_46
timestamp 1
transform 1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_60
timestamp 1
transform 1 0 6624 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_85
timestamp 1
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_93
timestamp 1
transform 1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_108
timestamp 1
transform 1 0 11040 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_117
timestamp 1636968456
transform 1 0 11868 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_129
timestamp 1
transform 1 0 12972 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_147
timestamp 1
transform 1 0 14628 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_9
timestamp 1
transform 1 0 1932 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_17
timestamp 1
transform 1 0 2668 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_41
timestamp 1
transform 1 0 4876 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_49
timestamp 1
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 1
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_65
timestamp 1
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_82
timestamp 1
transform 1 0 8648 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_88
timestamp 1
transform 1 0 9200 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_94
timestamp 1636968456
transform 1 0 9752 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_106
timestamp 1
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1636968456
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_125
timestamp 1
transform 1 0 12604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_129
timestamp 1
transform 1 0 12972 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_142
timestamp 1
transform 1 0 14168 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_150
timestamp 1
transform 1 0 14904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_169
timestamp 1
transform 1 0 16652 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_19
timestamp 1
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_29
timestamp 1
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_37
timestamp 1
transform 1 0 4508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_55
timestamp 1
transform 1 0 6164 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_63
timestamp 1
transform 1 0 6900 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 1
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_96
timestamp 1636968456
transform 1 0 9936 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_108
timestamp 1
transform 1 0 11040 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_115
timestamp 1
transform 1 0 11684 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_129
timestamp 1
transform 1 0 12972 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_135
timestamp 1
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_141
timestamp 1
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_150
timestamp 1
transform 1 0 14904 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_3
timestamp 1
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_26
timestamp 1
transform 1 0 3496 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_50
timestamp 1
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1636968456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1636968456
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_81
timestamp 1
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_90
timestamp 1
transform 1 0 9384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_103
timestamp 1
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_130
timestamp 1636968456
transform 1 0 13064 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_142
timestamp 1636968456
transform 1 0 14168 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_154
timestamp 1
transform 1 0 15272 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_160
timestamp 1
transform 1 0 15824 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_169
timestamp 1
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_3
timestamp 1
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_9
timestamp 1
transform 1 0 1932 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_20
timestamp 1
transform 1 0 2944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_24
timestamp 1
transform 1 0 3312 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_62
timestamp 1
transform 1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 1
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_116
timestamp 1636968456
transform 1 0 11776 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_128
timestamp 1
transform 1 0 12880 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_141
timestamp 1
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_156
timestamp 1
transform 1 0 15456 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_3
timestamp 1
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_21
timestamp 1
transform 1 0 3036 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1636968456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_39
timestamp 1
transform 1 0 4692 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_47
timestamp 1
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1636968456
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_80
timestamp 1
transform 1 0 8464 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_88
timestamp 1
transform 1 0 9200 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_118
timestamp 1
transform 1 0 11960 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_144
timestamp 1
transform 1 0 14352 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_152
timestamp 1
transform 1 0 15088 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_169
timestamp 1
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_3
timestamp 1
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_38
timestamp 1
transform 1 0 4600 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_55
timestamp 1
transform 1 0 6164 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_66
timestamp 1
transform 1 0 7176 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_76
timestamp 1
transform 1 0 8096 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1636968456
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_97
timestamp 1
transform 1 0 10028 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_105
timestamp 1
transform 1 0 10764 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_113
timestamp 1636968456
transform 1 0 11500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_125
timestamp 1
transform 1 0 12604 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_131
timestamp 1
transform 1 0 13156 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 1
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_147
timestamp 1
transform 1 0 14628 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_155
timestamp 1
transform 1 0 15364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_164
timestamp 1
transform 1 0 16192 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_173
timestamp 1
transform 1 0 17020 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 1
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_11
timestamp 1
transform 1 0 2116 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_22
timestamp 1636968456
transform 1 0 3128 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_34
timestamp 1
transform 1 0 4232 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_40
timestamp 1
transform 1 0 4784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_63
timestamp 1
transform 1 0 6900 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_67
timestamp 1
transform 1 0 7268 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_93
timestamp 1
transform 1 0 9660 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_101
timestamp 1
transform 1 0 10396 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_105
timestamp 1
transform 1 0 10764 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_118
timestamp 1636968456
transform 1 0 11960 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_130
timestamp 1
transform 1 0 13064 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_141
timestamp 1
transform 1 0 14076 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_145
timestamp 1
transform 1 0 14444 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_151
timestamp 1
transform 1 0 14996 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_169
timestamp 1
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_173
timestamp 1
transform 1 0 17020 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_3
timestamp 1
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_20
timestamp 1
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_96
timestamp 1636968456
transform 1 0 9936 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_108
timestamp 1
transform 1 0 11040 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_114
timestamp 1
transform 1 0 11592 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_122
timestamp 1
transform 1 0 12328 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_126
timestamp 1
transform 1 0 12696 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_141
timestamp 1
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_145
timestamp 1
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_151
timestamp 1636968456
transform 1 0 14996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_163
timestamp 1
transform 1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1636968456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_15
timestamp 1
transform 1 0 2484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_37
timestamp 1
transform 1 0 4508 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_48
timestamp 1
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_57
timestamp 1
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_61
timestamp 1
transform 1 0 6716 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_76
timestamp 1
transform 1 0 8096 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_80
timestamp 1
transform 1 0 8464 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_106
timestamp 1
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_118
timestamp 1636968456
transform 1 0 11960 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_130
timestamp 1
transform 1 0 13064 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_138
timestamp 1636968456
transform 1 0 13800 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_150
timestamp 1
transform 1 0 14904 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_158
timestamp 1
transform 1 0 15640 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_169
timestamp 1
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1636968456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1636968456
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_29
timestamp 1
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_37
timestamp 1
transform 1 0 4508 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_54
timestamp 1
transform 1 0 6072 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_62
timestamp 1
transform 1 0 6808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_85
timestamp 1
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_92
timestamp 1
transform 1 0 9568 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_98
timestamp 1
transform 1 0 10120 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_124
timestamp 1
transform 1 0 12512 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_135
timestamp 1
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_146
timestamp 1
transform 1 0 14536 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_150
timestamp 1
transform 1 0 14904 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1636968456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_15
timestamp 1
transform 1 0 2484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_30
timestamp 1
transform 1 0 3864 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_36
timestamp 1
transform 1 0 4416 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_44
timestamp 1636968456
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_65
timestamp 1
transform 1 0 7084 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_73
timestamp 1
transform 1 0 7820 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_81
timestamp 1
transform 1 0 8556 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_87
timestamp 1636968456
transform 1 0 9108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1636968456
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_125
timestamp 1
transform 1 0 12604 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_143
timestamp 1
transform 1 0 14260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_156
timestamp 1
transform 1 0 15456 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_173
timestamp 1
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_3
timestamp 1
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_11
timestamp 1
transform 1 0 2116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_29
timestamp 1
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_33
timestamp 1
transform 1 0 4140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_48
timestamp 1
transform 1 0 5520 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_75
timestamp 1
transform 1 0 8004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_85
timestamp 1
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_98
timestamp 1
transform 1 0 10120 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_118
timestamp 1
transform 1 0 11960 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_127
timestamp 1636968456
transform 1 0 12788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_141
timestamp 1
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_149
timestamp 1
transform 1 0 14812 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1636968456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_15
timestamp 1
transform 1 0 2484 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_30
timestamp 1
transform 1 0 3864 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_36
timestamp 1
transform 1 0 4416 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_44
timestamp 1
transform 1 0 5152 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_57
timestamp 1
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_72
timestamp 1636968456
transform 1 0 7728 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_84
timestamp 1636968456
transform 1 0 8832 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_96
timestamp 1
transform 1 0 9936 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_102
timestamp 1
transform 1 0 10488 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_108
timestamp 1
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_113
timestamp 1
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_121
timestamp 1
transform 1 0 12236 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_133
timestamp 1
transform 1 0 13340 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_141
timestamp 1
transform 1 0 14076 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_148
timestamp 1636968456
transform 1 0 14720 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_169
timestamp 1
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1636968456
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_15
timestamp 1
transform 1 0 2484 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_48
timestamp 1
transform 1 0 5520 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_76
timestamp 1
transform 1 0 8096 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_85
timestamp 1
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_91
timestamp 1
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_97
timestamp 1
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_107
timestamp 1636968456
transform 1 0 10948 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_119
timestamp 1
transform 1 0 12052 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_123
timestamp 1
transform 1 0 12420 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_130
timestamp 1
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_147
timestamp 1
transform 1 0 14628 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1636968456
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_15
timestamp 1
transform 1 0 2484 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_28
timestamp 1
transform 1 0 3680 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_34
timestamp 1
transform 1 0 4232 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_40
timestamp 1636968456
transform 1 0 4784 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_52
timestamp 1
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_57
timestamp 1
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_61
timestamp 1
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_74
timestamp 1
transform 1 0 7912 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_78
timestamp 1
transform 1 0 8280 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_90
timestamp 1
transform 1 0 9384 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_99
timestamp 1
transform 1 0 10212 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_106
timestamp 1
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_118
timestamp 1636968456
transform 1 0 11960 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_130
timestamp 1
transform 1 0 13064 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_138
timestamp 1
transform 1 0 13800 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_150
timestamp 1
transform 1 0 14904 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_159
timestamp 1
transform 1 0 15732 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_169
timestamp 1
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1636968456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1636968456
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1636968456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1636968456
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1636968456
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1636968456
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_90
timestamp 1636968456
transform 1 0 9384 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_102
timestamp 1
transform 1 0 10488 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_110
timestamp 1
transform 1 0 11224 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_117
timestamp 1
transform 1 0 11868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_126
timestamp 1
transform 1 0 12696 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1636968456
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_153
timestamp 1
transform 1 0 15180 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_170
timestamp 1
transform 1 0 16744 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1636968456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1636968456
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1636968456
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_39
timestamp 1
transform 1 0 4692 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_47
timestamp 1
transform 1 0 5428 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_63
timestamp 1
transform 1 0 6900 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_78
timestamp 1
transform 1 0 8280 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_86
timestamp 1
transform 1 0 9016 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_95
timestamp 1636968456
transform 1 0 9844 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_113
timestamp 1
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_123
timestamp 1
transform 1 0 12420 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_147
timestamp 1
transform 1 0 14628 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_169
timestamp 1
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1636968456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1636968456
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1636968456
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_41
timestamp 1
transform 1 0 4876 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_56
timestamp 1636968456
transform 1 0 6256 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_68
timestamp 1
transform 1 0 7360 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_72
timestamp 1
transform 1 0 7728 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_79
timestamp 1
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_85
timestamp 1
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_92
timestamp 1
transform 1 0 9568 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_104
timestamp 1
transform 1 0 10672 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_110
timestamp 1
transform 1 0 11224 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_126
timestamp 1636968456
transform 1 0 12696 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1636968456
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_153
timestamp 1
transform 1 0 15180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_157
timestamp 1
transform 1 0 15548 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1636968456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1636968456
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1636968456
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1636968456
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1636968456
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1636968456
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1636968456
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_93
timestamp 1
transform 1 0 9660 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_107
timestamp 1
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_113
timestamp 1
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_125
timestamp 1
transform 1 0 12604 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_129
timestamp 1
transform 1 0 12972 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_137
timestamp 1
transform 1 0 13708 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_162
timestamp 1
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_169
timestamp 1
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1636968456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1636968456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1636968456
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1636968456
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1636968456
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1636968456
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1636968456
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1636968456
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1636968456
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_121
timestamp 1
transform 1 0 12236 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_141
timestamp 1
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1636968456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1636968456
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1636968456
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1636968456
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1636968456
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1636968456
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1636968456
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1636968456
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_113
timestamp 1
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_157
timestamp 1
transform 1 0 15548 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_169
timestamp 1
transform 1 0 16652 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1636968456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1636968456
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1636968456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1636968456
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_53
timestamp 1
transform 1 0 5980 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_57
timestamp 1636968456
transform 1 0 6348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_69
timestamp 1636968456
transform 1 0 7452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_81
timestamp 1
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1636968456
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1636968456
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_109
timestamp 1
transform 1 0 11132 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_113
timestamp 1636968456
transform 1 0 11500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_125
timestamp 1
transform 1 0 12604 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_135
timestamp 1
transform 1 0 13524 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_147
timestamp 1636968456
transform 1 0 14628 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_159
timestamp 1
transform 1 0 15732 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_167
timestamp 1
transform 1 0 16468 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_169
timestamp 1
transform 1 0 16652 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_173
timestamp 1
transform 1 0 17020 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 15364 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform -1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 16560 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 16560 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform -1 0 16560 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform -1 0 16560 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform -1 0 16560 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 16560 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform -1 0 16560 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform -1 0 15640 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform -1 0 17020 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform -1 0 16560 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform -1 0 13892 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform -1 0 16560 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform -1 0 16560 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 15548 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform 1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform -1 0 6164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1
transform -1 0 16192 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap35
timestamp 1
transform -1 0 7360 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  max_cap36
timestamp 1
transform 1 0 9476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap39
timestamp 1
transform -1 0 7268 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap42
timestamp 1
transform -1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1
transform 1 0 16744 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1
transform 1 0 16744 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1
transform 1 0 16744 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1
transform 1 0 16376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1
transform 1 0 16744 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1
transform -1 0 13984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1
transform 1 0 16744 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1
transform -1 0 13524 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1
transform 1 0 16744 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1
transform 1 0 16744 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1
transform -1 0 14628 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1
transform 1 0 16744 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1
transform 1 0 16744 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1
transform 1 0 16744 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1
transform 1 0 16744 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1
transform -1 0 16560 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_29
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_30
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_31
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_32
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 17388 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_33
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_34
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 17388 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_35
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 17388 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_36
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 17388 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_37
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_38
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 17388 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_39
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 17388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_40
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 17388 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_41
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 17388 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_42
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 17388 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_43
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 17388 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_44
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 17388 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_45
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 17388 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_46
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 17388 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_47
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 17388 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_48
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 17388 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_49
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 17388 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_50
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 17388 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_51
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 17388 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_52
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 17388 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_53
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 17388 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_54
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 17388 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_55
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_56
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 17388 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_57
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 17388 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_64
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_65
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_66
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_67
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_68
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_69
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_70
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_71
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_72
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_73
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_74
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_75
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_77
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_78
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_80
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_81
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_83
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_85
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_86
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_89
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_90
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_92
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_93
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_94
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_95
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_96
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_97
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_98
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_99
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_100
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_101
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_102
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_103
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_104
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_105
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_106
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_107
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_108
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_109
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_110
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_111
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_112
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_113
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_114
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_115
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_116
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_117
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_118
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_119
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_120
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_121
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_122
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_123
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_124
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_125
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_126
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_127
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_128
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_129
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_130
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_131
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_132
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_133
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_134
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_135
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_136
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_137
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_138
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_139
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_140
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_141
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_142
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_143
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_144
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_145
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_146
timestamp 1
transform 1 0 6256 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_147
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_148
timestamp 1
transform 1 0 11408 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_149
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_150
timestamp 1
transform 1 0 16560 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire26
timestamp 1
transform -1 0 11316 0 1 4352
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 addr0[0]
port 0 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 addr0[1]
port 1 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 addr0[2]
port 2 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 addr0[3]
port 3 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 addr0[4]
port 4 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 addr0[5]
port 5 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 addr0[6]
port 6 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 clk0
port 7 nsew signal input
flabel metal3 s 17714 6808 18514 6928 0 FreeSans 480 0 0 0 cs0
port 8 nsew signal input
flabel metal3 s 17714 8848 18514 8968 0 FreeSans 480 0 0 0 dout0[0]
port 9 nsew signal output
flabel metal3 s 17714 14968 18514 15088 0 FreeSans 480 0 0 0 dout0[10]
port 10 nsew signal output
flabel metal3 s 17714 12928 18514 13048 0 FreeSans 480 0 0 0 dout0[11]
port 11 nsew signal output
flabel metal3 s 17714 9528 18514 9648 0 FreeSans 480 0 0 0 dout0[12]
port 12 nsew signal output
flabel metal3 s 17714 6128 18514 6248 0 FreeSans 480 0 0 0 dout0[13]
port 13 nsew signal output
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 dout0[14]
port 14 nsew signal output
flabel metal3 s 17714 5448 18514 5568 0 FreeSans 480 0 0 0 dout0[15]
port 15 nsew signal output
flabel metal2 s 12898 19858 12954 20658 0 FreeSans 224 90 0 0 dout0[1]
port 16 nsew signal output
flabel metal3 s 17714 10888 18514 11008 0 FreeSans 480 0 0 0 dout0[2]
port 17 nsew signal output
flabel metal3 s 17714 13608 18514 13728 0 FreeSans 480 0 0 0 dout0[3]
port 18 nsew signal output
flabel metal2 s 13542 19858 13598 20658 0 FreeSans 224 90 0 0 dout0[4]
port 19 nsew signal output
flabel metal3 s 17714 16328 18514 16448 0 FreeSans 480 0 0 0 dout0[5]
port 20 nsew signal output
flabel metal3 s 17714 11568 18514 11688 0 FreeSans 480 0 0 0 dout0[6]
port 21 nsew signal output
flabel metal3 s 17714 8168 18514 8288 0 FreeSans 480 0 0 0 dout0[7]
port 22 nsew signal output
flabel metal3 s 17714 15648 18514 15768 0 FreeSans 480 0 0 0 dout0[8]
port 23 nsew signal output
flabel metal3 s 17714 7488 18514 7608 0 FreeSans 480 0 0 0 dout0[9]
port 24 nsew signal output
flabel metal4 s 4208 2128 4528 18000 0 FreeSans 1920 90 0 0 vccd1
port 25 nsew power bidirectional
flabel metal4 s 4868 2128 5188 18000 0 FreeSans 1920 90 0 0 vssd1
port 26 nsew ground bidirectional
rlabel metal1 9246 17952 9246 17952 0 vccd1
rlabel metal1 9246 17408 9246 17408 0 vssd1
rlabel metal1 15762 5610 15762 5610 0 _000_
rlabel metal2 12558 16966 12558 16966 0 _001_
rlabel metal1 15762 11050 15762 11050 0 _002_
rlabel metal2 15686 14178 15686 14178 0 _003_
rlabel metal2 13662 16694 13662 16694 0 _004_
rlabel metal1 15394 16490 15394 16490 0 _005_
rlabel metal1 15762 12138 15762 12138 0 _006_
rlabel metal1 15860 7854 15860 7854 0 _007_
rlabel metal1 14756 16082 14756 16082 0 _008_
rlabel metal2 15778 6562 15778 6562 0 _009_
rlabel metal2 15778 15266 15778 15266 0 _010_
rlabel metal1 15931 13192 15931 13192 0 _011_
rlabel metal2 16146 9350 16146 9350 0 _012_
rlabel metal1 15762 4522 15762 4522 0 _013_
rlabel metal1 14214 2618 14214 2618 0 _014_
rlabel metal1 14750 3434 14750 3434 0 _015_
rlabel metal1 10948 12818 10948 12818 0 _016_
rlabel metal2 10442 15300 10442 15300 0 _017_
rlabel metal1 11914 12274 11914 12274 0 _018_
rlabel metal1 7774 15674 7774 15674 0 _019_
rlabel metal2 14674 11118 14674 11118 0 _020_
rlabel metal2 13018 9826 13018 9826 0 _021_
rlabel via1 12834 10421 12834 10421 0 _022_
rlabel metal1 13662 9894 13662 9894 0 _023_
rlabel metal1 11270 9962 11270 9962 0 _024_
rlabel metal1 13892 8942 13892 8942 0 _025_
rlabel metal1 14628 9146 14628 9146 0 _026_
rlabel metal2 14766 5916 14766 5916 0 _027_
rlabel metal1 8372 5678 8372 5678 0 _028_
rlabel metal1 7130 5678 7130 5678 0 _029_
rlabel metal1 13570 5610 13570 5610 0 _030_
rlabel metal1 9338 9554 9338 9554 0 _031_
rlabel metal1 13938 6256 13938 6256 0 _032_
rlabel metal2 13662 6358 13662 6358 0 _033_
rlabel metal1 13616 10574 13616 10574 0 _034_
rlabel metal1 13524 14994 13524 14994 0 _035_
rlabel metal1 4278 10744 4278 10744 0 _036_
rlabel metal1 7360 9146 7360 9146 0 _037_
rlabel metal1 4324 10506 4324 10506 0 _038_
rlabel metal1 6900 13294 6900 13294 0 _039_
rlabel metal1 10074 13906 10074 13906 0 _040_
rlabel metal1 13432 9554 13432 9554 0 _041_
rlabel metal1 14720 13906 14720 13906 0 _042_
rlabel metal1 11638 15470 11638 15470 0 _043_
rlabel metal1 12466 6936 12466 6936 0 _044_
rlabel metal2 12282 6052 12282 6052 0 _045_
rlabel metal2 8694 8296 8694 8296 0 _046_
rlabel metal1 11362 16150 11362 16150 0 _047_
rlabel metal2 13478 10846 13478 10846 0 _048_
rlabel metal1 13616 6834 13616 6834 0 _049_
rlabel metal2 11178 15334 11178 15334 0 _050_
rlabel metal2 7038 13770 7038 13770 0 _051_
rlabel metal2 8234 14586 8234 14586 0 _052_
rlabel metal1 6578 14960 6578 14960 0 _053_
rlabel metal1 12880 12274 12880 12274 0 _054_
rlabel metal1 13570 6698 13570 6698 0 _055_
rlabel metal1 13570 4590 13570 4590 0 _056_
rlabel metal1 8188 4590 8188 4590 0 _057_
rlabel metal1 7222 4624 7222 4624 0 _058_
rlabel metal1 9936 8942 9936 8942 0 _059_
rlabel metal1 8786 9554 8786 9554 0 _060_
rlabel metal1 12558 5236 12558 5236 0 _061_
rlabel via1 6298 5678 6298 5678 0 _062_
rlabel metal2 6394 5882 6394 5882 0 _063_
rlabel metal2 12742 5423 12742 5423 0 _064_
rlabel metal2 13754 4794 13754 4794 0 _065_
rlabel metal1 13938 14960 13938 14960 0 _066_
rlabel metal2 13570 5729 13570 5729 0 _067_
rlabel metal1 10764 4114 10764 4114 0 _068_
rlabel metal1 9936 10098 9936 10098 0 _069_
rlabel metal2 12098 5270 12098 5270 0 _070_
rlabel metal1 11316 4182 11316 4182 0 _071_
rlabel metal2 14122 14943 14122 14943 0 _072_
rlabel metal1 9384 11798 9384 11798 0 _073_
rlabel metal1 11638 10642 11638 10642 0 _074_
rlabel metal1 12696 15674 12696 15674 0 _075_
rlabel metal1 13478 4012 13478 4012 0 _076_
rlabel via2 6670 14909 6670 14909 0 _077_
rlabel metal2 6854 14790 6854 14790 0 _078_
rlabel metal1 5842 15436 5842 15436 0 _079_
rlabel metal1 11362 15436 11362 15436 0 _080_
rlabel metal1 12949 14586 12949 14586 0 _081_
rlabel metal1 9890 13362 9890 13362 0 _082_
rlabel metal2 10902 4386 10902 4386 0 _083_
rlabel metal1 14214 2414 14214 2414 0 _084_
rlabel via1 15410 15045 15410 15045 0 _085_
rlabel metal1 6348 12138 6348 12138 0 _086_
rlabel metal1 12006 5882 12006 5882 0 _087_
rlabel metal1 11454 5780 11454 5780 0 _088_
rlabel metal1 11224 13838 11224 13838 0 _089_
rlabel metal1 9568 4794 9568 4794 0 _090_
rlabel metal1 10396 5338 10396 5338 0 _091_
rlabel metal1 11362 5576 11362 5576 0 _092_
rlabel metal1 14214 5576 14214 5576 0 _093_
rlabel metal1 12466 10234 12466 10234 0 _094_
rlabel metal1 13018 11322 13018 11322 0 _095_
rlabel metal2 12558 13634 12558 13634 0 _096_
rlabel metal2 13018 13940 13018 13940 0 _097_
rlabel metal1 11454 14450 11454 14450 0 _098_
rlabel metal1 10626 14586 10626 14586 0 _099_
rlabel metal1 10166 9622 10166 9622 0 _100_
rlabel metal1 10902 9486 10902 9486 0 _101_
rlabel metal2 11454 7684 11454 7684 0 _102_
rlabel metal1 10396 14382 10396 14382 0 _103_
rlabel metal1 12052 14586 12052 14586 0 _104_
rlabel metal1 10350 9486 10350 9486 0 _105_
rlabel metal1 11454 14518 11454 14518 0 _106_
rlabel metal1 12880 14518 12880 14518 0 _107_
rlabel metal1 11454 8262 11454 8262 0 _108_
rlabel metal1 10948 7514 10948 7514 0 _109_
rlabel metal1 11638 8058 11638 8058 0 _110_
rlabel metal2 14398 10268 14398 10268 0 _111_
rlabel metal2 14214 13583 14214 13583 0 _112_
rlabel metal2 14122 6290 14122 6290 0 _113_
rlabel metal1 14536 11662 14536 11662 0 _114_
rlabel metal1 11316 13906 11316 13906 0 _115_
rlabel metal1 9706 12172 9706 12172 0 _116_
rlabel metal2 14490 11849 14490 11849 0 _117_
rlabel metal1 14996 11118 14996 11118 0 _118_
rlabel metal1 13432 14382 13432 14382 0 _119_
rlabel metal1 13892 13702 13892 13702 0 _120_
rlabel metal2 12466 13668 12466 13668 0 _121_
rlabel metal1 13846 10234 13846 10234 0 _122_
rlabel metal1 15134 13940 15134 13940 0 _123_
rlabel metal1 12650 15504 12650 15504 0 _124_
rlabel metal2 12282 15776 12282 15776 0 _125_
rlabel metal1 10258 16150 10258 16150 0 _126_
rlabel metal1 8924 13294 8924 13294 0 _127_
rlabel metal1 10304 8602 10304 8602 0 _128_
rlabel metal1 12834 6664 12834 6664 0 _129_
rlabel metal1 10212 14042 10212 14042 0 _130_
rlabel metal3 9913 15300 9913 15300 0 _131_
rlabel metal1 10810 15674 10810 15674 0 _132_
rlabel metal1 12834 16082 12834 16082 0 _133_
rlabel metal1 10810 10098 10810 10098 0 _134_
rlabel metal1 13662 11322 13662 11322 0 _135_
rlabel metal2 13754 11322 13754 11322 0 _136_
rlabel metal1 14444 13294 14444 13294 0 _137_
rlabel metal2 8050 13736 8050 13736 0 _138_
rlabel metal2 9338 13061 9338 13061 0 _139_
rlabel metal1 10212 12138 10212 12138 0 _140_
rlabel metal1 10902 12342 10902 12342 0 _141_
rlabel metal1 14536 12954 14536 12954 0 _142_
rlabel metal1 14766 11322 14766 11322 0 _143_
rlabel metal1 6486 12308 6486 12308 0 _144_
rlabel metal1 7038 13226 7038 13226 0 _145_
rlabel metal1 6716 12274 6716 12274 0 _146_
rlabel metal2 15042 11951 15042 11951 0 _147_
rlabel metal1 15272 11526 15272 11526 0 _148_
rlabel metal2 14398 7004 14398 7004 0 _149_
rlabel metal1 13018 10710 13018 10710 0 _150_
rlabel metal2 14582 10234 14582 10234 0 _151_
rlabel metal2 15042 8976 15042 8976 0 _152_
rlabel metal1 14950 6970 14950 6970 0 _153_
rlabel metal1 15318 8058 15318 8058 0 _154_
rlabel metal2 13294 13770 13294 13770 0 _155_
rlabel metal2 14306 14144 14306 14144 0 _156_
rlabel via2 12558 3723 12558 3723 0 _157_
rlabel metal1 13478 12954 13478 12954 0 _158_
rlabel metal1 14306 13430 14306 13430 0 _159_
rlabel metal2 9798 8670 9798 8670 0 _160_
rlabel metal2 12834 7582 12834 7582 0 _161_
rlabel metal1 12190 7276 12190 7276 0 _162_
rlabel metal1 11868 6970 11868 6970 0 _163_
rlabel metal1 12650 7480 12650 7480 0 _164_
rlabel metal1 15226 6324 15226 6324 0 _165_
rlabel metal1 9246 14994 9246 14994 0 _166_
rlabel metal1 14214 14824 14214 14824 0 _167_
rlabel metal1 13202 15096 13202 15096 0 _168_
rlabel metal1 14214 15028 14214 15028 0 _169_
rlabel metal1 14904 14994 14904 14994 0 _170_
rlabel metal1 10258 15912 10258 15912 0 _171_
rlabel metal1 10028 13498 10028 13498 0 _172_
rlabel metal2 8326 15878 8326 15878 0 _173_
rlabel metal1 14490 13940 14490 13940 0 _174_
rlabel metal2 15042 13498 15042 13498 0 _175_
rlabel metal2 13018 8738 13018 8738 0 _176_
rlabel metal1 13846 9146 13846 9146 0 _177_
rlabel metal1 15272 8942 15272 8942 0 _178_
rlabel metal1 13984 8466 13984 8466 0 _179_
rlabel metal1 13984 4590 13984 4590 0 _180_
rlabel metal1 15042 4556 15042 4556 0 _181_
rlabel metal1 16376 3706 16376 3706 0 _182_
rlabel metal2 7682 4386 7682 4386 0 _183_
rlabel metal1 2714 12172 2714 12172 0 _184_
rlabel metal1 10442 4080 10442 4080 0 _185_
rlabel metal1 6624 4250 6624 4250 0 _186_
rlabel metal1 2944 8806 2944 8806 0 _187_
rlabel metal1 10258 13294 10258 13294 0 _188_
rlabel metal1 6118 9894 6118 9894 0 _189_
rlabel metal1 5750 9962 5750 9962 0 _190_
rlabel metal1 5244 13906 5244 13906 0 _191_
rlabel metal1 6808 4114 6808 4114 0 _192_
rlabel via1 13478 8398 13478 8398 0 _193_
rlabel metal1 5060 8398 5060 8398 0 _194_
rlabel metal1 4324 8534 4324 8534 0 _195_
rlabel metal1 9844 9350 9844 9350 0 _196_
rlabel metal1 14214 11084 14214 11084 0 _197_
rlabel metal1 8602 13872 8602 13872 0 _198_
rlabel metal1 5522 5678 5522 5678 0 _199_
rlabel metal1 5842 5576 5842 5576 0 _200_
rlabel metal2 8418 14110 8418 14110 0 _201_
rlabel via1 12926 13141 12926 13141 0 _202_
rlabel metal2 9338 5729 9338 5729 0 _203_
rlabel metal1 4876 5270 4876 5270 0 _204_
rlabel via2 8510 5219 8510 5219 0 _205_
rlabel metal1 8096 7854 8096 7854 0 _206_
rlabel metal1 9246 5134 9246 5134 0 _207_
rlabel metal1 8786 5202 8786 5202 0 _208_
rlabel metal2 13294 6460 13294 6460 0 _209_
rlabel metal1 13984 7854 13984 7854 0 _210_
rlabel metal2 8970 14263 8970 14263 0 _211_
rlabel metal1 9568 6698 9568 6698 0 _212_
rlabel metal1 14030 8398 14030 8398 0 _213_
rlabel metal1 6118 5712 6118 5712 0 _214_
rlabel metal1 6946 8976 6946 8976 0 _215_
rlabel metal2 6762 8738 6762 8738 0 _216_
rlabel metal2 8970 8432 8970 8432 0 _217_
rlabel metal1 12696 14450 12696 14450 0 _218_
rlabel metal3 6417 13396 6417 13396 0 _219_
rlabel metal1 10166 7208 10166 7208 0 _220_
rlabel metal2 9982 8160 9982 8160 0 _221_
rlabel metal1 7682 6834 7682 6834 0 _222_
rlabel metal1 4462 6766 4462 6766 0 _223_
rlabel metal1 9752 14926 9752 14926 0 _224_
rlabel metal1 9982 7446 9982 7446 0 _225_
rlabel metal1 10442 7786 10442 7786 0 _226_
rlabel metal1 15134 7956 15134 7956 0 _227_
rlabel metal1 4048 13294 4048 13294 0 _228_
rlabel metal1 8004 13906 8004 13906 0 _229_
rlabel metal3 6578 12852 6578 12852 0 _230_
rlabel metal2 7314 12036 7314 12036 0 _231_
rlabel metal1 12558 13464 12558 13464 0 _232_
rlabel metal1 8234 8942 8234 8942 0 _233_
rlabel metal1 6302 12818 6302 12818 0 _234_
rlabel metal1 8648 12410 8648 12410 0 _235_
rlabel metal1 9154 11016 9154 11016 0 _236_
rlabel via1 8694 10438 8694 10438 0 _237_
rlabel metal2 9062 11934 9062 11934 0 _238_
rlabel metal1 13478 7888 13478 7888 0 _239_
rlabel metal1 10672 12818 10672 12818 0 _240_
rlabel metal3 1280 4148 1280 4148 0 addr0[0]
rlabel metal3 751 6188 751 6188 0 addr0[1]
rlabel metal3 1004 4828 1004 4828 0 addr0[2]
rlabel metal3 1280 5508 1280 5508 0 addr0[3]
rlabel metal2 10350 1588 10350 1588 0 addr0[4]
rlabel metal2 5842 1588 5842 1588 0 addr0[5]
rlabel metal2 9062 1588 9062 1588 0 addr0[6]
rlabel metal1 3036 4794 3036 4794 0 addr0_reg\[0\]
rlabel metal1 3312 7446 3312 7446 0 addr0_reg\[1\]
rlabel metal1 2944 5338 2944 5338 0 addr0_reg\[2\]
rlabel metal1 1978 7412 1978 7412 0 addr0_reg\[3\]
rlabel metal2 10166 4318 10166 4318 0 addr0_reg\[4\]
rlabel metal2 9154 3910 9154 3910 0 addr0_reg\[5\]
rlabel metal2 9982 3774 9982 3774 0 addr0_reg\[6\]
rlabel metal3 4638 17068 4638 17068 0 clk0
rlabel metal2 10350 9214 10350 9214 0 clknet_0_clk0
rlabel metal2 1426 3842 1426 3842 0 clknet_1_0__leaf_clk0
rlabel metal1 13386 17204 13386 17204 0 clknet_1_1__leaf_clk0
rlabel metal2 16146 7123 16146 7123 0 cs0
rlabel metal2 16974 8755 16974 8755 0 dout0[0]
rlabel metal2 16974 15079 16974 15079 0 dout0[10]
rlabel via2 16974 12971 16974 12971 0 dout0[11]
rlabel metal1 16560 9894 16560 9894 0 dout0[12]
rlabel via2 16974 6171 16974 6171 0 dout0[13]
rlabel metal2 13570 1520 13570 1520 0 dout0[14]
rlabel metal2 16974 5423 16974 5423 0 dout0[15]
rlabel metal1 13018 17850 13018 17850 0 dout0[1]
rlabel metal2 16974 10591 16974 10591 0 dout0[2]
rlabel via2 16974 13685 16974 13685 0 dout0[3]
rlabel metal1 13892 17850 13892 17850 0 dout0[4]
rlabel metal1 16744 16966 16744 16966 0 dout0[5]
rlabel metal1 17112 10778 17112 10778 0 dout0[6]
rlabel metal2 16974 7871 16974 7871 0 dout0[7]
rlabel metal2 16974 15793 16974 15793 0 dout0[8]
rlabel via2 16330 7531 16330 7531 0 dout0[9]
rlabel metal2 1702 4386 1702 4386 0 net1
rlabel metal1 16928 14994 16928 14994 0 net10
rlabel metal1 17112 12818 17112 12818 0 net11
rlabel metal2 16514 9180 16514 9180 0 net12
rlabel metal1 16928 4794 16928 4794 0 net13
rlabel metal1 14306 2482 14306 2482 0 net14
rlabel metal2 15778 4658 15778 4658 0 net15
rlabel metal2 13294 16796 13294 16796 0 net16
rlabel metal1 16560 10642 16560 10642 0 net17
rlabel metal2 16790 14076 16790 14076 0 net18
rlabel metal2 14766 17442 14766 17442 0 net19
rlabel metal1 1656 6426 1656 6426 0 net2
rlabel metal2 16790 16966 16790 16966 0 net20
rlabel metal1 16560 11730 16560 11730 0 net21
rlabel metal2 17066 8228 17066 8228 0 net22
rlabel metal1 15778 16218 15778 16218 0 net23
rlabel metal1 16790 6630 16790 6630 0 net24
rlabel metal1 15548 8874 15548 8874 0 net25
rlabel metal2 13570 4284 13570 4284 0 net26
rlabel via2 5014 8483 5014 8483 0 net27
rlabel metal1 7298 9350 7298 9350 0 net28
rlabel metal1 7038 9486 7038 9486 0 net29
rlabel metal1 1564 4250 1564 4250 0 net3
rlabel metal1 8004 10098 8004 10098 0 net30
rlabel metal2 2622 11832 2622 11832 0 net31
rlabel metal1 5152 13974 5152 13974 0 net32
rlabel metal1 7866 8976 7866 8976 0 net33
rlabel metal2 3450 14144 3450 14144 0 net34
rlabel metal1 7130 6834 7130 6834 0 net35
rlabel metal1 10074 4556 10074 4556 0 net36
rlabel metal2 8050 5287 8050 5287 0 net37
rlabel metal1 3404 12818 3404 12818 0 net38
rlabel metal2 8234 7905 8234 7905 0 net39
rlabel via1 1697 5678 1697 5678 0 net4
rlabel metal2 5382 7922 5382 7922 0 net40
rlabel metal2 3634 13056 3634 13056 0 net41
rlabel metal1 7682 12818 7682 12818 0 net42
rlabel metal1 7222 10030 7222 10030 0 net43
rlabel metal1 5612 8942 5612 8942 0 net44
rlabel metal1 8556 11050 8556 11050 0 net45
rlabel metal1 6670 5168 6670 5168 0 net46
rlabel metal1 11132 3434 11132 3434 0 net47
rlabel via1 2714 7973 2714 7973 0 net48
rlabel metal2 2714 9724 2714 9724 0 net49
rlabel metal1 10350 2618 10350 2618 0 net5
rlabel metal1 2254 7344 2254 7344 0 net50
rlabel metal1 2300 9690 2300 9690 0 net51
rlabel metal2 3450 8194 3450 8194 0 net52
rlabel metal2 2438 8738 2438 8738 0 net53
rlabel metal2 2714 7548 2714 7548 0 net54
rlabel metal2 2254 8738 2254 8738 0 net55
rlabel metal1 15410 13872 15410 13872 0 net56
rlabel metal1 15410 14994 15410 14994 0 net57
rlabel metal1 14628 2822 14628 2822 0 net58
rlabel metal1 15088 4114 15088 4114 0 net59
rlabel metal1 6302 2618 6302 2618 0 net6
rlabel metal1 15732 14994 15732 14994 0 net60
rlabel metal1 15686 13906 15686 13906 0 net61
rlabel metal2 15410 10948 15410 10948 0 net62
rlabel metal2 15410 12036 15410 12036 0 net63
rlabel metal2 15410 13124 15410 13124 0 net64
rlabel metal1 14996 16558 14996 16558 0 net65
rlabel metal1 15732 8466 15732 8466 0 net66
rlabel metal1 14306 16150 14306 16150 0 net67
rlabel metal1 16146 8942 16146 8942 0 net68
rlabel metal1 15732 6290 15732 6290 0 net69
rlabel metal1 8965 3026 8965 3026 0 net7
rlabel metal1 12880 16558 12880 16558 0 net70
rlabel metal2 15410 4420 15410 4420 0 net71
rlabel metal1 15594 5338 15594 5338 0 net72
rlabel metal1 13478 16116 13478 16116 0 net73
rlabel metal1 15410 2414 15410 2414 0 net8
rlabel metal1 16974 5882 16974 5882 0 net9
<< properties >>
string FIXED_BBOX 0 0 18514 20658
<< end >>
