* NGSPICE file created from cust_rom.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

.subckt cust_rom VGND VPWR addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6]
+ addr0[7] clk0 cs0 dout0[0] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15]
+ dout0[16] dout0[17] dout0[18] dout0[19] dout0[1] dout0[20] dout0[21] dout0[22] dout0[23]
+ dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[2] dout0[30] dout0[31]
+ dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9]
XTAP_TAPCELL_ROW_37_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1270_ _0539_ _0541_ _0546_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0985_ net116 net84 net82 net121 VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__a22o_2
X_1399_ net45 _0658_ _0666_ net165 net129 VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__o32a_1
Xfanout127 net128 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
Xfanout138 net4 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
Xfanout116 _0687_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__buf_2
XFILLER_0_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0770_ net135 net131 net133 net137 VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_59_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1253_ _0191_ _0193_ _0234_ _0405_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__or4_1
X_1322_ _0096_ _0193_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__or2_1
X_1184_ _0060_ _0228_ _0446_ _0466_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_19_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0968_ _0065_ _0259_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0899_ _0115_ _0185_ _0186_ _0187_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__or4_4
XFILLER_0_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0822_ net110 net92 net90 net100 VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__a22o_2
XFILLER_0_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0753_ _0040_ _0043_ _0044_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1236_ _0119_ _0199_ _0209_ _0514_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__or4_1
X_1305_ _0158_ _0576_ _0577_ _0578_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1167_ _0141_ _0205_ _0230_ _0248_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1098_ _0099_ _0102_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1021_ _0136_ _0142_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0805_ net84 net52 net49 net82 VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__a22o_4
X_0736_ net94 net92 net90 net96 VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__a22o_2
XFILLER_0_12_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1219_ _0166_ _0489_ _0497_ _0499_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold30 net23 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_5 _0097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1004_ _0069_ _0295_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__or2_2
XFILLER_0_44_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0719_ net124 net122 net120 net117 VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__a22o_2
XFILLER_0_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput20 net20 VGND VGND VPWR VPWR dout0[19] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput31 net31 VGND VGND VPWR VPWR dout0[29] sky130_fd_sc_hd__buf_2
XFILLER_0_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0984_ net122 net120 net117 net124 VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout128 net129 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_4
X_1398_ _0163_ _0659_ _0662_ _0665_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__or4_1
Xfanout139 net4 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__buf_1
Xfanout117 net118 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_49_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1252_ _0487_ _0489_ _0527_ _0529_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__or4_1
X_1321_ _0201_ _0231_ _0366_ _0548_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__or4_1
X_1183_ _0049_ _0389_ _0414_ _0459_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0967_ net60 net58 _0046_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0898_ _0185_ _0186_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__or2_2
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0752_ net84 net81 net78 net82 VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__a22o_2
XFILLER_0_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0821_ _0110_ net46 VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__or2_2
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1166_ _0069_ _0272_ _0297_ _0411_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__or4_1
X_1304_ _0165_ _0171_ _0219_ _0250_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__or4_1
X_1235_ _0090_ _0161_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1097_ net45 _0381_ _0384_ net151 net129 VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__o32a_1
XFILLER_0_30_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1020_ _0086_ _0310_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0804_ _0093_ _0094_ _0095_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__or3_1
X_0735_ net143 net141 net139 net145 VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1149_ net125 _0082_ _0431_ _0432_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1218_ _0068_ _0268_ _0307_ _0498_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold20 net28 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 net25 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_6 _0097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_7_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1003_ net68 net61 net58 net70 VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__a22o_2
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0718_ net136 net134 net130 net132 VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__nor4_1
XFILLER_0_57_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput32 net32 VGND VGND VPWR VPWR dout0[2] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_33_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput21 net21 VGND VGND VPWR VPWR dout0[1] sky130_fd_sc_hd__buf_2
Xoutput10 net10 VGND VGND VPWR VPWR dout0[0] sky130_fd_sc_hd__buf_2
XFILLER_0_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0983_ _0109_ _0274_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__or2_4
Xfanout129 net9 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1397_ _0430_ _0573_ _0663_ _0664_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1320_ _0074_ _0076_ _0221_ _0244_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__or4_1
X_1251_ _0069_ _0149_ _0297_ _0491_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__or4_1
X_1182_ _0252_ _0300_ _0406_ _0460_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_47_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0897_ _0115_ _0186_ _0187_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__or3_2
X_0966_ net114 net61 net58 net112 VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__a22o_2
XFILLER_0_27_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1449_ clknet_2_2__leaf_clk0 _0021_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_2_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0751_ net80 net69 net67 net78 VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__a22o_2
XFILLER_0_28_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0820_ _0702_ _0111_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1303_ _0180_ _0288_ _0305_ _0308_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1234_ _0107_ _0225_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__or2_1
X_1165_ _0149_ _0446_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__or2_1
X_1096_ _0370_ _0375_ _0382_ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0949_ _0239_ _0240_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0803_ net99 net60 net58 net103 VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__a22o_2
X_0734_ net145 net143 net141 net139 VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1079_ _0058_ _0171_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__or2_1
X_1148_ _0100_ _0194_ _0238_ _0314_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1217_ _0705_ _0711_ _0301_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__or3_1
XFILLER_0_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold21 net15 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 net24 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 net34 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_7 _0109_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1002_ _0696_ _0105_ _0290_ _0292_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_60_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0717_ net144 net140 net138 net142 VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_57_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput11 net11 VGND VGND VPWR VPWR dout0[10] sky130_fd_sc_hd__clkbuf_4
Xoutput22 net22 VGND VGND VPWR VPWR dout0[20] sky130_fd_sc_hd__buf_2
Xoutput33 net33 VGND VGND VPWR VPWR dout0[30] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0982_ net116 net69 net67 net121 VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__a22o_2
XFILLER_0_38_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout119 net120 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1396_ _0710_ _0131_ _0282_ _0285_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1181_ _0355_ _0457_ _0461_ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__or4_1
X_1250_ _0693_ _0221_ _0274_ _0285_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0896_ _0186_ _0187_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0965_ _0144_ _0216_ _0255_ _0256_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__or4_2
XFILLER_0_49_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1448_ clknet_2_3__leaf_clk0 _0020_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1379_ net43 _0643_ _0646_ net152 net127 VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_2_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0750_ net144 net142 net140 net138 VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__and4bb_1
Xfanout90 net91 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_2
X_1233_ _0094_ _0095_ _0261_ _0511_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__or4_1
X_1302_ _0101_ _0262_ _0574_ _0575_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1164_ _0057_ _0171_ _0246_ _0447_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__or4_1
X_1095_ _0240_ _0365_ _0368_ _0373_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__or4_1
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0948_ net80 net56 net54 net78 VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__a22o_2
XFILLER_0_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0879_ _0059_ _0170_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__or2_2
XFILLER_0_30_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0802_ net92 net60 net58 net90 VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__a22o_4
X_0733_ net104 net97 net95 net99 VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__a22o_2
XFILLER_0_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1216_ _0189_ _0371_ _0428_ _0490_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__or4_1
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1147_ _0140_ _0229_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__or2_1
X_1078_ _0189_ _0296_ _0297_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold22 net32 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 net22 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_8 _0167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ _0696_ _0292_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0716_ net130 net132 net136 net134 VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__and4b_1
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput12 net12 VGND VGND VPWR VPWR dout0[11] sky130_fd_sc_hd__buf_2
XFILLER_0_43_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput34 net34 VGND VGND VPWR VPWR dout0[31] sky130_fd_sc_hd__buf_2
XFILLER_0_31_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput23 net23 VGND VGND VPWR VPWR dout0[21] sky130_fd_sc_hd__buf_2
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0981_ _0093_ _0094_ _0095_ _0270_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__or4_2
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1395_ _0705_ _0203_ _0275_ _0277_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1180_ _0053_ _0275_ _0462_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__or3_1
XFILLER_0_54_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0964_ _0218_ _0224_ _0228_ _0231_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0895_ net119 net110 net100 net123 VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1447_ clknet_2_1__leaf_clk0 _0019_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1378_ _0425_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout80 _0038_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_2
Xfanout91 _0709_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
XFILLER_0_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1232_ _0693_ _0696_ _0130_ _0192_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__or4_1
X_1301_ _0076_ _0090_ _0181_ _0264_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__or4_1
X_1094_ _0169_ _0206_ _0371_ _0374_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__or4_1
X_1163_ net125 _0693_ _0073_ _0329_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__or4_1
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0947_ net103 net80 net78 net98 VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_15_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0878_ net67 net64 net62 net69 VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload0 clknet_2_0__leaf_clk0 VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_33_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0801_ net121 net58 _0702_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_21_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0732_ net136 net134 net130 net132 VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__and4b_1
X_1146_ _0707_ _0118_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1215_ _0235_ _0492_ _0494_ _0495_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_63_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1077_ _0236_ _0239_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__or2_1
Xhold12 net12 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 net10 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_9 _0167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1000_ net122 net117 _0046_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__o21ba_2
XTAP_TAPCELL_ROW_60_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0715_ net144 net138 net140 net142 VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1129_ _0105_ _0259_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput35 net35 VGND VGND VPWR VPWR dout0[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput24 net24 VGND VGND VPWR VPWR dout0[22] sky130_fd_sc_hd__buf_2
Xoutput13 net13 VGND VGND VPWR VPWR dout0[12] sky130_fd_sc_hd__buf_2
XFILLER_0_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0980_ _0093_ _0270_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_42_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1394_ _0149_ _0326_ _0660_ _0661_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0894_ net100 net85 net83 net110 VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__a22o_2
X_0963_ _0235_ _0243_ _0247_ _0254_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1377_ _0200_ _0228_ _0231_ _0644_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__or4_2
X_1446_ clknet_2_3__leaf_clk0 _0018_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout81 _0038_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout70 net73 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_2
Xfanout92 net93 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_24_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1162_ _0185_ _0186_ _0187_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__or3_2
X_1231_ net44 _0509_ _0510_ net154 net128 VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__o32a_1
X_1300_ _0088_ _0125_ _0134_ _0225_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1093_ _0377_ _0378_ _0379_ _0380_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_15_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0946_ _0236_ _0237_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__or2_1
X_0877_ _0122_ _0164_ _0166_ _0167_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__or4_1
XFILLER_0_55_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1429_ clknet_2_2__leaf_clk0 _0001_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_58_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload1 clknet_2_1__leaf_clk0 VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire105 _0698_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0800_ _0088_ _0089_ _0090_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__or3_1
X_0731_ _0701_ _0704_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1214_ _0049_ _0102_ _0270_ _0282_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__or4_1
X_1145_ _0064_ _0258_ _0259_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__or3_2
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1076_ net45 _0359_ _0364_ net169 net129 VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__o32a_1
XFILLER_0_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0929_ net123 net96 net94 net119 VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a22o_4
Xhold24 net35 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 net11 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0714_ net126 VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_27_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1059_ _0043_ _0220_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__or2_1
X_1128_ _0064_ _0068_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_11_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput36 net36 VGND VGND VPWR VPWR dout0[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput14 net14 VGND VGND VPWR VPWR dout0[13] sky130_fd_sc_hd__buf_2
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput25 net25 VGND VGND VPWR VPWR dout0[23] sky130_fd_sc_hd__buf_2
XFILLER_0_34_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1393_ _0102_ _0103_ _0241_ _0308_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__or4_1
XFILLER_0_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0893_ net110 net100 _0046_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__o21ba_1
X_0962_ _0117_ _0248_ _0249_ _0250_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1445_ clknet_2_2__leaf_clk0 _0017_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1376_ _0094_ _0137_ _0142_ _0270_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout93 _0708_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_2
Xfanout60 _0061_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout82 net83 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_4
X_1230_ _0306_ _0407_ _0445_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__or3_1
X_1092_ _0710_ _0121_ _0142_ _0250_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__or4_1
X_1161_ _0056_ _0065_ _0263_ _0444_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__or4_2
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0876_ _0166_ _0167_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__or2_1
X_0945_ net86 net80 _0702_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1428_ clknet_2_2__leaf_clk0 _0000_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfxtp_1
X_1359_ _0079_ _0159_ _0279_ _0617_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__or4_1
Xclkload2 clknet_2_3__leaf_clk0 VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire106 net107 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_29_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0730_ net111 net96 _0702_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1213_ _0288_ _0291_ _0493_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_63_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1075_ _0360_ _0361_ _0362_ _0363_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__or4_1
X_1144_ _0064_ _0258_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0928_ _0040_ _0219_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__or2_1
X_0859_ _0108_ _0115_ _0117_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold25 net30 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 net18 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1058_ _0711_ _0244_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__or2_1
X_1127_ _0137_ _0412_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_23_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput15 net15 VGND VGND VPWR VPWR dout0[14] sky130_fd_sc_hd__buf_2
Xoutput26 net26 VGND VGND VPWR VPWR dout0[24] sky130_fd_sc_hd__buf_2
Xoutput37 net37 VGND VGND VPWR VPWR dout0[5] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1392_ _0209_ _0230_ _0281_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0961_ _0117_ _0248_ _0249_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__or3_2
XFILLER_0_39_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0892_ _0079_ _0159_ _0173_ _0183_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1444_ clknet_2_3__leaf_clk0 _0016_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfxtp_1
X_1375_ _0526_ _0639_ _0641_ _0642_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout61 _0061_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout83 _0035_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_2
Xfanout94 _0706_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout50 net51 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1160_ _0040_ _0208_ _0210_ _0213_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__or4_1
X_1091_ _0076_ _0110_ _0178_ _0210_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0944_ net90 net80 net78 net92 VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__a22o_2
XFILLER_0_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0875_ net63 net56 net54 net64 VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1358_ _0234_ _0242_ _0458_ _0626_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__or4_1
X_1427_ _0647_ _0207_ _0257_ _0692_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__o31a_1
X_1289_ _0096_ _0243_ _0514_ _0563_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire107 net108 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_29_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1212_ _0040_ _0123_ _0212_ _0236_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1143_ _0181_ _0404_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__or2_1
X_1074_ _0068_ _0093_ _0104_ _0211_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0927_ net123 net81 net79 net119 VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0858_ _0705_ _0065_ _0113_ _0149_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__or4_1
X_0789_ net92 net80 net78 net91 VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__a22o_2
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold26 net16 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 net38 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1126_ _0136_ _0140_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1057_ net129 net167 net45 _0346_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_23_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput16 net16 VGND VGND VPWR VPWR dout0[15] sky130_fd_sc_hd__clkbuf_4
Xoutput38 net38 VGND VGND VPWR VPWR dout0[6] sky130_fd_sc_hd__buf_2
Xoutput27 net27 VGND VGND VPWR VPWR dout0[25] sky130_fd_sc_hd__buf_2
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_3__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_39_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ _0055_ _0253_ _0262_ _0332_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_36_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1391_ _0226_ _0473_ _0603_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_35_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0960_ _0117_ _0249_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0891_ _0177_ _0180_ _0182_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1443_ clknet_2_1__leaf_clk0 _0015_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfxtp_1
X_1374_ _0560_ _0605_ _0636_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_18_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout62 _0048_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout95 _0706_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout84 net85 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1090_ _0051_ _0065_ _0135_ _0271_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0943_ _0032_ _0033_ _0036_ _0232_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0874_ net63 net52 _0702_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__o21ba_4
XFILLER_0_15_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1426_ net126 net177 VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__or2_1
X_1357_ _0114_ _0122_ _0167_ _0197_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__or4_1
X_1288_ _0058_ _0129_ _0167_ _0202_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire108 net109 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1211_ _0469_ _0470_ _0487_ _0491_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__or4_1
X_1142_ _0052_ _0054_ _0162_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_63_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1073_ _0055_ _0079_ _0328_ _0356_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0926_ _0043_ _0044_ _0107_ _0217_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__or4_1
X_0857_ _0114_ _0121_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold16 net20 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold27 net33 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ _0201_ _0231_ _0273_ _0296_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__or4_1
X_0788_ net98 net80 net78 net103 VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__a22o_2
XFILLER_0_38_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1125_ _0232_ _0240_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__or2_1
X_1056_ _0331_ _0343_ _0345_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__or3_1
XFILLER_0_35_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput28 net28 VGND VGND VPWR VPWR dout0[26] sky130_fd_sc_hd__clkbuf_4
X_0909_ _0114_ _0121_ _0196_ _0197_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__or4_2
Xoutput17 net17 VGND VGND VPWR VPWR dout0[16] sky130_fd_sc_hd__buf_2
XFILLER_0_43_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput39 net39 VGND VGND VPWR VPWR dout0[7] sky130_fd_sc_hd__buf_2
XFILLER_0_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1108_ _0241_ _0386_ _0388_ _0391_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1039_ _0102_ _0103_ _0156_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__or3_1
XFILLER_0_63_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1390_ _0166_ _0489_ _0592_ _0656_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0890_ _0120_ _0181_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1442_ clknet_2_0__leaf_clk0 _0014_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfxtp_1
X_1373_ _0162_ _0203_ _0305_ _0640_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_18_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout63 _0048_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_2
Xfanout85 _0034_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_2
Xfanout96 _0703_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_4
Xfanout52 _0070_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_63_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0873_ _0122_ _0164_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__or2_1
X_0942_ _0032_ _0036_ _0232_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1425_ net126 net172 net42 _0691_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1356_ net128 net155 net44 _0625_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__o22a_1
X_1287_ _0275_ _0277_ _0559_ _0560_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1210_ net125 _0118_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__or2_2
X_1141_ _0221_ _0222_ _0244_ _0245_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__or4_1
X_1072_ _0347_ _0348_ _0355_ _0357_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0787_ _0075_ _0078_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__or2_2
X_0925_ net96 net94 _0046_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__o21ba_2
X_0856_ _0693_ _0696_ _0144_ _0147_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold28 net40 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold17 net31 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ net126 net146 net42 _0675_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__o22a_1
X_1339_ _0200_ _0385_ _0404_ _0412_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_26_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1055_ _0325_ _0334_ _0338_ _0344_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__or4_1
X_1124_ _0406_ _0407_ _0408_ _0409_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0908_ _0196_ _0197_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0839_ net114 net111 net101 net112 VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__a22o_2
Xoutput29 net29 VGND VGND VPWR VPWR dout0[27] sky130_fd_sc_hd__buf_2
XFILLER_0_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput18 net18 VGND VGND VPWR VPWR dout0[17] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_39_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1107_ _0208_ _0222_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__or2_1
X_1038_ _0089_ _0133_ _0141_ _0160_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_36_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1441_ clknet_2_3__leaf_clk0 _0013_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1372_ _0693_ _0052_ _0063_ _0104_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout86 _0713_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_2
Xfanout64 _0047_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_4
Xfanout42 net43 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
Xfanout97 _0703_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
Xfanout53 _0070_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_32_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0941_ _0032_ _0232_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0872_ net93 net64 net63 net91 VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__a22o_4
X_1355_ _0331_ _0619_ _0621_ _0624_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__or4_1
X_1424_ _0184_ _0207_ _0690_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__or3_1
X_1286_ net125 _0044_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1140_ _0252_ _0267_ _0424_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__or3_1
X_1071_ _0126_ _0286_ _0291_ _0358_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0924_ _0211_ _0213_ _0215_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0786_ _0072_ _0076_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0855_ _0068_ _0069_ _0118_ _0119_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold18 net41 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 net14 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__dlygate4sd3_1
X_1338_ _0097_ _0156_ _0416_ _0603_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__or4_1
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1407_ _0668_ _0671_ _0672_ _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__or4_1
X_1269_ _0337_ _0542_ _0543_ _0545_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_60_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1123_ _0696_ _0052_ _0054_ _0281_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__or4_1
X_1054_ _0326_ _0335_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__or2_1
X_0907_ _0197_ _0198_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput19 net19 VGND VGND VPWR VPWR dout0[18] sky130_fd_sc_hd__buf_2
X_0838_ net111 net70 net68 net101 VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__a22o_2
XFILLER_0_31_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0769_ net137 net131 net133 net135 VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1106_ _0198_ _0233_ _0296_ _0298_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__or4_1
XFILLER_0_63_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1037_ _0133_ _0141_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1440_ clknet_2_0__leaf_clk0 _0012_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfxtp_1
X_1371_ _0215_ _0308_ _0637_ _0638_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout65 net66 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout87 _0713_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_2
Xfanout98 _0700_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_2
Xfanout43 net44 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
Xfanout54 _0067_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0940_ net88 net69 net67 net86 VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0871_ _0056_ _0162_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__or2_1
X_1354_ _0175_ _0367_ _0622_ _0623_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__or4_1
X_1423_ _0108_ _0247_ _0269_ _0299_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__or4_1
X_1285_ _0098_ _0174_ _0473_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1070_ _0311_ _0351_ _0354_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0923_ net46 _0214_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0854_ _0037_ _0084_ _0101_ _0145_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0785_ _0075_ _0076_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1268_ _0431_ _0474_ _0475_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__or4_1
Xhold19 net19 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dlygate4sd3_1
X_1406_ _0226_ _0296_ _0308_ _0673_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__or4_1
X_1337_ _0514_ _0607_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__or2_1
X_1199_ _0476_ _0477_ _0480_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1122_ _0116_ _0251_ _0295_ _0299_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1053_ _0337_ _0340_ _0341_ _0342_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0906_ _0121_ _0196_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0837_ net124 net111 net101 net120 VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__a22o_2
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0768_ _0057_ _0058_ _0059_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__or3_2
XFILLER_0_47_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap51 _0071_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1105_ _0284_ _0290_ _0292_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__or3_1
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1036_ _0105_ _0179_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1019_ _0109_ _0274_ _0276_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__or3_1
XFILLER_0_63_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1370_ _0033_ _0036_ _0044_ _0222_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__or4_1
XFILLER_0_58_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout44 net45 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
Xfanout55 _0067_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout88 _0712_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
XFILLER_0_17_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout99 _0700_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0870_ _0088_ _0089_ _0090_ _0160_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__or4_2
XFILLER_0_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1422_ _0173_ net42 _0689_ net162 net126 VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__o32a_1
XPHY_EDGE_ROW_50_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1353_ _0081_ _0160_ _0196_ _0292_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__or4_1
X_1284_ _0075_ _0081_ _0082_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0999_ _0105_ _0290_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0922_ net96 net92 net90 net94 VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__a22o_2
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0853_ _0045_ _0060_ _0092_ _0106_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__or4_1
X_1405_ _0127_ _0188_ _0213_ _0275_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__or4_1
X_0784_ net93 net52 net49 net91 VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__a22o_2
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1267_ _0114_ _0130_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__or2_1
X_1198_ _0299_ _0478_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__or3_1
X_1336_ _0573_ _0602_ _0604_ _0605_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__or4_1
Xinput1 addr0[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1121_ _0274_ _0278_ _0286_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__or3_1
X_1052_ _0078_ _0176_ _0190_ _0227_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0836_ _0124_ _0127_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__or2_1
X_0767_ net113 net65 net62 net115 VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0905_ net103 net100 net98 net110 VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__a22o_2
XFILLER_0_28_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1319_ net129 net161 net45 _0591_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1035_ _0068_ _0253_ _0268_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__or3_1
X_1104_ _0236_ _0390_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_44_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0819_ net137 net135 net131 VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1018_ _0217_ _0244_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout89 _0712_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout67 _0042_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_4
Xfanout45 _0304_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_4
Xfanout78 _0039_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_2
Xfanout56 _0066_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1421_ _0072_ _0201_ _0216_ _0688_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__or4_1
X_1352_ _0107_ _0141_ _0142_ _0217_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__or4_1
X_1283_ net127 net153 net43 _0558_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0998_ net122 net57 net55 net116 VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__a22o_2
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0921_ _0110_ _0212_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_23_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0852_ _0138_ _0143_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__or2_1
X_0783_ net48 _0074_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__or2_2
X_1335_ _0710_ _0080_ _0123_ _0187_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__or4_1
X_1404_ _0177_ _0386_ _0604_ _0626_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__or4_1
X_1266_ _0113_ _0205_ _0290_ _0297_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__or4_1
X_1197_ _0051_ _0170_ _0194_ _0210_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput2 addr0[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_62_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1051_ _0261_ _0278_ _0288_ _0293_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__or4_1
X_1120_ _0209_ _0210_ _0405_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__or3_1
X_0904_ net100 net69 net67 net110 VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__a22o_2
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0835_ _0123_ _0125_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0766_ net83 net64 net62 net85 VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__a22o_4
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1318_ _0586_ _0587_ _0590_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1249_ _0040_ _0094_ _0272_ _0389_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_39_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1103_ _0043_ _0044_ _0219_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_36_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1034_ net126 net148 net42 _0324_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_44_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0818_ net95 net57 net55 net97 VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_10_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0749_ net144 net142 net138 net140 VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_54_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1017_ net125 _0043_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__or2_2
XFILLER_0_48_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout79 _0039_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_1
Xfanout68 _0042_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_2
Xfanout57 _0066_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1351_ _0408_ _0617_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__or3_1
X_1420_ _0183_ _0684_ _0685_ _0686_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__or4_1
X_1282_ _0549_ _0551_ _0552_ _0557_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0997_ _0085_ _0284_ _0288_ _0287_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__or4b_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0920_ net98 net96 net94 net103 VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0851_ _0139_ _0140_ _0141_ _0142_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0782_ net99 net53 net50 net104 VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__a22o_2
X_1265_ _0295_ _0327_ _0411_ _0412_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__or4_1
X_1403_ _0172_ _0243_ _0670_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__or3_1
X_1334_ _0087_ _0109_ _0277_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1196_ _0696_ _0074_ _0181_ _0201_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 addr0[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1050_ _0194_ _0205_ _0328_ _0339_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_38_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0834_ _0124_ _0125_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__or2_1
X_0903_ _0129_ _0191_ _0193_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0765_ net119 net65 net62 net123 VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__a22o_2
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1317_ _0083_ _0351_ _0588_ _0589_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_39_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1248_ _0240_ _0245_ _0501_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1179_ _0033_ _0098_ _0157_ _0167_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_30 _0244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1102_ _0044_ _0219_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__or2_2
XFILLER_0_17_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1033_ _0306_ _0315_ _0316_ _0323_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_36_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0817_ net117 net114 net112 net121 VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__a22o_2
X_0748_ net114 net81 net79 net112 VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__a22o_2
XFILLER_0_62_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1016_ _0097_ _0099_ _0198_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout69 net71 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_4
Xfanout58 net59 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_9_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1350_ _0072_ _0074_ _0365_ _0561_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__or4_1
X_1281_ _0370_ _0553_ _0554_ _0556_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0996_ _0086_ _0285_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__or2_2
XFILLER_0_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0850_ net119 net88 net86 net123 VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_11_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1402_ _0711_ _0208_ _0248_ _0669_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0781_ net136 net131 _0702_ net134 VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__nor4b_2
X_1264_ _0373_ _0405_ _0430_ _0540_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1333_ _0065_ _0258_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__or2_1
Xinput4 addr0[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_1195_ _0045_ _0128_ _0260_ _0373_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0979_ _0095_ _0270_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0902_ _0129_ _0192_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__or2_2
X_0833_ net112 net81 net79 net114 VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0764_ _0049_ _0050_ _0052_ _0053_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__or4_2
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1316_ _0043_ _0044_ _0209_ _0327_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1178_ _0705_ _0203_ _0458_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__or3_1
X_1247_ _0701_ _0202_ _0203_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_20 _0295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap66 _0047_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
Xmax_cap77 _0041_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1032_ _0317_ _0319_ _0321_ _0322_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1101_ _0109_ _0276_ _0288_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__or3_2
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0816_ net125 _0107_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__or2_2
XFILLER_0_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0747_ net136 net132 net130 net134 VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_12_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1015_ _0193_ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout59 _0062_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1280_ _0069_ _0074_ _0093_ _0555_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0995_ net136 net134 net133 _0702_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0780_ net55 net52 net49 net57 VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_11_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1401_ _0085_ _0157_ _0263_ _0270_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1194_ _0246_ _0457_ _0471_ _0472_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__or4_1
X_1332_ _0095_ _0264_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput5 addr0[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_1263_ _0158_ _0286_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0978_ net58 net56 net54 net60 VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__a22o_2
XFILLER_0_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0832_ net81 net79 _0046_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__o21ba_2
X_0901_ _0130_ _0131_ _0192_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__or3_2
X_0763_ _0049_ _0050_ _0053_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__or3_1
X_1315_ _0299_ _0387_ _0424_ _0513_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1177_ net125 _0133_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__or2_1
X_1246_ net44 _0519_ _0524_ net174 net128 VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__o32a_1
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_21 _0516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 _0167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1100_ _0068_ _0072_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_36_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1031_ _0135_ _0232_ _0284_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_44_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0815_ net115 net96 net94 net113 VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__a22o_2
X_0746_ net134 net130 net132 net136 VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__and4b_1
XFILLER_0_24_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1229_ _0504_ _0506_ _0508_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__or3_1
XFILLER_0_39_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_2__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_2__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1014_ _0704_ _0202_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_14_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0729_ net134 net132 net130 net136 VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_55_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout49 _0071_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0994_ _0085_ _0285_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__or2_2
XFILLER_0_49_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1331_ _0647_ _0251_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__or2_1
X_1400_ _0077_ _0163_ _0370_ _0392_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1193_ _0058_ _0122_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__or2_1
X_1262_ _0527_ _0535_ _0538_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__or3_1
Xinput6 addr0[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0977_ _0262_ _0265_ _0268_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ net111 net84 net82 net101 VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0831_ net119 net81 net79 net123 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0762_ _0050_ _0053_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__or2_2
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1314_ _0175_ _0354_ _0430_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1245_ _0515_ _0520_ _0523_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__or3_2
X_1176_ _0086_ _0094_ _0280_ _0282_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_11 _0196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_22 _0578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap46 _0112_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_1
X_1030_ _0052_ _0103_ _0170_ _0320_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0814_ _0102_ _0103_ _0104_ _0105_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__or4_1
XFILLER_0_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0745_ _0032_ _0033_ _0036_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1228_ _0336_ _0470_ _0501_ _0507_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1159_ _0117_ _0137_ _0217_ _0221_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__or4_1
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1013_ _0154_ _0155_ net42 net126 net168 VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__o32a_1
XFILLER_0_60_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0728_ net145 net143 net141 net139 VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__or4_4
XFILLER_0_62_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0993_ net116 net104 net99 net121 VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__a22o_2
XFILLER_0_41_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1261_ _0189_ _0228_ _0536_ _0537_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__or4_1
X_1330_ net127 net156 net43 _0601_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__o22a_1
X_1192_ _0107_ _0250_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__or2_1
Xinput7 addr0[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_62_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0976_ _0263_ _0266_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__or2_2
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1459_ clknet_2_2__leaf_clk0 _0031_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0830_ net98 net64 net63 net103 VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__a22o_2
XFILLER_0_28_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0761_ net85 net64 net62 net83 VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1244_ _0188_ _0231_ _0521_ _0522_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__or4_1
X_1313_ _0056_ _0243_ _0583_ _0585_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1175_ _0107_ _0217_ _0222_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__or3_1
X_0959_ _0117_ _0250_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_30_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_12 _0216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _0611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap47 net48 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0813_ net122 net70 net68 net116 VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__a22o_2
XFILLER_0_58_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0744_ net89 net84 net82 net87 VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1227_ _0116_ _0161_ _0300_ _0349_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__or4_1
X_1158_ net127 net147 net42 _0442_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1089_ _0126_ _0288_ _0366_ _0376_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_35_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_53_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1012_ _0184_ _0207_ _0257_ _0303_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__nor4_1
XFILLER_0_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_62_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0727_ net110 net103 net100 net98 VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0992_ _0693_ _0104_ _0280_ _0282_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__or4_2
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1260_ _0248_ _0249_ _0274_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__or3_1
X_1191_ _0185_ _0187_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__or2_2
Xinput8 addr0[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_62_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0975_ _0068_ _0264_ _0266_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__or3_2
XFILLER_0_27_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1389_ _0098_ _0176_ _0296_ _0297_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__or4_1
X_1458_ clknet_2_2__leaf_clk0 _0030_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0760_ net115 net65 net62 net113 VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__a22o_2
XFILLER_0_28_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1174_ _0089_ _0161_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1243_ _0086_ _0109_ _0292_ _0295_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__or4_1
X_1312_ _0085_ _0089_ _0229_ _0584_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__or4_1
XANTENNA_13 _0225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0958_ net87 net57 net55 net89 VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_30_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_24 _0615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0889_ net56 net52 net49 net54 VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__a22o_2
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap48 _0073_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0743_ net142 net140 net138 net144 VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__and4bb_1
X_0812_ net121 net103 net98 net116 VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__a22o_2
XFILLER_0_58_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1157_ _0435_ _0436_ _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_35_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1226_ _0138_ _0241_ _0254_ _0505_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1088_ _0043_ _0245_ _0369_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__or3_1
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1011_ _0269_ _0279_ _0289_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_6_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0726_ net144 net142 net140 net138 VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__and4b_1
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1209_ _0072_ _0075_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0991_ _0104_ _0282_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput9 cs0 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
X_1190_ _0113_ _0164_ _0166_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_62_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0974_ net70 net61 net59 net68 VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1457_ clknet_2_2__leaf_clk0 _0029_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1388_ net42 _0650_ _0655_ net149 net127 VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_25_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1311_ _0114_ _0197_ _0232_ _0245_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__or4_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1173_ net45 _0448_ _0456_ net173 net129 VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__o32a_1
X_1242_ _0214_ _0223_ _0244_ _0513_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_14 _0277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 _0654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0957_ net86 net69 net67 net88 VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_30_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0888_ _0178_ _0179_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0742_ net138 net140 net142 net144 VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__and4b_1
X_0811_ net119 net52 net49 net123 VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__a22o_2
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1156_ _0199_ _0437_ _0438_ _0440_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_35_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1087_ _0098_ _0176_ _0234_ _0367_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__or4_1
X_1225_ _0099_ _0127_ _0157_ _0179_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1010_ _0294_ _0301_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_6_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0725_ net137 net135 net133 net131 VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1208_ _0136_ _0250_ _0252_ _0488_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__or4_2
X_1139_ _0164_ _0167_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1 net29 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0990_ net116 net92 net90 net121 VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__a22o_2
XFILLER_0_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0973_ _0068_ _0264_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__or2_2
XFILLER_0_22_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1387_ _0649_ _0651_ _0653_ _0654_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__or4_1
X_1456_ clknet_2_2__leaf_clk0 _0028_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1241_ _0079_ _0253_ _0348_ _0413_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_22_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1310_ _0106_ _0273_ _0310_ _0332_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__or4_1
X_1172_ _0445_ _0450_ _0453_ _0455_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_15 _0280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _0707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0956_ net93 net88 net86 net91 VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__a22o_2
XFILLER_0_27_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0887_ net90 net52 net49 net92 VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__a22o_1
X_1439_ clknet_2_0__leaf_clk0 _0011_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_38_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0810_ net112 net53 net49 net114 VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__a22o_2
X_0741_ net123 net88 net86 net119 VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1224_ _0390_ _0458_ _0490_ _0503_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1155_ _0127_ _0389_ _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_35_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1086_ _0647_ net47 _0105_ _0274_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__or4_1
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0939_ _0123_ _0124_ _0125_ _0229_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__or4_4
XFILLER_0_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0724_ net144 net140 net138 net142 VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__nor4b_1
X_1207_ _0057_ _0058_ _0164_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_40_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1138_ net44 _0410_ _0423_ net160 net128 VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__o32a_1
X_1069_ _0097_ _0236_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 net39 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0972_ net104 net60 net58 net98 VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1386_ _0164_ _0166_ _0356_ _0550_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__or4_2
X_1455_ clknet_2_2__leaf_clk0 _0027_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1240_ _0512_ _0516_ _0517_ _0518_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__or4_1
X_1171_ _0084_ _0193_ _0290_ _0454_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__or4_1
XFILLER_0_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_27 _0707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_16 _0280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0955_ _0707_ _0710_ _0244_ _0245_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__or4_2
XFILLER_0_27_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0886_ net104 net53 net50 net99 VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__a22o_2
XFILLER_0_30_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1438_ clknet_2_1__leaf_clk0 _0010_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1369_ _0131_ _0192_ _0335_ _0415_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0740_ net114 net88 net86 net112 VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1154_ _0130_ _0156_ _0157_ _0214_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__or4_1
X_1223_ _0094_ _0270_ _0502_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__or3_1
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1085_ _0264_ _0268_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_35_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0938_ _0124_ _0229_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__or2_1
X_0869_ _0088_ _0160_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__or2_2
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire71 net72 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0723_ net137 net135 net131 net133 VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1206_ _0135_ _0141_ _0430_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__or3_1
X_1137_ _0417_ _0420_ _0421_ _0422_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__or4_2
X_1068_ _0107_ _0217_ _0221_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3 net21 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0971_ net91 net61 net58 net93 VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1454_ clknet_2_0__leaf_clk0 _0026_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1385_ _0704_ _0171_ _0203_ _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ _0275_ _0285_ _0405_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__or3_1
XFILLER_0_63_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0954_ _0711_ _0245_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__or2_1
XANTENNA_28 _0707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_17 _0291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0885_ _0097_ _0098_ _0099_ _0174_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__or4_1
X_1437_ clknet_2_1__leaf_clk0 _0009_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1299_ _0113_ _0214_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__or2_1
X_1368_ _0119_ _0180_ _0210_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1222_ _0104_ _0290_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__or2_1
X_1153_ _0696_ _0086_ _0104_ _0191_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__or4_1
X_1084_ _0263_ _0264_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_35_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0799_ _0089_ _0090_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__or2_2
X_0868_ net69 net65 net62 net67 VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__a22o_1
X_0937_ net83 net80 net78 net85 VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a22o_2
XFILLER_0_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire72 net77 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0722_ net122 net114 net112 net117 VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__a22o_4
X_1205_ net45 _0481_ _0486_ net158 net129 VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__o32a_1
XFILLER_0_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1136_ _0108_ _0220_ _0283_ _0372_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__or4_1
X_1067_ _0103_ _0156_ _0212_ _0214_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold4 net27 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1119_ _0120_ _0178_ _0179_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__or3_2
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_55_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0970_ _0063_ _0064_ _0258_ _0259_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__or4_4
XFILLER_0_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1453_ clknet_2_3__leaf_clk0 _0025_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfxtp_1
X_1384_ _0068_ _0069_ _0283_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_18 _0292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _0244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0953_ net97 net69 net67 net94 VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__a22o_2
XFILLER_0_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0884_ _0097_ _0174_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__or2_2
X_1436_ clknet_2_0__leaf_clk0 _0008_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dfxtp_1
X_1367_ net43 _0628_ _0635_ net176 net128 VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__o32a_1
XFILLER_0_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1298_ _0137_ _0140_ _0142_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__or3_2
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1221_ _0707_ _0237_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1152_ _0060_ _0203_ _0305_ _0430_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__or4_1
X_1083_ _0131_ _0192_ _0349_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__or3_1
XFILLER_0_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0936_ _0080_ _0081_ _0082_ _0225_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0867_ _0102_ _0103_ _0156_ _0157_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__or4_1
X_0798_ net91 net64 net62 net93 VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1419_ net125 _0696_ _0159_ _0370_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire73 net74 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0721_ net140 net138 net144 net142 VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__and4b_1
X_1204_ _0469_ _0482_ _0484_ _0485_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1135_ _0411_ _0414_ _0415_ _0416_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__or4_1
X_1066_ _0032_ _0164_ _0166_ _0240_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0919_ _0118_ _0119_ _0208_ _0210_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 net37 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_29_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap102 _0699_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1049_ _0115_ _0124_ _0137_ _0274_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__or4_1
X_1118_ _0120_ _0178_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1383_ _0190_ _0198_ _0388_ _0648_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__or4_1
X_1452_ clknet_2_3__leaf_clk0 _0024_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_19 _0295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0952_ net96 net57 net55 net94 VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__a22o_4
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0883_ _0100_ _0174_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1366_ _0627_ _0631_ _0634_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__or3_1
X_1435_ clknet_2_3__leaf_clk0 _0007_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1297_ net126 net159 net42 _0571_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__o22a_1
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1220_ net44 _0496_ _0500_ net157 net128 VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__o32a_1
X_1151_ _0077_ _0426_ _0428_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1082_ _0217_ _0221_ _0222_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__or3_2
XFILLER_0_55_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0935_ _0080_ _0225_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_43_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0866_ _0103_ _0157_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0797_ net103 net64 net63 net98 VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__a22o_2
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1349_ _0278_ _0286_ _0472_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1418_ _0083_ _0194_ _0283_ _0291_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire74 net75 VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_57_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0720_ net142 net138 net140 net144 VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1203_ _0272_ _0365_ _0460_ _0473_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__or4_1
X_1134_ _0128_ _0347_ _0418_ _0419_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1065_ _0204_ _0352_ _0353_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0849_ net89 net57 net55 net87 VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__a22o_2
XFILLER_0_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0918_ net112 net97 net95 net114 VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__a22o_2
XFILLER_0_59_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_1__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold6 net36 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1117_ net126 net150 net42 _0403_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_0_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1048_ _0220_ _0242_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1382_ _0391_ _0427_ _0512_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__or3_1
X_1451_ clknet_2_2__leaf_clk0 _0023_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0951_ _0236_ _0237_ _0239_ _0240_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0882_ net124 net53 net50 net120 VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__a22o_2
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1434_ clknet_2_3__leaf_clk0 _0006_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dfxtp_1
X_1365_ _0092_ _0313_ _0633_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__or3_1
X_1296_ _0562_ _0564_ _0567_ _0570_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_38_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1150_ _0425_ _0427_ _0433_ _0434_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1081_ _0088_ _0103_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0934_ _0082_ _0225_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__or2_1
X_0865_ net83 net52 net49 net85 VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__a22o_2
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0796_ net64 net56 net54 net63 VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__a22o_1
X_1417_ _0191_ _0273_ _0296_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1348_ _0091_ _0333_ _0372_ _0432_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__or4_1
X_1279_ _0130_ _0140_ _0166_ _0203_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire75 net76 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout140 net3 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_57_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1202_ _0204_ _0312_ _0483_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__or3_1
X_1064_ _0117_ _0131_ _0137_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__or3_1
X_1133_ _0057_ _0076_ _0097_ _0164_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0917_ _0118_ _0208_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__or2_2
XFILLER_0_43_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0848_ net89 net87 _0046_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0779_ net137 net130 net132 net135 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_59_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7 net26 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1047_ _0166_ _0221_ _0336_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__or3_1
XFILLER_0_48_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1116_ _0395_ _0400_ _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk0 clk0 VGND VGND VPWR VPWR clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1450_ clknet_2_0__leaf_clk0 _0022_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1381_ _0549_ _0559_ _0572_ _0602_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0950_ _0236_ _0237_ _0240_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__or3_1
X_0881_ _0056_ _0162_ _0169_ _0172_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__or4_2
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1433_ clknet_2_3__leaf_clk0 _0005_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_38_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1364_ _0063_ _0258_ _0292_ _0632_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__or4_1
X_1295_ _0301_ _0540_ _0568_ _0569_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__or4_1
XFILLER_0_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1080_ _0080_ _0226_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0933_ net78 net69 net67 net80 VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a22o_2
X_0795_ _0085_ _0086_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0864_ net68 net53 net50 net70 VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__a22o_4
X_1347_ _0129_ _0193_ _0525_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__or3_1
X_1416_ _0173_ net42 _0683_ net170 net126 VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__o32a_1
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1278_ _0369_ _0429_ _0491_ _0550_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__or4_1
Xwire76 _0041_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout141 net3 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__buf_1
Xfanout130 net131 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_57_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1201_ _0032_ _0036_ _0104_ _0105_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1063_ net125 _0186_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__or2_1
X_1132_ _0112_ _0185_ _0203_ _0237_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__or4_1
XFILLER_0_62_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0916_ net95 net69 net67 net97 VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__a22o_2
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0847_ _0702_ net89 VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__and2b_1
X_0778_ net135 net130 net132 net137 VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 net17 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1046_ net125 _0057_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__or2_1
X_1115_ _0392_ _0393_ _0401_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_0_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1029_ _0125_ _0137_ _0187_ _0212_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1380_ _0119_ _0209_ _0426_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__or3_1
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0880_ _0057_ _0058_ _0059_ _0170_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1432_ clknet_2_1__leaf_clk0 _0004_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1363_ _0058_ _0174_ _0214_ _0298_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_43_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1294_ _0696_ _0156_ _0280_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_52_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0932_ _0040_ _0219_ _0221_ _0222_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_43_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0863_ _0132_ _0146_ _0148_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0794_ net121 net92 net90 net116 VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__a22o_2
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1415_ _0636_ _0678_ _0680_ _0682_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__or4_1
X_1346_ net43 _0608_ _0616_ net175 net128 VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__o32a_1
X_1277_ _0135_ _0172_ _0232_ _0247_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout131 net8 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__buf_2
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout120 _0677_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout142 net2 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_57_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1200_ _0109_ _0277_ _0474_ _0475_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1062_ _0057_ _0171_ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_48_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1131_ _0135_ _0141_ _0368_ _0413_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0915_ _0195_ _0201_ _0206_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0846_ _0133_ _0134_ _0136_ _0137_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__or4_1
X_0777_ net113 net60 net59 net115 VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__a22o_4
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1329_ _0593_ _0595_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_3_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold9 net13 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1114_ _0100_ _0168_ _0387_ _0394_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__or4_1
X_1045_ _0049_ _0059_ _0069_ _0298_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_0_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0829_ net100 net56 net54 net110 VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__a22o_2
XFILLER_0_31_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1028_ _0051_ _0161_ _0318_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_34_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1431_ clknet_2_1__leaf_clk0 _0003_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dfxtp_1
X_1362_ _0051_ _0265_ _0629_ _0630_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1293_ _0049_ _0118_ _0120_ _0212_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__or4_1
XFILLER_0_58_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0931_ _0221_ _0222_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_43_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0862_ _0079_ _0096_ _0152_ _0153_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0793_ net116 net56 net54 net121 VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1276_ _0391_ _0409_ _0449_ _0548_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__or4_1
X_1414_ _0265_ _0268_ _0679_ _0681_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__or4_1
X_1345_ _0611_ _0612_ _0615_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout110 _0697_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_4
Xfanout121 _0667_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__buf_2
Xfanout143 net2 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__buf_1
Xfanout132 net133 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1130_ _0093_ _0170_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1061_ _0693_ _0280_ _0292_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0914_ _0705_ _0204_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__or2_1
X_0845_ net86 net84 net82 net88 VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__a22o_2
XFILLER_0_28_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0776_ net60 net56 net54 net59 VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__a22o_4
X_1259_ _0033_ _0052_ _0053_ _0089_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1328_ _0594_ _0596_ _0598_ _0599_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap118 _0687_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_1
X_1113_ _0352_ _0396_ _0397_ _0399_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__or4_2
X_1044_ _0121_ _0197_ _0332_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0759_ _0049_ _0050_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__or2_2
XFILLER_0_31_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0828_ net70 net53 net50 net68 VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_50_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1027_ _0036_ _0040_ _0080_ _0112_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1430_ clknet_2_1__leaf_clk0 _0002_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1292_ _0325_ _0516_ _0565_ _0566_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__or4_1
X_1361_ _0040_ _0121_ _0124_ _0245_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0861_ _0056_ _0109_ _0120_ _0122_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__or4_1
X_0930_ net96 net84 net82 net94 VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__a22o_4
X_0792_ _0082_ _0083_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1413_ _0182_ _0226_ _0278_ _0491_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1344_ _0078_ _0606_ _0613_ _0614_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__or4_2
X_1275_ _0267_ _0275_ _0285_ _0471_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout100 _0699_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_4
Xfanout111 _0697_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
Xfanout133 net7 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
Xfanout144 net1 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
Xfanout122 _0667_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_56_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1060_ _0693_ _0292_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0844_ net112 net88 net86 net114 VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__a22o_1
X_0913_ _0701_ _0202_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0775_ net143 net141 net139 net145 VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__and4b_1
X_1189_ _0082_ _0470_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__or2_1
X_1258_ _0281_ _0293_ _0385_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__or3_1
X_1327_ _0141_ _0203_ _0238_ _0262_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_19_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1112_ _0711_ _0057_ _0058_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__or4_1
X_1043_ _0707_ _0244_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0758_ net124 net65 net62 net120 VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_8_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0827_ net120 net97 net95 net124 VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__a22o_2
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1026_ _0078_ _0165_ _0265_ _0271_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1009_ _0069_ _0295_ _0297_ _0298_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__or4_2
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1360_ _0119_ _0208_ _0404_ _0561_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1291_ _0502_ _0544_ _0561_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0791_ _0080_ _0081_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_43_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0860_ _0711_ _0087_ _0150_ _0151_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1343_ _0157_ _0266_ _0297_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__or3_1
X_1412_ _0040_ _0350_ _0389_ _0525_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1274_ _0125_ _0229_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0989_ _0693_ _0280_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout101 net102 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout134 net135 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout123 net124 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_4
Xfanout112 net113 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_2
Xfanout145 net1 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__buf_1
XFILLER_0_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0912_ _0202_ _0203_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0843_ _0133_ _0134_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__or2_2
X_0774_ net141 net139 net145 net143 VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__and4bb_1
X_1326_ _0054_ _0178_ _0181_ _0597_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1188_ _0081_ _0225_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__or2_1
X_1257_ net44 _0530_ _0534_ net166 net128 VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_19_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap109 _0698_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1111_ _0088_ _0123_ _0136_ _0270_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__or4_1
X_1042_ net46 _0212_ _0214_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__or3_2
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0757_ net64 net62 _0046_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_24_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0826_ net94 net84 net82 net96 VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_8_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1309_ net43 _0580_ _0582_ net164 net127 VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_50_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1025_ _0260_ _0307_ _0313_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0809_ _0097_ _0098_ _0099_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 _0082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1008_ _0295_ _0298_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1290_ _0126_ _0309_ _0312_ _0429_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0790_ net78 net56 net54 net80 VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__a22o_4
XFILLER_0_11_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1342_ _0194_ _0205_ _0357_ _0488_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__or4_1
X_1273_ _0100_ _0178_ _0181_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__or3_1
X_1411_ _0115_ _0130_ _0131_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0988_ net121 net84 net82 net116 VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__a22o_2
Xfanout113 _0695_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_2
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout135 net6 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
Xfanout124 _0657_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__buf_2
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0911_ net110 net56 net54 net100 VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__a22o_4
X_0842_ net104 net89 net87 net99 VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0773_ _0063_ _0064_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__or2_2
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1256_ _0471_ _0525_ _0526_ _0533_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__or4_1
X_1325_ _0647_ _0082_ _0098_ _0156_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1187_ _0157_ _0174_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_19_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1110_ _0083_ _0102_ _0135_ _0156_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1041_ _0037_ _0182_ _0330_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0825_ net98 net88 net86 net103 VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__a22o_2
XFILLER_0_28_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0756_ net131 net133 net137 net135 VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__and4bb_1
X_1239_ _0178_ _0181_ _0336_ _0502_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1308_ _0195_ _0393_ _0501_ _0581_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__or4_1
XFILLER_0_62_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1024_ _0308_ _0309_ _0311_ _0314_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_64_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0808_ _0098_ _0099_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__or2_2
X_0739_ net132 net130 net134 net136 VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_27_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_2 _0082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1007_ _0297_ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1410_ _0077_ _0370_ _0676_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1272_ _0215_ _0248_ _0251_ _0283_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__or4_1
X_1341_ _0244_ _0245_ _0294_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0987_ _0273_ _0275_ _0278_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout103 net105 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_4
Xfanout125 _0647_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_4
Xfanout136 net137 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout114 net115 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__buf_2
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0772_ net123 net60 net59 net119 VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0841_ net90 net88 net87 net92 VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__a22o_2
X_0910_ net101 net93 net90 net111 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1186_ net45 _0464_ _0468_ net163 net129 VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__o32a_1
X_1324_ _0091_ _0171_ _0233_ _0349_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1255_ _0231_ _0528_ _0531_ _0532_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_45_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1040_ _0093_ _0094_ _0211_ _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0824_ _0114_ _0115_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0755_ net137 net135 net131 net133 VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1169_ _0091_ _0449_ _0451_ _0452_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__or4_1
X_1238_ _0168_ _0265_ _0305_ _0358_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__or4_1
X_1307_ _0054_ _0072_ _0074_ _0394_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1023_ _0069_ _0094_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0738_ net136 net134 net130 net132 VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0807_ net52 net49 _0046_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__o21ba_2
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_3 _0082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1006_ net119 net60 net59 net123 VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_32_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput40 net40 VGND VGND VPWR VPWR dout0[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1340_ _0338_ _0516_ _0609_ _0610_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__or4_1
XFILLER_0_64_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1271_ net129 net171 net45 _0547_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0986_ _0276_ _0277_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__or2_2
XFILLER_0_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout126 net128 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__buf_2
Xfanout115 _0694_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_2
Xfanout137 net5 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
Xfanout104 net106 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0840_ _0128_ _0129_ _0130_ _0131_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0771_ net84 net61 net58 net82 VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1323_ _0267_ _0390_ _0572_ _0592_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1185_ _0132_ _0334_ _0465_ _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__or4_1
X_1254_ _0051_ _0075_ _0213_ _0268_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0969_ _0258_ _0259_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0823_ net113 net110 net100 net115 VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__a22o_2
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0754_ net145 net143 net141 net139 VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__or4b_4
X_1306_ _0503_ _0572_ _0573_ _0579_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__or4_1
X_1168_ _0168_ _0176_ _0443_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1237_ _0037_ _0134_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__or2_2
X_1099_ _0704_ _0130_ _0131_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__or3_1
XFILLER_0_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_0__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_13_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1022_ _0248_ _0249_ _0312_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__or3_2
XFILLER_0_29_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0737_ _0707_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__or2_2
XFILLER_0_12_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0806_ net115 net52 net49 net113 VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__a22o_4
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_4 _0082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1005_ net83 net60 net59 net85 VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__a22o_2
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput41 net41 VGND VGND VPWR VPWR dout0[9] sky130_fd_sc_hd__clkbuf_4
Xoutput30 net30 VGND VGND VPWR VPWR dout0[28] sky130_fd_sc_hd__buf_2
XFILLER_0_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
.ends

