module cust_rom (clk0,
    cs0,
    addr0,
    dout0);
 input clk0;
 input cs0;
 input [6:0] addr0;
 output [15:0] dout0;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire \addr0_reg[0] ;
 wire \addr0_reg[1] ;
 wire \addr0_reg[2] ;
 wire \addr0_reg[3] ;
 wire \addr0_reg[4] ;
 wire \addr0_reg[5] ;
 wire \addr0_reg[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire clknet_0_clk0;
 wire clknet_1_0__leaf_clk0;
 wire clknet_1_1__leaf_clk0;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;

 sky130_fd_sc_hd__inv_2 _241_ (.A(net8),
    .Y(_182_));
 sky130_fd_sc_hd__and3_1 _242_ (.A(net47),
    .B(\addr0_reg[5] ),
    .C(\addr0_reg[6] ),
    .X(_183_));
 sky130_fd_sc_hd__and4bb_2 _243_ (.A_N(net51),
    .B_N(net55),
    .C(net53),
    .D(net49),
    .X(_184_));
 sky130_fd_sc_hd__nor2_1 _244_ (.A(net47),
    .B(\addr0_reg[5] ),
    .Y(_185_));
 sky130_fd_sc_hd__nor3b_1 _245_ (.A(net47),
    .B(\addr0_reg[5] ),
    .C_N(\addr0_reg[6] ),
    .Y(_186_));
 sky130_fd_sc_hd__and4bb_2 _246_ (.A_N(net49),
    .B_N(net55),
    .C(net53),
    .D(net51),
    .X(_187_));
 sky130_fd_sc_hd__a22o_1 _247_ (.A1(net45),
    .A2(_184_),
    .B1(net43),
    .B2(_187_),
    .X(_188_));
 sky130_fd_sc_hd__and4bb_2 _248_ (.A_N(net51),
    .B_N(net53),
    .C(net55),
    .D(net49),
    .X(_189_));
 sky130_fd_sc_hd__and4b_2 _249_ (.A_N(net49),
    .B(net53),
    .C(net55),
    .D(net51),
    .X(_190_));
 sky130_fd_sc_hd__a22o_1 _250_ (.A1(net46),
    .A2(_189_),
    .B1(_190_),
    .B2(net44),
    .X(_191_));
 sky130_fd_sc_hd__or4b_1 _251_ (.A(net50),
    .B(net52),
    .C(net54),
    .D_N(net48),
    .X(_192_));
 sky130_fd_sc_hd__o21ba_1 _252_ (.A1(net46),
    .A2(net44),
    .B1_N(_192_),
    .X(_193_));
 sky130_fd_sc_hd__and4b_2 _253_ (.A_N(net51),
    .B(net49),
    .C(net53),
    .D(net55),
    .X(_194_));
 sky130_fd_sc_hd__and4bb_2 _254_ (.A_N(net49),
    .B_N(net53),
    .C(net55),
    .D(net51),
    .X(_195_));
 sky130_fd_sc_hd__a22o_1 _255_ (.A1(net45),
    .A2(_194_),
    .B1(_195_),
    .B2(net43),
    .X(_196_));
 sky130_fd_sc_hd__or3_1 _256_ (.A(_188_),
    .B(_191_),
    .C(_196_),
    .X(_197_));
 sky130_fd_sc_hd__a22o_1 _257_ (.A1(net43),
    .A2(_194_),
    .B1(_195_),
    .B2(net45),
    .X(_198_));
 sky130_fd_sc_hd__nor4b_2 _258_ (.A(net48),
    .B(net52),
    .C(net54),
    .D_N(net50),
    .Y(_199_));
 sky130_fd_sc_hd__and4bb_2 _259_ (.A_N(net52),
    .B_N(net54),
    .C(net50),
    .D(net48),
    .X(_200_));
 sky130_fd_sc_hd__a22o_1 _260_ (.A1(net45),
    .A2(net42),
    .B1(_200_),
    .B2(net43),
    .X(_201_));
 sky130_fd_sc_hd__or2_1 _261_ (.A(_198_),
    .B(_201_),
    .X(_202_));
 sky130_fd_sc_hd__and3b_1 _262_ (.A_N(net47),
    .B(\addr0_reg[5] ),
    .C(\addr0_reg[6] ),
    .X(_203_));
 sky130_fd_sc_hd__nor4b_2 _263_ (.A(net50),
    .B(net48),
    .C(net52),
    .D_N(net54),
    .Y(_204_));
 sky130_fd_sc_hd__and3b_1 _264_ (.A_N(\addr0_reg[5] ),
    .B(\addr0_reg[6] ),
    .C(net47),
    .X(_205_));
 sky130_fd_sc_hd__and4_2 _265_ (.A(net50),
    .B(net48),
    .C(net52),
    .D(net54),
    .X(_206_));
 sky130_fd_sc_hd__a22o_1 _266_ (.A1(net40),
    .A2(net39),
    .B1(net37),
    .B2(_206_),
    .X(_207_));
 sky130_fd_sc_hd__nor4_1 _267_ (.A(net50),
    .B(net48),
    .C(net52),
    .D(net54),
    .Y(_208_));
 sky130_fd_sc_hd__a21o_1 _268_ (.A1(net40),
    .A2(_208_),
    .B1(_207_),
    .X(_209_));
 sky130_fd_sc_hd__or4_1 _269_ (.A(_193_),
    .B(_197_),
    .C(_202_),
    .D(_209_),
    .X(_210_));
 sky130_fd_sc_hd__a22o_1 _270_ (.A1(net44),
    .A2(_189_),
    .B1(_190_),
    .B2(net46),
    .X(_211_));
 sky130_fd_sc_hd__a22o_1 _271_ (.A1(_184_),
    .A2(net44),
    .B1(_187_),
    .B2(net46),
    .X(_212_));
 sky130_fd_sc_hd__or2_1 _272_ (.A(_211_),
    .B(_212_),
    .X(_213_));
 sky130_fd_sc_hd__a22oi_1 _273_ (.A1(_200_),
    .A2(net40),
    .B1(net37),
    .B2(_199_),
    .Y(_214_));
 sky130_fd_sc_hd__and4b_2 _274_ (.A_N(net52),
    .B(net54),
    .C(net50),
    .D(net48),
    .X(_215_));
 sky130_fd_sc_hd__and4bb_2 _275_ (.A_N(net50),
    .B_N(net48),
    .C(net52),
    .D(net54),
    .X(_216_));
 sky130_fd_sc_hd__a22o_1 _276_ (.A1(net40),
    .A2(_215_),
    .B1(_216_),
    .B2(net37),
    .X(_217_));
 sky130_fd_sc_hd__a221o_1 _277_ (.A1(_200_),
    .A2(net40),
    .B1(net37),
    .B2(_199_),
    .C1(_217_),
    .X(_218_));
 sky130_fd_sc_hd__a22o_1 _278_ (.A1(_187_),
    .A2(net41),
    .B1(net38),
    .B2(_184_),
    .X(_219_));
 sky130_fd_sc_hd__a22o_1 _279_ (.A1(_190_),
    .A2(net40),
    .B1(net37),
    .B2(_189_),
    .X(_220_));
 sky130_fd_sc_hd__or2_1 _280_ (.A(_219_),
    .B(_220_),
    .X(_221_));
 sky130_fd_sc_hd__and4b_2 _281_ (.A_N(net54),
    .B(net52),
    .C(net48),
    .D(net50),
    .X(_222_));
 sky130_fd_sc_hd__nor4b_2 _282_ (.A(net50),
    .B(net48),
    .C(net54),
    .D_N(net52),
    .Y(_223_));
 sky130_fd_sc_hd__a22o_1 _283_ (.A1(net40),
    .A2(_222_),
    .B1(_223_),
    .B2(net37),
    .X(_224_));
 sky130_fd_sc_hd__a22o_1 _284_ (.A1(net39),
    .A2(net37),
    .B1(_206_),
    .B2(net40),
    .X(_225_));
 sky130_fd_sc_hd__or2_1 _285_ (.A(_224_),
    .B(_225_),
    .X(_226_));
 sky130_fd_sc_hd__or4_1 _286_ (.A(_213_),
    .B(_218_),
    .C(_221_),
    .D(_226_),
    .X(_227_));
 sky130_fd_sc_hd__a22o_1 _287_ (.A1(_194_),
    .A2(net41),
    .B1(net38),
    .B2(_195_),
    .X(_228_));
 sky130_fd_sc_hd__a22o_1 _288_ (.A1(_184_),
    .A2(net41),
    .B1(net38),
    .B2(_187_),
    .X(_229_));
 sky130_fd_sc_hd__or2_1 _289_ (.A(_228_),
    .B(_229_),
    .X(_230_));
 sky130_fd_sc_hd__a22o_1 _290_ (.A1(_195_),
    .A2(net41),
    .B1(net38),
    .B2(_194_),
    .X(_231_));
 sky130_fd_sc_hd__a221o_1 _291_ (.A1(net38),
    .A2(_222_),
    .B1(net35),
    .B2(net41),
    .C1(_231_),
    .X(_232_));
 sky130_fd_sc_hd__a22o_1 _292_ (.A1(_189_),
    .A2(net40),
    .B1(net37),
    .B2(_190_),
    .X(_233_));
 sky130_fd_sc_hd__o21ba_1 _293_ (.A1(net40),
    .A2(net37),
    .B1_N(_192_),
    .X(_234_));
 sky130_fd_sc_hd__or2_1 _294_ (.A(_233_),
    .B(_234_),
    .X(_235_));
 sky130_fd_sc_hd__a22o_1 _295_ (.A1(net42),
    .A2(net41),
    .B1(net38),
    .B2(_200_),
    .X(_236_));
 sky130_fd_sc_hd__a22o_1 _296_ (.A1(net37),
    .A2(_215_),
    .B1(_216_),
    .B2(net41),
    .X(_237_));
 sky130_fd_sc_hd__or2_1 _297_ (.A(_236_),
    .B(_237_),
    .X(_238_));
 sky130_fd_sc_hd__or4_1 _298_ (.A(_230_),
    .B(_232_),
    .C(_235_),
    .D(_238_),
    .X(_239_));
 sky130_fd_sc_hd__a22o_1 _299_ (.A1(net45),
    .A2(_215_),
    .B1(_216_),
    .B2(net43),
    .X(_240_));
 sky130_fd_sc_hd__a22o_1 _300_ (.A1(net43),
    .A2(net39),
    .B1(_206_),
    .B2(net45),
    .X(_016_));
 sky130_fd_sc_hd__or2_1 _301_ (.A(_240_),
    .B(_016_),
    .X(_017_));
 sky130_fd_sc_hd__a22o_1 _302_ (.A1(net43),
    .A2(net42),
    .B1(_200_),
    .B2(net45),
    .X(_018_));
 sky130_fd_sc_hd__a22o_1 _303_ (.A1(net45),
    .A2(_222_),
    .B1(net35),
    .B2(net43),
    .X(_019_));
 sky130_fd_sc_hd__or4_1 _304_ (.A(_240_),
    .B(_016_),
    .C(_018_),
    .D(_019_),
    .X(_020_));
 sky130_fd_sc_hd__a22o_1 _305_ (.A1(net43),
    .A2(_222_),
    .B1(net35),
    .B2(net45),
    .X(_021_));
 sky130_fd_sc_hd__a22o_1 _306_ (.A1(net43),
    .A2(_215_),
    .B1(_216_),
    .B2(net45),
    .X(_022_));
 sky130_fd_sc_hd__or2_1 _307_ (.A(_021_),
    .B(_022_),
    .X(_023_));
 sky130_fd_sc_hd__a22o_1 _308_ (.A1(net46),
    .A2(_204_),
    .B1(_206_),
    .B2(net44),
    .X(_024_));
 sky130_fd_sc_hd__and3_1 _309_ (.A(\addr0_reg[4] ),
    .B(\addr0_reg[6] ),
    .C(net36),
    .X(_025_));
 sky130_fd_sc_hd__or4_1 _310_ (.A(_020_),
    .B(_023_),
    .C(_024_),
    .D(_025_),
    .X(_026_));
 sky130_fd_sc_hd__o41a_1 _311_ (.A1(_210_),
    .A2(_227_),
    .A3(_239_),
    .A4(_026_),
    .B1(net8),
    .X(_027_));
 sky130_fd_sc_hd__nor3b_1 _312_ (.A(net47),
    .B(\addr0_reg[6] ),
    .C_N(\addr0_reg[5] ),
    .Y(_028_));
 sky130_fd_sc_hd__nor3b_1 _313_ (.A(\addr0_reg[5] ),
    .B(\addr0_reg[6] ),
    .C_N(net47),
    .Y(_029_));
 sky130_fd_sc_hd__a22o_1 _314_ (.A1(_199_),
    .A2(net33),
    .B1(net31),
    .B2(_200_),
    .X(_030_));
 sky130_fd_sc_hd__a22o_1 _315_ (.A1(_216_),
    .A2(net33),
    .B1(net31),
    .B2(_215_),
    .X(_031_));
 sky130_fd_sc_hd__a22o_1 _316_ (.A1(_223_),
    .A2(net33),
    .B1(net31),
    .B2(_222_),
    .X(_032_));
 sky130_fd_sc_hd__a22o_1 _317_ (.A1(net39),
    .A2(net33),
    .B1(net31),
    .B2(_206_),
    .X(_033_));
 sky130_fd_sc_hd__or2_1 _318_ (.A(_032_),
    .B(_033_),
    .X(_034_));
 sky130_fd_sc_hd__or4_2 _319_ (.A(_030_),
    .B(_031_),
    .C(_032_),
    .D(_033_),
    .X(_035_));
 sky130_fd_sc_hd__a22o_1 _320_ (.A1(_187_),
    .A2(net34),
    .B1(net32),
    .B2(_184_),
    .X(_036_));
 sky130_fd_sc_hd__o21ba_1 _321_ (.A1(net33),
    .A2(net31),
    .B1_N(_192_),
    .X(_037_));
 sky130_fd_sc_hd__a22o_1 _322_ (.A1(_195_),
    .A2(net34),
    .B1(net32),
    .B2(_194_),
    .X(_038_));
 sky130_fd_sc_hd__a22o_1 _323_ (.A1(_190_),
    .A2(net34),
    .B1(net32),
    .B2(_189_),
    .X(_039_));
 sky130_fd_sc_hd__or2_1 _324_ (.A(_036_),
    .B(_038_),
    .X(_040_));
 sky130_fd_sc_hd__or4_1 _325_ (.A(_036_),
    .B(_037_),
    .C(_038_),
    .D(_039_),
    .X(_041_));
 sky130_fd_sc_hd__or2_1 _326_ (.A(_035_),
    .B(_041_),
    .X(_042_));
 sky130_fd_sc_hd__a22o_1 _327_ (.A1(_222_),
    .A2(net33),
    .B1(net31),
    .B2(_223_),
    .X(_043_));
 sky130_fd_sc_hd__a22o_1 _328_ (.A1(_215_),
    .A2(net33),
    .B1(net31),
    .B2(_216_),
    .X(_044_));
 sky130_fd_sc_hd__and3b_1 _329_ (.A_N(\addr0_reg[6] ),
    .B(net36),
    .C(net47),
    .X(_045_));
 sky130_fd_sc_hd__a22o_1 _330_ (.A1(_206_),
    .A2(net33),
    .B1(net31),
    .B2(_204_),
    .X(_046_));
 sky130_fd_sc_hd__or2_1 _331_ (.A(_045_),
    .B(_046_),
    .X(_047_));
 sky130_fd_sc_hd__or3_1 _332_ (.A(_043_),
    .B(_044_),
    .C(_046_),
    .X(_048_));
 sky130_fd_sc_hd__or4_1 _333_ (.A(_043_),
    .B(_044_),
    .C(_045_),
    .D(_046_),
    .X(_049_));
 sky130_fd_sc_hd__a22o_1 _334_ (.A1(_200_),
    .A2(net34),
    .B1(net32),
    .B2(net42),
    .X(_050_));
 sky130_fd_sc_hd__a22o_1 _335_ (.A1(_194_),
    .A2(net34),
    .B1(net32),
    .B2(_195_),
    .X(_051_));
 sky130_fd_sc_hd__or2_1 _336_ (.A(_050_),
    .B(_051_),
    .X(_052_));
 sky130_fd_sc_hd__a22o_1 _337_ (.A1(_184_),
    .A2(net33),
    .B1(net31),
    .B2(_187_),
    .X(_053_));
 sky130_fd_sc_hd__a22o_1 _338_ (.A1(_189_),
    .A2(net33),
    .B1(net31),
    .B2(_190_),
    .X(_054_));
 sky130_fd_sc_hd__or4_2 _339_ (.A(_050_),
    .B(_051_),
    .C(_053_),
    .D(_054_),
    .X(_055_));
 sky130_fd_sc_hd__nor4_1 _340_ (.A(_035_),
    .B(_041_),
    .C(_049_),
    .D(_055_),
    .Y(_056_));
 sky130_fd_sc_hd__and3b_1 _341_ (.A_N(\addr0_reg[6] ),
    .B(\addr0_reg[5] ),
    .C(net47),
    .X(_057_));
 sky130_fd_sc_hd__nor3_1 _342_ (.A(net47),
    .B(\addr0_reg[5] ),
    .C(\addr0_reg[6] ),
    .Y(_058_));
 sky130_fd_sc_hd__a22o_1 _343_ (.A1(net42),
    .A2(net30),
    .B1(net28),
    .B2(_200_),
    .X(_059_));
 sky130_fd_sc_hd__a22o_1 _344_ (.A1(_216_),
    .A2(net29),
    .B1(net27),
    .B2(_215_),
    .X(_060_));
 sky130_fd_sc_hd__or2_1 _345_ (.A(_059_),
    .B(_060_),
    .X(_061_));
 sky130_fd_sc_hd__a22oi_1 _346_ (.A1(_204_),
    .A2(net29),
    .B1(net27),
    .B2(_206_),
    .Y(_062_));
 sky130_fd_sc_hd__a22oi_1 _347_ (.A1(_223_),
    .A2(net29),
    .B1(net27),
    .B2(_222_),
    .Y(_063_));
 sky130_fd_sc_hd__nand2_1 _348_ (.A(_062_),
    .B(_063_),
    .Y(_064_));
 sky130_fd_sc_hd__nor2_1 _349_ (.A(_061_),
    .B(_064_),
    .Y(_065_));
 sky130_fd_sc_hd__a22o_1 _350_ (.A1(_187_),
    .A2(net30),
    .B1(net28),
    .B2(_184_),
    .X(_066_));
 sky130_fd_sc_hd__a22o_1 _351_ (.A1(_195_),
    .A2(net29),
    .B1(net27),
    .B2(_194_),
    .X(_067_));
 sky130_fd_sc_hd__or2_1 _352_ (.A(_066_),
    .B(_067_),
    .X(_068_));
 sky130_fd_sc_hd__a22o_1 _353_ (.A1(_206_),
    .A2(net29),
    .B1(net27),
    .B2(_204_),
    .X(_069_));
 sky130_fd_sc_hd__a22o_1 _354_ (.A1(_190_),
    .A2(net29),
    .B1(net27),
    .B2(_189_),
    .X(_070_));
 sky130_fd_sc_hd__o21ba_1 _355_ (.A1(net29),
    .A2(net27),
    .B1_N(_192_),
    .X(_071_));
 sky130_fd_sc_hd__or2_1 _356_ (.A(_070_),
    .B(_071_),
    .X(_072_));
 sky130_fd_sc_hd__a22o_1 _357_ (.A1(_184_),
    .A2(net30),
    .B1(net28),
    .B2(_187_),
    .X(_073_));
 sky130_fd_sc_hd__a22o_1 _358_ (.A1(_189_),
    .A2(net30),
    .B1(net28),
    .B2(_190_),
    .X(_074_));
 sky130_fd_sc_hd__or2_1 _359_ (.A(_073_),
    .B(_074_),
    .X(_075_));
 sky130_fd_sc_hd__nor2_1 _360_ (.A(_072_),
    .B(_075_),
    .Y(_076_));
 sky130_fd_sc_hd__a22o_1 _361_ (.A1(_222_),
    .A2(net29),
    .B1(net27),
    .B2(_223_),
    .X(_077_));
 sky130_fd_sc_hd__a22o_1 _362_ (.A1(_215_),
    .A2(net29),
    .B1(net27),
    .B2(_216_),
    .X(_078_));
 sky130_fd_sc_hd__a22o_1 _363_ (.A1(_194_),
    .A2(net30),
    .B1(net28),
    .B2(_195_),
    .X(_079_));
 sky130_fd_sc_hd__a22o_1 _364_ (.A1(_200_),
    .A2(net30),
    .B1(net28),
    .B2(net42),
    .X(_080_));
 sky130_fd_sc_hd__or2_1 _365_ (.A(_079_),
    .B(_080_),
    .X(_081_));
 sky130_fd_sc_hd__or4_2 _366_ (.A(_077_),
    .B(_078_),
    .C(_079_),
    .D(_080_),
    .X(_082_));
 sky130_fd_sc_hd__a2111oi_1 _367_ (.A1(_185_),
    .A2(net36),
    .B1(_068_),
    .C1(_069_),
    .D1(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__a41oi_1 _368_ (.A1(_056_),
    .A2(_065_),
    .A3(_076_),
    .A4(net26),
    .B1(net56),
    .Y(_084_));
 sky130_fd_sc_hd__or2_2 _369_ (.A(_027_),
    .B(_084_),
    .X(_085_));
 sky130_fd_sc_hd__nand2_1 _370_ (.A(_214_),
    .B(_062_),
    .Y(_086_));
 sky130_fd_sc_hd__or3_1 _371_ (.A(_224_),
    .B(_070_),
    .C(_086_),
    .X(_087_));
 sky130_fd_sc_hd__or4_1 _372_ (.A(_032_),
    .B(_037_),
    .C(_043_),
    .D(_055_),
    .X(_088_));
 sky130_fd_sc_hd__or2_1 _373_ (.A(_198_),
    .B(_079_),
    .X(_089_));
 sky130_fd_sc_hd__a2111o_1 _374_ (.A1(\addr0_reg[4] ),
    .A2(net36),
    .B1(_219_),
    .C1(_024_),
    .D1(_196_),
    .X(_090_));
 sky130_fd_sc_hd__or4_1 _375_ (.A(_213_),
    .B(_030_),
    .C(_031_),
    .D(_090_),
    .X(_091_));
 sky130_fd_sc_hd__or4_1 _376_ (.A(_040_),
    .B(_068_),
    .C(_089_),
    .D(_091_),
    .X(_092_));
 sky130_fd_sc_hd__or4_1 _377_ (.A(_239_),
    .B(_087_),
    .C(_088_),
    .D(_092_),
    .X(_093_));
 sky130_fd_sc_hd__a22o_1 _378_ (.A1(net72),
    .A2(net56),
    .B1(net25),
    .B2(_093_),
    .X(_000_));
 sky130_fd_sc_hd__or2_1 _379_ (.A(_059_),
    .B(_064_),
    .X(_094_));
 sky130_fd_sc_hd__or2_1 _380_ (.A(_220_),
    .B(_236_),
    .X(_095_));
 sky130_fd_sc_hd__or3_1 _381_ (.A(_234_),
    .B(_019_),
    .C(_095_),
    .X(_096_));
 sky130_fd_sc_hd__or4_1 _382_ (.A(_230_),
    .B(_232_),
    .C(_094_),
    .D(_096_),
    .X(_097_));
 sky130_fd_sc_hd__or2_1 _383_ (.A(_050_),
    .B(_054_),
    .X(_098_));
 sky130_fd_sc_hd__or2_1 _384_ (.A(_039_),
    .B(_077_),
    .X(_099_));
 sky130_fd_sc_hd__or2_1 _385_ (.A(_031_),
    .B(_036_),
    .X(_100_));
 sky130_fd_sc_hd__or2_1 _386_ (.A(_068_),
    .B(_071_),
    .X(_101_));
 sky130_fd_sc_hd__or2_1 _387_ (.A(_021_),
    .B(_025_),
    .X(_102_));
 sky130_fd_sc_hd__or2_1 _388_ (.A(_201_),
    .B(_211_),
    .X(_103_));
 sky130_fd_sc_hd__or3_1 _389_ (.A(_098_),
    .B(_099_),
    .C(_103_),
    .X(_104_));
 sky130_fd_sc_hd__or4_1 _390_ (.A(_193_),
    .B(_196_),
    .C(_224_),
    .D(_100_),
    .X(_105_));
 sky130_fd_sc_hd__or3_1 _391_ (.A(_101_),
    .B(_102_),
    .C(_105_),
    .X(_106_));
 sky130_fd_sc_hd__or3_1 _392_ (.A(_097_),
    .B(_104_),
    .C(_106_),
    .X(_107_));
 sky130_fd_sc_hd__a22o_1 _393_ (.A1(net56),
    .A2(net70),
    .B1(net25),
    .B2(_107_),
    .X(_001_));
 sky130_fd_sc_hd__or4_1 _394_ (.A(_240_),
    .B(_018_),
    .C(_069_),
    .D(_073_),
    .X(_108_));
 sky130_fd_sc_hd__or3_1 _395_ (.A(_207_),
    .B(_220_),
    .C(_046_),
    .X(_109_));
 sky130_fd_sc_hd__or3_1 _396_ (.A(_226_),
    .B(_102_),
    .C(_109_),
    .X(_110_));
 sky130_fd_sc_hd__or3_1 _397_ (.A(_082_),
    .B(_108_),
    .C(_110_),
    .X(_111_));
 sky130_fd_sc_hd__or4_1 _398_ (.A(_229_),
    .B(_235_),
    .C(_040_),
    .D(_052_),
    .X(_112_));
 sky130_fd_sc_hd__or2_1 _399_ (.A(_030_),
    .B(_067_),
    .X(_113_));
 sky130_fd_sc_hd__or4_1 _400_ (.A(_031_),
    .B(_033_),
    .C(_072_),
    .D(_113_),
    .X(_114_));
 sky130_fd_sc_hd__or2_1 _401_ (.A(_024_),
    .B(_059_),
    .X(_115_));
 sky130_fd_sc_hd__a221o_1 _402_ (.A1(net38),
    .A2(_222_),
    .B1(net35),
    .B2(net41),
    .C1(_212_),
    .X(_116_));
 sky130_fd_sc_hd__or4_1 _403_ (.A(_188_),
    .B(_016_),
    .C(_115_),
    .D(_116_),
    .X(_117_));
 sky130_fd_sc_hd__or4_1 _404_ (.A(_111_),
    .B(_112_),
    .C(_114_),
    .D(_117_),
    .X(_118_));
 sky130_fd_sc_hd__a22o_1 _405_ (.A1(net57),
    .A2(net62),
    .B1(net25),
    .B2(_118_),
    .X(_002_));
 sky130_fd_sc_hd__or2_1 _406_ (.A(_066_),
    .B(_072_),
    .X(_119_));
 sky130_fd_sc_hd__or3_1 _407_ (.A(_218_),
    .B(_081_),
    .C(_119_),
    .X(_120_));
 sky130_fd_sc_hd__or4_1 _408_ (.A(_188_),
    .B(_198_),
    .C(_017_),
    .D(_100_),
    .X(_121_));
 sky130_fd_sc_hd__or4_1 _409_ (.A(_025_),
    .B(_033_),
    .C(_048_),
    .D(_054_),
    .X(_122_));
 sky130_fd_sc_hd__or4_1 _410_ (.A(_097_),
    .B(_120_),
    .C(_121_),
    .D(_122_),
    .X(_123_));
 sky130_fd_sc_hd__a22o_1 _411_ (.A1(net56),
    .A2(net61),
    .B1(net25),
    .B2(_123_),
    .X(_003_));
 sky130_fd_sc_hd__or3_1 _412_ (.A(_043_),
    .B(_050_),
    .C(_080_),
    .X(_124_));
 sky130_fd_sc_hd__or3_1 _413_ (.A(_072_),
    .B(_075_),
    .C(_124_),
    .X(_125_));
 sky130_fd_sc_hd__or3_1 _414_ (.A(_202_),
    .B(_053_),
    .C(_054_),
    .X(_126_));
 sky130_fd_sc_hd__or2_1 _415_ (.A(_191_),
    .B(_228_),
    .X(_127_));
 sky130_fd_sc_hd__or2_1 _416_ (.A(_196_),
    .B(_225_),
    .X(_128_));
 sky130_fd_sc_hd__or2_1 _417_ (.A(_237_),
    .B(_025_),
    .X(_129_));
 sky130_fd_sc_hd__or4_1 _418_ (.A(_040_),
    .B(_127_),
    .C(_128_),
    .D(_129_),
    .X(_130_));
 sky130_fd_sc_hd__or4_1 _419_ (.A(_207_),
    .B(_212_),
    .C(_217_),
    .D(_032_),
    .X(_131_));
 sky130_fd_sc_hd__or4_1 _420_ (.A(_017_),
    .B(_064_),
    .C(_130_),
    .D(_131_),
    .X(_132_));
 sky130_fd_sc_hd__or4_1 _421_ (.A(_096_),
    .B(_125_),
    .C(_126_),
    .D(_132_),
    .X(_133_));
 sky130_fd_sc_hd__a22o_1 _422_ (.A1(net57),
    .A2(net73),
    .B1(net25),
    .B2(_133_),
    .X(_004_));
 sky130_fd_sc_hd__or4_1 _423_ (.A(_036_),
    .B(_037_),
    .C(_069_),
    .D(_078_),
    .X(_134_));
 sky130_fd_sc_hd__or3_1 _424_ (.A(_034_),
    .B(_095_),
    .C(_134_),
    .X(_135_));
 sky130_fd_sc_hd__or2_1 _425_ (.A(_231_),
    .B(_023_),
    .X(_136_));
 sky130_fd_sc_hd__or3_1 _426_ (.A(_048_),
    .B(_135_),
    .C(_136_),
    .X(_137_));
 sky130_fd_sc_hd__a221o_1 _427_ (.A1(net39),
    .A2(net29),
    .B1(net27),
    .B2(_206_),
    .C1(_080_),
    .X(_138_));
 sky130_fd_sc_hd__or4_1 _428_ (.A(_052_),
    .B(_103_),
    .C(_129_),
    .D(_138_),
    .X(_139_));
 sky130_fd_sc_hd__or4_1 _429_ (.A(_233_),
    .B(_019_),
    .C(_053_),
    .D(_060_),
    .X(_140_));
 sky130_fd_sc_hd__or4_1 _430_ (.A(_197_),
    .B(_101_),
    .C(_139_),
    .D(_140_),
    .X(_141_));
 sky130_fd_sc_hd__or2_1 _431_ (.A(_137_),
    .B(_141_),
    .X(_142_));
 sky130_fd_sc_hd__a22o_1 _432_ (.A1(net57),
    .A2(net65),
    .B1(_085_),
    .B2(_142_),
    .X(_005_));
 sky130_fd_sc_hd__or3_1 _433_ (.A(_197_),
    .B(_049_),
    .C(_136_),
    .X(_143_));
 sky130_fd_sc_hd__or4_1 _434_ (.A(_053_),
    .B(_054_),
    .C(_077_),
    .D(_078_),
    .X(_144_));
 sky130_fd_sc_hd__or4_1 _435_ (.A(_201_),
    .B(_219_),
    .C(_234_),
    .D(_016_),
    .X(_145_));
 sky130_fd_sc_hd__or4_1 _436_ (.A(_039_),
    .B(_051_),
    .C(_080_),
    .D(_145_),
    .X(_146_));
 sky130_fd_sc_hd__or4_1 _437_ (.A(_086_),
    .B(_116_),
    .C(_144_),
    .D(_146_),
    .X(_147_));
 sky130_fd_sc_hd__or3_1 _438_ (.A(_114_),
    .B(_143_),
    .C(_147_),
    .X(_148_));
 sky130_fd_sc_hd__a22o_1 _439_ (.A1(net56),
    .A2(net63),
    .B1(_085_),
    .B2(_148_),
    .X(_006_));
 sky130_fd_sc_hd__or2_1 _440_ (.A(_229_),
    .B(_051_),
    .X(_149_));
 sky130_fd_sc_hd__or4_1 _441_ (.A(_231_),
    .B(_234_),
    .C(_054_),
    .D(_079_),
    .X(_150_));
 sky130_fd_sc_hd__or4_1 _442_ (.A(_193_),
    .B(_022_),
    .C(_034_),
    .D(_150_),
    .X(_151_));
 sky130_fd_sc_hd__or3_1 _443_ (.A(_020_),
    .B(_094_),
    .C(_151_),
    .X(_152_));
 sky130_fd_sc_hd__or4_1 _444_ (.A(_075_),
    .B(_113_),
    .C(_129_),
    .D(_149_),
    .X(_153_));
 sky130_fd_sc_hd__or3_1 _445_ (.A(_227_),
    .B(_152_),
    .C(_153_),
    .X(_154_));
 sky130_fd_sc_hd__a22o_1 _446_ (.A1(net56),
    .A2(net66),
    .B1(net25),
    .B2(_154_),
    .X(_007_));
 sky130_fd_sc_hd__or3_1 _447_ (.A(_089_),
    .B(_098_),
    .C(_115_),
    .X(_155_));
 sky130_fd_sc_hd__or3_1 _448_ (.A(_188_),
    .B(_193_),
    .C(_074_),
    .X(_156_));
 sky130_fd_sc_hd__or4_1 _449_ (.A(_212_),
    .B(_031_),
    .C(_045_),
    .D(_070_),
    .X(_157_));
 sky130_fd_sc_hd__or4_1 _450_ (.A(_230_),
    .B(_018_),
    .C(_019_),
    .D(_157_),
    .X(_158_));
 sky130_fd_sc_hd__or4_1 _451_ (.A(_137_),
    .B(_155_),
    .C(_156_),
    .D(_158_),
    .X(_159_));
 sky130_fd_sc_hd__a22o_1 _452_ (.A1(net57),
    .A2(net67),
    .B1(_085_),
    .B2(_159_),
    .X(_008_));
 sky130_fd_sc_hd__or4_1 _453_ (.A(_233_),
    .B(_037_),
    .C(_038_),
    .D(_046_),
    .X(_160_));
 sky130_fd_sc_hd__or4_1 _454_ (.A(_191_),
    .B(_193_),
    .C(_221_),
    .D(_160_),
    .X(_161_));
 sky130_fd_sc_hd__or4_1 _455_ (.A(_061_),
    .B(_089_),
    .C(_102_),
    .D(_149_),
    .X(_162_));
 sky130_fd_sc_hd__or4_1 _456_ (.A(_035_),
    .B(_044_),
    .C(_066_),
    .D(_077_),
    .X(_163_));
 sky130_fd_sc_hd__or4_1 _457_ (.A(_087_),
    .B(_108_),
    .C(_162_),
    .D(_163_),
    .X(_164_));
 sky130_fd_sc_hd__or2_1 _458_ (.A(_161_),
    .B(_164_),
    .X(_165_));
 sky130_fd_sc_hd__a22o_1 _459_ (.A1(net56),
    .A2(net69),
    .B1(net25),
    .B2(_165_),
    .X(_009_));
 sky130_fd_sc_hd__or4_1 _460_ (.A(_217_),
    .B(_021_),
    .C(_024_),
    .D(_060_),
    .X(_166_));
 sky130_fd_sc_hd__or4_1 _461_ (.A(_202_),
    .B(_211_),
    .C(_224_),
    .D(_166_),
    .X(_167_));
 sky130_fd_sc_hd__or4_1 _462_ (.A(_017_),
    .B(_047_),
    .C(_081_),
    .D(_099_),
    .X(_168_));
 sky130_fd_sc_hd__or4_1 _463_ (.A(_035_),
    .B(_066_),
    .C(_112_),
    .D(_168_),
    .X(_169_));
 sky130_fd_sc_hd__or3_1 _464_ (.A(_156_),
    .B(_167_),
    .C(_169_),
    .X(_170_));
 sky130_fd_sc_hd__a22o_1 _465_ (.A1(net57),
    .A2(net60),
    .B1(_085_),
    .B2(_170_),
    .X(_010_));
 sky130_fd_sc_hd__or2_1 _466_ (.A(_047_),
    .B(_064_),
    .X(_171_));
 sky130_fd_sc_hd__or3_1 _467_ (.A(_188_),
    .B(_016_),
    .C(_127_),
    .X(_172_));
 sky130_fd_sc_hd__or4_1 _468_ (.A(_224_),
    .B(_019_),
    .C(_022_),
    .D(_078_),
    .X(_173_));
 sky130_fd_sc_hd__or4_1 _469_ (.A(_126_),
    .B(_171_),
    .C(_172_),
    .D(_173_),
    .X(_174_));
 sky130_fd_sc_hd__or3_1 _470_ (.A(_042_),
    .B(_120_),
    .C(_174_),
    .X(_175_));
 sky130_fd_sc_hd__a22o_1 _471_ (.A1(net57),
    .A2(net64),
    .B1(net25),
    .B2(_175_),
    .X(_011_));
 sky130_fd_sc_hd__or4_1 _472_ (.A(_202_),
    .B(_043_),
    .C(_044_),
    .D(_075_),
    .X(_176_));
 sky130_fd_sc_hd__or4_1 _473_ (.A(_055_),
    .B(_119_),
    .C(_128_),
    .D(_176_),
    .X(_177_));
 sky130_fd_sc_hd__or3_1 _474_ (.A(_026_),
    .B(_042_),
    .C(_177_),
    .X(_178_));
 sky130_fd_sc_hd__a22o_1 _475_ (.A1(net56),
    .A2(net68),
    .B1(net25),
    .B2(_178_),
    .X(_012_));
 sky130_fd_sc_hd__or3_1 _476_ (.A(_193_),
    .B(_197_),
    .C(_067_),
    .X(_179_));
 sky130_fd_sc_hd__nor3_1 _477_ (.A(_213_),
    .B(_020_),
    .C(_179_),
    .Y(_180_));
 sky130_fd_sc_hd__nand3_1 _478_ (.A(_056_),
    .B(_065_),
    .C(_180_),
    .Y(_181_));
 sky130_fd_sc_hd__a22o_1 _479_ (.A1(net56),
    .A2(net71),
    .B1(net25),
    .B2(_181_),
    .X(_013_));
 sky130_fd_sc_hd__o21ba_1 _480_ (.A1(net8),
    .A2(net58),
    .B1_N(_084_),
    .X(_014_));
 sky130_fd_sc_hd__a21o_1 _481_ (.A1(net56),
    .A2(net59),
    .B1(_027_),
    .X(_015_));
 sky130_fd_sc_hd__dfxtp_1 _482_ (.CLK(clknet_1_0__leaf_clk0),
    .D(net1),
    .Q(\addr0_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _483_ (.CLK(clknet_1_0__leaf_clk0),
    .D(net2),
    .Q(\addr0_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _484_ (.CLK(clknet_1_0__leaf_clk0),
    .D(net3),
    .Q(\addr0_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _485_ (.CLK(clknet_1_0__leaf_clk0),
    .D(net4),
    .Q(\addr0_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _486_ (.CLK(clknet_1_0__leaf_clk0),
    .D(net5),
    .Q(\addr0_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _487_ (.CLK(clknet_1_0__leaf_clk0),
    .D(net6),
    .Q(\addr0_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _488_ (.CLK(clknet_1_0__leaf_clk0),
    .D(net7),
    .Q(\addr0_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _489_ (.CLK(clknet_1_0__leaf_clk0),
    .D(_000_),
    .Q(net9));
 sky130_fd_sc_hd__dfxtp_1 _490_ (.CLK(clknet_1_1__leaf_clk0),
    .D(_001_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_1 _491_ (.CLK(clknet_1_1__leaf_clk0),
    .D(_002_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_1 _492_ (.CLK(clknet_1_1__leaf_clk0),
    .D(_003_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_1 _493_ (.CLK(clknet_1_1__leaf_clk0),
    .D(_004_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_1 _494_ (.CLK(clknet_1_1__leaf_clk0),
    .D(_005_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_1 _495_ (.CLK(clknet_1_1__leaf_clk0),
    .D(_006_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_1 _496_ (.CLK(clknet_1_0__leaf_clk0),
    .D(_007_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_1 _497_ (.CLK(clknet_1_1__leaf_clk0),
    .D(_008_),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_1 _498_ (.CLK(clknet_1_0__leaf_clk0),
    .D(_009_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_1 _499_ (.CLK(clknet_1_1__leaf_clk0),
    .D(_010_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_1 _500_ (.CLK(clknet_1_1__leaf_clk0),
    .D(_011_),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_1 _501_ (.CLK(clknet_1_1__leaf_clk0),
    .D(_012_),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_1 _502_ (.CLK(clknet_1_0__leaf_clk0),
    .D(_013_),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_1 _503_ (.CLK(clknet_1_0__leaf_clk0),
    .D(_014_),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_1 _504_ (.CLK(clknet_1_0__leaf_clk0),
    .D(_015_),
    .Q(net15));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_150 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(addr0[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(addr0[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(addr0[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(addr0[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(addr0[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(addr0[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(addr0[6]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(cs0),
    .X(net8));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(dout0[0]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(dout0[10]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(dout0[11]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(dout0[12]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(dout0[13]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(dout0[14]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(dout0[15]));
 sky130_fd_sc_hd__clkbuf_4 output16 (.A(net16),
    .X(dout0[1]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(dout0[2]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(dout0[3]));
 sky130_fd_sc_hd__clkbuf_4 output19 (.A(net19),
    .X(dout0[4]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(dout0[5]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(dout0[6]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(dout0[7]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(dout0[8]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(dout0[9]));
 sky130_fd_sc_hd__buf_2 fanout25 (.A(_085_),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 wire26 (.A(_083_),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(_058_),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 fanout28 (.A(_058_),
    .X(net28));
 sky130_fd_sc_hd__buf_2 fanout29 (.A(_057_),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 fanout30 (.A(_057_),
    .X(net30));
 sky130_fd_sc_hd__buf_2 fanout31 (.A(_029_),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout32 (.A(_029_),
    .X(net32));
 sky130_fd_sc_hd__buf_2 fanout33 (.A(_028_),
    .X(net33));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout34 (.A(_028_),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 max_cap35 (.A(_223_),
    .X(net35));
 sky130_fd_sc_hd__buf_1 max_cap36 (.A(_208_),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(_205_),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 fanout38 (.A(_205_),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 max_cap39 (.A(_204_),
    .X(net39));
 sky130_fd_sc_hd__buf_2 fanout40 (.A(_203_),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 fanout41 (.A(_203_),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 max_cap42 (.A(_199_),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 fanout44 (.A(_186_),
    .X(net44));
 sky130_fd_sc_hd__buf_2 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 fanout46 (.A(_183_),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 fanout47 (.A(\addr0_reg[4] ),
    .X(net47));
 sky130_fd_sc_hd__buf_2 fanout48 (.A(\addr0_reg[3] ),
    .X(net48));
 sky130_fd_sc_hd__buf_1 fanout49 (.A(\addr0_reg[3] ),
    .X(net49));
 sky130_fd_sc_hd__buf_2 fanout50 (.A(\addr0_reg[2] ),
    .X(net50));
 sky130_fd_sc_hd__buf_1 fanout51 (.A(\addr0_reg[2] ),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 fanout52 (.A(\addr0_reg[1] ),
    .X(net52));
 sky130_fd_sc_hd__buf_1 fanout53 (.A(\addr0_reg[1] ),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 fanout54 (.A(\addr0_reg[0] ),
    .X(net54));
 sky130_fd_sc_hd__buf_1 fanout55 (.A(\addr0_reg[0] ),
    .X(net55));
 sky130_fd_sc_hd__buf_2 fanout56 (.A(_182_),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 fanout57 (.A(_182_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk0 (.A(clk0),
    .X(clknet_0_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_1_0__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_1_1__leaf_clk0));
 sky130_fd_sc_hd__clkinv_2 clkload0 (.A(clknet_1_1__leaf_clk0));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net14),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net15),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net10),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net18),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net17),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net21),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net11),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net20),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net22),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net23),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net12),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net24),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net16),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net13),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net9),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net19),
    .X(net73));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_173 ();
endmodule
