VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rom7
  CLASS BLOCK ;
  FOREIGN rom7 ;
  ORIGIN 0.000 0.000 ;
  SIZE 260.000 BY 260.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 247.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 247.760 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 247.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 247.760 ;
    END
  END VPWR
  PIN addr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 37.440 260.000 38.040 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 40.840 260.000 41.440 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 256.000 44.240 260.000 44.840 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 47.640 260.000 48.240 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 51.040 260.000 51.640 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 54.440 260.000 55.040 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END addr0[8]
  PIN clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END clk0
  PIN dout0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 102.040 260.000 102.640 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 61.240 260.000 61.840 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 105.440 260.000 106.040 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 136.040 260.000 136.640 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 122.450 256.000 122.730 260.000 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 190.440 260.000 191.040 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 173.970 256.000 174.250 260.000 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 183.630 256.000 183.910 260.000 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 199.730 256.000 200.010 260.000 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 148.210 256.000 148.490 260.000 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 96.690 256.000 96.970 260.000 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 116.010 256.000 116.290 260.000 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 109.570 256.000 109.850 260.000 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 80.590 256.000 80.870 260.000 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 70.930 256.000 71.210 260.000 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 64.490 256.000 64.770 260.000 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 256.000 158.150 260.000 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.000 17.040 260.000 17.640 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END dout0[31]
  PIN dout0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 132.640 260.000 133.240 ;
    END
  END dout0[3]
  PIN dout0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END dout0[4]
  PIN dout0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END dout0[5]
  PIN dout0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END dout0[9]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 254.570 247.710 ;
      LAYER li1 ;
        RECT 5.520 10.795 254.380 247.605 ;
      LAYER met1 ;
        RECT 2.370 10.640 254.380 249.180 ;
      LAYER met2 ;
        RECT 2.390 255.720 64.210 256.770 ;
        RECT 65.050 255.720 70.650 256.770 ;
        RECT 71.490 255.720 80.310 256.770 ;
        RECT 81.150 255.720 96.410 256.770 ;
        RECT 97.250 255.720 109.290 256.770 ;
        RECT 110.130 255.720 115.730 256.770 ;
        RECT 116.570 255.720 122.170 256.770 ;
        RECT 123.010 255.720 147.930 256.770 ;
        RECT 148.770 255.720 157.590 256.770 ;
        RECT 158.430 255.720 173.690 256.770 ;
        RECT 174.530 255.720 183.350 256.770 ;
        RECT 184.190 255.720 199.450 256.770 ;
        RECT 200.290 255.720 252.910 256.770 ;
        RECT 2.390 4.280 252.910 255.720 ;
        RECT 2.390 4.000 51.330 4.280 ;
        RECT 52.170 4.000 54.550 4.280 ;
        RECT 55.390 4.000 57.770 4.280 ;
        RECT 58.610 4.000 131.830 4.280 ;
        RECT 132.670 4.000 189.790 4.280 ;
        RECT 190.630 4.000 234.870 4.280 ;
        RECT 235.710 4.000 252.910 4.280 ;
      LAYER met3 ;
        RECT 2.365 232.240 256.000 251.425 ;
        RECT 4.400 230.840 256.000 232.240 ;
        RECT 2.365 218.640 256.000 230.840 ;
        RECT 4.400 217.240 256.000 218.640 ;
        RECT 2.365 215.240 256.000 217.240 ;
        RECT 4.400 213.840 256.000 215.240 ;
        RECT 2.365 198.240 256.000 213.840 ;
        RECT 4.400 196.840 256.000 198.240 ;
        RECT 2.365 191.440 256.000 196.840 ;
        RECT 2.365 190.040 255.600 191.440 ;
        RECT 2.365 160.840 256.000 190.040 ;
        RECT 4.400 159.440 256.000 160.840 ;
        RECT 2.365 154.040 256.000 159.440 ;
        RECT 4.400 152.640 256.000 154.040 ;
        RECT 2.365 137.040 256.000 152.640 ;
        RECT 2.365 135.640 255.600 137.040 ;
        RECT 2.365 133.640 256.000 135.640 ;
        RECT 4.400 132.240 255.600 133.640 ;
        RECT 2.365 120.040 256.000 132.240 ;
        RECT 4.400 118.640 256.000 120.040 ;
        RECT 2.365 113.240 256.000 118.640 ;
        RECT 4.400 111.840 256.000 113.240 ;
        RECT 2.365 106.440 256.000 111.840 ;
        RECT 2.365 105.040 255.600 106.440 ;
        RECT 2.365 103.040 256.000 105.040 ;
        RECT 2.365 101.640 255.600 103.040 ;
        RECT 2.365 99.640 256.000 101.640 ;
        RECT 4.400 98.240 256.000 99.640 ;
        RECT 2.365 75.840 256.000 98.240 ;
        RECT 4.400 74.440 256.000 75.840 ;
        RECT 2.365 62.240 256.000 74.440 ;
        RECT 2.365 60.840 255.600 62.240 ;
        RECT 2.365 55.440 256.000 60.840 ;
        RECT 2.365 54.040 255.600 55.440 ;
        RECT 2.365 52.040 256.000 54.040 ;
        RECT 2.365 50.640 255.600 52.040 ;
        RECT 2.365 48.640 256.000 50.640 ;
        RECT 2.365 47.240 255.600 48.640 ;
        RECT 2.365 45.240 256.000 47.240 ;
        RECT 2.365 43.840 255.600 45.240 ;
        RECT 2.365 41.840 256.000 43.840 ;
        RECT 2.365 40.440 255.600 41.840 ;
        RECT 2.365 38.440 256.000 40.440 ;
        RECT 2.365 37.040 255.600 38.440 ;
        RECT 2.365 18.040 256.000 37.040 ;
        RECT 2.365 16.640 255.600 18.040 ;
        RECT 2.365 10.715 256.000 16.640 ;
      LAYER met4 ;
        RECT 3.055 248.160 244.425 251.425 ;
        RECT 3.055 17.855 20.640 248.160 ;
        RECT 23.040 17.855 23.940 248.160 ;
        RECT 26.340 17.855 174.240 248.160 ;
        RECT 176.640 17.855 177.540 248.160 ;
        RECT 179.940 17.855 244.425 248.160 ;
  END
END rom7
END LIBRARY

