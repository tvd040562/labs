assign table1[0] = 32'h00000000;
assign table1[1] = 32'hff36f170;
assign table1[2] = 32'hfe6deaa1;
assign table1[3] = 32'hfda4f351;
assign table1[4] = 32'hfcdc1342;
assign table1[5] = 32'hfc135231;
assign table1[6] = 32'hfb4ab7db;
assign table1[7] = 32'hfa824bfd;
assign table1[8] = 32'hf9ba1651;
assign table1[9] = 32'hf8f21e8e;
assign table1[10] = 32'hf82a6c6a;
assign table1[11] = 32'hf7630799;
assign table1[12] = 32'hf69bf7c9;
assign table1[13] = 32'hf5d544a7;
assign table1[14] = 32'hf50ef5de;
assign table1[15] = 32'hf4491311;
assign table1[16] = 32'hf383a3e2;
assign table1[17] = 32'hf2beafed;
assign table1[18] = 32'hf1fa3ecb;
assign table1[19] = 32'hf136580d;
assign table1[20] = 32'hf0730342;
assign table1[21] = 32'hefb047f2;
assign table1[22] = 32'heeee2d9d;
assign table1[23] = 32'hee2cbbc1;
assign table1[24] = 32'hed6bf9d1;
assign table1[25] = 32'hecabef3d;
assign table1[26] = 32'hebeca36c;
assign table1[27] = 32'heb2e1dbe;
assign table1[28] = 32'hea70658a;
assign table1[29] = 32'he9b38223;
assign table1[30] = 32'he8f77acf;
assign table1[31] = 32'he83c56cf;
assign table1[32] = 32'he7821d59;
assign table1[33] = 32'he6c8d59c;
assign table1[34] = 32'he61086bc;
assign table1[35] = 32'he55937d5;
assign table1[36] = 32'he4a2eff6;
assign table1[37] = 32'he3edb628;
assign table1[38] = 32'he3399167;
assign table1[39] = 32'he28688a4;
assign table1[40] = 32'he1d4a2c8;
assign table1[41] = 32'he123e6ad;
assign table1[42] = 32'he0745b24;
assign table1[43] = 32'hdfc606f1;
assign table1[44] = 32'hdf18f0ce;
assign table1[45] = 32'hde6d1f65;
assign table1[46] = 32'hddc29958;
assign table1[47] = 32'hdd196538;
assign table1[48] = 32'hdc71898d;
assign table1[49] = 32'hdbcb0cce;
assign table1[50] = 32'hdb25f566;
assign table1[51] = 32'hda8249b4;
assign table1[52] = 32'hd9e01006;
assign table1[53] = 32'hd93f4e9e;
assign table1[54] = 32'hd8a00bae;
assign table1[55] = 32'hd8024d59;
assign table1[56] = 32'hd76619b6;
assign table1[57] = 32'hd6cb76c9;
assign table1[58] = 32'hd6326a88;
assign table1[59] = 32'hd59afadb;
assign table1[60] = 32'hd5052d97;
assign table1[61] = 32'hd4710883;
assign table1[62] = 32'hd3de9156;
assign table1[63] = 32'hd34dcdb4;
assign table1[64] = 32'hd2bec333;
assign table1[65] = 32'hd2317756;
assign table1[66] = 32'hd1a5ef90;
assign table1[67] = 32'hd11c3142;
assign table1[68] = 32'hd09441bb;
assign table1[69] = 32'hd00e2639;
assign table1[70] = 32'hcf89e3e8;
assign table1[71] = 32'hcf077fe1;
assign table1[72] = 32'hce86ff2a;
assign table1[73] = 32'hce0866b8;
assign table1[74] = 32'hcd8bbb6d;
assign table1[75] = 32'hcd110216;
assign table1[76] = 32'hcc983f70;
assign table1[77] = 32'hcc217822;
assign table1[78] = 32'hcbacb0bf;
assign table1[79] = 32'hcb39edca;
assign table1[80] = 32'hcac933ae;
assign table1[81] = 32'hca5a86c4;
assign table1[82] = 32'hc9edeb50;
assign table1[83] = 32'hc9836582;
assign table1[84] = 32'hc91af976;
assign table1[85] = 32'hc8b4ab32;
assign table1[86] = 32'hc8507ea7;
assign table1[87] = 32'hc7ee77b3;
assign table1[88] = 32'hc78e9a1d;
assign table1[89] = 32'hc730e997;
assign table1[90] = 32'hc6d569be;
assign table1[91] = 32'hc67c1e18;
assign table1[92] = 32'hc6250a18;
assign table1[93] = 32'hc5d03118;
assign table1[94] = 32'hc57d965d;
assign table1[95] = 32'hc52d3d18;
assign table1[96] = 32'hc4df2862;
assign table1[97] = 32'hc4935b3c;
assign table1[98] = 32'hc449d892;
assign table1[99] = 32'hc402a33c;
assign table1[100] = 32'hc3bdbdf6;
assign table1[101] = 32'hc37b2b6a;
assign table1[102] = 32'hc33aee27;
assign table1[103] = 32'hc2fd08a9;
assign table1[104] = 32'hc2c17d52;
assign table1[105] = 32'hc2884e6e;
assign table1[106] = 32'hc2517e31;
assign table1[107] = 32'hc21d0eb8;
assign table1[108] = 32'hc1eb0209;
assign table1[109] = 32'hc1bb5a11;
assign table1[110] = 32'hc18e18a7;
assign table1[111] = 32'hc1633f8a;
assign table1[112] = 32'hc13ad060;
assign table1[113] = 32'hc114ccb9;
assign table1[114] = 32'hc0f1360b;
assign table1[115] = 32'hc0d00db6;
assign table1[116] = 32'hc0b15502;
assign table1[117] = 32'hc0950d1d;
assign table1[118] = 32'hc07b371e;
assign table1[119] = 32'hc063d405;
assign table1[120] = 32'hc04ee4b8;
assign table1[121] = 32'hc03c6a07;
assign table1[122] = 32'hc02c64a6;
assign table1[123] = 32'hc01ed535;
assign table1[124] = 32'hc013bc39;
assign table1[125] = 32'hc00b1a20;
assign table1[126] = 32'hc004ef3f;
assign table1[127] = 32'hc0013bd3;
assign table1[128] = 32'hc0000000;
assign table1[129] = 32'hc0013bd3;
assign table1[130] = 32'hc004ef3f;
assign table1[131] = 32'hc00b1a20;
assign table1[132] = 32'hc013bc39;
assign table1[133] = 32'hc01ed535;
assign table1[134] = 32'hc02c64a6;
assign table1[135] = 32'hc03c6a07;
assign table1[136] = 32'hc04ee4b8;
assign table1[137] = 32'hc063d405;
assign table1[138] = 32'hc07b371e;
assign table1[139] = 32'hc0950d1d;
assign table1[140] = 32'hc0b15502;
assign table1[141] = 32'hc0d00db6;
assign table1[142] = 32'hc0f1360b;
assign table1[143] = 32'hc114ccb9;
assign table1[144] = 32'hc13ad060;
assign table1[145] = 32'hc1633f8a;
assign table1[146] = 32'hc18e18a7;
assign table1[147] = 32'hc1bb5a11;
assign table1[148] = 32'hc1eb0209;
assign table1[149] = 32'hc21d0eb8;
assign table1[150] = 32'hc2517e31;
assign table1[151] = 32'hc2884e6e;
assign table1[152] = 32'hc2c17d52;
assign table1[153] = 32'hc2fd08a9;
assign table1[154] = 32'hc33aee27;
assign table1[155] = 32'hc37b2b6a;
assign table1[156] = 32'hc3bdbdf6;
assign table1[157] = 32'hc402a33c;
assign table1[158] = 32'hc449d892;
assign table1[159] = 32'hc4935b3c;
assign table1[160] = 32'hc4df2862;
assign table1[161] = 32'hc52d3d18;
assign table1[162] = 32'hc57d965d;
assign table1[163] = 32'hc5d03118;
assign table1[164] = 32'hc6250a18;
assign table1[165] = 32'hc67c1e18;
assign table1[166] = 32'hc6d569be;
assign table1[167] = 32'hc730e997;
assign table1[168] = 32'hc78e9a1d;
assign table1[169] = 32'hc7ee77b3;
assign table1[170] = 32'hc8507ea7;
assign table1[171] = 32'hc8b4ab32;
assign table1[172] = 32'hc91af976;
assign table1[173] = 32'hc9836582;
assign table1[174] = 32'hc9edeb50;
assign table1[175] = 32'hca5a86c4;
assign table1[176] = 32'hcac933ae;
assign table1[177] = 32'hcb39edca;
assign table1[178] = 32'hcbacb0bf;
assign table1[179] = 32'hcc217822;
assign table1[180] = 32'hcc983f70;
assign table1[181] = 32'hcd110216;
assign table1[182] = 32'hcd8bbb6d;
assign table1[183] = 32'hce0866b8;
assign table1[184] = 32'hce86ff2a;
assign table1[185] = 32'hcf077fe1;
assign table1[186] = 32'hcf89e3e8;
assign table1[187] = 32'hd00e2639;
assign table1[188] = 32'hd09441bb;
assign table1[189] = 32'hd11c3142;
assign table1[190] = 32'hd1a5ef90;
assign table1[191] = 32'hd2317756;
assign table1[192] = 32'hd2bec333;
assign table1[193] = 32'hd34dcdb4;
assign table1[194] = 32'hd3de9156;
assign table1[195] = 32'hd4710883;
assign table1[196] = 32'hd5052d97;
assign table1[197] = 32'hd59afadb;
assign table1[198] = 32'hd6326a88;
assign table1[199] = 32'hd6cb76c9;
assign table1[200] = 32'hd76619b6;
assign table1[201] = 32'hd8024d59;
assign table1[202] = 32'hd8a00bae;
assign table1[203] = 32'hd93f4e9e;
assign table1[204] = 32'hd9e01006;
assign table1[205] = 32'hda8249b4;
assign table1[206] = 32'hdb25f566;
assign table1[207] = 32'hdbcb0cce;
assign table1[208] = 32'hdc71898d;
assign table1[209] = 32'hdd196538;
assign table1[210] = 32'hddc29958;
assign table1[211] = 32'hde6d1f65;
assign table1[212] = 32'hdf18f0ce;
assign table1[213] = 32'hdfc606f1;
assign table1[214] = 32'he0745b24;
assign table1[215] = 32'he123e6ad;
assign table1[216] = 32'he1d4a2c8;
assign table1[217] = 32'he28688a4;
assign table1[218] = 32'he3399167;
assign table1[219] = 32'he3edb628;
assign table1[220] = 32'he4a2eff6;
assign table1[221] = 32'he55937d5;
assign table1[222] = 32'he61086bc;
assign table1[223] = 32'he6c8d59c;
assign table1[224] = 32'he7821d59;
assign table1[225] = 32'he83c56cf;
assign table1[226] = 32'he8f77acf;
assign table1[227] = 32'he9b38223;
assign table1[228] = 32'hea70658a;
assign table1[229] = 32'heb2e1dbe;
assign table1[230] = 32'hebeca36c;
assign table1[231] = 32'hecabef3d;
assign table1[232] = 32'hed6bf9d1;
assign table1[233] = 32'hee2cbbc1;
assign table1[234] = 32'heeee2d9d;
assign table1[235] = 32'hefb047f2;
assign table1[236] = 32'hf0730342;
assign table1[237] = 32'hf136580d;
assign table1[238] = 32'hf1fa3ecb;
assign table1[239] = 32'hf2beafed;
assign table1[240] = 32'hf383a3e2;
assign table1[241] = 32'hf4491311;
assign table1[242] = 32'hf50ef5de;
assign table1[243] = 32'hf5d544a7;
assign table1[244] = 32'hf69bf7c9;
assign table1[245] = 32'hf7630799;
assign table1[246] = 32'hf82a6c6a;
assign table1[247] = 32'hf8f21e8e;
assign table1[248] = 32'hf9ba1651;
assign table1[249] = 32'hfa824bfd;
assign table1[250] = 32'hfb4ab7db;
assign table1[251] = 32'hfc135231;
assign table1[252] = 32'hfcdc1342;
assign table1[253] = 32'hfda4f351;
assign table1[254] = 32'hfe6deaa1;
assign table1[255] = 32'hff36f170;
