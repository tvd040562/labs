VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rom6
  CLASS BLOCK ;
  FOREIGN rom6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 260.000 BY 260.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 247.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 247.760 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 247.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 247.760 ;
    END
  END VPWR
  PIN addr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 37.440 260.000 38.040 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 40.840 260.000 41.440 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 44.240 260.000 44.840 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 256.000 47.640 260.000 48.240 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 256.000 51.040 260.000 51.640 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 54.440 260.000 55.040 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 215.830 256.000 216.110 260.000 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 212.610 256.000 212.890 260.000 ;
    END
  END addr0[8]
  PIN clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END clk0
  PIN dout0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 156.440 260.000 157.040 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 95.240 260.000 95.840 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 122.440 260.000 123.040 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 190.070 256.000 190.350 260.000 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 105.440 260.000 106.040 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 200.640 260.000 201.240 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 167.530 256.000 167.810 260.000 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 187.040 260.000 187.640 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 180.410 256.000 180.690 260.000 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 122.450 256.000 122.730 260.000 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 103.130 256.000 103.410 260.000 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 70.930 256.000 71.210 260.000 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 87.030 256.000 87.310 260.000 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 51.610 256.000 51.890 260.000 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 256.000 55.110 260.000 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.000 210.840 260.000 211.440 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.000 241.440 260.000 242.040 ;
    END
  END dout0[31]
  PIN dout0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 99.910 256.000 100.190 260.000 ;
    END
  END dout0[3]
  PIN dout0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 256.000 98.640 260.000 99.240 ;
    END
  END dout0[4]
  PIN dout0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END dout0[5]
  PIN dout0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END dout0[9]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 254.570 247.710 ;
      LAYER li1 ;
        RECT 5.520 10.795 254.380 247.605 ;
      LAYER met1 ;
        RECT 1.910 10.240 257.070 249.860 ;
      LAYER met2 ;
        RECT 1.930 255.720 51.330 256.770 ;
        RECT 52.170 255.720 54.550 256.770 ;
        RECT 55.390 255.720 70.650 256.770 ;
        RECT 71.490 255.720 86.750 256.770 ;
        RECT 87.590 255.720 99.630 256.770 ;
        RECT 100.470 255.720 102.850 256.770 ;
        RECT 103.690 255.720 122.170 256.770 ;
        RECT 123.010 255.720 167.250 256.770 ;
        RECT 168.090 255.720 180.130 256.770 ;
        RECT 180.970 255.720 189.790 256.770 ;
        RECT 190.630 255.720 212.330 256.770 ;
        RECT 213.170 255.720 215.550 256.770 ;
        RECT 216.390 255.720 257.050 256.770 ;
        RECT 1.930 4.280 257.050 255.720 ;
        RECT 1.930 4.000 83.530 4.280 ;
        RECT 84.370 4.000 167.250 4.280 ;
        RECT 168.090 4.000 199.450 4.280 ;
        RECT 200.290 4.000 257.050 4.280 ;
      LAYER met3 ;
        RECT 1.905 242.440 257.075 250.740 ;
        RECT 1.905 241.040 255.600 242.440 ;
        RECT 1.905 228.840 257.075 241.040 ;
        RECT 4.400 227.440 257.075 228.840 ;
        RECT 1.905 218.640 257.075 227.440 ;
        RECT 4.400 217.240 257.075 218.640 ;
        RECT 1.905 211.840 257.075 217.240 ;
        RECT 1.905 210.440 255.600 211.840 ;
        RECT 1.905 208.440 257.075 210.440 ;
        RECT 4.400 207.040 257.075 208.440 ;
        RECT 1.905 201.640 257.075 207.040 ;
        RECT 1.905 200.240 255.600 201.640 ;
        RECT 1.905 188.040 257.075 200.240 ;
        RECT 1.905 186.640 255.600 188.040 ;
        RECT 1.905 160.840 257.075 186.640 ;
        RECT 4.400 159.440 257.075 160.840 ;
        RECT 1.905 157.440 257.075 159.440 ;
        RECT 1.905 156.040 255.600 157.440 ;
        RECT 1.905 140.440 257.075 156.040 ;
        RECT 4.400 139.040 257.075 140.440 ;
        RECT 1.905 137.040 257.075 139.040 ;
        RECT 4.400 135.640 257.075 137.040 ;
        RECT 1.905 126.840 257.075 135.640 ;
        RECT 4.400 125.440 257.075 126.840 ;
        RECT 1.905 123.440 257.075 125.440 ;
        RECT 1.905 122.040 255.600 123.440 ;
        RECT 1.905 106.440 257.075 122.040 ;
        RECT 4.400 105.040 255.600 106.440 ;
        RECT 1.905 99.640 257.075 105.040 ;
        RECT 1.905 98.240 255.600 99.640 ;
        RECT 1.905 96.240 257.075 98.240 ;
        RECT 4.400 94.840 255.600 96.240 ;
        RECT 1.905 82.640 257.075 94.840 ;
        RECT 4.400 81.240 257.075 82.640 ;
        RECT 1.905 75.840 257.075 81.240 ;
        RECT 4.400 74.440 257.075 75.840 ;
        RECT 1.905 62.240 257.075 74.440 ;
        RECT 4.400 60.840 257.075 62.240 ;
        RECT 1.905 55.440 257.075 60.840 ;
        RECT 1.905 54.040 255.600 55.440 ;
        RECT 1.905 52.040 257.075 54.040 ;
        RECT 1.905 50.640 255.600 52.040 ;
        RECT 1.905 48.640 257.075 50.640 ;
        RECT 1.905 47.240 255.600 48.640 ;
        RECT 1.905 45.240 257.075 47.240 ;
        RECT 1.905 43.840 255.600 45.240 ;
        RECT 1.905 41.840 257.075 43.840 ;
        RECT 1.905 40.440 255.600 41.840 ;
        RECT 1.905 38.440 257.075 40.440 ;
        RECT 1.905 37.040 255.600 38.440 ;
        RECT 1.905 8.335 257.075 37.040 ;
      LAYER met4 ;
        RECT 3.055 248.160 246.265 250.745 ;
        RECT 3.055 10.240 20.640 248.160 ;
        RECT 23.040 10.240 23.940 248.160 ;
        RECT 26.340 10.240 174.240 248.160 ;
        RECT 176.640 10.240 177.540 248.160 ;
        RECT 179.940 10.240 246.265 248.160 ;
        RECT 3.055 8.335 246.265 10.240 ;
  END
END rom6
END LIBRARY

