logic [0:(ROM_DEPTH/2)-1] [DATA_WIDTH-1:0] table1 = {
32'h00000000,
32'h00c90e90,
32'h0192155f,
32'h025b0caf,
32'h0323ecbe,
32'h03ecadcf,
32'h04b54825,
32'h057db403,
32'h0645e9af,
32'h070de172,
32'h07d59396,
32'h089cf867,
32'h09640837,
32'h0a2abb59,
32'h0af10a22,
32'h0bb6ecef,
32'h0c7c5c1e,
32'h0d415013,
32'h0e05c135,
32'h0ec9a7f3,
32'h0f8cfcbe,
32'h104fb80e,
32'h1111d263,
32'h11d3443f,
32'h1294062f,
32'h135410c3,
32'h14135c94,
32'h14d1e242,
32'h158f9a76,
32'h164c7ddd,
32'h17088531,
32'h17c3a931,
32'h187de2a7,
32'h19372a64,
32'h19ef7944,
32'h1aa6c82b,
32'h1b5d100a,
32'h1c1249d8,
32'h1cc66e99,
32'h1d79775c,
32'h1e2b5d38,
32'h1edc1953,
32'h1f8ba4dc,
32'h2039f90f,
32'h20e70f32,
32'h2192e09b,
32'h223d66a8,
32'h22e69ac8,
32'h238e7673,
32'h2434f332,
32'h24da0a9a,
32'h257db64c,
32'h261feffa,
32'h26c0b162,
32'h275ff452,
32'h27fdb2a7,
32'h2899e64a,
32'h29348937,
32'h29cd9578,
32'h2a650525,
32'h2afad269,
32'h2b8ef77d,
32'h2c216eaa,
32'h2cb2324c,
32'h2d413ccd,
32'h2dce88aa,
32'h2e5a1070,
32'h2ee3cebe,
32'h2f6bbe45,
32'h2ff1d9c7,
32'h30761c18,
32'h30f8801f,
32'h317900d6,
32'h31f79948,
32'h32744493,
32'h32eefdea,
32'h3367c090,
32'h33de87de,
32'h34534f41,
32'h34c61236,
32'h3536cc52,
32'h35a5793c,
32'h361214b0,
32'h367c9a7e,
32'h36e5068a,
32'h374b54ce,
32'h37af8159,
32'h3811884d,
32'h387165e3,
32'h38cf1669,
32'h392a9642,
32'h3983e1e8,
32'h39daf5e8,
32'h3a2fcee8,
32'h3a8269a3,
32'h3ad2c2e8,
32'h3b20d79e,
32'h3b6ca4c4,
32'h3bb6276e,
32'h3bfd5cc4,
32'h3c42420a,
32'h3c84d496,
32'h3cc511d9,
32'h3d02f757,
32'h3d3e82ae,
32'h3d77b192,
32'h3dae81cf,
32'h3de2f148,
32'h3e14fdf7,
32'h3e44a5ef,
32'h3e71e759,
32'h3e9cc076,
32'h3ec52fa0,
32'h3eeb3347,
32'h3f0ec9f5,
32'h3f2ff24a,
32'h3f4eaafe,
32'h3f6af2e3,
32'h3f84c8e2,
32'h3f9c2bfb,
32'h3fb11b48,
32'h3fc395f9,
32'h3fd39b5a,
32'h3fe12acb,
32'h3fec43c7,
32'h3ff4e5e0,
32'h3ffb10c1,
32'h3ffec42d,
32'h40000000,
32'h3ffec42d,
32'h3ffb10c1,
32'h3ff4e5e0,
32'h3fec43c7,
32'h3fe12acb,
32'h3fd39b5a,
32'h3fc395f9,
32'h3fb11b48,
32'h3f9c2bfb,
32'h3f84c8e2,
32'h3f6af2e3,
32'h3f4eaafe,
32'h3f2ff24a,
32'h3f0ec9f5,
32'h3eeb3347,
32'h3ec52fa0,
32'h3e9cc076,
32'h3e71e759,
32'h3e44a5ef,
32'h3e14fdf7,
32'h3de2f148,
32'h3dae81cf,
32'h3d77b192,
32'h3d3e82ae,
32'h3d02f757,
32'h3cc511d9,
32'h3c84d496,
32'h3c42420a,
32'h3bfd5cc4,
32'h3bb6276e,
32'h3b6ca4c4,
32'h3b20d79e,
32'h3ad2c2e8,
32'h3a8269a3,
32'h3a2fcee8,
32'h39daf5e8,
32'h3983e1e8,
32'h392a9642,
32'h38cf1669,
32'h387165e3,
32'h3811884d,
32'h37af8159,
32'h374b54ce,
32'h36e5068a,
32'h367c9a7e,
32'h361214b0,
32'h35a5793c,
32'h3536cc52,
32'h34c61236,
32'h34534f41,
32'h33de87de,
32'h3367c090,
32'h32eefdea,
32'h32744493,
32'h31f79948,
32'h317900d6,
32'h30f8801f,
32'h30761c18,
32'h2ff1d9c7,
32'h2f6bbe45,
32'h2ee3cebe,
32'h2e5a1070,
32'h2dce88aa,
32'h2d413ccd,
32'h2cb2324c,
32'h2c216eaa,
32'h2b8ef77d,
32'h2afad269,
32'h2a650525,
32'h29cd9578,
32'h29348937,
32'h2899e64a,
32'h27fdb2a7,
32'h275ff452,
32'h26c0b162,
32'h261feffa,
32'h257db64c,
32'h24da0a9a,
32'h2434f332,
32'h238e7673,
32'h22e69ac8,
32'h223d66a8,
32'h2192e09b,
32'h20e70f32,
32'h2039f90f,
32'h1f8ba4dc,
32'h1edc1953,
32'h1e2b5d38,
32'h1d79775c,
32'h1cc66e99,
32'h1c1249d8,
32'h1b5d100a,
32'h1aa6c82b,
32'h19ef7944,
32'h19372a64,
32'h187de2a7,
32'h17c3a931,
32'h17088531,
32'h164c7ddd,
32'h158f9a76,
32'h14d1e242,
32'h14135c94,
32'h135410c3,
32'h1294062f,
32'h11d3443f,
32'h1111d263,
32'h104fb80e,
32'h0f8cfcbe,
32'h0ec9a7f3,
32'h0e05c135,
32'h0d415013,
32'h0c7c5c1e,
32'h0bb6ecef,
32'h0af10a22,
32'h0a2abb59,
32'h09640837,
32'h089cf867,
32'h07d59396,
32'h070de172,
32'h0645e9af,
32'h057db403,
32'h04b54825,
32'h03ecadcf,
32'h0323ecbe,
32'h025b0caf,
32'h0192155f,
32'h00c90e90
};
