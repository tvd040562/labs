logic [0:ROM_DEPTH-1] [DATA_WIDTH-1:0] table_ = {
32'hd2bec333,
32'hd2d08c33,
32'hd2e25c2b,
32'hd2f43318,
32'hd30610f7,
32'hd317f5c6,
32'hd329e181,
32'hd33bd427,
32'hd34dcdb4,
32'hd35fce26,
32'hd371d579,
32'hd383e3ab,
32'hd395f8ba,
32'hd3a814a2,
32'hd3ba3760,
32'hd3cc60f2,
32'hd3de9156,
32'hd3f0c887,
32'hd4030684,
32'hd4154b4a,
32'hd42796d5,
32'hd439e923,
32'hd44c4232,
32'hd45ea1fd,
32'hd4710883,
32'hd48375c1,
32'hd495e9b3,
32'hd4a86458,
32'hd4bae5ab,
32'hd4cd6dab,
32'hd4dffc54,
32'hd4f291a4,
32'hd5052d97,
32'hd517d02b,
32'hd52a795d,
32'hd53d292a,
32'hd54fdf8f,
32'hd5629c89,
32'hd5756016,
32'hd5882a32,
32'hd59afadb,
32'hd5add20d,
32'hd5c0afc6,
32'hd5d39403,
32'hd5e67ec1,
32'hd5f96ffd,
32'hd60c67b4,
32'hd61f65e4,
32'hd6326a88,
32'hd645759f,
32'hd6588725,
32'hd66b9f18,
32'hd67ebd74,
32'hd691e237,
32'hd6a50d5d,
32'hd6b83ee4,
32'hd6cb76c9,
32'hd6deb508,
32'hd6f1f99f,
32'hd705448b,
32'hd71895c9,
32'hd72bed55,
32'hd73f4b2e,
32'hd752af4f,
32'hd76619b6,
32'hd7798a60,
32'hd78d014a,
32'hd7a07e70,
32'hd7b401d1,
32'hd7c78b68,
32'hd7db1b34,
32'hd7eeb130,
32'hd8024d59,
32'hd815efae,
32'hd829982b,
32'hd83d46cc,
32'hd850fb8e,
32'hd864b670,
32'hd878776d,
32'hd88c3e83,
32'hd8a00bae,
32'hd8b3deeb,
32'hd8c7b838,
32'hd8db9792,
32'hd8ef7cf4,
32'hd903685d,
32'hd91759c9,
32'hd92b5135,
32'hd93f4e9e,
32'hd9535201,
32'hd9675b5a,
32'hd97b6aa8,
32'hd98f7fe6,
32'hd9a39b11,
32'hd9b7bc27,
32'hd9cbe325,
32'hd9e01006,
32'hd9f442c9,
32'hda087b69,
32'hda1cb9e5,
32'hda30fe38,
32'hda454860,
32'hda599859,
32'hda6dee21,
32'hda8249b4,
32'hda96ab0f,
32'hdaab122f,
32'hdabf7f11,
32'hdad3f1b1,
32'hdae86a0d,
32'hdafce821,
32'hdb116beb,
32'hdb25f566,
32'hdb3a8491,
32'hdb4f1967,
32'hdb63b3e5,
32'hdb785409,
32'hdb8cf9cf,
32'hdba1a534,
32'hdbb65634,
32'hdbcb0cce,
32'hdbdfc8fc,
32'hdbf48abd,
32'hdc09520d,
32'hdc1e1ee9,
32'hdc32f14d,
32'hdc47c936,
32'hdc5ca6a2,
32'hdc71898d,
32'hdc8671f3,
32'hdc9b5fd2,
32'hdcb05326,
32'hdcc54bec,
32'hdcda4a21,
32'hdcef4dc2,
32'hdd0456ca,
32'hdd196538,
32'hdd2e7908,
32'hdd439236,
32'hdd58b0c0,
32'hdd6dd4a2,
32'hdd82fdd8,
32'hdd982c60,
32'hddad6036,
32'hddc29958,
32'hddd7d7c1,
32'hdded1b6e,
32'hde02645d,
32'hde17b28a,
32'hde2d05f1,
32'hde425e8f,
32'hde57bc62,
32'hde6d1f65,
32'hde828796,
32'hde97f4f1,
32'hdead6773,
32'hdec2df18,
32'hded85bdd,
32'hdeedddc0,
32'hdf0364bc,
32'hdf18f0ce,
32'hdf2e81f3,
32'hdf441828,
32'hdf59b369,
32'hdf6f53b3,
32'hdf84f902,
32'hdf9aa354,
32'hdfb052a5,
32'hdfc606f1,
32'hdfdbc036,
32'hdff17e70,
32'he007419b,
32'he01d09b4,
32'he032d6b8,
32'he048a8a4,
32'he05e7f74,
32'he0745b24,
32'he08a3bb2,
32'he0a0211a,
32'he0b60b58,
32'he0cbfa6a,
32'he0e1ee4b,
32'he0f7e6f9,
32'he10de470,
32'he123e6ad,
32'he139edac,
32'he14ff96a,
32'he16609e3,
32'he17c1f15,
32'he19238fb,
32'he1a85793,
32'he1be7ad8,
32'he1d4a2c8,
32'he1eacf5f,
32'he2010099,
32'he2173674,
32'he22d70eb,
32'he243affc,
32'he259f3a3,
32'he2703bdc,
32'he28688a4,
32'he29cd9f8,
32'he2b32fd4,
32'he2c98a35,
32'he2dfe917,
32'he2f64c77,
32'he30cb451,
32'he32320a2,
32'he3399167,
32'he350069b,
32'he366803c,
32'he37cfe47,
32'he39380b6,
32'he3aa0788,
32'he3c092b9,
32'he3d72245,
32'he3edb628,
32'he4044e60,
32'he41aeae8,
32'he4318bbe,
32'he44830dd,
32'he45eda43,
32'he47587eb,
32'he48c39d3,
32'he4a2eff6,
32'he4b9aa52,
32'he4d068e2,
32'he4e72ba4,
32'he4fdf294,
32'he514bdad,
32'he52b8cee,
32'he5426051,
32'he55937d5,
32'he5701374,
32'he586f32c,
32'he59dd6f9,
32'he5b4bed8,
32'he5cbaac5,
32'he5e29abc,
32'he5f98ebb,
32'he61086bc,
32'he62782be,
32'he63e82bc,
32'he65586b3,
32'he66c8e9f,
32'he6839a7c,
32'he69aaa48,
32'he6b1bdff,
32'he6c8d59c,
32'he6dff11d,
32'he6f7107e,
32'he70e33bb,
32'he7255ad1,
32'he73c85bc,
32'he753b479,
32'he76ae704,
32'he7821d59,
32'he7995776,
32'he7b09555,
32'he7c7d6f4,
32'he7df1c50,
32'he7f66564,
32'he80db22d,
32'he82502a7,
32'he83c56cf,
32'he853aea1,
32'he86b0a1a,
32'he8826936,
32'he899cbf1,
32'he8b13248,
32'he8c89c37,
32'he8e009ba,
32'he8f77acf,
32'he90eef71,
32'he926679c,
32'he93de34e,
32'he9556282,
32'he96ce535,
32'he9846b63,
32'he99bf509,
32'he9b38223,
32'he9cb12ad,
32'he9e2a6a3,
32'he9fa3e03,
32'hea11d8c8,
32'hea2976ef,
32'hea411874,
32'hea58bd54,
32'hea70658a,
32'hea881114,
32'hea9fbfed,
32'heab77212,
32'heacf277f,
32'heae6e031,
32'heafe9c24,
32'heb165b54,
32'heb2e1dbe,
32'heb45e35d,
32'heb5dac2f,
32'heb75782f,
32'heb8d475b,
32'heba519ad,
32'hebbcef23,
32'hebd4c7ba,
32'hebeca36c,
32'hec048237,
32'hec1c6417,
32'hec344908,
32'hec4c3106,
32'hec641c0e,
32'hec7c0a1d,
32'hec93fb2e,
32'hecabef3d,
32'hecc3e648,
32'hecdbe04a,
32'hecf3dd3f,
32'hed0bdd25,
32'hed23dff7,
32'hed3be5b1,
32'hed53ee51,
32'hed6bf9d1,
32'hed84082f,
32'hed9c1967,
32'hedb42d74,
32'hedcc4454,
32'hede45e03,
32'hedfc7a7c,
32'hee1499bd,
32'hee2cbbc1,
32'hee44e084,
32'hee5d0804,
32'hee75323c,
32'hee8d5f29,
32'heea58ec6,
32'heebdc110,
32'heed5f604,
32'heeee2d9d,
32'hef0667d9,
32'hef1ea4b2,
32'hef36e426,
32'hef4f2630,
32'hef676ace,
32'hef7fb1fa,
32'hef97fbb2,
32'hefb047f2,
32'hefc896b5,
32'hefe0e7f9,
32'heff93bba,
32'hf01191f3,
32'hf029eaa1,
32'hf04245c0,
32'hf05aa34c,
32'hf0730342,
32'hf08b659f,
32'hf0a3ca5d,
32'hf0bc317a,
32'hf0d49af1,
32'hf0ed06bf,
32'hf10574e0,
32'hf11de551,
32'hf136580d,
32'hf14ecd11,
32'hf1674459,
32'hf17fbde2,
32'hf19839a6,
32'hf1b0b7a4,
32'hf1c937d6,
32'hf1e1ba3a,
32'hf1fa3ecb,
32'hf212c585,
32'hf22b4e66,
32'hf243d968,
32'hf25c6688,
32'hf274f5c3,
32'hf28d8715,
32'hf2a61a7a,
32'hf2beafed,
32'hf2d7476c,
32'hf2efe0f2,
32'hf3087c7d,
32'hf3211a07,
32'hf339b98d,
32'hf3525b0b,
32'hf36afe7e,
32'hf383a3e2,
32'hf39c4b32,
32'hf3b4f46c,
32'hf3cd9f8b,
32'hf3e64c8c,
32'hf3fefb6a,
32'hf417ac22,
32'hf4305eb0,
32'hf4491311,
32'hf461c940,
32'hf47a8139,
32'hf4933afa,
32'hf4abf67e,
32'hf4c4b3c0,
32'hf4dd72be,
32'hf4f63374,
32'hf50ef5de,
32'hf527b9f7,
32'hf5407fbd,
32'hf559472b,
32'hf572103d,
32'hf58adaf0,
32'hf5a3a740,
32'hf5bc7529,
32'hf5d544a7,
32'hf5ee15b7,
32'hf606e854,
32'hf61fbc7b,
32'hf6389228,
32'hf6516956,
32'hf66a4203,
32'hf6831c2b,
32'hf69bf7c9,
32'hf6b4d4d9,
32'hf6cdb359,
32'hf6e69344,
32'hf6ff7496,
32'hf718574b,
32'hf7313b60,
32'hf74a20d0,
32'hf7630799,
32'hf77befb5,
32'hf794d922,
32'hf7adc3db,
32'hf7c6afdc,
32'hf7df9d22,
32'hf7f88ba9,
32'hf8117b6d,
32'hf82a6c6a,
32'hf8435e9d,
32'hf85c5201,
32'hf8754692,
32'hf88e3c4d,
32'hf8a7332e,
32'hf8c02b31,
32'hf8d92452,
32'hf8f21e8e,
32'hf90b19e0,
32'hf9241645,
32'hf93d13b8,
32'hf9561237,
32'hf96f11bc,
32'hf9881245,
32'hf9a113cd,
32'hf9ba1651,
32'hf9d319cc,
32'hf9ec1e3b,
32'hfa05239a,
32'hfa1e29e5,
32'hfa373119,
32'hfa503930,
32'hfa694229,
32'hfa824bfd,
32'hfa9b56ab,
32'hfab4622d,
32'hfacd6e81,
32'hfae67ba2,
32'hfaff898c,
32'hfb18983b,
32'hfb31a7ac,
32'hfb4ab7db,
32'hfb63c8c4,
32'hfb7cda63,
32'hfb95ecb4,
32'hfbaeffb3,
32'hfbc8135c,
32'hfbe127ac,
32'hfbfa3c9f,
32'hfc135231,
32'hfc2c685d,
32'hfc457f21,
32'hfc5e9678,
32'hfc77ae5e,
32'hfc90c6cf,
32'hfca9dfc8,
32'hfcc2f945,
32'hfcdc1342,
32'hfcf52dbb,
32'hfd0e48ab,
32'hfd276410,
32'hfd407fe6,
32'hfd599c28,
32'hfd72b8d2,
32'hfd8bd5e1,
32'hfda4f351,
32'hfdbe111e,
32'hfdd72f45,
32'hfdf04dc0,
32'hfe096c8d,
32'hfe228ba7,
32'hfe3bab0b,
32'hfe54cab5,
32'hfe6deaa1,
32'hfe870aca,
32'hfea02b2e,
32'hfeb94bc8,
32'hfed26c94,
32'hfeeb8d8f,
32'hff04aeb5,
32'hff1dd001,
32'hff36f170,
32'hff5012fe,
32'hff6934a8,
32'hff825668,
32'hff9b783c,
32'hffb49a1f,
32'hffcdbc0f,
32'hffe6de05
};
