VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_256byte_1rw1r_32x64_8
   CLASS BLOCK ;
   SIZE 370.18 BY 261.11 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  100.54 0.0 100.92 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  106.38 0.0 106.76 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  112.22 0.0 112.6 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  118.06 0.0 118.44 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  123.9 0.0 124.28 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  129.74 0.0 130.12 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  135.58 0.0 135.96 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  141.42 0.0 141.8 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  147.26 0.0 147.64 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  153.1 0.0 153.48 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  158.94 0.0 159.32 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  164.78 0.0 165.16 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  170.62 0.0 171.0 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  176.46 0.0 176.84 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  182.3 0.0 182.68 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  188.14 0.0 188.52 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  193.98 0.0 194.36 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  199.82 0.0 200.2 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  205.66 0.0 206.04 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  211.5 0.0 211.88 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  217.34 0.0 217.72 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  223.18 0.0 223.56 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  229.02 0.0 229.4 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  234.86 0.0 235.24 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  240.7 0.0 241.08 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  246.54 0.0 246.92 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  252.38 0.0 252.76 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  258.22 0.0 258.6 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  264.06 0.0 264.44 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  269.9 0.0 270.28 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  275.74 0.0 276.12 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  281.58 0.0 281.96 0.38 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 109.585 0.38 109.965 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 117.985 0.38 118.365 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 123.85 0.38 124.23 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 132.35 0.38 132.73 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 137.99 0.38 138.37 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 146.49 0.38 146.87 ;
      END
   END addr0[5]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  369.8 72.47 370.18 72.85 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  369.8 63.97 370.18 64.35 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  307.76 0.0 308.14 0.38 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  304.785 0.0 305.165 0.38 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  305.475 0.0 305.855 0.38 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  306.22 0.0 306.6 0.38 ;
      END
   END addr1[5]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 16.73 0.38 17.11 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  369.8 245.86 370.18 246.24 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 25.23 0.38 25.61 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  31.1 0.0 31.48 0.38 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  339.54 260.73 339.92 261.11 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  77.18 0.0 77.56 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  83.02 0.0 83.4 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  88.86 0.0 89.24 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  94.7 0.0 95.08 0.38 ;
      END
   END wmask0[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  137.685 0.0 138.065 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  142.11 0.0 142.49 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  143.925 0.0 144.305 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  147.95 0.0 148.33 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  148.785 0.0 149.165 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  153.815 0.0 154.195 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.025 0.0 155.405 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  160.0 0.0 160.38 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  162.645 0.0 163.025 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.295 0.0 166.675 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.505 0.0 167.885 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.535 0.0 172.915 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  173.745 0.0 174.125 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.775 0.0 179.155 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  179.985 0.0 180.365 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.96 0.0 185.34 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  186.285 0.0 186.665 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.255 0.0 191.635 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.175 0.0 192.555 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.495 0.0 197.875 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  200.51 0.0 200.89 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.735 0.0 204.115 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  206.35 0.0 206.73 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  209.695 0.0 210.075 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  212.565 0.0 212.945 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  215.535 0.0 215.915 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  218.03 0.0 218.41 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  220.515 0.0 220.895 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  223.87 0.0 224.25 0.38 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  229.71 0.0 230.09 0.38 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  231.285 0.0 231.665 0.38 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  235.68 0.0 236.06 0.38 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  136.365 260.73 136.745 261.11 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  141.335 260.73 141.715 261.11 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  142.605 260.73 142.985 261.11 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  147.575 260.73 147.955 261.11 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  148.845 260.73 149.225 261.11 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  153.815 260.73 154.195 261.11 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.085 260.73 155.465 261.11 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  160.055 260.73 160.435 261.11 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  161.325 260.73 161.705 261.11 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.295 260.73 166.675 261.11 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.565 260.73 167.945 261.11 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.535 260.73 172.915 261.11 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  173.805 260.73 174.185 261.11 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.775 260.73 179.155 261.11 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.045 260.73 180.425 261.11 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  185.015 260.73 185.395 261.11 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  186.285 260.73 186.665 261.11 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.255 260.73 191.635 261.11 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.525 260.73 192.905 261.11 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.495 260.73 197.875 261.11 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  198.765 260.73 199.145 261.11 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.735 260.73 204.115 261.11 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.005 260.73 205.385 261.11 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  209.975 260.73 210.355 261.11 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  211.245 260.73 211.625 261.11 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.215 260.73 216.595 261.11 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.485 260.73 217.865 261.11 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  222.455 260.73 222.835 261.11 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  223.725 260.73 224.105 261.11 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  228.695 260.73 229.075 261.11 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  229.965 260.73 230.345 261.11 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  234.935 260.73 235.315 261.11 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  0.0 0.0 1.74 261.11 ;
         LAYER met3 ;
         RECT  0.0 259.37 370.18 261.11 ;
         LAYER met4 ;
         RECT  368.44 0.0 370.18 261.11 ;
         LAYER met3 ;
         RECT  0.0 0.0 370.18 1.74 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  3.48 255.89 366.7 257.63 ;
         LAYER met4 ;
         RECT  3.48 3.48 5.22 257.63 ;
         LAYER met4 ;
         RECT  364.96 3.48 366.7 257.63 ;
         LAYER met3 ;
         RECT  3.48 3.48 366.7 5.22 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 369.56 260.49 ;
   LAYER  met2 ;
      RECT  0.62 0.62 369.56 260.49 ;
   LAYER  met3 ;
      RECT  0.98 108.985 369.56 110.565 ;
      RECT  0.62 110.565 0.98 117.385 ;
      RECT  0.62 118.965 0.98 123.25 ;
      RECT  0.62 124.83 0.98 131.75 ;
      RECT  0.62 133.33 0.98 137.39 ;
      RECT  0.62 138.97 0.98 145.89 ;
      RECT  0.98 71.87 369.2 73.45 ;
      RECT  0.98 73.45 369.2 108.985 ;
      RECT  369.2 73.45 369.56 108.985 ;
      RECT  369.2 64.95 369.56 71.87 ;
      RECT  0.98 110.565 369.2 245.26 ;
      RECT  0.98 245.26 369.2 246.84 ;
      RECT  369.2 110.565 369.56 245.26 ;
      RECT  0.62 17.71 0.98 24.63 ;
      RECT  0.62 26.21 0.98 108.985 ;
      RECT  0.62 147.47 0.98 258.77 ;
      RECT  369.2 246.84 369.56 258.77 ;
      RECT  369.2 2.34 369.56 63.37 ;
      RECT  0.62 2.34 0.98 16.13 ;
      RECT  0.98 246.84 2.88 255.29 ;
      RECT  0.98 255.29 2.88 258.23 ;
      RECT  0.98 258.23 2.88 258.77 ;
      RECT  2.88 246.84 367.3 255.29 ;
      RECT  2.88 258.23 367.3 258.77 ;
      RECT  367.3 246.84 369.2 255.29 ;
      RECT  367.3 255.29 369.2 258.23 ;
      RECT  367.3 258.23 369.2 258.77 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 71.87 ;
      RECT  2.88 2.34 367.3 2.88 ;
      RECT  2.88 5.82 367.3 71.87 ;
      RECT  367.3 2.34 369.2 2.88 ;
      RECT  367.3 2.88 369.2 5.82 ;
      RECT  367.3 5.82 369.2 71.87 ;
   LAYER  met4 ;
      RECT  99.94 0.98 101.52 260.49 ;
      RECT  101.52 0.62 105.78 0.98 ;
      RECT  107.36 0.62 111.62 0.98 ;
      RECT  113.2 0.62 117.46 0.98 ;
      RECT  119.04 0.62 123.3 0.98 ;
      RECT  124.88 0.62 129.14 0.98 ;
      RECT  130.72 0.62 134.98 0.98 ;
      RECT  241.68 0.62 245.94 0.98 ;
      RECT  247.52 0.62 251.78 0.98 ;
      RECT  253.36 0.62 257.62 0.98 ;
      RECT  259.2 0.62 263.46 0.98 ;
      RECT  265.04 0.62 269.3 0.98 ;
      RECT  270.88 0.62 275.14 0.98 ;
      RECT  276.72 0.62 280.98 0.98 ;
      RECT  282.56 0.62 304.185 0.98 ;
      RECT  101.52 0.98 338.94 260.13 ;
      RECT  338.94 0.98 340.52 260.13 ;
      RECT  32.08 0.62 76.58 0.98 ;
      RECT  78.16 0.62 82.42 0.98 ;
      RECT  84.0 0.62 88.26 0.98 ;
      RECT  89.84 0.62 94.1 0.98 ;
      RECT  95.68 0.62 99.94 0.98 ;
      RECT  136.56 0.62 137.085 0.98 ;
      RECT  138.665 0.62 140.82 0.98 ;
      RECT  143.09 0.62 143.325 0.98 ;
      RECT  144.905 0.62 146.66 0.98 ;
      RECT  149.765 0.62 152.5 0.98 ;
      RECT  156.005 0.62 158.34 0.98 ;
      RECT  160.98 0.62 162.045 0.98 ;
      RECT  163.625 0.62 164.18 0.98 ;
      RECT  168.485 0.62 170.02 0.98 ;
      RECT  171.6 0.62 171.935 0.98 ;
      RECT  174.725 0.62 175.86 0.98 ;
      RECT  177.44 0.62 178.175 0.98 ;
      RECT  180.965 0.62 181.7 0.98 ;
      RECT  183.28 0.62 184.36 0.98 ;
      RECT  187.265 0.62 187.54 0.98 ;
      RECT  189.12 0.62 190.655 0.98 ;
      RECT  193.155 0.62 193.38 0.98 ;
      RECT  194.96 0.62 196.895 0.98 ;
      RECT  198.475 0.62 199.22 0.98 ;
      RECT  201.49 0.62 203.135 0.98 ;
      RECT  204.715 0.62 205.06 0.98 ;
      RECT  207.33 0.62 209.095 0.98 ;
      RECT  210.675 0.62 210.9 0.98 ;
      RECT  213.545 0.62 214.935 0.98 ;
      RECT  216.515 0.62 216.74 0.98 ;
      RECT  219.01 0.62 219.915 0.98 ;
      RECT  221.495 0.62 222.58 0.98 ;
      RECT  224.85 0.62 228.42 0.98 ;
      RECT  232.265 0.62 234.26 0.98 ;
      RECT  236.66 0.62 240.1 0.98 ;
      RECT  101.52 260.13 135.765 260.49 ;
      RECT  137.345 260.13 140.735 260.49 ;
      RECT  143.585 260.13 146.975 260.49 ;
      RECT  149.825 260.13 153.215 260.49 ;
      RECT  156.065 260.13 159.455 260.49 ;
      RECT  162.305 260.13 165.695 260.49 ;
      RECT  168.545 260.13 171.935 260.49 ;
      RECT  174.785 260.13 178.175 260.49 ;
      RECT  181.025 260.13 184.415 260.49 ;
      RECT  187.265 260.13 190.655 260.49 ;
      RECT  193.505 260.13 196.895 260.49 ;
      RECT  199.745 260.13 203.135 260.49 ;
      RECT  205.985 260.13 209.375 260.49 ;
      RECT  212.225 260.13 215.615 260.49 ;
      RECT  218.465 260.13 221.855 260.49 ;
      RECT  224.705 260.13 228.095 260.49 ;
      RECT  230.945 260.13 234.335 260.49 ;
      RECT  235.915 260.13 338.94 260.49 ;
      RECT  2.34 0.62 30.5 0.98 ;
      RECT  308.74 0.62 367.84 0.98 ;
      RECT  340.52 260.13 367.84 260.49 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 258.23 ;
      RECT  2.34 258.23 2.88 260.49 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 258.23 5.82 260.49 ;
      RECT  5.82 0.98 99.94 2.88 ;
      RECT  5.82 2.88 99.94 258.23 ;
      RECT  5.82 258.23 99.94 260.49 ;
      RECT  340.52 0.98 364.36 2.88 ;
      RECT  340.52 2.88 364.36 258.23 ;
      RECT  340.52 258.23 364.36 260.13 ;
      RECT  364.36 0.98 367.3 2.88 ;
      RECT  364.36 258.23 367.3 260.13 ;
      RECT  367.3 0.98 367.84 2.88 ;
      RECT  367.3 2.88 367.84 258.23 ;
      RECT  367.3 258.23 367.84 260.13 ;
   END
END    sky130_sram_256byte_1rw1r_32x64_8
END    LIBRARY
