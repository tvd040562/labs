magic
tech sky130A
magscale 1 2
timestamp 1727679568
<< viali >>
rect 19441 31433 19475 31467
rect 22201 31433 22235 31467
rect 25421 31433 25455 31467
rect 16865 31365 16899 31399
rect 23305 31365 23339 31399
rect 17233 31297 17267 31331
rect 19349 31297 19383 31331
rect 21925 31297 21959 31331
rect 23673 31297 23707 31331
rect 25329 31297 25363 31331
rect 21649 30345 21683 30379
rect 17417 30209 17451 30243
rect 17684 30209 17718 30243
rect 19441 30209 19475 30243
rect 20536 30209 20570 30243
rect 22385 30209 22419 30243
rect 22753 30209 22787 30243
rect 20269 30141 20303 30175
rect 18797 30073 18831 30107
rect 21833 30073 21867 30107
rect 18889 30005 18923 30039
rect 22569 30005 22603 30039
rect 9137 29801 9171 29835
rect 10333 29801 10367 29835
rect 15945 29801 15979 29835
rect 18705 29801 18739 29835
rect 20729 29801 20763 29835
rect 23397 29801 23431 29835
rect 9505 29733 9539 29767
rect 10241 29733 10275 29767
rect 17325 29665 17359 29699
rect 17969 29665 18003 29699
rect 22017 29665 22051 29699
rect 24041 29665 24075 29699
rect 3157 29597 3191 29631
rect 3249 29597 3283 29631
rect 9321 29597 9355 29631
rect 9689 29597 9723 29631
rect 10057 29597 10091 29631
rect 10517 29597 10551 29631
rect 10609 29597 10643 29631
rect 18153 29597 18187 29631
rect 18521 29597 18555 29631
rect 20913 29597 20947 29631
rect 21281 29597 21315 29631
rect 21925 29597 21959 29631
rect 25789 29597 25823 29631
rect 17080 29529 17114 29563
rect 18337 29529 18371 29563
rect 18429 29529 18463 29563
rect 21005 29529 21039 29563
rect 21097 29529 21131 29563
rect 22284 29529 22318 29563
rect 25522 29529 25556 29563
rect 2973 29461 3007 29495
rect 3433 29461 3467 29495
rect 10793 29461 10827 29495
rect 17417 29461 17451 29495
rect 21741 29461 21775 29495
rect 23489 29461 23523 29495
rect 24409 29461 24443 29495
rect 3709 29257 3743 29291
rect 9137 29257 9171 29291
rect 9689 29257 9723 29291
rect 10517 29257 10551 29291
rect 12817 29257 12851 29291
rect 15945 29257 15979 29291
rect 16313 29257 16347 29291
rect 22477 29257 22511 29291
rect 24501 29257 24535 29291
rect 16865 29189 16899 29223
rect 16957 29189 16991 29223
rect 22109 29189 22143 29223
rect 24133 29189 24167 29223
rect 24225 29189 24259 29223
rect 1409 29121 1443 29155
rect 2513 29121 2547 29155
rect 2973 29121 3007 29155
rect 3157 29121 3191 29155
rect 3525 29121 3559 29155
rect 3985 29121 4019 29155
rect 4261 29121 4295 29155
rect 4445 29121 4479 29155
rect 4721 29121 4755 29155
rect 5181 29121 5215 29155
rect 5273 29121 5307 29155
rect 7205 29121 7239 29155
rect 7481 29121 7515 29155
rect 7757 29121 7791 29155
rect 8033 29121 8067 29155
rect 8861 29121 8895 29155
rect 8953 29121 8987 29155
rect 9413 29121 9447 29155
rect 9873 29121 9907 29155
rect 9965 29121 9999 29155
rect 10425 29121 10459 29155
rect 10701 29121 10735 29155
rect 10793 29121 10827 29155
rect 11069 29121 11103 29155
rect 11713 29121 11747 29155
rect 12173 29121 12207 29155
rect 12265 29121 12299 29155
rect 12725 29121 12759 29155
rect 13001 29121 13035 29155
rect 16129 29121 16163 29155
rect 16681 29121 16715 29155
rect 17049 29121 17083 29155
rect 17969 29121 18003 29155
rect 18245 29121 18279 29155
rect 20177 29121 20211 29155
rect 21925 29121 21959 29155
rect 22201 29121 22235 29155
rect 22293 29121 22327 29155
rect 23489 29121 23523 29155
rect 23949 29121 23983 29155
rect 24317 29121 24351 29155
rect 24593 29121 24627 29155
rect 25237 29121 25271 29155
rect 2697 28985 2731 29019
rect 7021 28985 7055 29019
rect 7573 28985 7607 29019
rect 7849 28985 7883 29019
rect 11253 28985 11287 29019
rect 12449 28985 12483 29019
rect 17233 28985 17267 29019
rect 18153 28985 18187 29019
rect 1593 28917 1627 28951
rect 2789 28917 2823 28951
rect 3341 28917 3375 28951
rect 3801 28917 3835 28951
rect 4077 28917 4111 28951
rect 4629 28917 4663 28951
rect 4905 28917 4939 28951
rect 4997 28917 5031 28951
rect 5457 28917 5491 28951
rect 7297 28917 7331 28951
rect 8677 28917 8711 28951
rect 9229 28917 9263 28951
rect 10149 28917 10183 28951
rect 10241 28917 10275 28951
rect 10977 28917 11011 28951
rect 11529 28917 11563 28951
rect 11989 28917 12023 28951
rect 12541 28917 12575 28951
rect 18429 28917 18463 28951
rect 20361 28917 20395 28951
rect 23673 28917 23707 28951
rect 2973 28713 3007 28747
rect 3985 28713 4019 28747
rect 6101 28713 6135 28747
rect 12541 28713 12575 28747
rect 13553 28713 13587 28747
rect 16497 28713 16531 28747
rect 19901 28713 19935 28747
rect 23213 28713 23247 28747
rect 23765 28713 23799 28747
rect 2789 28645 2823 28679
rect 5365 28645 5399 28679
rect 8493 28645 8527 28679
rect 9505 28645 9539 28679
rect 11897 28645 11931 28679
rect 13277 28645 13311 28679
rect 14381 28645 14415 28679
rect 3157 28577 3191 28611
rect 4905 28577 4939 28611
rect 5733 28577 5767 28611
rect 5825 28577 5859 28611
rect 5917 28577 5951 28611
rect 19901 28577 19935 28611
rect 20269 28577 20303 28611
rect 1409 28509 1443 28543
rect 1676 28509 1710 28543
rect 3341 28509 3375 28543
rect 3801 28509 3835 28543
rect 4261 28509 4295 28543
rect 4353 28509 4387 28543
rect 5641 28509 5675 28543
rect 6837 28509 6871 28543
rect 6929 28509 6963 28543
rect 7205 28509 7239 28543
rect 7665 28509 7699 28543
rect 8033 28509 8067 28543
rect 8309 28509 8343 28543
rect 8585 28509 8619 28543
rect 8953 28509 8987 28543
rect 9345 28509 9379 28543
rect 9781 28509 9815 28543
rect 10241 28509 10275 28543
rect 10517 28509 10551 28543
rect 10793 28509 10827 28543
rect 10885 28509 10919 28543
rect 11345 28509 11379 28543
rect 11529 28509 11563 28543
rect 11713 28509 11747 28543
rect 11989 28509 12023 28543
rect 12357 28509 12391 28543
rect 12633 28509 12667 28543
rect 12817 28509 12851 28543
rect 12909 28509 12943 28543
rect 13001 28509 13035 28543
rect 13461 28509 13495 28543
rect 13737 28509 13771 28543
rect 14289 28509 14323 28543
rect 14565 28509 14599 28543
rect 16313 28509 16347 28543
rect 17969 28509 18003 28543
rect 18337 28509 18371 28543
rect 20009 28509 20043 28543
rect 20545 28509 20579 28543
rect 23213 28509 23247 28543
rect 23397 28509 23431 28543
rect 23765 28509 23799 28543
rect 23949 28509 23983 28543
rect 2881 28441 2915 28475
rect 5365 28441 5399 28475
rect 9137 28441 9171 28475
rect 9229 28441 9263 28475
rect 10701 28441 10735 28475
rect 11621 28441 11655 28475
rect 12173 28441 12207 28475
rect 12265 28441 12299 28475
rect 15853 28441 15887 28475
rect 16037 28441 16071 28475
rect 17325 28441 17359 28475
rect 17509 28441 17543 28475
rect 18153 28441 18187 28475
rect 19717 28441 19751 28475
rect 3525 28373 3559 28407
rect 4077 28373 4111 28407
rect 4537 28373 4571 28407
rect 4629 28373 4663 28407
rect 4813 28373 4847 28407
rect 6653 28373 6687 28407
rect 7113 28373 7147 28407
rect 7389 28373 7423 28407
rect 7849 28373 7883 28407
rect 8217 28373 8251 28407
rect 8769 28373 8803 28407
rect 9965 28373 9999 28407
rect 10425 28373 10459 28407
rect 11069 28373 11103 28407
rect 13185 28373 13219 28407
rect 14105 28373 14139 28407
rect 16221 28373 16255 28407
rect 17693 28373 17727 28407
rect 17785 28373 17819 28407
rect 18521 28373 18555 28407
rect 20177 28373 20211 28407
rect 23581 28373 23615 28407
rect 24133 28373 24167 28407
rect 2789 28169 2823 28203
rect 5365 28169 5399 28203
rect 6009 28169 6043 28203
rect 8217 28169 8251 28203
rect 8493 28169 8527 28203
rect 11345 28169 11379 28203
rect 12725 28169 12759 28203
rect 15393 28169 15427 28203
rect 3341 28101 3375 28135
rect 3985 28101 4019 28135
rect 4445 28101 4479 28135
rect 4905 28101 4939 28135
rect 8769 28101 8803 28135
rect 8861 28101 8895 28135
rect 11897 28101 11931 28135
rect 13737 28101 13771 28135
rect 23305 28101 23339 28135
rect 25605 28101 25639 28135
rect 1676 28033 1710 28067
rect 3550 28033 3584 28067
rect 5457 28033 5491 28067
rect 5733 28033 5767 28067
rect 6193 28033 6227 28067
rect 6377 28033 6411 28067
rect 6561 28033 6595 28067
rect 6653 28033 6687 28067
rect 6745 28033 6779 28067
rect 7021 28033 7055 28067
rect 7205 28033 7239 28067
rect 7481 28033 7515 28067
rect 7757 28033 7791 28067
rect 8033 28033 8067 28067
rect 8309 28033 8343 28067
rect 8585 28033 8619 28067
rect 8953 28033 8987 28067
rect 9505 28033 9539 28067
rect 9781 28033 9815 28067
rect 10057 28033 10091 28067
rect 10149 28033 10183 28067
rect 10333 28033 10367 28067
rect 10609 28023 10643 28057
rect 10793 28033 10827 28067
rect 10885 28033 10919 28067
rect 11161 28033 11195 28067
rect 11621 28033 11655 28067
rect 11805 28033 11839 28067
rect 11989 28033 12023 28067
rect 12449 28033 12483 28067
rect 12541 28033 12575 28067
rect 13001 28033 13035 28067
rect 14013 28033 14047 28067
rect 14657 28033 14691 28067
rect 14841 28033 14875 28067
rect 15025 28033 15059 28067
rect 15209 28033 15243 28067
rect 17877 28033 17911 28067
rect 18245 28033 18279 28067
rect 19533 28033 19567 28067
rect 19809 28033 19843 28067
rect 20177 28033 20211 28067
rect 22017 28033 22051 28067
rect 22293 28033 22327 28067
rect 22569 28033 22603 28067
rect 23581 28033 23615 28067
rect 24869 28033 24903 28067
rect 25145 28033 25179 28067
rect 1409 27965 1443 27999
rect 3065 27965 3099 27999
rect 3433 27965 3467 27999
rect 4537 27965 4571 27999
rect 5641 27965 5675 27999
rect 7665 27965 7699 27999
rect 13829 27965 13863 27999
rect 16957 27965 16991 27999
rect 17233 27965 17267 27999
rect 18337 27965 18371 27999
rect 19717 27965 19751 27999
rect 20453 27965 20487 27999
rect 22109 27965 22143 27999
rect 23489 27965 23523 27999
rect 24961 27965 24995 27999
rect 3985 27897 4019 27931
rect 4905 27897 4939 27931
rect 5917 27897 5951 27931
rect 9137 27897 9171 27931
rect 9873 27897 9907 27931
rect 18061 27897 18095 27931
rect 21833 27897 21867 27931
rect 22385 27897 22419 27931
rect 23765 27897 23799 27931
rect 3709 27829 3743 27863
rect 4721 27829 4755 27863
rect 6929 27829 6963 27863
rect 7941 27829 7975 27863
rect 9321 27829 9355 27863
rect 9597 27829 9631 27863
rect 11069 27829 11103 27863
rect 12173 27829 12207 27863
rect 12265 27829 12299 27863
rect 12817 27829 12851 27863
rect 13921 27829 13955 27863
rect 14197 27829 14231 27863
rect 14565 27829 14599 27863
rect 18245 27829 18279 27863
rect 18613 27829 18647 27863
rect 19809 27829 19843 27863
rect 19993 27829 20027 27863
rect 22293 27829 22327 27863
rect 23397 27829 23431 27863
rect 25145 27829 25179 27863
rect 25329 27829 25363 27863
rect 25513 27829 25547 27863
rect 1593 27625 1627 27659
rect 7297 27625 7331 27659
rect 7389 27625 7423 27659
rect 9689 27625 9723 27659
rect 14565 27625 14599 27659
rect 15209 27625 15243 27659
rect 16037 27625 16071 27659
rect 16773 27625 16807 27659
rect 18889 27625 18923 27659
rect 20453 27625 20487 27659
rect 22477 27625 22511 27659
rect 23673 27625 23707 27659
rect 24225 27625 24259 27659
rect 25605 27625 25639 27659
rect 2237 27557 2271 27591
rect 3525 27557 3559 27591
rect 3985 27557 4019 27591
rect 4905 27557 4939 27591
rect 5641 27557 5675 27591
rect 6377 27557 6411 27591
rect 7665 27557 7699 27591
rect 8217 27557 8251 27591
rect 11253 27557 11287 27591
rect 12357 27557 12391 27591
rect 13001 27557 13035 27591
rect 15577 27557 15611 27591
rect 16313 27557 16347 27591
rect 22753 27557 22787 27591
rect 23765 27557 23799 27591
rect 2513 27489 2547 27523
rect 2605 27489 2639 27523
rect 2881 27489 2915 27523
rect 3249 27489 3283 27523
rect 3366 27489 3400 27523
rect 4445 27489 4479 27523
rect 5365 27489 5399 27523
rect 16037 27489 16071 27523
rect 16865 27489 16899 27523
rect 18797 27489 18831 27523
rect 19257 27489 19291 27523
rect 19533 27489 19567 27523
rect 22385 27489 22419 27523
rect 25789 27489 25823 27523
rect 1409 27421 1443 27455
rect 2421 27421 2455 27455
rect 2697 27421 2731 27455
rect 4537 27421 4571 27455
rect 6009 27421 6043 27455
rect 6101 27421 6135 27455
rect 6561 27421 6595 27455
rect 6837 27421 6871 27455
rect 7113 27421 7147 27455
rect 7573 27421 7607 27455
rect 7849 27421 7883 27455
rect 8125 27421 8159 27455
rect 8401 27421 8435 27455
rect 8585 27421 8619 27455
rect 9137 27421 9171 27455
rect 9413 27421 9447 27455
rect 9505 27421 9539 27455
rect 9781 27421 9815 27455
rect 10149 27421 10183 27455
rect 10609 27421 10643 27455
rect 10977 27421 11011 27455
rect 11437 27421 11471 27455
rect 11529 27421 11563 27455
rect 11805 27421 11839 27455
rect 11989 27421 12023 27455
rect 12173 27421 12207 27455
rect 12449 27421 12483 27455
rect 12633 27421 12667 27455
rect 12817 27421 12851 27455
rect 13277 27421 13311 27455
rect 14289 27421 14323 27455
rect 14381 27421 14415 27455
rect 14565 27421 14599 27455
rect 15025 27421 15059 27455
rect 15301 27421 15335 27455
rect 15393 27421 15427 27455
rect 15945 27421 15979 27455
rect 16497 27421 16531 27455
rect 17049 27421 17083 27455
rect 17325 27421 17359 27455
rect 17785 27421 17819 27455
rect 18705 27421 18739 27455
rect 20361 27421 20395 27455
rect 20453 27421 20487 27455
rect 22569 27421 22603 27455
rect 23949 27421 23983 27455
rect 24041 27421 24075 27455
rect 25605 27421 25639 27455
rect 25881 27421 25915 27455
rect 3157 27353 3191 27387
rect 3985 27353 4019 27387
rect 4905 27353 4939 27387
rect 5457 27353 5491 27387
rect 9321 27353 9355 27387
rect 9965 27353 9999 27387
rect 10057 27353 10091 27387
rect 10793 27353 10827 27387
rect 10885 27353 10919 27387
rect 12081 27353 12115 27387
rect 12725 27353 12759 27387
rect 15117 27353 15151 27387
rect 16773 27353 16807 27387
rect 20177 27353 20211 27387
rect 22293 27353 22327 27387
rect 24225 27353 24259 27387
rect 26617 27353 26651 27387
rect 26801 27353 26835 27387
rect 4721 27285 4755 27319
rect 5825 27285 5859 27319
rect 6285 27285 6319 27319
rect 7021 27285 7055 27319
rect 7941 27285 7975 27319
rect 8769 27285 8803 27319
rect 10333 27285 10367 27319
rect 11161 27285 11195 27319
rect 11713 27285 11747 27319
rect 13093 27285 13127 27319
rect 14105 27285 14139 27319
rect 14749 27285 14783 27319
rect 14841 27285 14875 27319
rect 16681 27285 16715 27319
rect 17233 27285 17267 27319
rect 17509 27285 17543 27319
rect 17601 27285 17635 27319
rect 19073 27285 19107 27319
rect 20637 27285 20671 27319
rect 26065 27285 26099 27319
rect 26985 27285 27019 27319
rect 3985 27081 4019 27115
rect 4629 27081 4663 27115
rect 4997 27081 5031 27115
rect 6561 27081 6595 27115
rect 7205 27081 7239 27115
rect 10609 27081 10643 27115
rect 14381 27081 14415 27115
rect 14933 27081 14967 27115
rect 28273 27081 28307 27115
rect 6837 27013 6871 27047
rect 7573 27013 7607 27047
rect 8953 27013 8987 27047
rect 10149 27013 10183 27047
rect 14473 27013 14507 27047
rect 17325 27013 17359 27047
rect 18521 27013 18555 27047
rect 23489 27013 23523 27047
rect 31217 27013 31251 27047
rect 2053 26945 2087 26979
rect 2329 26945 2363 26979
rect 2881 26945 2915 26979
rect 2973 26945 3007 26979
rect 3249 26945 3283 26979
rect 3525 26945 3559 26979
rect 3801 26945 3835 26979
rect 4077 26945 4111 26979
rect 4445 26945 4479 26979
rect 4721 26945 4755 26979
rect 5206 26945 5240 26979
rect 5549 26945 5583 26979
rect 5825 26945 5859 26979
rect 6377 26945 6411 26979
rect 6653 26945 6687 26979
rect 6929 26945 6963 26979
rect 7021 26945 7055 26979
rect 7297 26945 7331 26979
rect 7481 26945 7515 26979
rect 7665 26945 7699 26979
rect 7941 26945 7975 26979
rect 8125 26945 8159 26979
rect 8217 26945 8251 26979
rect 8309 26945 8343 26979
rect 8861 26945 8895 26979
rect 9045 26945 9079 26979
rect 9229 26945 9263 26979
rect 9321 26945 9355 26979
rect 9505 26945 9539 26979
rect 9597 26945 9631 26979
rect 9689 26945 9723 26979
rect 9965 26945 9999 26979
rect 10241 26945 10275 26979
rect 10333 26945 10367 26979
rect 10793 26945 10827 26979
rect 11069 26945 11103 26979
rect 13093 26945 13127 26979
rect 13284 26945 13318 26979
rect 13461 26945 13495 26979
rect 13553 26945 13587 26979
rect 14013 26945 14047 26979
rect 14197 26945 14231 26979
rect 14749 26945 14783 26979
rect 16405 26945 16439 26979
rect 16865 26945 16899 26979
rect 17601 26945 17635 26979
rect 18337 26945 18371 26979
rect 18797 26945 18831 26979
rect 19625 26945 19659 26979
rect 19717 26945 19751 26979
rect 22477 26945 22511 26979
rect 22661 26945 22695 26979
rect 23305 26945 23339 26979
rect 23581 26945 23615 26979
rect 24961 26945 24995 26979
rect 25145 26945 25179 26979
rect 25237 26945 25271 26979
rect 25605 26945 25639 26979
rect 25881 26945 25915 26979
rect 26985 26945 27019 26979
rect 27261 26945 27295 26979
rect 28641 26945 28675 26979
rect 30941 26945 30975 26979
rect 31125 26945 31159 26979
rect 31309 26945 31343 26979
rect 32505 26945 32539 26979
rect 2605 26877 2639 26911
rect 2789 26877 2823 26911
rect 3065 26877 3099 26911
rect 5089 26877 5123 26911
rect 13829 26877 13863 26911
rect 14565 26877 14599 26911
rect 17417 26877 17451 26911
rect 18705 26877 18739 26911
rect 19533 26877 19567 26911
rect 25697 26877 25731 26911
rect 2237 26809 2271 26843
rect 2513 26809 2547 26843
rect 3709 26809 3743 26843
rect 17049 26809 17083 26843
rect 18981 26809 19015 26843
rect 19257 26809 19291 26843
rect 25421 26809 25455 26843
rect 3433 26741 3467 26775
rect 4261 26741 4295 26775
rect 5365 26741 5399 26775
rect 5733 26741 5767 26775
rect 6009 26741 6043 26775
rect 7849 26741 7883 26775
rect 8493 26741 8527 26775
rect 8677 26741 8711 26775
rect 9873 26741 9907 26775
rect 10517 26741 10551 26775
rect 10885 26741 10919 26775
rect 13001 26741 13035 26775
rect 13553 26741 13587 26775
rect 13737 26741 13771 26775
rect 14473 26741 14507 26775
rect 16221 26741 16255 26775
rect 17417 26741 17451 26775
rect 17785 26741 17819 26775
rect 19533 26741 19567 26775
rect 19901 26741 19935 26775
rect 22845 26741 22879 26775
rect 23121 26741 23155 26775
rect 23765 26741 23799 26775
rect 25237 26741 25271 26775
rect 25697 26741 25731 26775
rect 26065 26741 26099 26775
rect 27169 26741 27203 26775
rect 27445 26741 27479 26775
rect 28457 26741 28491 26775
rect 31493 26741 31527 26775
rect 32321 26741 32355 26775
rect 2789 26537 2823 26571
rect 4905 26537 4939 26571
rect 5457 26537 5491 26571
rect 7849 26537 7883 26571
rect 8125 26537 8159 26571
rect 13645 26537 13679 26571
rect 15025 26537 15059 26571
rect 15209 26537 15243 26571
rect 16037 26537 16071 26571
rect 18153 26537 18187 26571
rect 23121 26537 23155 26571
rect 26617 26537 26651 26571
rect 26985 26537 27019 26571
rect 27629 26537 27663 26571
rect 27905 26537 27939 26571
rect 28365 26537 28399 26571
rect 31861 26537 31895 26571
rect 3893 26469 3927 26503
rect 5181 26469 5215 26503
rect 6101 26469 6135 26503
rect 6653 26469 6687 26503
rect 7573 26469 7607 26503
rect 11161 26469 11195 26503
rect 13921 26469 13955 26503
rect 16497 26469 16531 26503
rect 21649 26469 21683 26503
rect 23581 26469 23615 26503
rect 28733 26469 28767 26503
rect 3341 26401 3375 26435
rect 4353 26401 4387 26435
rect 14841 26401 14875 26435
rect 18061 26401 18095 26435
rect 18429 26401 18463 26435
rect 23029 26401 23063 26435
rect 23213 26401 23247 26435
rect 26893 26401 26927 26435
rect 28365 26401 28399 26435
rect 1409 26333 1443 26367
rect 2973 26333 3007 26367
rect 4445 26333 4479 26367
rect 4721 26333 4755 26367
rect 4997 26333 5031 26367
rect 5273 26333 5307 26367
rect 5549 26333 5583 26367
rect 5733 26333 5767 26367
rect 5825 26333 5859 26367
rect 5917 26333 5951 26367
rect 6377 26333 6411 26367
rect 6837 26333 6871 26367
rect 7021 26333 7055 26367
rect 7389 26333 7423 26367
rect 7665 26333 7699 26367
rect 7941 26333 7975 26367
rect 8953 26333 8987 26367
rect 9229 26333 9263 26367
rect 9873 26333 9907 26367
rect 10333 26333 10367 26367
rect 11345 26333 11379 26367
rect 11713 26333 11747 26367
rect 11805 26333 11839 26367
rect 12173 26333 12207 26367
rect 13461 26333 13495 26367
rect 13737 26333 13771 26367
rect 15025 26333 15059 26367
rect 16221 26333 16255 26367
rect 16313 26333 16347 26367
rect 18153 26333 18187 26367
rect 18613 26333 18647 26367
rect 18797 26333 18831 26367
rect 21373 26333 21407 26367
rect 21833 26333 21867 26367
rect 23121 26333 23155 26367
rect 23397 26333 23431 26367
rect 26801 26333 26835 26367
rect 27537 26333 27571 26367
rect 27629 26333 27663 26367
rect 27721 26333 27755 26367
rect 28273 26333 28307 26367
rect 28549 26333 28583 26367
rect 31585 26333 31619 26367
rect 32505 26333 32539 26367
rect 1676 26265 1710 26299
rect 3458 26265 3492 26299
rect 3893 26265 3927 26299
rect 7205 26265 7239 26299
rect 7297 26265 7331 26299
rect 11437 26265 11471 26299
rect 11529 26265 11563 26299
rect 11989 26265 12023 26299
rect 12081 26265 12115 26299
rect 14749 26265 14783 26299
rect 16037 26265 16071 26299
rect 17877 26265 17911 26299
rect 21189 26265 21223 26299
rect 21557 26265 21591 26299
rect 27077 26265 27111 26299
rect 3249 26197 3283 26231
rect 3617 26197 3651 26231
rect 4629 26197 4663 26231
rect 6561 26197 6595 26231
rect 9137 26197 9171 26231
rect 9413 26197 9447 26231
rect 10057 26197 10091 26231
rect 10149 26197 10183 26231
rect 12357 26197 12391 26231
rect 18337 26197 18371 26231
rect 27261 26197 27295 26231
rect 30941 26197 30975 26231
rect 1593 25993 1627 26027
rect 3065 25993 3099 26027
rect 3525 25993 3559 26027
rect 4721 25993 4755 26027
rect 5917 25993 5951 26027
rect 7021 25993 7055 26027
rect 8677 25993 8711 26027
rect 9413 25993 9447 26027
rect 9873 25993 9907 26027
rect 20177 25993 20211 26027
rect 30205 25993 30239 26027
rect 3249 25925 3283 25959
rect 3801 25925 3835 25959
rect 5273 25925 5307 25959
rect 8953 25925 8987 25959
rect 10609 25925 10643 25959
rect 29837 25925 29871 25959
rect 29929 25925 29963 25959
rect 30542 25925 30576 25959
rect 1409 25857 1443 25891
rect 2881 25857 2915 25891
rect 3157 25857 3191 25891
rect 3709 25857 3743 25891
rect 4077 25857 4111 25891
rect 4537 25857 4571 25891
rect 4813 25857 4847 25891
rect 5089 25857 5123 25891
rect 5365 25857 5399 25891
rect 5457 25857 5491 25891
rect 5733 25857 5767 25891
rect 6009 25857 6043 25891
rect 6377 25857 6411 25891
rect 6561 25857 6595 25891
rect 6653 25857 6687 25891
rect 6745 25857 6779 25891
rect 7205 25857 7239 25891
rect 7297 25857 7331 25891
rect 8217 25857 8251 25891
rect 8493 25857 8527 25891
rect 8769 25857 8803 25891
rect 9045 25857 9079 25891
rect 9137 25857 9171 25891
rect 9597 25857 9631 25891
rect 9689 25857 9723 25891
rect 10425 25857 10459 25891
rect 10701 25857 10735 25891
rect 10793 25857 10827 25891
rect 13185 25857 13219 25891
rect 13461 25857 13495 25891
rect 16773 25857 16807 25891
rect 16957 25857 16991 25891
rect 18153 25857 18187 25891
rect 18337 25857 18371 25891
rect 19441 25857 19475 25891
rect 19717 25857 19751 25891
rect 19901 25857 19935 25891
rect 19993 25857 20027 25891
rect 20269 25857 20303 25891
rect 20453 25857 20487 25891
rect 21005 25857 21039 25891
rect 21281 25857 21315 25891
rect 21833 25857 21867 25891
rect 22017 25857 22051 25891
rect 23397 25857 23431 25891
rect 23581 25857 23615 25891
rect 23673 25857 23707 25891
rect 24041 25857 24075 25891
rect 29653 25857 29687 25891
rect 30021 25857 30055 25891
rect 32229 25857 32263 25891
rect 3893 25789 3927 25823
rect 30297 25789 30331 25823
rect 3433 25721 3467 25755
rect 6193 25721 6227 25755
rect 6929 25721 6963 25755
rect 9321 25721 9355 25755
rect 19625 25721 19659 25755
rect 20637 25721 20671 25755
rect 22201 25721 22235 25755
rect 23949 25721 23983 25755
rect 31677 25721 31711 25755
rect 3801 25653 3835 25687
rect 4261 25653 4295 25687
rect 4997 25653 5031 25687
rect 5641 25653 5675 25687
rect 7481 25653 7515 25687
rect 8401 25653 8435 25687
rect 10977 25653 11011 25687
rect 13001 25653 13035 25687
rect 13277 25653 13311 25687
rect 19349 25653 19383 25687
rect 19993 25653 20027 25687
rect 20269 25653 20303 25687
rect 21189 25653 21223 25687
rect 21465 25653 21499 25687
rect 21833 25653 21867 25687
rect 23213 25653 23247 25687
rect 23673 25653 23707 25687
rect 24225 25653 24259 25687
rect 32413 25653 32447 25687
rect 2789 25449 2823 25483
rect 6469 25449 6503 25483
rect 6745 25449 6779 25483
rect 10333 25449 10367 25483
rect 12817 25449 12851 25483
rect 13645 25449 13679 25483
rect 16773 25449 16807 25483
rect 17049 25449 17083 25483
rect 17417 25449 17451 25483
rect 19625 25449 19659 25483
rect 20545 25449 20579 25483
rect 21373 25449 21407 25483
rect 22753 25449 22787 25483
rect 23673 25449 23707 25483
rect 24225 25449 24259 25483
rect 25053 25449 25087 25483
rect 25513 25449 25547 25483
rect 25973 25449 26007 25483
rect 26341 25449 26375 25483
rect 29561 25449 29595 25483
rect 29929 25449 29963 25483
rect 32505 25449 32539 25483
rect 4077 25381 4111 25415
rect 5457 25381 5491 25415
rect 9597 25381 9631 25415
rect 12633 25381 12667 25415
rect 13277 25381 13311 25415
rect 16957 25381 16991 25415
rect 19257 25381 19291 25415
rect 20729 25381 20763 25415
rect 21005 25381 21039 25415
rect 21649 25381 21683 25415
rect 13461 25313 13495 25347
rect 20361 25313 20395 25347
rect 25145 25313 25179 25347
rect 25789 25313 25823 25347
rect 26525 25313 26559 25347
rect 31125 25313 31159 25347
rect 1409 25245 1443 25279
rect 3065 25245 3099 25279
rect 3157 25245 3191 25279
rect 3617 25245 3651 25279
rect 3893 25245 3927 25279
rect 4169 25245 4203 25279
rect 4445 25245 4479 25279
rect 5273 25245 5307 25279
rect 5733 25245 5767 25279
rect 5825 25245 5859 25279
rect 6101 25245 6135 25279
rect 6193 25245 6227 25279
rect 6653 25245 6687 25279
rect 6929 25245 6963 25279
rect 8953 25245 8987 25279
rect 9137 25245 9171 25279
rect 9413 25245 9447 25279
rect 9689 25245 9723 25279
rect 9873 25245 9907 25279
rect 10057 25245 10091 25279
rect 10517 25245 10551 25279
rect 10793 25245 10827 25279
rect 10977 25245 11011 25279
rect 11069 25245 11103 25279
rect 11437 25245 11471 25279
rect 11621 25245 11655 25279
rect 11713 25245 11747 25279
rect 11805 25245 11839 25279
rect 12081 25245 12115 25279
rect 12357 25245 12391 25279
rect 12449 25245 12483 25279
rect 13001 25245 13035 25279
rect 13093 25245 13127 25279
rect 13645 25245 13679 25279
rect 14473 25245 14507 25279
rect 15945 25245 15979 25279
rect 16589 25245 16623 25279
rect 16681 25245 16715 25279
rect 17233 25245 17267 25279
rect 17417 25245 17451 25279
rect 17693 25245 17727 25279
rect 17785 25245 17819 25279
rect 18061 25245 18095 25279
rect 19441 25245 19475 25279
rect 19625 25245 19659 25279
rect 20269 25245 20303 25279
rect 20545 25245 20579 25279
rect 20821 25245 20855 25279
rect 21281 25245 21315 25279
rect 21373 25245 21407 25279
rect 21925 25245 21959 25279
rect 22937 25245 22971 25279
rect 23213 25245 23247 25279
rect 23949 25245 23983 25279
rect 24041 25245 24075 25279
rect 25329 25245 25363 25279
rect 25973 25245 26007 25279
rect 26617 25245 26651 25279
rect 29561 25245 29595 25279
rect 29653 25245 29687 25279
rect 31033 25245 31067 25279
rect 31392 25245 31426 25279
rect 1676 25177 1710 25211
rect 6009 25177 6043 25211
rect 9965 25177 9999 25211
rect 12265 25177 12299 25211
rect 12817 25177 12851 25211
rect 13369 25177 13403 25211
rect 16129 25177 16163 25211
rect 16313 25177 16347 25211
rect 24225 25177 24259 25211
rect 25053 25177 25087 25211
rect 25697 25177 25731 25211
rect 26341 25177 26375 25211
rect 2881 25109 2915 25143
rect 3341 25109 3375 25143
rect 3433 25109 3467 25143
rect 4353 25109 4387 25143
rect 4629 25109 4663 25143
rect 5549 25109 5583 25143
rect 6377 25109 6411 25143
rect 10241 25109 10275 25143
rect 11253 25109 11287 25143
rect 11989 25109 12023 25143
rect 13829 25109 13863 25143
rect 14289 25109 14323 25143
rect 16405 25109 16439 25143
rect 17509 25109 17543 25143
rect 17969 25109 18003 25143
rect 18245 25109 18279 25143
rect 22109 25109 22143 25143
rect 23121 25109 23155 25143
rect 23397 25109 23431 25143
rect 23765 25109 23799 25143
rect 26157 25109 26191 25143
rect 26801 25109 26835 25143
rect 30849 25109 30883 25143
rect 2053 24905 2087 24939
rect 3525 24905 3559 24939
rect 3985 24905 4019 24939
rect 16681 24905 16715 24939
rect 21373 24905 21407 24939
rect 22753 24905 22787 24939
rect 23765 24905 23799 24939
rect 27997 24905 28031 24939
rect 2789 24837 2823 24871
rect 3341 24837 3375 24871
rect 5549 24837 5583 24871
rect 7205 24837 7239 24871
rect 17969 24837 18003 24871
rect 22017 24837 22051 24871
rect 1869 24769 1903 24803
rect 2145 24769 2179 24803
rect 2421 24769 2455 24803
rect 3801 24769 3835 24803
rect 4077 24769 4111 24803
rect 5181 24769 5215 24803
rect 5365 24769 5399 24803
rect 5641 24769 5675 24803
rect 5733 24769 5767 24803
rect 6193 24769 6227 24803
rect 7021 24769 7055 24803
rect 7297 24769 7331 24803
rect 7389 24769 7423 24803
rect 8309 24769 8343 24803
rect 8493 24769 8527 24803
rect 8769 24769 8803 24803
rect 9229 24793 9263 24827
rect 9321 24769 9355 24803
rect 9597 24769 9631 24803
rect 11529 24769 11563 24803
rect 11713 24769 11747 24803
rect 11805 24769 11839 24803
rect 11897 24769 11931 24803
rect 12817 24769 12851 24803
rect 13277 24769 13311 24803
rect 13461 24769 13495 24803
rect 14105 24769 14139 24803
rect 14381 24769 14415 24803
rect 14841 24769 14875 24803
rect 15025 24769 15059 24803
rect 16865 24769 16899 24803
rect 16957 24769 16991 24803
rect 17141 24769 17175 24803
rect 17601 24769 17635 24803
rect 17785 24769 17819 24803
rect 18153 24769 18187 24803
rect 18337 24769 18371 24803
rect 18429 24769 18463 24803
rect 18981 24769 19015 24803
rect 19165 24769 19199 24803
rect 19257 24769 19291 24803
rect 19901 24769 19935 24803
rect 20177 24769 20211 24803
rect 20453 24769 20487 24803
rect 20729 24769 20763 24803
rect 21189 24769 21223 24803
rect 21465 24793 21499 24827
rect 22201 24769 22235 24803
rect 22477 24769 22511 24803
rect 22569 24769 22603 24803
rect 23305 24769 23339 24803
rect 23397 24769 23431 24803
rect 23489 24769 23523 24803
rect 23857 24769 23891 24803
rect 24041 24769 24075 24803
rect 27537 24769 27571 24803
rect 27813 24769 27847 24803
rect 28181 24769 28215 24803
rect 28457 24769 28491 24803
rect 30205 24769 30239 24803
rect 31861 24769 31895 24803
rect 32229 24769 32263 24803
rect 3249 24701 3283 24735
rect 4353 24701 4387 24735
rect 14289 24701 14323 24735
rect 20269 24701 20303 24735
rect 20821 24701 20855 24735
rect 23213 24701 23247 24735
rect 24225 24701 24259 24735
rect 28365 24701 28399 24735
rect 30481 24701 30515 24735
rect 2329 24633 2363 24667
rect 2789 24633 2823 24667
rect 4997 24633 5031 24667
rect 5917 24633 5951 24667
rect 6009 24633 6043 24667
rect 9045 24633 9079 24667
rect 13093 24633 13127 24667
rect 13645 24633 13679 24667
rect 18613 24633 18647 24667
rect 21097 24633 21131 24667
rect 21833 24633 21867 24667
rect 22293 24633 22327 24667
rect 22937 24633 22971 24667
rect 27721 24633 27755 24667
rect 28641 24633 28675 24667
rect 2605 24565 2639 24599
rect 7573 24565 7607 24599
rect 8953 24565 8987 24599
rect 9505 24565 9539 24599
rect 9781 24565 9815 24599
rect 12081 24565 12115 24599
rect 13001 24565 13035 24599
rect 14381 24565 14415 24599
rect 14565 24565 14599 24599
rect 14657 24565 14691 24599
rect 17141 24565 17175 24599
rect 18245 24565 18279 24599
rect 19257 24565 19291 24599
rect 19441 24565 19475 24599
rect 20085 24565 20119 24599
rect 20177 24565 20211 24599
rect 20637 24565 20671 24599
rect 20729 24565 20763 24599
rect 21649 24565 21683 24599
rect 23305 24565 23339 24599
rect 23397 24565 23431 24599
rect 28181 24565 28215 24599
rect 31309 24565 31343 24599
rect 32413 24565 32447 24599
rect 1593 24361 1627 24395
rect 2145 24361 2179 24395
rect 3617 24361 3651 24395
rect 5365 24361 5399 24395
rect 6377 24361 6411 24395
rect 8769 24361 8803 24395
rect 11069 24361 11103 24395
rect 11345 24361 11379 24395
rect 20729 24361 20763 24395
rect 21097 24361 21131 24395
rect 23857 24361 23891 24395
rect 25329 24361 25363 24395
rect 25697 24361 25731 24395
rect 28089 24361 28123 24395
rect 28181 24361 28215 24395
rect 2881 24293 2915 24327
rect 3893 24293 3927 24327
rect 4629 24293 4663 24327
rect 9505 24293 9539 24327
rect 10793 24293 10827 24327
rect 29837 24293 29871 24327
rect 31493 24293 31527 24327
rect 2329 24225 2363 24259
rect 2421 24225 2455 24259
rect 3433 24225 3467 24259
rect 4353 24225 4387 24259
rect 21005 24225 21039 24259
rect 27997 24225 28031 24259
rect 28273 24225 28307 24259
rect 32137 24225 32171 24259
rect 1409 24157 1443 24191
rect 1869 24157 1903 24191
rect 2513 24157 2547 24191
rect 2605 24157 2639 24191
rect 4721 24157 4755 24191
rect 4997 24157 5031 24191
rect 5457 24157 5491 24191
rect 5733 24157 5767 24191
rect 6009 24157 6043 24191
rect 6101 24157 6135 24191
rect 6561 24157 6595 24191
rect 6929 24157 6963 24191
rect 7113 24157 7147 24191
rect 7205 24157 7239 24191
rect 7297 24157 7331 24191
rect 8585 24157 8619 24191
rect 8953 24157 8987 24191
rect 9229 24157 9263 24191
rect 9321 24157 9355 24191
rect 9597 24157 9631 24191
rect 9873 24157 9907 24191
rect 9965 24157 9999 24191
rect 10241 24157 10275 24191
rect 10425 24157 10459 24191
rect 10517 24157 10551 24191
rect 10609 24157 10643 24191
rect 10885 24157 10919 24191
rect 11161 24157 11195 24191
rect 21097 24157 21131 24191
rect 21465 24157 21499 24191
rect 21741 24157 21775 24191
rect 22845 24157 22879 24191
rect 25329 24157 25363 24191
rect 25421 24157 25455 24191
rect 27813 24157 27847 24191
rect 28181 24157 28215 24191
rect 28825 24157 28859 24191
rect 29009 24157 29043 24191
rect 29193 24157 29227 24191
rect 30021 24157 30055 24191
rect 30113 24157 30147 24191
rect 2881 24089 2915 24123
rect 3893 24089 3927 24123
rect 5089 24089 5123 24123
rect 5206 24089 5240 24123
rect 5917 24089 5951 24123
rect 9137 24089 9171 24123
rect 9781 24089 9815 24123
rect 11989 24089 12023 24123
rect 12173 24089 12207 24123
rect 21649 24089 21683 24123
rect 23581 24089 23615 24123
rect 23765 24089 23799 24123
rect 28089 24089 28123 24123
rect 29101 24089 29135 24123
rect 30380 24089 30414 24123
rect 2053 24021 2087 24055
rect 3341 24021 3375 24055
rect 4445 24021 4479 24055
rect 5641 24021 5675 24055
rect 6285 24021 6319 24055
rect 7481 24021 7515 24055
rect 10149 24021 10183 24055
rect 11805 24021 11839 24055
rect 21281 24021 21315 24055
rect 21925 24021 21959 24055
rect 23029 24021 23063 24055
rect 27629 24021 27663 24055
rect 28549 24021 28583 24055
rect 29377 24021 29411 24055
rect 31585 24021 31619 24055
rect 2973 23817 3007 23851
rect 3065 23817 3099 23851
rect 3893 23817 3927 23851
rect 4169 23817 4203 23851
rect 6009 23817 6043 23851
rect 10977 23817 11011 23851
rect 12081 23817 12115 23851
rect 12357 23817 12391 23851
rect 13001 23817 13035 23851
rect 24593 23817 24627 23851
rect 30481 23817 30515 23851
rect 31953 23817 31987 23851
rect 3433 23749 3467 23783
rect 10609 23749 10643 23783
rect 11805 23749 11839 23783
rect 15209 23749 15243 23783
rect 17969 23749 18003 23783
rect 24317 23749 24351 23783
rect 30818 23749 30852 23783
rect 2697 23681 2731 23715
rect 2789 23681 2823 23715
rect 3249 23681 3283 23715
rect 4445 23681 4479 23715
rect 4537 23681 4571 23715
rect 5089 23681 5123 23715
rect 5181 23681 5215 23715
rect 5641 23681 5675 23715
rect 5917 23681 5951 23715
rect 6193 23681 6227 23715
rect 6561 23681 6595 23715
rect 8769 23681 8803 23715
rect 8953 23681 8987 23715
rect 9045 23681 9079 23715
rect 9137 23681 9171 23715
rect 10425 23681 10459 23715
rect 10701 23681 10735 23715
rect 10793 23681 10827 23715
rect 11529 23681 11563 23715
rect 11713 23681 11747 23715
rect 11897 23681 11931 23715
rect 12173 23681 12207 23715
rect 12541 23681 12575 23715
rect 12725 23681 12759 23715
rect 13185 23681 13219 23715
rect 13829 23681 13863 23715
rect 14013 23681 14047 23715
rect 14289 23681 14323 23715
rect 15025 23681 15059 23715
rect 15669 23681 15703 23715
rect 16681 23681 16715 23715
rect 16865 23681 16899 23715
rect 18245 23681 18279 23715
rect 19717 23681 19751 23715
rect 22017 23681 22051 23715
rect 22937 23681 22971 23715
rect 24041 23681 24075 23715
rect 24409 23681 24443 23715
rect 26065 23681 26099 23715
rect 29929 23681 29963 23715
rect 30113 23681 30147 23715
rect 30205 23681 30239 23715
rect 30297 23681 30331 23715
rect 30573 23681 30607 23715
rect 32229 23681 32263 23715
rect 3985 23613 4019 23647
rect 4353 23613 4387 23647
rect 4629 23613 4663 23647
rect 17049 23613 17083 23647
rect 18153 23613 18187 23647
rect 24133 23613 24167 23647
rect 26157 23613 26191 23647
rect 2513 23545 2547 23579
rect 3433 23545 3467 23579
rect 6377 23545 6411 23579
rect 13645 23545 13679 23579
rect 15485 23545 15519 23579
rect 23121 23545 23155 23579
rect 4813 23477 4847 23511
rect 4905 23477 4939 23511
rect 5365 23477 5399 23511
rect 5457 23477 5491 23511
rect 5733 23477 5767 23511
rect 9321 23477 9355 23511
rect 12909 23477 12943 23511
rect 14105 23477 14139 23511
rect 15393 23477 15427 23511
rect 18245 23477 18279 23511
rect 18429 23477 18463 23511
rect 19901 23477 19935 23511
rect 22201 23477 22235 23511
rect 23857 23477 23891 23511
rect 24041 23477 24075 23511
rect 26065 23477 26099 23511
rect 26433 23477 26467 23511
rect 32413 23477 32447 23511
rect 2145 23273 2179 23307
rect 4353 23273 4387 23307
rect 6009 23273 6043 23307
rect 7113 23273 7147 23307
rect 14105 23273 14139 23307
rect 16221 23273 16255 23307
rect 16405 23273 16439 23307
rect 17785 23273 17819 23307
rect 18705 23273 18739 23307
rect 20085 23273 20119 23307
rect 21741 23273 21775 23307
rect 24685 23273 24719 23307
rect 25789 23273 25823 23307
rect 25973 23273 26007 23307
rect 26433 23273 26467 23307
rect 26893 23273 26927 23307
rect 28641 23273 28675 23307
rect 2605 23205 2639 23239
rect 2881 23205 2915 23239
rect 10977 23205 11011 23239
rect 14565 23205 14599 23239
rect 19901 23205 19935 23239
rect 24869 23205 24903 23239
rect 4077 23137 4111 23171
rect 17969 23137 18003 23171
rect 18521 23137 18555 23171
rect 24593 23137 24627 23171
rect 26525 23137 26559 23171
rect 28825 23137 28859 23171
rect 31125 23137 31159 23171
rect 2329 23069 2363 23103
rect 2421 23069 2455 23103
rect 2697 23069 2731 23103
rect 2973 23069 3007 23103
rect 3249 23069 3283 23103
rect 3893 23069 3927 23103
rect 3985 23069 4019 23103
rect 4169 23069 4203 23103
rect 4629 23069 4663 23103
rect 4905 23069 4939 23103
rect 5089 23069 5123 23103
rect 5365 23069 5399 23103
rect 5457 23069 5491 23103
rect 5825 23069 5859 23103
rect 6285 23069 6319 23103
rect 6561 23069 6595 23103
rect 6745 23069 6779 23103
rect 6837 23069 6871 23103
rect 6929 23069 6963 23103
rect 7205 23069 7239 23103
rect 7481 23069 7515 23103
rect 7573 23069 7607 23103
rect 7849 23069 7883 23103
rect 8125 23069 8159 23103
rect 8217 23069 8251 23103
rect 10793 23069 10827 23103
rect 11069 23069 11103 23103
rect 11345 23069 11379 23103
rect 12357 23069 12391 23103
rect 12633 23069 12667 23103
rect 14289 23069 14323 23103
rect 14381 23069 14415 23103
rect 16037 23069 16071 23103
rect 16221 23069 16255 23103
rect 18061 23069 18095 23103
rect 18429 23069 18463 23103
rect 18705 23069 18739 23103
rect 20085 23069 20119 23103
rect 20177 23069 20211 23103
rect 21741 23069 21775 23103
rect 21833 23069 21867 23103
rect 22477 23069 22511 23103
rect 23121 23069 23155 23103
rect 23305 23069 23339 23103
rect 24409 23069 24443 23103
rect 24685 23069 24719 23103
rect 25697 23069 25731 23103
rect 25789 23069 25823 23103
rect 26433 23069 26467 23103
rect 26709 23069 26743 23103
rect 28641 23069 28675 23103
rect 28917 23069 28951 23103
rect 31033 23069 31067 23103
rect 5641 23001 5675 23035
rect 5733 23001 5767 23035
rect 7389 23001 7423 23035
rect 8033 23001 8067 23035
rect 11529 23001 11563 23035
rect 14105 23001 14139 23035
rect 17601 23001 17635 23035
rect 17785 23001 17819 23035
rect 20361 23001 20395 23035
rect 20453 23001 20487 23035
rect 20637 23001 20671 23035
rect 20821 23001 20855 23035
rect 21557 23001 21591 23035
rect 22293 23001 22327 23035
rect 22661 23001 22695 23035
rect 24961 23001 24995 23035
rect 25513 23001 25547 23035
rect 29561 23001 29595 23035
rect 29745 23001 29779 23035
rect 31392 23001 31426 23035
rect 3157 22933 3191 22967
rect 3433 22933 3467 22967
rect 4445 22933 4479 22967
rect 5181 22933 5215 22967
rect 6101 22933 6135 22967
rect 7757 22933 7791 22967
rect 8401 22933 8435 22967
rect 11253 22933 11287 22967
rect 11713 22933 11747 22967
rect 18245 22933 18279 22967
rect 18889 22933 18923 22967
rect 22017 22933 22051 22967
rect 22109 22933 22143 22967
rect 22753 22933 22787 22967
rect 22937 22933 22971 22967
rect 29101 22933 29135 22967
rect 29929 22933 29963 22967
rect 30389 22933 30423 22967
rect 32505 22933 32539 22967
rect 2789 22729 2823 22763
rect 3249 22729 3283 22763
rect 3525 22729 3559 22763
rect 6193 22729 6227 22763
rect 7205 22729 7239 22763
rect 7481 22729 7515 22763
rect 11115 22729 11149 22763
rect 12541 22729 12575 22763
rect 13185 22729 13219 22763
rect 19073 22729 19107 22763
rect 19349 22729 19383 22763
rect 20545 22729 20579 22763
rect 25421 22729 25455 22763
rect 30297 22729 30331 22763
rect 3366 22661 3400 22695
rect 3985 22661 4019 22695
rect 4721 22661 4755 22695
rect 6561 22661 6595 22695
rect 9873 22661 9907 22695
rect 12725 22661 12759 22695
rect 16037 22661 16071 22695
rect 21005 22661 21039 22695
rect 30021 22661 30055 22695
rect 30634 22661 30668 22695
rect 1676 22593 1710 22627
rect 2881 22593 2915 22627
rect 4102 22593 4136 22627
rect 4629 22593 4663 22627
rect 4813 22593 4847 22627
rect 4997 22593 5031 22627
rect 5181 22593 5215 22627
rect 5632 22597 5666 22631
rect 5733 22617 5767 22651
rect 6009 22593 6043 22627
rect 6377 22593 6411 22627
rect 6653 22593 6687 22627
rect 6745 22593 6779 22627
rect 7021 22593 7055 22627
rect 7297 22593 7331 22627
rect 7573 22593 7607 22627
rect 8585 22593 8619 22627
rect 8769 22593 8803 22627
rect 8861 22593 8895 22627
rect 8977 22593 9011 22627
rect 10057 22593 10091 22627
rect 10241 22593 10275 22627
rect 11805 22593 11839 22627
rect 11897 22593 11931 22627
rect 12081 22593 12115 22627
rect 12357 22593 12391 22627
rect 13001 22593 13035 22627
rect 16313 22593 16347 22627
rect 17601 22593 17635 22627
rect 18889 22593 18923 22627
rect 19165 22593 19199 22627
rect 19441 22593 19475 22627
rect 19809 22593 19843 22627
rect 20085 22593 20119 22627
rect 20729 22593 20763 22627
rect 20821 22593 20855 22627
rect 21833 22593 21867 22627
rect 22109 22593 22143 22627
rect 22845 22593 22879 22627
rect 25053 22593 25087 22627
rect 25237 22593 25271 22627
rect 27629 22593 27663 22627
rect 27813 22593 27847 22627
rect 29745 22593 29779 22627
rect 29929 22593 29963 22627
rect 30113 22593 30147 22627
rect 32229 22593 32263 22627
rect 1409 22525 1443 22559
rect 3157 22525 3191 22559
rect 3617 22525 3651 22559
rect 3893 22525 3927 22559
rect 9689 22525 9723 22559
rect 11345 22525 11379 22559
rect 12817 22525 12851 22559
rect 16129 22525 16163 22559
rect 19901 22525 19935 22559
rect 21925 22525 21959 22559
rect 30389 22525 30423 22559
rect 4261 22457 4295 22491
rect 5457 22457 5491 22491
rect 5917 22457 5951 22491
rect 9137 22457 9171 22491
rect 10425 22457 10459 22491
rect 12265 22457 12299 22491
rect 4445 22389 4479 22423
rect 5365 22389 5399 22423
rect 6929 22389 6963 22423
rect 7757 22389 7791 22423
rect 11529 22389 11563 22423
rect 11805 22389 11839 22423
rect 12725 22389 12759 22423
rect 16221 22389 16255 22423
rect 16497 22389 16531 22423
rect 17785 22389 17819 22423
rect 19625 22389 19659 22423
rect 19809 22389 19843 22423
rect 20269 22389 20303 22423
rect 20453 22389 20487 22423
rect 20913 22389 20947 22423
rect 21833 22389 21867 22423
rect 22293 22389 22327 22423
rect 23029 22389 23063 22423
rect 27813 22389 27847 22423
rect 27997 22389 28031 22423
rect 31769 22389 31803 22423
rect 32413 22389 32447 22423
rect 2237 22185 2271 22219
rect 5641 22185 5675 22219
rect 8493 22185 8527 22219
rect 13369 22185 13403 22219
rect 21097 22185 21131 22219
rect 22109 22185 22143 22219
rect 22937 22185 22971 22219
rect 24041 22185 24075 22219
rect 25789 22185 25823 22219
rect 31493 22185 31527 22219
rect 4353 22117 4387 22151
rect 5917 22117 5951 22151
rect 9597 22117 9631 22151
rect 17141 22117 17175 22151
rect 19717 22117 19751 22151
rect 4077 22049 4111 22083
rect 4169 22049 4203 22083
rect 11161 22049 11195 22083
rect 11989 22049 12023 22083
rect 15393 22049 15427 22083
rect 22753 22049 22787 22083
rect 25881 22049 25915 22083
rect 32505 22049 32539 22083
rect 2053 21981 2087 22015
rect 2513 21981 2547 22015
rect 2605 21981 2639 22015
rect 2881 21981 2915 22015
rect 3341 21981 3375 22015
rect 3433 21981 3467 22015
rect 3893 21981 3927 22015
rect 3985 21981 4019 22015
rect 4629 21981 4663 22015
rect 4721 21981 4755 22015
rect 4997 21981 5031 22015
rect 5457 21981 5491 22015
rect 5733 21981 5767 22015
rect 6009 21981 6043 22015
rect 6837 21981 6871 22015
rect 7113 21981 7147 22015
rect 7205 21981 7239 22015
rect 8309 21981 8343 22015
rect 8585 21981 8619 22015
rect 8953 21981 8987 22015
rect 9137 21981 9171 22015
rect 9413 21981 9447 22015
rect 10241 21981 10275 22015
rect 10885 21981 10919 22015
rect 11621 21981 11655 22015
rect 11897 21997 11931 22031
rect 12265 21981 12299 22015
rect 13553 21981 13587 22015
rect 13645 21981 13679 22015
rect 15209 21981 15243 22015
rect 16957 21981 16991 22015
rect 17509 21981 17543 22015
rect 17785 21981 17819 22015
rect 18981 21981 19015 22015
rect 21281 21981 21315 22015
rect 22109 21981 22143 22015
rect 22201 21981 22235 22015
rect 22385 21981 22419 22015
rect 22661 21981 22695 22015
rect 22937 21981 22971 22015
rect 23949 21981 23983 22015
rect 24041 21981 24075 22015
rect 26065 21981 26099 22015
rect 30941 21981 30975 22015
rect 31309 21981 31343 22015
rect 31861 21981 31895 22015
rect 7021 21913 7055 21947
rect 10057 21913 10091 21947
rect 11437 21913 11471 21947
rect 13369 21913 13403 21947
rect 15025 21913 15059 21947
rect 17325 21913 17359 21947
rect 21005 21913 21039 21947
rect 23765 21913 23799 21947
rect 25789 21913 25823 21947
rect 31125 21913 31159 21947
rect 31217 21913 31251 21947
rect 2329 21845 2363 21879
rect 2789 21845 2823 21879
rect 3065 21845 3099 21879
rect 3157 21845 3191 21879
rect 3617 21845 3651 21879
rect 4445 21845 4479 21879
rect 4905 21845 4939 21879
rect 5181 21845 5215 21879
rect 6193 21845 6227 21879
rect 7389 21845 7423 21879
rect 8769 21845 8803 21879
rect 9873 21845 9907 21879
rect 11253 21845 11287 21879
rect 11713 21845 11747 21879
rect 13829 21845 13863 21879
rect 17693 21845 17727 21879
rect 17969 21845 18003 21879
rect 21925 21845 21959 21879
rect 23121 21845 23155 21879
rect 24225 21845 24259 21879
rect 26249 21845 26283 21879
rect 2789 21641 2823 21675
rect 3341 21641 3375 21675
rect 3709 21641 3743 21675
rect 4537 21641 4571 21675
rect 5917 21641 5951 21675
rect 7849 21641 7883 21675
rect 9229 21641 9263 21675
rect 13553 21641 13587 21675
rect 17233 21641 17267 21675
rect 19165 21641 19199 21675
rect 19717 21641 19751 21675
rect 27629 21641 27663 21675
rect 28641 21641 28675 21675
rect 29193 21641 29227 21675
rect 31953 21641 31987 21675
rect 3157 21573 3191 21607
rect 3249 21573 3283 21607
rect 3617 21573 3651 21607
rect 3985 21573 4019 21607
rect 6745 21573 6779 21607
rect 10241 21573 10275 21607
rect 16773 21573 16807 21607
rect 20637 21573 20671 21607
rect 23949 21573 23983 21607
rect 24501 21573 24535 21607
rect 28089 21573 28123 21607
rect 1409 21505 1443 21539
rect 1665 21505 1699 21539
rect 2973 21505 3007 21539
rect 4077 21505 4111 21539
rect 4353 21505 4387 21539
rect 4629 21505 4663 21539
rect 5089 21505 5123 21539
rect 5365 21505 5399 21539
rect 5457 21505 5491 21539
rect 5733 21505 5767 21539
rect 6009 21505 6043 21539
rect 6561 21505 6595 21539
rect 6837 21505 6871 21539
rect 6929 21505 6963 21539
rect 7205 21505 7239 21539
rect 7389 21505 7423 21539
rect 7665 21505 7699 21539
rect 7941 21505 7975 21539
rect 9045 21505 9079 21539
rect 9321 21505 9355 21539
rect 9505 21505 9539 21539
rect 9965 21505 9999 21539
rect 10793 21505 10827 21539
rect 10977 21505 11011 21539
rect 11161 21505 11195 21539
rect 11713 21505 11747 21539
rect 11897 21505 11931 21539
rect 13001 21505 13035 21539
rect 13093 21505 13127 21539
rect 13369 21505 13403 21539
rect 14841 21505 14875 21539
rect 16129 21505 16163 21539
rect 16313 21505 16347 21539
rect 17049 21505 17083 21539
rect 17601 21505 17635 21539
rect 17877 21505 17911 21539
rect 17969 21505 18003 21539
rect 18245 21505 18279 21539
rect 18705 21505 18739 21539
rect 18981 21505 19015 21539
rect 19257 21505 19291 21539
rect 19533 21505 19567 21539
rect 19993 21505 20027 21539
rect 20085 21505 20119 21539
rect 20361 21505 20395 21539
rect 20913 21505 20947 21539
rect 24225 21505 24259 21539
rect 24777 21505 24811 21539
rect 26985 21505 27019 21539
rect 27261 21505 27295 21539
rect 27813 21505 27847 21539
rect 28181 21505 28215 21539
rect 28457 21505 28491 21539
rect 28733 21505 28767 21539
rect 29009 21505 29043 21539
rect 30573 21505 30607 21539
rect 30840 21505 30874 21539
rect 32229 21505 32263 21539
rect 3893 21437 3927 21471
rect 9689 21437 9723 21471
rect 10149 21437 10183 21471
rect 12725 21437 12759 21471
rect 13185 21437 13219 21471
rect 16957 21437 16991 21471
rect 17785 21437 17819 21471
rect 18797 21437 18831 21471
rect 19441 21437 19475 21471
rect 20177 21437 20211 21471
rect 20729 21437 20763 21471
rect 24041 21437 24075 21471
rect 24685 21437 24719 21471
rect 27077 21437 27111 21471
rect 27905 21437 27939 21471
rect 28273 21437 28307 21471
rect 28825 21437 28859 21471
rect 4905 21369 4939 21403
rect 9781 21369 9815 21403
rect 12081 21369 12115 21403
rect 16497 21369 16531 21403
rect 20545 21369 20579 21403
rect 24961 21369 24995 21403
rect 3525 21301 3559 21335
rect 3801 21301 3835 21335
rect 4261 21301 4295 21335
rect 4813 21301 4847 21335
rect 5181 21301 5215 21335
rect 5641 21301 5675 21335
rect 6193 21301 6227 21335
rect 7113 21301 7147 21335
rect 8125 21301 8159 21335
rect 10241 21301 10275 21335
rect 11345 21301 11379 21335
rect 13369 21301 13403 21335
rect 14657 21301 14691 21335
rect 16865 21301 16899 21335
rect 17417 21301 17451 21335
rect 17693 21301 17727 21335
rect 18153 21301 18187 21335
rect 18429 21301 18463 21335
rect 18981 21301 19015 21335
rect 19533 21301 19567 21335
rect 19809 21301 19843 21335
rect 20269 21301 20303 21335
rect 20821 21301 20855 21335
rect 21097 21301 21131 21335
rect 23857 21301 23891 21335
rect 24225 21301 24259 21335
rect 24409 21301 24443 21335
rect 24501 21301 24535 21335
rect 26985 21301 27019 21335
rect 27445 21301 27479 21335
rect 28089 21301 28123 21335
rect 28273 21301 28307 21335
rect 28733 21301 28767 21335
rect 32413 21301 32447 21335
rect 2237 21097 2271 21131
rect 2513 21097 2547 21131
rect 4537 21097 4571 21131
rect 9965 21097 9999 21131
rect 12173 21097 12207 21131
rect 12633 21097 12667 21131
rect 12817 21097 12851 21131
rect 14749 21097 14783 21131
rect 14933 21097 14967 21131
rect 21557 21097 21591 21131
rect 22017 21097 22051 21131
rect 25789 21097 25823 21131
rect 25881 21097 25915 21131
rect 27169 21097 27203 21131
rect 31309 21097 31343 21131
rect 1961 21029 1995 21063
rect 2697 21029 2731 21063
rect 5641 21029 5675 21063
rect 8769 21029 8803 21063
rect 10057 21029 10091 21063
rect 26249 21029 26283 21063
rect 32321 21029 32355 21063
rect 10425 20961 10459 20995
rect 12265 20961 12299 20995
rect 21649 20961 21683 20995
rect 27353 20961 27387 20995
rect 32229 20961 32263 20995
rect 1501 20893 1535 20927
rect 1777 20893 1811 20927
rect 2053 20893 2087 20927
rect 2329 20893 2363 20927
rect 3985 20893 4019 20927
rect 4169 20893 4203 20927
rect 4353 20893 4387 20927
rect 4721 20893 4755 20927
rect 4813 20893 4847 20927
rect 5181 20893 5215 20927
rect 5457 20893 5491 20927
rect 5733 20893 5767 20927
rect 6101 20893 6135 20927
rect 8217 20893 8251 20927
rect 8585 20893 8619 20927
rect 9413 20893 9447 20927
rect 9781 20893 9815 20927
rect 10241 20893 10275 20927
rect 12081 20893 12115 20927
rect 12449 20893 12483 20927
rect 12909 20893 12943 20927
rect 13093 20893 13127 20927
rect 14473 20893 14507 20927
rect 14657 20893 14691 20927
rect 14749 20893 14783 20927
rect 20177 20889 20211 20923
rect 21833 20893 21867 20927
rect 25605 20893 25639 20927
rect 25881 20893 25915 20927
rect 26065 20893 26099 20927
rect 27169 20893 27203 20927
rect 27445 20893 27479 20927
rect 30757 20893 30791 20927
rect 30941 20893 30975 20927
rect 31125 20893 31159 20927
rect 31585 20893 31619 20927
rect 32505 20893 32539 20927
rect 2697 20825 2731 20859
rect 4077 20825 4111 20859
rect 4997 20825 5031 20859
rect 5089 20825 5123 20859
rect 5917 20825 5951 20859
rect 6009 20825 6043 20859
rect 8401 20825 8435 20859
rect 8493 20825 8527 20859
rect 9597 20825 9631 20859
rect 9689 20825 9723 20859
rect 12173 20825 12207 20859
rect 21557 20825 21591 20859
rect 31033 20825 31067 20859
rect 1685 20757 1719 20791
rect 3157 20757 3191 20791
rect 3249 20757 3283 20791
rect 3433 20757 3467 20791
rect 3801 20757 3835 20791
rect 5365 20757 5399 20791
rect 6285 20757 6319 20791
rect 13277 20757 13311 20791
rect 20361 20757 20395 20791
rect 26985 20757 27019 20791
rect 27629 20757 27663 20791
rect 2421 20553 2455 20587
rect 3709 20553 3743 20587
rect 5733 20553 5767 20587
rect 18429 20553 18463 20587
rect 21281 20553 21315 20587
rect 30389 20553 30423 20587
rect 2538 20485 2572 20519
rect 2881 20485 2915 20519
rect 3433 20485 3467 20519
rect 5365 20485 5399 20519
rect 8125 20485 8159 20519
rect 8217 20485 8251 20519
rect 10977 20485 11011 20519
rect 13829 20485 13863 20519
rect 14565 20485 14599 20519
rect 15485 20485 15519 20519
rect 15945 20485 15979 20519
rect 17969 20485 18003 20519
rect 20821 20485 20855 20519
rect 22753 20485 22787 20519
rect 30849 20485 30883 20519
rect 30941 20485 30975 20519
rect 1777 20417 1811 20451
rect 2053 20417 2087 20451
rect 3893 20417 3927 20451
rect 3985 20417 4019 20451
rect 4445 20417 4479 20451
rect 4721 20417 4755 20451
rect 5089 20417 5123 20451
rect 5181 20417 5215 20451
rect 5457 20417 5491 20451
rect 5549 20417 5583 20451
rect 5825 20417 5859 20451
rect 7941 20417 7975 20451
rect 8309 20417 8343 20451
rect 10517 20417 10551 20451
rect 10793 20417 10827 20451
rect 11161 20417 11195 20451
rect 11529 20417 11563 20451
rect 11713 20417 11747 20451
rect 11805 20417 11839 20451
rect 12265 20417 12299 20451
rect 12357 20417 12391 20451
rect 14105 20417 14139 20451
rect 15301 20417 15335 20451
rect 15761 20417 15795 20451
rect 16681 20417 16715 20451
rect 16865 20417 16899 20451
rect 16957 20417 16991 20451
rect 18245 20417 18279 20451
rect 18889 20417 18923 20451
rect 19993 20417 20027 20451
rect 20269 20417 20303 20451
rect 21097 20417 21131 20451
rect 22569 20417 22603 20451
rect 24225 20417 24259 20451
rect 24501 20417 24535 20451
rect 30021 20417 30055 20451
rect 30665 20417 30699 20451
rect 31033 20417 31067 20451
rect 31309 20417 31343 20451
rect 32229 20417 32263 20451
rect 2329 20349 2363 20383
rect 3341 20349 3375 20383
rect 14013 20349 14047 20383
rect 14381 20349 14415 20383
rect 18153 20349 18187 20383
rect 18981 20349 19015 20383
rect 20085 20349 20119 20383
rect 20913 20349 20947 20383
rect 24317 20349 24351 20383
rect 30113 20349 30147 20383
rect 31953 20349 31987 20383
rect 1961 20281 1995 20315
rect 2697 20281 2731 20315
rect 2881 20281 2915 20315
rect 4261 20281 4295 20315
rect 4537 20281 4571 20315
rect 11989 20281 12023 20315
rect 12081 20281 12115 20315
rect 12541 20281 12575 20315
rect 17141 20281 17175 20315
rect 19257 20281 19291 20315
rect 20453 20281 20487 20315
rect 3617 20213 3651 20247
rect 4169 20213 4203 20247
rect 4905 20213 4939 20247
rect 6009 20213 6043 20247
rect 8493 20213 8527 20247
rect 10701 20213 10735 20247
rect 11529 20213 11563 20247
rect 14013 20213 14047 20247
rect 14289 20213 14323 20247
rect 15669 20213 15703 20247
rect 16129 20213 16163 20247
rect 16681 20213 16715 20247
rect 17785 20213 17819 20247
rect 17969 20213 18003 20247
rect 18797 20213 18831 20247
rect 18889 20213 18923 20247
rect 20269 20213 20303 20247
rect 20821 20213 20855 20247
rect 22937 20213 22971 20247
rect 24409 20213 24443 20247
rect 24685 20213 24719 20247
rect 30021 20213 30055 20247
rect 31217 20213 31251 20247
rect 32413 20213 32447 20247
rect 3433 20009 3467 20043
rect 5641 20009 5675 20043
rect 8217 20009 8251 20043
rect 9413 20009 9447 20043
rect 13737 20009 13771 20043
rect 14657 20009 14691 20043
rect 14841 20009 14875 20043
rect 16497 20009 16531 20043
rect 16957 20009 16991 20043
rect 20729 20009 20763 20043
rect 20913 20009 20947 20043
rect 24409 20009 24443 20043
rect 24777 20009 24811 20043
rect 26065 20009 26099 20043
rect 26525 20009 26559 20043
rect 26801 20009 26835 20043
rect 27905 20009 27939 20043
rect 27997 20009 28031 20043
rect 29561 20009 29595 20043
rect 30205 20009 30239 20043
rect 30573 20009 30607 20043
rect 30849 20009 30883 20043
rect 32505 20009 32539 20043
rect 2789 19941 2823 19975
rect 3801 19941 3835 19975
rect 5549 19941 5583 19975
rect 29929 19941 29963 19975
rect 1409 19873 1443 19907
rect 10241 19873 10275 19907
rect 12265 19873 12299 19907
rect 13645 19873 13679 19907
rect 14473 19873 14507 19907
rect 24501 19873 24535 19907
rect 26249 19873 26283 19907
rect 26709 19873 26743 19907
rect 28089 19873 28123 19907
rect 30297 19873 30331 19907
rect 2973 19805 3007 19839
rect 3065 19805 3099 19839
rect 3157 19805 3191 19839
rect 3249 19805 3283 19839
rect 3985 19805 4019 19839
rect 4353 19805 4387 19839
rect 4629 19805 4663 19839
rect 4721 19805 4755 19839
rect 4997 19805 5031 19839
rect 5365 19805 5399 19839
rect 5825 19805 5859 19839
rect 6101 19805 6135 19839
rect 6377 19805 6411 19839
rect 6469 19805 6503 19839
rect 7021 19805 7055 19839
rect 7297 19805 7331 19839
rect 7389 19805 7423 19839
rect 7665 19805 7699 19839
rect 8401 19805 8435 19839
rect 8953 19805 8987 19839
rect 9229 19805 9263 19839
rect 9413 19805 9447 19839
rect 10057 19805 10091 19839
rect 10517 19781 10551 19815
rect 11989 19805 12023 19839
rect 13461 19805 13495 19839
rect 13737 19805 13771 19839
rect 14105 19805 14139 19839
rect 14657 19805 14691 19839
rect 16681 19805 16715 19839
rect 16773 19805 16807 19839
rect 16957 19805 16991 19839
rect 20913 19805 20947 19839
rect 21097 19805 21131 19839
rect 24409 19805 24443 19839
rect 25789 19805 25823 19839
rect 26065 19805 26099 19839
rect 26341 19805 26375 19839
rect 26617 19805 26651 19839
rect 26893 19805 26927 19839
rect 27997 19805 28031 19839
rect 29561 19805 29595 19839
rect 29653 19805 29687 19839
rect 30205 19805 30239 19839
rect 30665 19805 30699 19839
rect 31125 19805 31159 19839
rect 31381 19805 31415 19839
rect 1676 19737 1710 19771
rect 4537 19737 4571 19771
rect 5181 19737 5215 19771
rect 5273 19737 5307 19771
rect 6285 19737 6319 19771
rect 7205 19737 7239 19771
rect 7941 19737 7975 19771
rect 8125 19737 8159 19771
rect 8585 19737 8619 19771
rect 9873 19737 9907 19771
rect 14381 19737 14415 19771
rect 28457 19737 28491 19771
rect 28641 19737 28675 19771
rect 30021 19737 30055 19771
rect 4905 19669 4939 19703
rect 6653 19669 6687 19703
rect 7573 19669 7607 19703
rect 7849 19669 7883 19703
rect 9137 19669 9171 19703
rect 9597 19669 9631 19703
rect 10333 19669 10367 19703
rect 13921 19669 13955 19703
rect 14289 19669 14323 19703
rect 25973 19669 26007 19703
rect 27077 19669 27111 19703
rect 28365 19669 28399 19703
rect 28825 19669 28859 19703
rect 1593 19465 1627 19499
rect 4537 19465 4571 19499
rect 11529 19465 11563 19499
rect 13645 19465 13679 19499
rect 16221 19465 16255 19499
rect 20637 19465 20671 19499
rect 24133 19465 24167 19499
rect 24869 19465 24903 19499
rect 26617 19465 26651 19499
rect 29377 19465 29411 19499
rect 30297 19465 30331 19499
rect 32413 19465 32447 19499
rect 7573 19397 7607 19431
rect 11989 19397 12023 19431
rect 14105 19397 14139 19431
rect 15025 19397 15059 19431
rect 15768 19397 15802 19431
rect 19809 19397 19843 19431
rect 28917 19397 28951 19431
rect 30849 19397 30883 19431
rect 30941 19397 30975 19431
rect 1409 19329 1443 19363
rect 4077 19329 4111 19363
rect 4445 19329 4479 19363
rect 4721 19329 4755 19363
rect 5273 19313 5307 19347
rect 11713 19329 11747 19363
rect 11897 19329 11931 19363
rect 12265 19329 12299 19363
rect 13369 19329 13403 19363
rect 13829 19329 13863 19363
rect 14013 19329 14047 19363
rect 14289 19329 14323 19363
rect 14749 19329 14783 19363
rect 15209 19329 15243 19363
rect 15317 19329 15351 19363
rect 15945 19329 15979 19363
rect 16037 19329 16071 19363
rect 19993 19329 20027 19363
rect 20269 19329 20303 19363
rect 22753 19329 22787 19363
rect 23673 19329 23707 19363
rect 23857 19329 23891 19363
rect 23949 19329 23983 19363
rect 24409 19329 24443 19363
rect 24593 19329 24627 19363
rect 24685 19329 24719 19363
rect 25605 19329 25639 19363
rect 25789 19329 25823 19363
rect 25881 19329 25915 19363
rect 26157 19329 26191 19363
rect 26341 19329 26375 19363
rect 26433 19329 26467 19363
rect 27721 19329 27755 19363
rect 29101 19329 29135 19363
rect 29193 19329 29227 19363
rect 30113 19329 30147 19363
rect 30573 19329 30607 19363
rect 30665 19329 30699 19363
rect 31033 19329 31067 19363
rect 31309 19329 31343 19363
rect 32229 19329 32263 19363
rect 12173 19261 12207 19295
rect 14565 19261 14599 19295
rect 15669 19261 15703 19295
rect 20361 19261 20395 19295
rect 27813 19261 27847 19295
rect 31953 19261 31987 19295
rect 5089 19193 5123 19227
rect 12449 19193 12483 19227
rect 13553 19193 13587 19227
rect 14933 19193 14967 19227
rect 15485 19193 15519 19227
rect 16313 19193 16347 19227
rect 30389 19193 30423 19227
rect 3893 19125 3927 19159
rect 4261 19125 4295 19159
rect 7665 19125 7699 19159
rect 11897 19125 11931 19159
rect 12265 19125 12299 19159
rect 14473 19125 14507 19159
rect 15117 19125 15151 19159
rect 15761 19125 15795 19159
rect 20177 19125 20211 19159
rect 20269 19125 20303 19159
rect 22937 19125 22971 19159
rect 23949 19125 23983 19159
rect 24409 19125 24443 19159
rect 25881 19125 25915 19159
rect 26065 19125 26099 19159
rect 26341 19125 26375 19159
rect 27813 19125 27847 19159
rect 28089 19125 28123 19159
rect 29193 19125 29227 19159
rect 31217 19125 31251 19159
rect 2789 18921 2823 18955
rect 6837 18921 6871 18955
rect 7941 18921 7975 18955
rect 9229 18921 9263 18955
rect 9965 18921 9999 18955
rect 10241 18921 10275 18955
rect 10517 18921 10551 18955
rect 11621 18921 11655 18955
rect 12081 18921 12115 18955
rect 12633 18921 12667 18955
rect 14565 18921 14599 18955
rect 17233 18921 17267 18955
rect 19257 18921 19291 18955
rect 21281 18921 21315 18955
rect 21465 18921 21499 18955
rect 21833 18921 21867 18955
rect 22109 18921 22143 18955
rect 22477 18921 22511 18955
rect 23029 18921 23063 18955
rect 23765 18921 23799 18955
rect 24133 18921 24167 18955
rect 24961 18921 24995 18955
rect 30757 18921 30791 18955
rect 32505 18921 32539 18955
rect 8309 18853 8343 18887
rect 9689 18853 9723 18887
rect 17693 18853 17727 18887
rect 19717 18853 19751 18887
rect 1409 18785 1443 18819
rect 8033 18785 8067 18819
rect 9321 18785 9355 18819
rect 9873 18785 9907 18819
rect 11713 18785 11747 18819
rect 17141 18785 17175 18819
rect 17325 18785 17359 18819
rect 19349 18785 19383 18819
rect 21741 18785 21775 18819
rect 22201 18785 22235 18819
rect 22845 18785 22879 18819
rect 23305 18785 23339 18819
rect 31125 18785 31159 18819
rect 3341 18717 3375 18751
rect 3433 18717 3467 18751
rect 3985 18717 4019 18751
rect 4261 18717 4295 18751
rect 4445 18717 4479 18751
rect 5365 18717 5399 18751
rect 5917 18717 5951 18751
rect 6101 18717 6135 18751
rect 6377 18717 6411 18751
rect 6653 18717 6687 18751
rect 7021 18717 7055 18751
rect 7481 18717 7515 18751
rect 7941 18717 7975 18751
rect 9505 18717 9539 18751
rect 10057 18717 10091 18751
rect 10333 18717 10367 18751
rect 10609 18717 10643 18751
rect 11345 18717 11379 18751
rect 11529 18717 11563 18751
rect 11937 18717 11971 18751
rect 12357 18717 12391 18751
rect 12817 18717 12851 18751
rect 14197 18717 14231 18751
rect 16957 18717 16991 18751
rect 17509 18717 17543 18751
rect 17785 18717 17819 18751
rect 19533 18717 19567 18751
rect 21097 18717 21131 18751
rect 21281 18717 21315 18751
rect 21833 18717 21867 18751
rect 22109 18717 22143 18751
rect 22661 18717 22695 18751
rect 23029 18717 23063 18751
rect 23765 18717 23799 18751
rect 23857 18717 23891 18751
rect 24961 18717 24995 18751
rect 25145 18717 25179 18751
rect 29101 18717 29135 18751
rect 29285 18717 29319 18751
rect 30573 18717 30607 18751
rect 31033 18717 31067 18751
rect 31381 18717 31415 18751
rect 1676 18649 1710 18683
rect 7205 18649 7239 18683
rect 7297 18649 7331 18683
rect 9229 18649 9263 18683
rect 9781 18649 9815 18683
rect 11610 18649 11644 18683
rect 12541 18649 12575 18683
rect 14381 18649 14415 18683
rect 14657 18649 14691 18683
rect 17233 18649 17267 18683
rect 19257 18649 19291 18683
rect 21557 18649 21591 18683
rect 22753 18649 22787 18683
rect 23489 18649 23523 18683
rect 23673 18649 23707 18683
rect 24869 18649 24903 18683
rect 3157 18581 3191 18615
rect 3617 18581 3651 18615
rect 3801 18581 3835 18615
rect 5181 18581 5215 18615
rect 6561 18581 6595 18615
rect 7665 18581 7699 18615
rect 10793 18581 10827 18615
rect 12173 18581 12207 18615
rect 16773 18581 16807 18615
rect 17969 18581 18003 18615
rect 22017 18581 22051 18615
rect 23213 18581 23247 18615
rect 25329 18581 25363 18615
rect 29193 18581 29227 18615
rect 30849 18581 30883 18615
rect 2421 18377 2455 18411
rect 3525 18377 3559 18411
rect 3617 18377 3651 18411
rect 7297 18377 7331 18411
rect 9413 18377 9447 18411
rect 12173 18377 12207 18411
rect 12541 18377 12575 18411
rect 23857 18377 23891 18411
rect 28365 18377 28399 18411
rect 30481 18377 30515 18411
rect 31953 18377 31987 18411
rect 2881 18309 2915 18343
rect 2973 18309 3007 18343
rect 5089 18309 5123 18343
rect 9781 18309 9815 18343
rect 16957 18309 16991 18343
rect 19165 18309 19199 18343
rect 23673 18309 23707 18343
rect 2605 18241 2639 18275
rect 2697 18241 2731 18275
rect 3111 18241 3145 18275
rect 3341 18241 3375 18275
rect 3801 18241 3835 18275
rect 4353 18241 4387 18275
rect 4813 18241 4847 18275
rect 4997 18241 5031 18275
rect 5181 18241 5215 18275
rect 7481 18241 7515 18275
rect 7757 18241 7791 18275
rect 7849 18241 7883 18275
rect 9597 18241 9631 18275
rect 12357 18241 12391 18275
rect 13461 18265 13495 18299
rect 14565 18241 14599 18275
rect 14841 18241 14875 18275
rect 15393 18241 15427 18275
rect 17233 18241 17267 18275
rect 18889 18241 18923 18275
rect 18981 18241 19015 18275
rect 23489 18241 23523 18275
rect 26433 18241 26467 18275
rect 27905 18241 27939 18275
rect 28181 18241 28215 18275
rect 29745 18241 29779 18275
rect 29929 18241 29963 18275
rect 30297 18241 30331 18275
rect 30573 18241 30607 18275
rect 30840 18241 30874 18275
rect 32229 18241 32263 18275
rect 7573 18173 7607 18207
rect 14289 18173 14323 18207
rect 14657 18173 14691 18207
rect 17049 18173 17083 18207
rect 27997 18173 28031 18207
rect 3249 18105 3283 18139
rect 8033 18105 8067 18139
rect 17417 18105 17451 18139
rect 4169 18037 4203 18071
rect 5365 18037 5399 18071
rect 7665 18037 7699 18071
rect 13645 18037 13679 18071
rect 14381 18037 14415 18071
rect 14841 18037 14875 18071
rect 15209 18037 15243 18071
rect 17233 18037 17267 18071
rect 18705 18037 18739 18071
rect 19165 18037 19199 18071
rect 27905 18037 27939 18071
rect 30113 18037 30147 18071
rect 32413 18037 32447 18071
rect 2697 17833 2731 17867
rect 12449 17833 12483 17867
rect 14105 17833 14139 17867
rect 14657 17833 14691 17867
rect 15117 17833 15151 17867
rect 17325 17833 17359 17867
rect 21833 17833 21867 17867
rect 22937 17833 22971 17867
rect 23397 17833 23431 17867
rect 26249 17833 26283 17867
rect 26801 17833 26835 17867
rect 27261 17833 27295 17867
rect 30849 17833 30883 17867
rect 31493 17833 31527 17867
rect 4537 17765 4571 17799
rect 7573 17765 7607 17799
rect 9965 17765 9999 17799
rect 12633 17765 12667 17799
rect 13553 17765 13587 17799
rect 14841 17765 14875 17799
rect 12265 17697 12299 17731
rect 13461 17697 13495 17731
rect 14473 17697 14507 17731
rect 17417 17697 17451 17731
rect 21925 17697 21959 17731
rect 23029 17697 23063 17731
rect 26157 17697 26191 17731
rect 26433 17697 26467 17731
rect 26985 17697 27019 17731
rect 32229 17697 32263 17731
rect 2881 17629 2915 17663
rect 3157 17629 3191 17663
rect 3433 17629 3467 17663
rect 3985 17629 4019 17663
rect 4169 17629 4203 17663
rect 4353 17629 4387 17663
rect 4813 17629 4847 17663
rect 5089 17629 5123 17663
rect 5549 17629 5583 17663
rect 5825 17629 5859 17663
rect 7757 17629 7791 17663
rect 9781 17629 9815 17663
rect 10057 17629 10091 17663
rect 10517 17629 10551 17663
rect 12449 17629 12483 17663
rect 12725 17629 12759 17663
rect 13277 17629 13311 17663
rect 13737 17629 13771 17663
rect 14289 17629 14323 17663
rect 14657 17629 14691 17663
rect 15025 17629 15059 17663
rect 15117 17629 15151 17663
rect 17325 17629 17359 17663
rect 19993 17629 20027 17663
rect 20821 17629 20855 17663
rect 22109 17629 22143 17663
rect 22937 17629 22971 17663
rect 23213 17629 23247 17663
rect 26525 17629 26559 17663
rect 27077 17629 27111 17663
rect 28733 17629 28767 17663
rect 28917 17629 28951 17663
rect 30665 17629 30699 17663
rect 30941 17629 30975 17663
rect 31217 17629 31251 17663
rect 31309 17629 31343 17663
rect 31677 17629 31711 17663
rect 4261 17561 4295 17595
rect 12173 17561 12207 17595
rect 13093 17561 13127 17595
rect 13921 17561 13955 17595
rect 14381 17561 14415 17595
rect 20177 17561 20211 17595
rect 20637 17561 20671 17595
rect 21833 17561 21867 17595
rect 24409 17561 24443 17595
rect 26249 17561 26283 17595
rect 26801 17561 26835 17595
rect 31125 17561 31159 17595
rect 2973 17493 3007 17527
rect 3249 17493 3283 17527
rect 4629 17493 4663 17527
rect 4905 17493 4939 17527
rect 5365 17493 5399 17527
rect 5641 17493 5675 17527
rect 10241 17493 10275 17527
rect 10333 17493 10367 17527
rect 12909 17493 12943 17527
rect 15393 17493 15427 17527
rect 17693 17493 17727 17527
rect 19809 17493 19843 17527
rect 20453 17493 20487 17527
rect 22293 17493 22327 17527
rect 26709 17493 26743 17527
rect 28549 17493 28583 17527
rect 5825 17289 5859 17323
rect 7113 17289 7147 17323
rect 10609 17289 10643 17323
rect 15117 17289 15151 17323
rect 18153 17289 18187 17323
rect 24685 17289 24719 17323
rect 27445 17289 27479 17323
rect 28641 17289 28675 17323
rect 2605 17221 2639 17255
rect 4445 17221 4479 17255
rect 4537 17221 4571 17255
rect 5457 17221 5491 17255
rect 7389 17221 7423 17255
rect 9321 17221 9355 17255
rect 10057 17221 10091 17255
rect 10149 17221 10183 17255
rect 12265 17221 12299 17255
rect 16681 17221 16715 17255
rect 22569 17221 22603 17255
rect 25605 17221 25639 17255
rect 28181 17221 28215 17255
rect 28917 17221 28951 17255
rect 2421 17153 2455 17187
rect 2697 17153 2731 17187
rect 2789 17153 2823 17187
rect 4261 17153 4295 17187
rect 4629 17153 4663 17187
rect 5273 17153 5307 17187
rect 5549 17153 5583 17187
rect 5641 17153 5675 17187
rect 6377 17153 6411 17187
rect 6561 17153 6595 17187
rect 6653 17153 6687 17187
rect 6929 17153 6963 17187
rect 7205 17153 7239 17187
rect 7481 17153 7515 17187
rect 7573 17153 7607 17187
rect 7849 17153 7883 17187
rect 8125 17153 8159 17187
rect 9505 17153 9539 17187
rect 9781 17153 9815 17187
rect 10333 17153 10367 17187
rect 10425 17153 10459 17187
rect 10885 17153 10919 17187
rect 11069 17153 11103 17187
rect 11161 17153 11195 17187
rect 11713 17153 11747 17187
rect 11989 17153 12023 17187
rect 12541 17153 12575 17187
rect 13921 17153 13955 17187
rect 14749 17153 14783 17187
rect 21925 17153 21959 17187
rect 22109 17153 22143 17187
rect 22201 17153 22235 17187
rect 22753 17153 22787 17187
rect 24225 17153 24259 17187
rect 24409 17153 24443 17187
rect 24501 17153 24535 17187
rect 25789 17153 25823 17187
rect 26985 17153 27019 17187
rect 27169 17153 27203 17187
rect 27261 17153 27295 17187
rect 27629 17153 27663 17187
rect 27905 17153 27939 17187
rect 28457 17153 28491 17187
rect 28733 17153 28767 17187
rect 30573 17153 30607 17187
rect 30840 17153 30874 17187
rect 32229 17153 32263 17187
rect 8033 17085 8067 17119
rect 9965 17085 9999 17119
rect 11897 17085 11931 17119
rect 12357 17085 12391 17119
rect 14841 17085 14875 17119
rect 22845 17085 22879 17119
rect 27721 17085 27755 17119
rect 28273 17085 28307 17119
rect 4813 17017 4847 17051
rect 9597 17017 9631 17051
rect 11345 17017 11379 17051
rect 14105 17017 14139 17051
rect 22385 17017 22419 17051
rect 25973 17017 26007 17051
rect 31953 17017 31987 17051
rect 32413 17017 32447 17051
rect 2973 16949 3007 16983
rect 6469 16949 6503 16983
rect 6837 16949 6871 16983
rect 7757 16949 7791 16983
rect 8125 16949 8159 16983
rect 8309 16949 8343 16983
rect 9137 16949 9171 16983
rect 9781 16949 9815 16983
rect 10149 16949 10183 16983
rect 10885 16949 10919 16983
rect 11713 16949 11747 16983
rect 12173 16949 12207 16983
rect 12265 16949 12299 16983
rect 12725 16949 12759 16983
rect 14749 16949 14783 16983
rect 21925 16949 21959 16983
rect 22753 16949 22787 16983
rect 23121 16949 23155 16983
rect 24041 16949 24075 16983
rect 24501 16949 24535 16983
rect 26985 16949 27019 16983
rect 27629 16949 27663 16983
rect 28089 16949 28123 16983
rect 28181 16949 28215 16983
rect 29101 16949 29135 16983
rect 8033 16745 8067 16779
rect 8401 16745 8435 16779
rect 9965 16745 9999 16779
rect 12817 16745 12851 16779
rect 13277 16745 13311 16779
rect 15761 16745 15795 16779
rect 16037 16745 16071 16779
rect 16497 16745 16531 16779
rect 16681 16745 16715 16779
rect 17141 16745 17175 16779
rect 17969 16745 18003 16779
rect 18705 16745 18739 16779
rect 20361 16745 20395 16779
rect 25421 16745 25455 16779
rect 25697 16745 25731 16779
rect 28089 16745 28123 16779
rect 28365 16745 28399 16779
rect 28733 16745 28767 16779
rect 29009 16745 29043 16779
rect 31585 16745 31619 16779
rect 14933 16677 14967 16711
rect 8309 16609 8343 16643
rect 15577 16609 15611 16643
rect 16773 16609 16807 16643
rect 17325 16609 17359 16643
rect 18521 16609 18555 16643
rect 20177 16609 20211 16643
rect 25329 16609 25363 16643
rect 27997 16609 28031 16643
rect 28733 16609 28767 16643
rect 29101 16609 29135 16643
rect 32321 16609 32355 16643
rect 1409 16541 1443 16575
rect 2697 16541 2731 16575
rect 2973 16541 3007 16575
rect 3065 16541 3099 16575
rect 4353 16541 4387 16575
rect 4629 16541 4663 16575
rect 4721 16541 4755 16575
rect 5365 16541 5399 16575
rect 5549 16541 5583 16575
rect 5733 16541 5767 16575
rect 8401 16541 8435 16575
rect 9505 16541 9539 16575
rect 12817 16541 12851 16575
rect 13001 16541 13035 16575
rect 13461 16541 13495 16575
rect 14749 16541 14783 16575
rect 15209 16541 15243 16575
rect 15393 16541 15427 16575
rect 15761 16541 15795 16575
rect 16681 16541 16715 16575
rect 17417 16541 17451 16575
rect 17969 16541 18003 16575
rect 18061 16541 18095 16575
rect 18705 16541 18739 16575
rect 20085 16541 20119 16575
rect 25513 16541 25547 16575
rect 27905 16541 27939 16575
rect 28181 16541 28215 16575
rect 28825 16541 28859 16575
rect 29009 16541 29043 16575
rect 31033 16541 31067 16575
rect 31401 16541 31435 16575
rect 31769 16541 31803 16575
rect 2881 16473 2915 16507
rect 4537 16473 4571 16507
rect 5641 16473 5675 16507
rect 10149 16473 10183 16507
rect 10333 16473 10367 16507
rect 13645 16473 13679 16507
rect 15025 16473 15059 16507
rect 15485 16473 15519 16507
rect 16221 16473 16255 16507
rect 16405 16473 16439 16507
rect 16957 16473 16991 16507
rect 17141 16473 17175 16507
rect 18429 16473 18463 16507
rect 20361 16473 20395 16507
rect 25237 16473 25271 16507
rect 31217 16473 31251 16507
rect 31309 16473 31343 16507
rect 1593 16405 1627 16439
rect 3249 16405 3283 16439
rect 4905 16405 4939 16439
rect 5917 16405 5951 16439
rect 9689 16405 9723 16439
rect 13185 16405 13219 16439
rect 15945 16405 15979 16439
rect 17601 16405 17635 16439
rect 18337 16405 18371 16439
rect 18889 16405 18923 16439
rect 19901 16405 19935 16439
rect 28457 16405 28491 16439
rect 29377 16405 29411 16439
rect 4169 16201 4203 16235
rect 10517 16201 10551 16235
rect 13001 16201 13035 16235
rect 20453 16201 20487 16235
rect 23489 16201 23523 16235
rect 25881 16201 25915 16235
rect 30205 16201 30239 16235
rect 2881 16133 2915 16167
rect 6009 16133 6043 16167
rect 6653 16133 6687 16167
rect 8493 16133 8527 16167
rect 12541 16133 12575 16167
rect 19809 16133 19843 16167
rect 19993 16133 20027 16167
rect 22845 16133 22879 16167
rect 30941 16133 30975 16167
rect 2605 16065 2639 16099
rect 2789 16065 2823 16099
rect 2973 16065 3007 16099
rect 4353 16065 4387 16099
rect 4537 16065 4571 16099
rect 6837 16065 6871 16099
rect 7021 16065 7055 16099
rect 8677 16065 8711 16099
rect 8861 16065 8895 16099
rect 10701 16065 10735 16099
rect 10793 16065 10827 16099
rect 10977 16065 11011 16099
rect 11253 16065 11287 16099
rect 12817 16065 12851 16099
rect 15290 16065 15324 16099
rect 15485 16065 15519 16099
rect 15577 16065 15611 16099
rect 20269 16065 20303 16099
rect 20545 16065 20579 16099
rect 20729 16065 20763 16099
rect 20821 16065 20855 16099
rect 23121 16065 23155 16099
rect 23581 16065 23615 16099
rect 25513 16065 25547 16099
rect 25697 16065 25731 16099
rect 26433 16065 26467 16099
rect 29745 16065 29779 16099
rect 30021 16065 30055 16099
rect 30573 16065 30607 16099
rect 30665 16065 30699 16099
rect 30849 16065 30883 16099
rect 31033 16065 31067 16099
rect 31309 16065 31343 16099
rect 31953 16065 31987 16099
rect 32229 16065 32263 16099
rect 7205 15997 7239 16031
rect 12725 15997 12759 16031
rect 20085 15997 20119 16031
rect 22937 15997 22971 16031
rect 23673 15997 23707 16031
rect 26525 15997 26559 16031
rect 29837 15997 29871 16031
rect 4721 15929 4755 15963
rect 6469 15929 6503 15963
rect 15761 15929 15795 15963
rect 26801 15929 26835 15963
rect 3157 15861 3191 15895
rect 6101 15861 6135 15895
rect 10701 15861 10735 15895
rect 11161 15861 11195 15895
rect 12541 15861 12575 15895
rect 15577 15861 15611 15895
rect 19993 15861 20027 15895
rect 20545 15861 20579 15895
rect 21005 15861 21039 15895
rect 22845 15861 22879 15895
rect 23305 15861 23339 15895
rect 23581 15861 23615 15895
rect 23949 15861 23983 15895
rect 25513 15861 25547 15895
rect 26341 15861 26375 15895
rect 26433 15861 26467 15895
rect 29745 15861 29779 15895
rect 30389 15861 30423 15895
rect 31217 15861 31251 15895
rect 32413 15861 32447 15895
rect 3985 15657 4019 15691
rect 5457 15657 5491 15691
rect 6745 15657 6779 15691
rect 13737 15657 13771 15691
rect 15025 15657 15059 15691
rect 15209 15657 15243 15691
rect 16405 15657 16439 15691
rect 16773 15657 16807 15691
rect 21925 15657 21959 15691
rect 22385 15657 22419 15691
rect 22477 15657 22511 15691
rect 23029 15657 23063 15691
rect 27261 15657 27295 15691
rect 29653 15657 29687 15691
rect 30205 15657 30239 15691
rect 30573 15657 30607 15691
rect 32505 15657 32539 15691
rect 9597 15589 9631 15623
rect 10241 15589 10275 15623
rect 10609 15589 10643 15623
rect 15485 15589 15519 15623
rect 27445 15589 27479 15623
rect 30113 15589 30147 15623
rect 4353 15521 4387 15555
rect 14841 15521 14875 15555
rect 16497 15521 16531 15555
rect 22201 15521 22235 15555
rect 23121 15521 23155 15555
rect 27077 15521 27111 15555
rect 29837 15521 29871 15555
rect 30297 15521 30331 15555
rect 31125 15521 31159 15555
rect 3433 15453 3467 15487
rect 3893 15453 3927 15487
rect 4629 15453 4663 15487
rect 5273 15453 5307 15487
rect 6285 15453 6319 15487
rect 6561 15453 6595 15487
rect 6653 15453 6687 15487
rect 6837 15453 6871 15487
rect 6929 15453 6963 15487
rect 9781 15453 9815 15487
rect 10057 15453 10091 15487
rect 10425 15453 10459 15487
rect 10793 15453 10827 15487
rect 10885 15453 10919 15487
rect 15025 15453 15059 15487
rect 15301 15453 15335 15487
rect 15577 15453 15611 15487
rect 16405 15453 16439 15487
rect 22109 15453 22143 15487
rect 22845 15453 22879 15487
rect 23305 15453 23339 15487
rect 25513 15453 25547 15487
rect 27261 15453 27295 15487
rect 27905 15453 27939 15487
rect 29653 15453 29687 15487
rect 29929 15453 29963 15487
rect 30205 15453 30239 15487
rect 31381 15453 31415 15487
rect 13369 15385 13403 15419
rect 13553 15385 13587 15419
rect 14749 15385 14783 15419
rect 19993 15385 20027 15419
rect 20177 15385 20211 15419
rect 22385 15385 22419 15419
rect 22661 15385 22695 15419
rect 23029 15385 23063 15419
rect 25329 15385 25363 15419
rect 26985 15385 27019 15419
rect 28089 15385 28123 15419
rect 3617 15317 3651 15351
rect 7113 15317 7147 15351
rect 9873 15317 9907 15351
rect 11069 15317 11103 15351
rect 15761 15317 15795 15351
rect 20361 15317 20395 15351
rect 23489 15317 23523 15351
rect 25697 15317 25731 15351
rect 28273 15317 28307 15351
rect 2881 15113 2915 15147
rect 3893 15113 3927 15147
rect 8125 15113 8159 15147
rect 9137 15113 9171 15147
rect 10609 15113 10643 15147
rect 17969 15113 18003 15147
rect 23857 15113 23891 15147
rect 26065 15113 26099 15147
rect 32413 15113 32447 15147
rect 10057 15045 10091 15079
rect 13553 15045 13587 15079
rect 14013 15045 14047 15079
rect 21005 15045 21039 15079
rect 23397 15045 23431 15079
rect 27905 15045 27939 15079
rect 2237 14977 2271 15011
rect 2421 14977 2455 15011
rect 2697 14977 2731 15011
rect 2973 14977 3007 15011
rect 3157 14977 3191 15011
rect 3433 14977 3467 15011
rect 3709 14977 3743 15011
rect 4353 14977 4387 15011
rect 4629 14977 4663 15011
rect 4905 14977 4939 15011
rect 5181 14977 5215 15011
rect 7941 14977 7975 15011
rect 8309 14977 8343 15011
rect 8401 14977 8435 15011
rect 8585 14977 8619 15011
rect 8677 14977 8711 15011
rect 8953 14977 8987 15011
rect 9229 14977 9263 15011
rect 9413 14977 9447 15011
rect 9689 14977 9723 15011
rect 10333 14977 10367 15011
rect 10793 14977 10827 15011
rect 10885 14977 10919 15011
rect 11069 14977 11103 15011
rect 12081 14977 12115 15011
rect 13737 14977 13771 15011
rect 14289 14977 14323 15011
rect 14565 14977 14599 15011
rect 17325 14977 17359 15011
rect 17417 14977 17451 15011
rect 17693 14977 17727 15011
rect 17785 14977 17819 15011
rect 18429 14977 18463 15011
rect 18889 14977 18923 15011
rect 19349 14977 19383 15011
rect 19717 14977 19751 15011
rect 21189 14977 21223 15011
rect 21373 14977 21407 15011
rect 23673 14977 23707 15011
rect 25697 14977 25731 15011
rect 28089 14977 28123 15011
rect 30573 14977 30607 15011
rect 31033 14977 31067 15011
rect 31401 14977 31435 15011
rect 32229 14977 32263 15011
rect 4537 14909 4571 14943
rect 5457 14909 5491 14943
rect 6377 14909 6411 14943
rect 6653 14909 6687 14943
rect 10149 14909 10183 14943
rect 11989 14909 12023 14943
rect 14105 14909 14139 14943
rect 18521 14909 18555 14943
rect 23489 14909 23523 14943
rect 25789 14909 25823 14943
rect 31125 14909 31159 14943
rect 18797 14841 18831 14875
rect 19073 14841 19107 14875
rect 19165 14841 19199 14875
rect 30757 14841 30791 14875
rect 3617 14773 3651 14807
rect 4169 14773 4203 14807
rect 4629 14773 4663 14807
rect 5089 14773 5123 14807
rect 7757 14773 7791 14807
rect 8585 14773 8619 14807
rect 8861 14773 8895 14807
rect 9873 14773 9907 14807
rect 10057 14773 10091 14807
rect 10517 14773 10551 14807
rect 10885 14773 10919 14807
rect 11713 14773 11747 14807
rect 12081 14773 12115 14807
rect 13921 14773 13955 14807
rect 14289 14773 14323 14807
rect 14473 14773 14507 14807
rect 14749 14773 14783 14807
rect 17049 14773 17083 14807
rect 17417 14773 17451 14807
rect 17509 14773 17543 14807
rect 18429 14773 18463 14807
rect 19901 14773 19935 14807
rect 23673 14773 23707 14807
rect 25697 14773 25731 14807
rect 28273 14773 28307 14807
rect 30849 14773 30883 14807
rect 1593 14569 1627 14603
rect 4077 14569 4111 14603
rect 4261 14569 4295 14603
rect 5457 14569 5491 14603
rect 5733 14569 5767 14603
rect 6101 14569 6135 14603
rect 6561 14569 6595 14603
rect 7389 14569 7423 14603
rect 7849 14569 7883 14603
rect 9413 14569 9447 14603
rect 9873 14569 9907 14603
rect 9965 14569 9999 14603
rect 11253 14569 11287 14603
rect 11621 14569 11655 14603
rect 13369 14569 13403 14603
rect 15853 14569 15887 14603
rect 16497 14569 16531 14603
rect 16773 14569 16807 14603
rect 17509 14569 17543 14603
rect 18613 14569 18647 14603
rect 19625 14569 19659 14603
rect 22109 14569 22143 14603
rect 23581 14569 23615 14603
rect 24685 14569 24719 14603
rect 25053 14569 25087 14603
rect 28825 14569 28859 14603
rect 30297 14569 30331 14603
rect 30389 14569 30423 14603
rect 30665 14569 30699 14603
rect 31217 14569 31251 14603
rect 4997 14501 5031 14535
rect 6009 14501 6043 14535
rect 7021 14501 7055 14535
rect 9321 14501 9355 14535
rect 10701 14501 10735 14535
rect 11529 14501 11563 14535
rect 12081 14501 12115 14535
rect 12173 14501 12207 14535
rect 16313 14501 16347 14535
rect 19993 14501 20027 14535
rect 22017 14501 22051 14535
rect 23949 14501 23983 14535
rect 25697 14501 25731 14535
rect 28549 14501 28583 14535
rect 3893 14433 3927 14467
rect 5641 14433 5675 14467
rect 6193 14433 6227 14467
rect 6929 14433 6963 14467
rect 7573 14433 7607 14467
rect 7941 14433 7975 14467
rect 9597 14433 9631 14467
rect 10057 14433 10091 14467
rect 11253 14433 11287 14467
rect 11713 14433 11747 14467
rect 13461 14433 13495 14467
rect 17325 14433 17359 14467
rect 18429 14433 18463 14467
rect 20453 14433 20487 14467
rect 28641 14433 28675 14467
rect 29009 14433 29043 14467
rect 31953 14433 31987 14467
rect 1409 14365 1443 14399
rect 3801 14365 3835 14399
rect 4077 14365 4111 14399
rect 4721 14365 4755 14399
rect 5181 14365 5215 14399
rect 5273 14365 5307 14399
rect 5549 14365 5583 14399
rect 5825 14365 5859 14399
rect 6377 14365 6411 14399
rect 6745 14365 6779 14399
rect 7205 14365 7239 14399
rect 7665 14365 7699 14399
rect 8217 14365 8251 14399
rect 9137 14365 9171 14399
rect 9689 14365 9723 14399
rect 10241 14365 10275 14399
rect 11161 14365 11195 14399
rect 11897 14365 11931 14399
rect 12357 14365 12391 14399
rect 13369 14365 13403 14399
rect 15853 14365 15887 14399
rect 16037 14365 16071 14399
rect 16129 14365 16163 14399
rect 16405 14365 16439 14399
rect 16497 14365 16531 14399
rect 17509 14365 17543 14399
rect 18613 14365 18647 14399
rect 19625 14365 19659 14399
rect 19809 14365 19843 14399
rect 20085 14365 20119 14399
rect 20269 14365 20303 14399
rect 23581 14365 23615 14399
rect 23673 14365 23707 14399
rect 24685 14365 24719 14399
rect 24777 14365 24811 14399
rect 25513 14365 25547 14399
rect 28181 14365 28215 14399
rect 29101 14365 29135 14399
rect 30113 14365 30147 14399
rect 30573 14365 30607 14399
rect 30849 14365 30883 14399
rect 30941 14365 30975 14399
rect 31401 14365 31435 14399
rect 31677 14365 31711 14399
rect 5457 14297 5491 14331
rect 6101 14297 6135 14331
rect 7389 14297 7423 14331
rect 9413 14297 9447 14331
rect 9965 14297 9999 14331
rect 10885 14297 10919 14331
rect 11069 14297 11103 14331
rect 11621 14297 11655 14331
rect 15393 14297 15427 14331
rect 15577 14297 15611 14331
rect 17233 14297 17267 14331
rect 18337 14297 18371 14331
rect 21465 14297 21499 14331
rect 21649 14297 21683 14331
rect 21925 14297 21959 14331
rect 22293 14297 22327 14331
rect 24961 14297 24995 14331
rect 25237 14297 25271 14331
rect 25421 14297 25455 14331
rect 28365 14297 28399 14331
rect 28825 14297 28859 14331
rect 4905 14229 4939 14263
rect 10425 14229 10459 14263
rect 13737 14229 13771 14263
rect 15761 14229 15795 14263
rect 17693 14229 17727 14263
rect 18797 14229 18831 14263
rect 21833 14229 21867 14263
rect 22201 14229 22235 14263
rect 24501 14229 24535 14263
rect 29285 14229 29319 14263
rect 31125 14229 31159 14263
rect 3709 14025 3743 14059
rect 3985 14025 4019 14059
rect 6009 14025 6043 14059
rect 7297 14025 7331 14059
rect 9505 14025 9539 14059
rect 11345 14025 11379 14059
rect 12449 14025 12483 14059
rect 13185 14025 13219 14059
rect 13461 14025 13495 14059
rect 13553 14025 13587 14059
rect 14657 14025 14691 14059
rect 21097 14025 21131 14059
rect 21189 14025 21223 14059
rect 24317 14025 24351 14059
rect 27905 14025 27939 14059
rect 30113 14025 30147 14059
rect 31953 14025 31987 14059
rect 32413 14025 32447 14059
rect 5549 13957 5583 13991
rect 7757 13957 7791 13991
rect 9045 13957 9079 13991
rect 11989 13957 12023 13991
rect 15117 13957 15151 13991
rect 23857 13957 23891 13991
rect 2697 13889 2731 13923
rect 3525 13889 3559 13923
rect 3801 13889 3835 13923
rect 4077 13889 4111 13923
rect 4537 13889 4571 13923
rect 5825 13889 5859 13923
rect 7481 13889 7515 13923
rect 8677 13889 8711 13923
rect 8769 13889 8803 13923
rect 9321 13889 9355 13923
rect 9781 13889 9815 13923
rect 9873 13889 9907 13923
rect 10333 13889 10367 13923
rect 11161 13889 11195 13923
rect 11713 13889 11747 13923
rect 12265 13889 12299 13923
rect 12725 13889 12759 13923
rect 12909 13889 12943 13923
rect 13001 13889 13035 13923
rect 13277 13889 13311 13923
rect 13737 13889 13771 13923
rect 14841 13889 14875 13923
rect 15393 13889 15427 13923
rect 18613 13889 18647 13923
rect 18705 13889 18739 13923
rect 18889 13889 18923 13923
rect 19073 13889 19107 13923
rect 20637 13889 20671 13923
rect 20913 13889 20947 13923
rect 21373 13889 21407 13923
rect 21465 13889 21499 13923
rect 22017 13889 22051 13923
rect 22201 13889 22235 13923
rect 22293 13889 22327 13923
rect 22569 13889 22603 13923
rect 24133 13889 24167 13923
rect 26341 13889 26375 13923
rect 26617 13889 26651 13923
rect 26985 13889 27019 13923
rect 27169 13889 27203 13923
rect 27261 13889 27295 13923
rect 27537 13889 27571 13923
rect 27629 13889 27663 13923
rect 29653 13889 29687 13923
rect 29837 13889 29871 13923
rect 29929 13889 29963 13923
rect 30205 13889 30239 13923
rect 30389 13889 30423 13923
rect 30840 13889 30874 13923
rect 32229 13889 32263 13923
rect 5641 13821 5675 13855
rect 6929 13821 6963 13855
rect 7205 13821 7239 13855
rect 7573 13821 7607 13855
rect 9229 13821 9263 13855
rect 12173 13821 12207 13855
rect 15025 13821 15059 13855
rect 20821 13821 20855 13855
rect 22661 13821 22695 13855
rect 23949 13821 23983 13855
rect 26525 13821 26559 13855
rect 29469 13821 29503 13855
rect 30573 13821 30607 13855
rect 9597 13753 9631 13787
rect 11897 13753 11931 13787
rect 21649 13753 21683 13787
rect 22937 13753 22971 13787
rect 30297 13753 30331 13787
rect 2513 13685 2547 13719
rect 4261 13685 4295 13719
rect 4353 13685 4387 13719
rect 5825 13685 5859 13719
rect 7481 13685 7515 13719
rect 8493 13685 8527 13719
rect 8953 13685 8987 13719
rect 9045 13685 9079 13719
rect 10057 13685 10091 13719
rect 10149 13685 10183 13719
rect 11989 13685 12023 13719
rect 13001 13685 13035 13719
rect 14933 13685 14967 13719
rect 15209 13685 15243 13719
rect 18337 13685 18371 13719
rect 18521 13685 18555 13719
rect 20729 13685 20763 13719
rect 21833 13685 21867 13719
rect 22293 13685 22327 13719
rect 22477 13685 22511 13719
rect 22569 13685 22603 13719
rect 24133 13685 24167 13719
rect 26341 13685 26375 13719
rect 26801 13685 26835 13719
rect 27169 13685 27203 13719
rect 27445 13685 27479 13719
rect 27721 13685 27755 13719
rect 29929 13685 29963 13719
rect 2329 13481 2363 13515
rect 3617 13481 3651 13515
rect 8125 13481 8159 13515
rect 9597 13481 9631 13515
rect 11253 13481 11287 13515
rect 13277 13481 13311 13515
rect 14473 13481 14507 13515
rect 18153 13481 18187 13515
rect 18337 13481 18371 13515
rect 20453 13481 20487 13515
rect 21005 13481 21039 13515
rect 28273 13481 28307 13515
rect 28733 13481 28767 13515
rect 29285 13481 29319 13515
rect 31493 13481 31527 13515
rect 7278 13413 7312 13447
rect 7389 13413 7423 13447
rect 12725 13413 12759 13447
rect 20913 13413 20947 13447
rect 26433 13413 26467 13447
rect 28457 13413 28491 13447
rect 28825 13413 28859 13447
rect 6193 13345 6227 13379
rect 7481 13345 7515 13379
rect 13093 13345 13127 13379
rect 17969 13345 18003 13379
rect 20545 13345 20579 13379
rect 26157 13345 26191 13379
rect 32229 13345 32263 13379
rect 2513 13277 2547 13311
rect 3433 13277 3467 13311
rect 3801 13277 3835 13311
rect 3985 13277 4019 13311
rect 4169 13277 4203 13311
rect 4629 13277 4663 13311
rect 5825 13277 5859 13311
rect 6101 13277 6135 13311
rect 6469 13277 6503 13311
rect 9045 13277 9079 13311
rect 9321 13277 9355 13311
rect 9413 13277 9447 13311
rect 11437 13277 11471 13311
rect 12909 13277 12943 13311
rect 13277 13277 13311 13311
rect 14289 13277 14323 13311
rect 15117 13277 15151 13311
rect 15301 13277 15335 13311
rect 18153 13277 18187 13311
rect 20177 13277 20211 13311
rect 20729 13277 20763 13311
rect 21005 13277 21039 13311
rect 21189 13277 21223 13311
rect 24409 13277 24443 13311
rect 26249 13277 26283 13311
rect 26433 13277 26467 13311
rect 27813 13277 27847 13311
rect 27905 13277 27939 13311
rect 28273 13277 28307 13311
rect 28549 13277 28583 13311
rect 28917 13277 28951 13311
rect 29009 13277 29043 13311
rect 30941 13277 30975 13311
rect 31217 13277 31251 13311
rect 31309 13277 31343 13311
rect 31677 13277 31711 13311
rect 2697 13209 2731 13243
rect 4077 13209 4111 13243
rect 7113 13209 7147 13243
rect 7849 13209 7883 13243
rect 8033 13209 8067 13243
rect 9229 13209 9263 13243
rect 13001 13209 13035 13243
rect 14105 13209 14139 13243
rect 15485 13209 15519 13243
rect 17877 13209 17911 13243
rect 20453 13209 20487 13243
rect 31125 13209 31159 13243
rect 4353 13141 4387 13175
rect 4445 13141 4479 13175
rect 13461 13141 13495 13175
rect 20361 13141 20395 13175
rect 21373 13141 21407 13175
rect 27629 13141 27663 13175
rect 6377 12937 6411 12971
rect 15393 12937 15427 12971
rect 23857 12937 23891 12971
rect 27629 12937 27663 12971
rect 30389 12937 30423 12971
rect 3525 12869 3559 12903
rect 4629 12869 4663 12903
rect 8677 12869 8711 12903
rect 11529 12869 11563 12903
rect 14933 12869 14967 12903
rect 15669 12869 15703 12903
rect 16773 12869 16807 12903
rect 19901 12869 19935 12903
rect 20269 12869 20303 12903
rect 24225 12869 24259 12903
rect 25789 12869 25823 12903
rect 28181 12869 28215 12903
rect 3249 12801 3283 12835
rect 3341 12801 3375 12835
rect 3617 12801 3651 12835
rect 3801 12801 3835 12835
rect 3985 12801 4019 12835
rect 4813 12801 4847 12835
rect 4997 12801 5031 12835
rect 5273 12801 5307 12835
rect 5549 12801 5583 12835
rect 5917 12801 5951 12835
rect 6101 12801 6135 12835
rect 6561 12801 6595 12835
rect 6837 12801 6871 12835
rect 7389 12801 7423 12835
rect 8401 12801 8435 12835
rect 8861 12801 8895 12835
rect 8953 12801 8987 12835
rect 9505 12801 9539 12835
rect 9781 12801 9815 12835
rect 11052 12801 11086 12835
rect 11345 12801 11379 12835
rect 11805 12801 11839 12835
rect 12357 12801 12391 12835
rect 15209 12801 15243 12835
rect 15485 12801 15519 12835
rect 15945 12801 15979 12835
rect 16221 12801 16255 12835
rect 17049 12801 17083 12835
rect 17325 12801 17359 12835
rect 18613 12801 18647 12835
rect 18705 12801 18739 12835
rect 20085 12801 20119 12835
rect 22017 12801 22051 12835
rect 22201 12801 22235 12835
rect 23397 12801 23431 12835
rect 24041 12801 24075 12835
rect 24317 12801 24351 12835
rect 24777 12801 24811 12835
rect 24869 12801 24903 12835
rect 26065 12801 26099 12835
rect 27169 12801 27203 12835
rect 27445 12801 27479 12835
rect 28457 12801 28491 12835
rect 30297 12801 30331 12835
rect 31697 12801 31731 12835
rect 31953 12801 31987 12835
rect 32505 12801 32539 12835
rect 6653 12733 6687 12767
rect 7113 12733 7147 12767
rect 11253 12733 11287 12767
rect 11713 12733 11747 12767
rect 15025 12733 15059 12767
rect 15853 12733 15887 12767
rect 16129 12733 16163 12767
rect 16865 12733 16899 12767
rect 23489 12733 23523 12767
rect 25881 12733 25915 12767
rect 27261 12733 27295 12767
rect 28273 12733 28307 12767
rect 3065 12665 3099 12699
rect 5089 12665 5123 12699
rect 5733 12665 5767 12699
rect 8585 12665 8619 12699
rect 11989 12665 12023 12699
rect 17509 12665 17543 12699
rect 24501 12665 24535 12699
rect 26249 12665 26283 12699
rect 30573 12665 30607 12699
rect 32321 12665 32355 12699
rect 3525 12597 3559 12631
rect 5365 12597 5399 12631
rect 6745 12597 6779 12631
rect 8953 12597 8987 12631
rect 9137 12597 9171 12631
rect 9321 12597 9355 12631
rect 9597 12597 9631 12631
rect 10885 12597 10919 12631
rect 11161 12597 11195 12631
rect 11529 12597 11563 12631
rect 12173 12597 12207 12631
rect 15117 12597 15151 12631
rect 16221 12597 16255 12631
rect 16405 12597 16439 12631
rect 16865 12597 16899 12631
rect 17233 12597 17267 12631
rect 18613 12597 18647 12631
rect 18981 12597 19015 12631
rect 22109 12597 22143 12631
rect 22385 12597 22419 12631
rect 23489 12597 23523 12631
rect 23765 12597 23799 12631
rect 24593 12597 24627 12631
rect 25053 12597 25087 12631
rect 25789 12597 25823 12631
rect 27169 12597 27203 12631
rect 28457 12597 28491 12631
rect 28641 12597 28675 12631
rect 3065 12393 3099 12427
rect 3157 12393 3191 12427
rect 6101 12393 6135 12427
rect 9413 12393 9447 12427
rect 11345 12393 11379 12427
rect 11897 12393 11931 12427
rect 16405 12393 16439 12427
rect 16773 12393 16807 12427
rect 21925 12393 21959 12427
rect 22661 12393 22695 12427
rect 23673 12393 23707 12427
rect 24409 12393 24443 12427
rect 24961 12393 24995 12427
rect 25421 12393 25455 12427
rect 25605 12393 25639 12427
rect 25973 12393 26007 12427
rect 26893 12393 26927 12427
rect 27077 12393 27111 12427
rect 27997 12393 28031 12427
rect 30113 12393 30147 12427
rect 5273 12325 5307 12359
rect 17233 12325 17267 12359
rect 24869 12325 24903 12359
rect 11713 12257 11747 12291
rect 16865 12257 16899 12291
rect 21925 12257 21959 12291
rect 22477 12257 22511 12291
rect 24501 12257 24535 12291
rect 25053 12257 25087 12291
rect 27813 12257 27847 12291
rect 29929 12257 29963 12291
rect 30205 12257 30239 12291
rect 2421 12189 2455 12223
rect 2513 12189 2547 12223
rect 2881 12189 2915 12223
rect 3341 12189 3375 12223
rect 3617 12189 3651 12223
rect 4721 12189 4755 12223
rect 4997 12189 5031 12223
rect 5113 12189 5147 12223
rect 5365 12189 5399 12223
rect 5549 12189 5583 12223
rect 5825 12189 5859 12223
rect 6285 12189 6319 12223
rect 6745 12189 6779 12223
rect 6929 12189 6963 12223
rect 7205 12189 7239 12223
rect 8033 12189 8067 12223
rect 9144 12189 9178 12223
rect 9321 12189 9355 12223
rect 9413 12189 9447 12223
rect 11161 12189 11195 12223
rect 11897 12189 11931 12223
rect 16221 12189 16255 12223
rect 17049 12189 17083 12223
rect 17969 12189 18003 12223
rect 18245 12189 18279 12223
rect 19257 12189 19291 12223
rect 22109 12189 22143 12223
rect 22661 12189 22695 12223
rect 23857 12189 23891 12223
rect 24041 12189 24075 12223
rect 24685 12189 24719 12223
rect 25237 12189 25271 12223
rect 25697 12189 25731 12223
rect 25789 12189 25823 12223
rect 26709 12189 26743 12223
rect 26801 12189 26835 12223
rect 27997 12189 28031 12223
rect 30113 12189 30147 12223
rect 30941 12189 30975 12223
rect 31309 12189 31343 12223
rect 31677 12189 31711 12223
rect 32229 12189 32263 12223
rect 2697 12121 2731 12155
rect 2789 12121 2823 12155
rect 4905 12121 4939 12155
rect 6009 12121 6043 12155
rect 6561 12121 6595 12155
rect 7849 12121 7883 12155
rect 11621 12121 11655 12155
rect 16773 12121 16807 12155
rect 19441 12121 19475 12155
rect 19625 12121 19659 12155
rect 21833 12121 21867 12155
rect 22385 12121 22419 12155
rect 24409 12121 24443 12155
rect 24961 12121 24995 12155
rect 25513 12121 25547 12155
rect 27721 12121 27755 12155
rect 31125 12121 31159 12155
rect 31217 12121 31251 12155
rect 2237 12053 2271 12087
rect 3433 12053 3467 12087
rect 8217 12053 8251 12087
rect 9597 12053 9631 12087
rect 12081 12053 12115 12087
rect 22293 12053 22327 12087
rect 22845 12053 22879 12087
rect 28181 12053 28215 12087
rect 30481 12053 30515 12087
rect 31493 12053 31527 12087
rect 3249 11849 3283 11883
rect 4261 11849 4295 11883
rect 7021 11849 7055 11883
rect 7481 11849 7515 11883
rect 9229 11849 9263 11883
rect 10885 11849 10919 11883
rect 11161 11849 11195 11883
rect 17141 11849 17175 11883
rect 17509 11849 17543 11883
rect 17969 11849 18003 11883
rect 19073 11849 19107 11883
rect 20729 11849 20763 11883
rect 21005 11849 21039 11883
rect 31953 11849 31987 11883
rect 6929 11781 6963 11815
rect 8217 11781 8251 11815
rect 14749 11781 14783 11815
rect 15209 11781 15243 11815
rect 18153 11781 18187 11815
rect 19901 11781 19935 11815
rect 24133 11781 24167 11815
rect 29561 11781 29595 11815
rect 30840 11781 30874 11815
rect 2789 11713 2823 11747
rect 3065 11713 3099 11747
rect 3525 11713 3559 11747
rect 3801 11713 3835 11747
rect 4169 11713 4203 11747
rect 4445 11713 4479 11747
rect 4629 11713 4663 11747
rect 5181 11713 5215 11747
rect 5457 11713 5491 11747
rect 6169 11713 6203 11747
rect 6561 11713 6595 11747
rect 7297 11713 7331 11747
rect 8769 11713 8803 11747
rect 9045 11713 9079 11747
rect 10609 11713 10643 11747
rect 10701 11713 10735 11747
rect 10977 11713 11011 11747
rect 11529 11713 11563 11747
rect 11805 11713 11839 11747
rect 12173 11713 12207 11747
rect 12357 11713 12391 11747
rect 12909 11713 12943 11747
rect 13185 11713 13219 11747
rect 14473 11713 14507 11747
rect 14841 11713 14875 11747
rect 15025 11713 15059 11747
rect 16681 11713 16715 11747
rect 16957 11713 16991 11747
rect 17693 11713 17727 11747
rect 18429 11713 18463 11747
rect 18705 11713 18739 11747
rect 19717 11713 19751 11747
rect 20361 11713 20395 11747
rect 20545 11713 20579 11747
rect 20821 11713 20855 11747
rect 23949 11713 23983 11747
rect 28457 11713 28491 11747
rect 28641 11713 28675 11747
rect 28733 11713 28767 11747
rect 29837 11713 29871 11747
rect 32229 11713 32263 11747
rect 8953 11645 8987 11679
rect 11621 11645 11655 11679
rect 13001 11645 13035 11679
rect 14657 11645 14691 11679
rect 16865 11645 16899 11679
rect 18245 11645 18279 11679
rect 18797 11645 18831 11679
rect 29653 11645 29687 11679
rect 30573 11645 30607 11679
rect 3617 11577 3651 11611
rect 4813 11577 4847 11611
rect 8493 11577 8527 11611
rect 12541 11577 12575 11611
rect 32413 11577 32447 11611
rect 2973 11509 3007 11543
rect 3341 11509 3375 11543
rect 3985 11509 4019 11543
rect 4997 11509 5031 11543
rect 5273 11509 5307 11543
rect 6009 11509 6043 11543
rect 6745 11509 6779 11543
rect 8677 11509 8711 11543
rect 9045 11509 9079 11543
rect 10425 11509 10459 11543
rect 11529 11509 11563 11543
rect 11989 11509 12023 11543
rect 12173 11509 12207 11543
rect 12909 11509 12943 11543
rect 13369 11509 13403 11543
rect 14289 11509 14323 11543
rect 14749 11509 14783 11543
rect 16773 11509 16807 11543
rect 18153 11509 18187 11543
rect 18613 11509 18647 11543
rect 18705 11509 18739 11543
rect 20085 11509 20119 11543
rect 23765 11509 23799 11543
rect 28457 11509 28491 11543
rect 28917 11509 28951 11543
rect 29837 11509 29871 11543
rect 30021 11509 30055 11543
rect 1593 11305 1627 11339
rect 4721 11305 4755 11339
rect 7665 11305 7699 11339
rect 10517 11305 10551 11339
rect 10885 11305 10919 11339
rect 11069 11305 11103 11339
rect 11897 11305 11931 11339
rect 14473 11305 14507 11339
rect 14933 11305 14967 11339
rect 15301 11305 15335 11339
rect 16037 11305 16071 11339
rect 20453 11305 20487 11339
rect 21005 11305 21039 11339
rect 21189 11305 21223 11339
rect 22201 11305 22235 11339
rect 23857 11305 23891 11339
rect 25697 11305 25731 11339
rect 26249 11305 26283 11339
rect 26801 11305 26835 11339
rect 28089 11305 28123 11339
rect 32229 11305 32263 11339
rect 3157 11237 3191 11271
rect 4077 11237 4111 11271
rect 7113 11237 7147 11271
rect 7941 11237 7975 11271
rect 10057 11237 10091 11271
rect 16313 11237 16347 11271
rect 20913 11237 20947 11271
rect 22385 11237 22419 11271
rect 26065 11237 26099 11271
rect 26709 11237 26743 11271
rect 27169 11237 27203 11271
rect 30757 11237 30791 11271
rect 7573 11169 7607 11203
rect 10333 11169 10367 11203
rect 10701 11169 10735 11203
rect 14565 11169 14599 11203
rect 20545 11169 20579 11203
rect 23673 11169 23707 11203
rect 26433 11169 26467 11203
rect 1409 11101 1443 11135
rect 1961 11101 1995 11135
rect 2145 11101 2179 11135
rect 2237 11101 2271 11135
rect 2329 11101 2363 11135
rect 2605 11101 2639 11135
rect 2881 11101 2915 11135
rect 2973 11101 3007 11135
rect 3433 11101 3467 11135
rect 3893 11101 3927 11135
rect 4169 11101 4203 11135
rect 4537 11101 4571 11135
rect 4997 11101 5031 11135
rect 5089 11101 5123 11135
rect 5365 11101 5399 11135
rect 5457 11101 5491 11135
rect 5917 11101 5951 11135
rect 6377 11101 6411 11135
rect 6561 11101 6595 11135
rect 6837 11101 6871 11135
rect 6929 11101 6963 11135
rect 7205 11101 7239 11135
rect 7757 11101 7791 11135
rect 8309 11101 8343 11135
rect 8585 11101 8619 11135
rect 10241 11101 10275 11135
rect 10517 11101 10551 11135
rect 10609 11101 10643 11135
rect 10885 11101 10919 11135
rect 14473 11101 14507 11135
rect 14749 11101 14783 11135
rect 15301 11101 15335 11135
rect 15485 11101 15519 11135
rect 16221 11101 16255 11135
rect 16497 11101 16531 11135
rect 17233 11101 17267 11135
rect 17417 11101 17451 11135
rect 20729 11101 20763 11135
rect 21281 11101 21315 11135
rect 21373 11101 21407 11135
rect 22017 11101 22051 11135
rect 22201 11101 22235 11135
rect 22661 11101 22695 11135
rect 23581 11101 23615 11135
rect 23857 11101 23891 11135
rect 25697 11101 25731 11135
rect 25789 11101 25823 11135
rect 26249 11101 26283 11135
rect 26525 11101 26559 11135
rect 26801 11101 26835 11135
rect 26893 11101 26927 11135
rect 30205 11101 30239 11135
rect 30389 11101 30423 11135
rect 30573 11101 30607 11135
rect 30849 11101 30883 11135
rect 31105 11101 31139 11135
rect 2789 11033 2823 11067
rect 4353 11033 4387 11067
rect 4445 11033 4479 11067
rect 5273 11033 5307 11067
rect 6745 11033 6779 11067
rect 7481 11033 7515 11067
rect 8125 11033 8159 11067
rect 11805 11033 11839 11067
rect 17601 11033 17635 11067
rect 20453 11033 20487 11067
rect 27721 11033 27755 11067
rect 27905 11033 27939 11067
rect 30481 11033 30515 11067
rect 2513 10965 2547 10999
rect 3617 10965 3651 10999
rect 4813 10965 4847 10999
rect 5641 10965 5675 10999
rect 6101 10965 6135 10999
rect 6285 10965 6319 10999
rect 7389 10965 7423 10999
rect 8401 10965 8435 10999
rect 15669 10965 15703 10999
rect 22477 10965 22511 10999
rect 24041 10965 24075 10999
rect 4721 10761 4755 10795
rect 6929 10761 6963 10795
rect 7481 10761 7515 10795
rect 11897 10761 11931 10795
rect 13093 10761 13127 10795
rect 18061 10761 18095 10795
rect 19441 10761 19475 10795
rect 20637 10761 20671 10795
rect 22201 10761 22235 10795
rect 22845 10761 22879 10795
rect 24409 10761 24443 10795
rect 25145 10761 25179 10795
rect 25973 10761 26007 10795
rect 27537 10761 27571 10795
rect 27997 10761 28031 10795
rect 28457 10761 28491 10795
rect 31309 10761 31343 10795
rect 4261 10693 4295 10727
rect 6561 10693 6595 10727
rect 7021 10693 7055 10727
rect 7573 10693 7607 10727
rect 9229 10693 9263 10727
rect 9413 10693 9447 10727
rect 12633 10693 12667 10727
rect 15853 10693 15887 10727
rect 18981 10693 19015 10727
rect 19986 10693 20020 10727
rect 21097 10693 21131 10727
rect 23949 10693 23983 10727
rect 24685 10693 24719 10727
rect 25513 10693 25547 10727
rect 4077 10625 4111 10659
rect 4353 10625 4387 10659
rect 4445 10625 4479 10659
rect 4905 10625 4939 10659
rect 4997 10625 5031 10659
rect 5457 10625 5491 10659
rect 5891 10629 5925 10663
rect 6009 10629 6043 10663
rect 6377 10625 6411 10659
rect 6653 10625 6687 10659
rect 6769 10625 6803 10659
rect 7297 10625 7331 10659
rect 7757 10625 7791 10659
rect 9689 10625 9723 10659
rect 11529 10625 11563 10659
rect 11713 10625 11747 10659
rect 11989 10625 12023 10659
rect 12909 10625 12943 10659
rect 14289 10625 14323 10659
rect 14565 10625 14599 10659
rect 16129 10625 16163 10659
rect 16957 10625 16991 10659
rect 17141 10625 17175 10659
rect 17601 10625 17635 10659
rect 17693 10625 17727 10659
rect 19257 10625 19291 10659
rect 19717 10625 19751 10659
rect 20085 10625 20119 10659
rect 20545 10625 20579 10659
rect 20821 10625 20855 10659
rect 21281 10625 21315 10659
rect 21465 10625 21499 10659
rect 21833 10625 21867 10659
rect 22017 10625 22051 10659
rect 22385 10625 22419 10659
rect 22661 10625 22695 10659
rect 22937 10625 22971 10659
rect 23489 10625 23523 10659
rect 24133 10625 24167 10659
rect 24225 10625 24259 10659
rect 24961 10625 24995 10659
rect 25789 10625 25823 10659
rect 26065 10625 26099 10659
rect 27077 10625 27111 10659
rect 27353 10625 27387 10659
rect 27629 10625 27663 10659
rect 27813 10625 27847 10659
rect 28089 10625 28123 10659
rect 28273 10625 28307 10659
rect 30389 10625 30423 10659
rect 30481 10625 30515 10659
rect 30941 10625 30975 10659
rect 31033 10625 31067 10659
rect 32229 10625 32263 10659
rect 7113 10557 7147 10591
rect 9045 10557 9079 10591
rect 12725 10557 12759 10591
rect 14381 10557 14415 10591
rect 16037 10557 16071 10591
rect 17785 10557 17819 10591
rect 19073 10557 19107 10591
rect 19901 10557 19935 10591
rect 20913 10557 20947 10591
rect 22477 10557 22511 10591
rect 23029 10557 23063 10591
rect 23581 10557 23615 10591
rect 24777 10557 24811 10591
rect 25605 10557 25639 10591
rect 26157 10557 26191 10591
rect 27169 10557 27203 10591
rect 31953 10557 31987 10591
rect 4629 10489 4663 10523
rect 5273 10489 5307 10523
rect 14749 10489 14783 10523
rect 17325 10489 17359 10523
rect 21649 10489 21683 10523
rect 23305 10489 23339 10523
rect 23857 10489 23891 10523
rect 26433 10489 26467 10523
rect 30757 10489 30791 10523
rect 5181 10421 5215 10455
rect 5733 10421 5767 10455
rect 6193 10421 6227 10455
rect 7297 10421 7331 10455
rect 7941 10421 7975 10455
rect 9505 10421 9539 10455
rect 12173 10421 12207 10455
rect 12909 10421 12943 10455
rect 14289 10421 14323 10455
rect 15853 10421 15887 10455
rect 16313 10421 16347 10455
rect 16773 10421 16807 10455
rect 17417 10421 17451 10455
rect 17785 10421 17819 10455
rect 19257 10421 19291 10455
rect 19533 10421 19567 10455
rect 19901 10421 19935 10455
rect 20269 10421 20303 10455
rect 20361 10421 20395 10455
rect 21097 10421 21131 10455
rect 21281 10421 21315 10455
rect 22661 10421 22695 10455
rect 22937 10421 22971 10455
rect 23489 10421 23523 10455
rect 23949 10421 23983 10455
rect 24961 10421 24995 10455
rect 25605 10421 25639 10455
rect 26249 10421 26283 10455
rect 27077 10421 27111 10455
rect 30205 10421 30239 10455
rect 30665 10421 30699 10455
rect 31217 10421 31251 10455
rect 32413 10421 32447 10455
rect 6009 10217 6043 10251
rect 9137 10217 9171 10251
rect 9597 10217 9631 10251
rect 9689 10217 9723 10251
rect 10793 10217 10827 10251
rect 15577 10217 15611 10251
rect 16037 10217 16071 10251
rect 16957 10217 16991 10251
rect 17417 10217 17451 10251
rect 19993 10217 20027 10251
rect 22477 10217 22511 10251
rect 24685 10217 24719 10251
rect 27721 10217 27755 10251
rect 29653 10217 29687 10251
rect 3617 10149 3651 10183
rect 4353 10149 4387 10183
rect 6469 10149 6503 10183
rect 7113 10149 7147 10183
rect 15761 10149 15795 10183
rect 22109 10149 22143 10183
rect 10885 10081 10919 10115
rect 15393 10081 15427 10115
rect 17141 10081 17175 10115
rect 19625 10081 19659 10115
rect 24501 10081 24535 10115
rect 27721 10081 27755 10115
rect 29653 10081 29687 10115
rect 31861 10081 31895 10115
rect 3433 10013 3467 10047
rect 3801 10013 3835 10047
rect 4077 10013 4111 10047
rect 4169 10013 4203 10047
rect 5365 10013 5399 10047
rect 5917 10013 5951 10047
rect 6193 10013 6227 10047
rect 6285 10013 6319 10047
rect 6929 10013 6963 10047
rect 7757 10013 7791 10047
rect 9321 10013 9355 10047
rect 9413 10013 9447 10047
rect 9873 10013 9907 10047
rect 10793 10013 10827 10047
rect 11069 10013 11103 10047
rect 15577 10013 15611 10047
rect 15853 10013 15887 10047
rect 16405 10013 16439 10047
rect 16865 10013 16899 10047
rect 17233 10013 17267 10047
rect 18521 10013 18555 10047
rect 19257 10013 19291 10047
rect 19814 10007 19848 10041
rect 19993 10013 20027 10047
rect 22293 10013 22327 10047
rect 22385 10013 22419 10047
rect 22569 10013 22603 10047
rect 24409 10013 24443 10047
rect 24685 10013 24719 10047
rect 27537 10013 27571 10047
rect 29561 10013 29595 10047
rect 29837 10013 29871 10047
rect 30205 10013 30239 10047
rect 30573 10013 30607 10047
rect 31493 10013 31527 10047
rect 31585 10013 31619 10047
rect 32505 10013 32539 10047
rect 3985 9945 4019 9979
rect 9597 9945 9631 9979
rect 15301 9945 15335 9979
rect 16957 9945 16991 9979
rect 19441 9945 19475 9979
rect 27169 9945 27203 9979
rect 27813 9945 27847 9979
rect 30389 9945 30423 9979
rect 30481 9945 30515 9979
rect 30849 9945 30883 9979
rect 5549 9877 5583 9911
rect 5733 9877 5767 9911
rect 7573 9877 7607 9911
rect 11253 9877 11287 9911
rect 16589 9877 16623 9911
rect 16681 9877 16715 9911
rect 18337 9877 18371 9911
rect 20177 9877 20211 9911
rect 24869 9877 24903 9911
rect 27353 9877 27387 9911
rect 30021 9877 30055 9911
rect 30757 9877 30791 9911
rect 31769 9877 31803 9911
rect 4537 9673 4571 9707
rect 6837 9673 6871 9707
rect 8769 9673 8803 9707
rect 10701 9673 10735 9707
rect 11069 9673 11103 9707
rect 12449 9673 12483 9707
rect 16497 9673 16531 9707
rect 18613 9673 18647 9707
rect 20085 9673 20119 9707
rect 31585 9673 31619 9707
rect 3617 9605 3651 9639
rect 4261 9605 4295 9639
rect 5549 9605 5583 9639
rect 5641 9605 5675 9639
rect 7205 9605 7239 9639
rect 8493 9605 8527 9639
rect 25237 9605 25271 9639
rect 29745 9605 29779 9639
rect 29837 9605 29871 9639
rect 3065 9537 3099 9571
rect 3341 9537 3375 9571
rect 3525 9537 3559 9571
rect 3709 9537 3743 9571
rect 3985 9537 4019 9571
rect 4169 9537 4203 9571
rect 4353 9537 4387 9571
rect 5273 9537 5307 9571
rect 5365 9537 5399 9571
rect 5733 9537 5767 9571
rect 6001 9541 6035 9575
rect 6377 9537 6411 9571
rect 6653 9537 6687 9571
rect 6929 9537 6963 9571
rect 7113 9537 7147 9571
rect 7297 9537 7331 9571
rect 7573 9537 7607 9571
rect 7757 9537 7791 9571
rect 7849 9537 7883 9571
rect 7941 9537 7975 9571
rect 8217 9537 8251 9571
rect 8401 9537 8435 9571
rect 8585 9537 8619 9571
rect 10057 9537 10091 9571
rect 10149 9537 10183 9571
rect 10333 9537 10367 9571
rect 10425 9537 10459 9571
rect 10517 9537 10551 9571
rect 10977 9537 11011 9571
rect 11253 9537 11287 9571
rect 11989 9537 12023 9571
rect 12265 9537 12299 9571
rect 12817 9537 12851 9571
rect 13093 9537 13127 9571
rect 13369 9537 13403 9571
rect 13553 9537 13587 9571
rect 13829 9537 13863 9571
rect 14013 9537 14047 9571
rect 16037 9537 16071 9571
rect 16313 9537 16347 9571
rect 17785 9537 17819 9571
rect 17969 9537 18003 9571
rect 18245 9537 18279 9571
rect 18429 9537 18463 9571
rect 19441 9537 19475 9571
rect 19901 9537 19935 9571
rect 20913 9537 20947 9571
rect 21097 9537 21131 9571
rect 21465 9537 21499 9571
rect 21925 9537 21959 9571
rect 22201 9537 22235 9571
rect 23029 9537 23063 9571
rect 24961 9537 24995 9571
rect 26341 9537 26375 9571
rect 29561 9537 29595 9571
rect 29929 9537 29963 9571
rect 30461 9537 30495 9571
rect 31953 9537 31987 9571
rect 32505 9537 32539 9571
rect 8953 9469 8987 9503
rect 9229 9469 9263 9503
rect 13001 9469 13035 9503
rect 16129 9469 16163 9503
rect 19533 9469 19567 9503
rect 21281 9469 21315 9503
rect 22109 9469 22143 9503
rect 22937 9469 22971 9503
rect 25053 9469 25087 9503
rect 30205 9469 30239 9503
rect 3249 9401 3283 9435
rect 5089 9401 5123 9435
rect 8125 9401 8159 9435
rect 10793 9401 10827 9435
rect 12173 9401 12207 9435
rect 13277 9401 13311 9435
rect 19809 9401 19843 9435
rect 22661 9401 22695 9435
rect 24777 9401 24811 9435
rect 30113 9401 30147 9435
rect 32321 9401 32355 9435
rect 3893 9333 3927 9367
rect 5917 9333 5951 9367
rect 6193 9333 6227 9367
rect 6561 9333 6595 9367
rect 7481 9333 7515 9367
rect 9873 9333 9907 9367
rect 13001 9333 13035 9367
rect 13553 9333 13587 9367
rect 14197 9333 14231 9367
rect 16313 9333 16347 9367
rect 18153 9333 18187 9367
rect 19441 9333 19475 9367
rect 21649 9333 21683 9367
rect 22201 9333 22235 9367
rect 22385 9333 22419 9367
rect 22569 9333 22603 9367
rect 22845 9333 22879 9367
rect 24593 9333 24627 9367
rect 25237 9333 25271 9367
rect 26525 9333 26559 9367
rect 31769 9333 31803 9367
rect 3617 9129 3651 9163
rect 5549 9129 5583 9163
rect 6837 9129 6871 9163
rect 8953 9129 8987 9163
rect 9137 9129 9171 9163
rect 12541 9129 12575 9163
rect 12725 9129 12759 9163
rect 14565 9129 14599 9163
rect 17417 9129 17451 9163
rect 18613 9129 18647 9163
rect 21925 9129 21959 9163
rect 22109 9129 22143 9163
rect 25605 9129 25639 9163
rect 25973 9129 26007 9163
rect 26157 9129 26191 9163
rect 26617 9129 26651 9163
rect 26985 9129 27019 9163
rect 27721 9129 27755 9163
rect 28089 9129 28123 9163
rect 29285 9129 29319 9163
rect 32505 9129 32539 9163
rect 4905 9061 4939 9095
rect 6193 9061 6227 9095
rect 14749 9061 14783 9095
rect 11621 8993 11655 9027
rect 12357 8993 12391 9027
rect 18521 8993 18555 9027
rect 26341 8993 26375 9027
rect 27721 8993 27755 9027
rect 3433 8925 3467 8959
rect 3985 8925 4019 8959
rect 4077 8925 4111 8959
rect 4445 8925 4479 8959
rect 4721 8925 4755 8959
rect 4997 8925 5031 8959
rect 5365 8925 5399 8959
rect 5641 8925 5675 8959
rect 6009 8925 6043 8959
rect 6285 8925 6319 8959
rect 6469 8925 6503 8959
rect 6561 8925 6595 8959
rect 6653 8925 6687 8959
rect 7297 8925 7331 8959
rect 7573 8925 7607 8959
rect 8033 8925 8067 8959
rect 9137 8925 9171 8959
rect 9229 8925 9263 8959
rect 11345 8925 11379 8959
rect 12541 8925 12575 8959
rect 14105 8925 14139 8959
rect 14381 8925 14415 8959
rect 14565 8925 14599 8959
rect 17141 8925 17175 8959
rect 17601 8925 17635 8959
rect 18429 8925 18463 8959
rect 18705 8925 18739 8959
rect 22109 8925 22143 8959
rect 22201 8925 22235 8959
rect 22396 8925 22430 8959
rect 25513 8925 25547 8959
rect 25697 8925 25731 8959
rect 25789 8925 25823 8959
rect 26426 8925 26460 8959
rect 26893 8925 26927 8959
rect 26985 8925 27019 8959
rect 27905 8925 27939 8959
rect 28365 8925 28399 8959
rect 29101 8925 29135 8959
rect 31125 8925 31159 8959
rect 4261 8857 4295 8891
rect 4353 8857 4387 8891
rect 5181 8857 5215 8891
rect 5273 8857 5307 8891
rect 5825 8857 5859 8891
rect 5917 8857 5951 8891
rect 9413 8857 9447 8891
rect 12265 8857 12299 8891
rect 17785 8857 17819 8891
rect 26157 8857 26191 8891
rect 26709 8857 26743 8891
rect 27629 8857 27663 8891
rect 28917 8857 28951 8891
rect 31370 8857 31404 8891
rect 3801 8789 3835 8823
rect 4629 8789 4663 8823
rect 7481 8789 7515 8823
rect 7757 8789 7791 8823
rect 7849 8789 7883 8823
rect 16957 8789 16991 8823
rect 17325 8789 17359 8823
rect 18889 8789 18923 8823
rect 25329 8789 25363 8823
rect 27169 8789 27203 8823
rect 28181 8789 28215 8823
rect 4077 8585 4111 8619
rect 4629 8585 4663 8619
rect 9413 8585 9447 8619
rect 11345 8585 11379 8619
rect 11897 8585 11931 8619
rect 12541 8585 12575 8619
rect 14013 8585 14047 8619
rect 15485 8585 15519 8619
rect 16865 8585 16899 8619
rect 17325 8585 17359 8619
rect 20085 8585 20119 8619
rect 20729 8585 20763 8619
rect 24685 8585 24719 8619
rect 5457 8517 5491 8551
rect 7389 8517 7423 8551
rect 9689 8517 9723 8551
rect 10425 8517 10459 8551
rect 10977 8517 11011 8551
rect 11069 8517 11103 8551
rect 12081 8517 12115 8551
rect 14933 8517 14967 8551
rect 23489 8517 23523 8551
rect 24225 8517 24259 8551
rect 30849 8517 30883 8551
rect 30941 8517 30975 8551
rect 4261 8449 4295 8483
rect 4445 8449 4479 8483
rect 5273 8449 5307 8483
rect 5549 8449 5583 8483
rect 5641 8449 5675 8483
rect 5917 8449 5951 8483
rect 7205 8449 7239 8483
rect 7481 8449 7515 8483
rect 7573 8449 7607 8483
rect 8033 8449 8067 8483
rect 8309 8449 8343 8483
rect 8585 8449 8619 8483
rect 8769 8449 8803 8483
rect 8861 8449 8895 8483
rect 8953 8449 8987 8483
rect 9229 8449 9263 8483
rect 9505 8449 9539 8483
rect 9781 8449 9815 8483
rect 9873 8449 9907 8483
rect 10195 8449 10229 8483
rect 10333 8449 10367 8483
rect 10517 8449 10551 8483
rect 10793 8449 10827 8483
rect 11161 8449 11195 8483
rect 11529 8449 11563 8483
rect 11713 8449 11747 8483
rect 12265 8449 12299 8483
rect 12357 8449 12391 8483
rect 12725 8449 12759 8483
rect 12817 8449 12851 8483
rect 13553 8449 13587 8483
rect 13829 8449 13863 8483
rect 15117 8449 15151 8483
rect 15209 8449 15243 8483
rect 15669 8449 15703 8483
rect 15761 8449 15795 8483
rect 15945 8449 15979 8483
rect 16681 8449 16715 8483
rect 16957 8449 16991 8483
rect 17509 8449 17543 8483
rect 17693 8449 17727 8483
rect 20294 8449 20328 8483
rect 20545 8449 20579 8483
rect 23673 8449 23707 8483
rect 23949 8449 23983 8483
rect 24501 8449 24535 8483
rect 29745 8449 29779 8483
rect 30665 8449 30699 8483
rect 31033 8449 31067 8483
rect 31309 8449 31343 8483
rect 31953 8449 31987 8483
rect 32229 8449 32263 8483
rect 13737 8381 13771 8415
rect 17049 8381 17083 8415
rect 20453 8381 20487 8415
rect 23765 8381 23799 8415
rect 24317 8381 24351 8415
rect 29837 8381 29871 8415
rect 7757 8313 7791 8347
rect 9137 8313 9171 8347
rect 10701 8313 10735 8347
rect 13001 8313 13035 8347
rect 15393 8313 15427 8347
rect 17877 8313 17911 8347
rect 24133 8313 24167 8347
rect 30113 8313 30147 8347
rect 32413 8313 32447 8347
rect 5825 8245 5859 8279
rect 6101 8245 6135 8279
rect 8217 8245 8251 8279
rect 8493 8245 8527 8279
rect 10057 8245 10091 8279
rect 11529 8245 11563 8279
rect 12173 8245 12207 8279
rect 13553 8245 13587 8279
rect 14933 8245 14967 8279
rect 15945 8245 15979 8279
rect 16957 8245 16991 8279
rect 17509 8245 17543 8279
rect 20269 8245 20303 8279
rect 23765 8245 23799 8279
rect 24225 8245 24259 8279
rect 29929 8245 29963 8279
rect 31217 8245 31251 8279
rect 8585 8041 8619 8075
rect 8953 8041 8987 8075
rect 11253 8041 11287 8075
rect 11713 8041 11747 8075
rect 13185 8041 13219 8075
rect 14657 8041 14691 8075
rect 14841 8041 14875 8075
rect 16681 8041 16715 8075
rect 17141 8041 17175 8075
rect 19533 8041 19567 8075
rect 20085 8041 20119 8075
rect 21741 8041 21775 8075
rect 22201 8041 22235 8075
rect 22845 8041 22879 8075
rect 25789 8041 25823 8075
rect 32505 8041 32539 8075
rect 17601 7973 17635 8007
rect 22109 7973 22143 8007
rect 29377 7973 29411 8007
rect 14565 7905 14599 7939
rect 16865 7905 16899 7939
rect 19349 7905 19383 7939
rect 19901 7905 19935 7939
rect 21833 7905 21867 7939
rect 25881 7905 25915 7939
rect 6193 7837 6227 7871
rect 6469 7837 6503 7871
rect 6561 7837 6595 7871
rect 8401 7837 8435 7871
rect 9137 7837 9171 7871
rect 9229 7837 9263 7871
rect 9321 7837 9355 7871
rect 9505 7837 9539 7871
rect 11437 7837 11471 7871
rect 11529 7837 11563 7871
rect 12725 7837 12759 7871
rect 13001 7837 13035 7871
rect 14473 7837 14507 7871
rect 16221 7837 16255 7871
rect 16957 7837 16991 7871
rect 17233 7837 17267 7871
rect 19533 7837 19567 7871
rect 20085 7837 20119 7871
rect 21741 7837 21775 7871
rect 22201 7837 22235 7871
rect 22293 7837 22327 7871
rect 22661 7837 22695 7871
rect 22753 7837 22787 7871
rect 26065 7837 26099 7871
rect 28825 7837 28859 7871
rect 29193 7837 29227 7871
rect 29561 7837 29595 7871
rect 31125 7837 31159 7871
rect 31381 7837 31415 7871
rect 6377 7769 6411 7803
rect 16037 7769 16071 7803
rect 16681 7769 16715 7803
rect 17417 7769 17451 7803
rect 19257 7769 19291 7803
rect 19809 7769 19843 7803
rect 25789 7769 25823 7803
rect 29009 7769 29043 7803
rect 29101 7769 29135 7803
rect 29806 7769 29840 7803
rect 6745 7701 6779 7735
rect 12909 7701 12943 7735
rect 16405 7701 16439 7735
rect 19717 7701 19751 7735
rect 20269 7701 20303 7735
rect 22569 7701 22603 7735
rect 23029 7701 23063 7735
rect 26249 7701 26283 7735
rect 30941 7701 30975 7735
rect 6929 7497 6963 7531
rect 7205 7497 7239 7531
rect 7849 7497 7883 7531
rect 8493 7497 8527 7531
rect 13461 7497 13495 7531
rect 16313 7497 16347 7531
rect 21925 7497 21959 7531
rect 24317 7497 24351 7531
rect 26249 7497 26283 7531
rect 30113 7497 30147 7531
rect 4077 7429 4111 7463
rect 4169 7429 4203 7463
rect 5825 7429 5859 7463
rect 6561 7429 6595 7463
rect 6653 7429 6687 7463
rect 7481 7429 7515 7463
rect 13369 7429 13403 7463
rect 19349 7429 19383 7463
rect 22109 7429 22143 7463
rect 23857 7429 23891 7463
rect 28089 7429 28123 7463
rect 3893 7361 3927 7395
rect 4261 7361 4295 7395
rect 4537 7361 4571 7395
rect 4721 7361 4755 7395
rect 4813 7361 4847 7395
rect 4905 7361 4939 7395
rect 5365 7361 5399 7395
rect 5641 7361 5675 7395
rect 5917 7361 5951 7395
rect 6009 7361 6043 7395
rect 6377 7361 6411 7395
rect 6745 7361 6779 7395
rect 7021 7361 7055 7395
rect 7297 7361 7331 7395
rect 7573 7361 7607 7395
rect 7665 7361 7699 7395
rect 7941 7361 7975 7395
rect 8125 7361 8159 7395
rect 8217 7361 8251 7395
rect 8309 7361 8343 7395
rect 8585 7361 8619 7395
rect 8769 7361 8803 7395
rect 8861 7361 8895 7395
rect 8953 7361 8987 7395
rect 9229 7361 9263 7395
rect 9413 7361 9447 7395
rect 9505 7361 9539 7395
rect 9597 7361 9631 7395
rect 9873 7361 9907 7395
rect 10425 7361 10459 7395
rect 12541 7361 12575 7395
rect 12817 7361 12851 7395
rect 13185 7361 13219 7395
rect 13645 7361 13679 7395
rect 16497 7361 16531 7395
rect 22385 7361 22419 7395
rect 24133 7361 24167 7395
rect 25881 7361 25915 7395
rect 25973 7361 26007 7395
rect 27813 7361 27847 7395
rect 31953 7361 31987 7395
rect 32137 7361 32171 7395
rect 12357 7293 12391 7327
rect 12633 7293 12667 7327
rect 22293 7293 22327 7327
rect 24041 7293 24075 7327
rect 27905 7293 27939 7327
rect 30757 7293 30791 7327
rect 4445 7225 4479 7259
rect 5089 7225 5123 7259
rect 5181 7225 5215 7259
rect 9781 7225 9815 7259
rect 10057 7225 10091 7259
rect 27629 7225 27663 7259
rect 6193 7157 6227 7191
rect 9137 7157 9171 7191
rect 10609 7157 10643 7191
rect 12817 7157 12851 7191
rect 13001 7157 13035 7191
rect 22109 7157 22143 7191
rect 22569 7157 22603 7191
rect 24133 7157 24167 7191
rect 26065 7157 26099 7191
rect 27813 7157 27847 7191
rect 31309 7157 31343 7191
rect 32321 7157 32355 7191
rect 4721 6953 4755 6987
rect 7849 6953 7883 6987
rect 9597 6953 9631 6987
rect 10517 6953 10551 6987
rect 13001 6953 13035 6987
rect 13645 6953 13679 6987
rect 17969 6953 18003 6987
rect 18521 6953 18555 6987
rect 20361 6953 20395 6987
rect 22201 6953 22235 6987
rect 22569 6953 22603 6987
rect 26433 6953 26467 6987
rect 32505 6953 32539 6987
rect 13829 6885 13863 6919
rect 10333 6817 10367 6851
rect 11713 6817 11747 6851
rect 13553 6817 13587 6851
rect 18429 6817 18463 6851
rect 20269 6817 20303 6851
rect 24777 6817 24811 6851
rect 31125 6817 31159 6851
rect 4905 6749 4939 6783
rect 7665 6749 7699 6783
rect 9321 6749 9355 6783
rect 9413 6749 9447 6783
rect 10517 6749 10551 6783
rect 10885 6749 10919 6783
rect 11161 6749 11195 6783
rect 11437 6749 11471 6783
rect 12817 6749 12851 6783
rect 13461 6749 13495 6783
rect 15209 6749 15243 6783
rect 15853 6765 15887 6799
rect 16221 6749 16255 6783
rect 17785 6749 17819 6783
rect 18245 6749 18279 6783
rect 18797 6749 18831 6783
rect 20085 6749 20119 6783
rect 20361 6749 20395 6783
rect 22477 6749 22511 6783
rect 22569 6749 22603 6783
rect 24409 6749 24443 6783
rect 26433 6749 26467 6783
rect 26525 6749 26559 6783
rect 30481 6749 30515 6783
rect 30757 6749 30791 6783
rect 30849 6749 30883 6783
rect 9597 6681 9631 6715
rect 10241 6681 10275 6715
rect 15393 6681 15427 6715
rect 15577 6681 15611 6715
rect 16037 6681 16071 6715
rect 17601 6681 17635 6715
rect 18521 6681 18555 6715
rect 22293 6681 22327 6715
rect 24593 6681 24627 6715
rect 30665 6681 30699 6715
rect 31370 6681 31404 6715
rect 9137 6613 9171 6647
rect 10701 6613 10735 6647
rect 11069 6613 11103 6647
rect 11345 6613 11379 6647
rect 15669 6613 15703 6647
rect 16405 6613 16439 6647
rect 18061 6613 18095 6647
rect 18613 6613 18647 6647
rect 18981 6613 19015 6647
rect 20545 6613 20579 6647
rect 22753 6613 22787 6647
rect 26801 6613 26835 6647
rect 31033 6613 31067 6647
rect 14565 6409 14599 6443
rect 15761 6409 15795 6443
rect 18613 6409 18647 6443
rect 22293 6409 22327 6443
rect 22753 6409 22787 6443
rect 23397 6409 23431 6443
rect 26617 6409 26651 6443
rect 32413 6409 32447 6443
rect 19901 6341 19935 6375
rect 20913 6341 20947 6375
rect 24869 6341 24903 6375
rect 10609 6273 10643 6307
rect 10793 6273 10827 6307
rect 11529 6273 11563 6307
rect 14197 6295 14231 6329
rect 15393 6273 15427 6307
rect 15577 6273 15611 6307
rect 17049 6273 17083 6307
rect 17325 6273 17359 6307
rect 17601 6273 17635 6307
rect 17877 6273 17911 6307
rect 18889 6273 18923 6307
rect 18981 6273 19015 6307
rect 19257 6273 19291 6307
rect 20177 6273 20211 6307
rect 21097 6273 21131 6307
rect 21833 6273 21867 6307
rect 22109 6273 22143 6307
rect 22385 6273 22419 6307
rect 23213 6273 23247 6307
rect 23489 6273 23523 6307
rect 25053 6273 25087 6307
rect 25329 6273 25363 6307
rect 25421 6273 25455 6307
rect 25973 6273 26007 6307
rect 26157 6273 26191 6307
rect 26341 6273 26375 6307
rect 26433 6273 26467 6307
rect 32229 6273 32263 6307
rect 11621 6205 11655 6239
rect 14289 6205 14323 6239
rect 17233 6205 17267 6239
rect 19993 6205 20027 6239
rect 21281 6205 21315 6239
rect 21925 6205 21959 6239
rect 22477 6205 22511 6239
rect 19073 6137 19107 6171
rect 10977 6069 11011 6103
rect 11713 6069 11747 6103
rect 11897 6069 11931 6103
rect 14197 6069 14231 6103
rect 17049 6069 17083 6103
rect 17509 6069 17543 6103
rect 17785 6069 17819 6103
rect 18061 6069 18095 6103
rect 18981 6069 19015 6103
rect 20085 6069 20119 6103
rect 20361 6069 20395 6103
rect 22109 6069 22143 6103
rect 22385 6069 22419 6103
rect 23673 6069 23707 6103
rect 25237 6069 25271 6103
rect 25329 6069 25363 6103
rect 25697 6069 25731 6103
rect 26157 6069 26191 6103
rect 6837 5865 6871 5899
rect 13553 5865 13587 5899
rect 18245 5865 18279 5899
rect 18705 5865 18739 5899
rect 23029 5865 23063 5899
rect 23489 5865 23523 5899
rect 23949 5865 23983 5899
rect 9229 5797 9263 5831
rect 17325 5729 17359 5763
rect 18337 5729 18371 5763
rect 23673 5729 23707 5763
rect 7389 5661 7423 5695
rect 8125 5661 8159 5695
rect 8585 5661 8619 5695
rect 9045 5661 9079 5695
rect 18521 5661 18555 5695
rect 23397 5661 23431 5695
rect 23765 5661 23799 5695
rect 6929 5593 6963 5627
rect 7113 5593 7147 5627
rect 13185 5593 13219 5627
rect 13369 5593 13403 5627
rect 16957 5593 16991 5627
rect 17141 5593 17175 5627
rect 18245 5593 18279 5627
rect 23213 5593 23247 5627
rect 23489 5593 23523 5627
rect 7205 5525 7239 5559
rect 8309 5525 8343 5559
rect 8401 5525 8435 5559
rect 8677 5321 8711 5355
rect 12081 5321 12115 5355
rect 23121 5321 23155 5355
rect 8217 5253 8251 5287
rect 11621 5253 11655 5287
rect 18061 5253 18095 5287
rect 23857 5253 23891 5287
rect 24685 5253 24719 5287
rect 8493 5185 8527 5219
rect 11897 5185 11931 5219
rect 14473 5185 14507 5219
rect 14565 5185 14599 5219
rect 14841 5185 14875 5219
rect 18337 5185 18371 5219
rect 23581 5185 23615 5219
rect 23765 5185 23799 5219
rect 23949 5185 23983 5219
rect 24409 5185 24443 5219
rect 24501 5185 24535 5219
rect 24777 5185 24811 5219
rect 24869 5185 24903 5219
rect 25145 5185 25179 5219
rect 8401 5117 8435 5151
rect 11713 5117 11747 5151
rect 18153 5117 18187 5151
rect 25697 5117 25731 5151
rect 14197 5049 14231 5083
rect 14657 5049 14691 5083
rect 18521 5049 18555 5083
rect 8401 4981 8435 5015
rect 11621 4981 11655 5015
rect 14565 4981 14599 5015
rect 18061 4981 18095 5015
rect 24133 4981 24167 5015
rect 24225 4981 24259 5015
rect 25053 4981 25087 5015
rect 12357 4777 12391 4811
rect 14565 4777 14599 4811
rect 14749 4777 14783 4811
rect 16129 4777 16163 4811
rect 16313 4777 16347 4811
rect 12633 4709 12667 4743
rect 13001 4709 13035 4743
rect 22845 4709 22879 4743
rect 23765 4709 23799 4743
rect 24409 4709 24443 4743
rect 12265 4641 12299 4675
rect 15945 4641 15979 4675
rect 9965 4573 9999 4607
rect 10149 4573 10183 4607
rect 10333 4573 10367 4607
rect 12173 4573 12207 4607
rect 12449 4573 12483 4607
rect 12817 4573 12851 4607
rect 14381 4573 14415 4607
rect 14565 4573 14599 4607
rect 15853 4573 15887 4607
rect 16129 4573 16163 4607
rect 19809 4573 19843 4607
rect 20821 4573 20855 4607
rect 21189 4573 21223 4607
rect 22293 4573 22327 4607
rect 22477 4573 22511 4607
rect 22661 4573 22695 4607
rect 23029 4573 23063 4607
rect 23581 4573 23615 4607
rect 23949 4573 23983 4607
rect 24225 4573 24259 4607
rect 24593 4573 24627 4607
rect 24869 4573 24903 4607
rect 25125 4573 25159 4607
rect 21005 4505 21039 4539
rect 21097 4505 21131 4539
rect 22569 4505 22603 4539
rect 19257 4437 19291 4471
rect 21373 4437 21407 4471
rect 24041 4437 24075 4471
rect 26249 4437 26283 4471
rect 18889 4233 18923 4267
rect 21557 4233 21591 4267
rect 25329 4233 25363 4267
rect 16937 4097 16971 4131
rect 20002 4097 20036 4131
rect 20269 4097 20303 4131
rect 22201 4097 22235 4131
rect 22468 4097 22502 4131
rect 23857 4097 23891 4131
rect 24124 4097 24158 4131
rect 16681 4029 16715 4063
rect 20913 4029 20947 4063
rect 25881 4029 25915 4063
rect 18245 3961 18279 3995
rect 18061 3893 18095 3927
rect 23581 3893 23615 3927
rect 25237 3893 25271 3927
rect 16773 3621 16807 3655
rect 18797 3621 18831 3655
rect 17509 3553 17543 3587
rect 21925 3553 21959 3587
rect 16221 3485 16255 3519
rect 16405 3485 16439 3519
rect 16589 3485 16623 3519
rect 16865 3485 16899 3519
rect 18245 3485 18279 3519
rect 18521 3485 18555 3519
rect 18613 3485 18647 3519
rect 21658 3485 21692 3519
rect 16497 3417 16531 3451
rect 18429 3417 18463 3451
rect 20545 3349 20579 3383
rect 17785 2397 17819 2431
rect 19717 2397 19751 2431
rect 21373 2397 21407 2431
rect 22937 2397 22971 2431
rect 24869 2397 24903 2431
rect 25881 2397 25915 2431
rect 29745 2397 29779 2431
rect 17601 2261 17635 2295
rect 19533 2261 19567 2295
rect 21557 2261 21591 2295
rect 22753 2261 22787 2295
rect 24685 2261 24719 2295
rect 26065 2261 26099 2295
<< metal1 >>
rect 1104 31578 32844 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 32844 31578
rect 1104 31504 32844 31526
rect 18690 31424 18696 31476
rect 18748 31464 18754 31476
rect 19429 31467 19487 31473
rect 19429 31464 19441 31467
rect 18748 31436 19441 31464
rect 18748 31424 18754 31436
rect 19429 31433 19441 31436
rect 19475 31433 19487 31467
rect 19429 31427 19487 31433
rect 21266 31424 21272 31476
rect 21324 31464 21330 31476
rect 22189 31467 22247 31473
rect 22189 31464 22201 31467
rect 21324 31436 22201 31464
rect 21324 31424 21330 31436
rect 22189 31433 22201 31436
rect 22235 31433 22247 31467
rect 22189 31427 22247 31433
rect 25130 31424 25136 31476
rect 25188 31464 25194 31476
rect 25409 31467 25467 31473
rect 25409 31464 25421 31467
rect 25188 31436 25421 31464
rect 25188 31424 25194 31436
rect 25409 31433 25421 31436
rect 25455 31433 25467 31467
rect 25409 31427 25467 31433
rect 16758 31356 16764 31408
rect 16816 31396 16822 31408
rect 16853 31399 16911 31405
rect 16853 31396 16865 31399
rect 16816 31368 16865 31396
rect 16816 31356 16822 31368
rect 16853 31365 16865 31368
rect 16899 31365 16911 31399
rect 16853 31359 16911 31365
rect 23198 31356 23204 31408
rect 23256 31396 23262 31408
rect 23293 31399 23351 31405
rect 23293 31396 23305 31399
rect 23256 31368 23305 31396
rect 23256 31356 23262 31368
rect 23293 31365 23305 31368
rect 23339 31365 23351 31399
rect 23293 31359 23351 31365
rect 17126 31288 17132 31340
rect 17184 31328 17190 31340
rect 17221 31331 17279 31337
rect 17221 31328 17233 31331
rect 17184 31300 17233 31328
rect 17184 31288 17190 31300
rect 17221 31297 17233 31300
rect 17267 31297 17279 31331
rect 17221 31291 17279 31297
rect 19334 31288 19340 31340
rect 19392 31288 19398 31340
rect 21910 31288 21916 31340
rect 21968 31288 21974 31340
rect 23658 31288 23664 31340
rect 23716 31288 23722 31340
rect 25314 31288 25320 31340
rect 25372 31288 25378 31340
rect 1104 31034 32844 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 32844 31034
rect 1104 30960 32844 30982
rect 13446 30744 13452 30796
rect 13504 30784 13510 30796
rect 26970 30784 26976 30796
rect 13504 30756 26976 30784
rect 13504 30744 13510 30756
rect 26970 30744 26976 30756
rect 27028 30744 27034 30796
rect 18506 30716 18512 30728
rect 2746 30688 18512 30716
rect 1302 30540 1308 30592
rect 1360 30580 1366 30592
rect 2746 30580 2774 30688
rect 18506 30676 18512 30688
rect 18564 30676 18570 30728
rect 14826 30608 14832 30660
rect 14884 30648 14890 30660
rect 32306 30648 32312 30660
rect 14884 30620 32312 30648
rect 14884 30608 14890 30620
rect 32306 30608 32312 30620
rect 32364 30608 32370 30660
rect 1360 30552 2774 30580
rect 1360 30540 1366 30552
rect 14090 30540 14096 30592
rect 14148 30580 14154 30592
rect 28258 30580 28264 30592
rect 14148 30552 28264 30580
rect 14148 30540 14154 30552
rect 28258 30540 28264 30552
rect 28316 30540 28322 30592
rect 1104 30490 32844 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 32844 30490
rect 1104 30416 32844 30438
rect 6086 30336 6092 30388
rect 6144 30376 6150 30388
rect 14090 30376 14096 30388
rect 6144 30348 14096 30376
rect 6144 30336 6150 30348
rect 14090 30336 14096 30348
rect 14148 30336 14154 30388
rect 21637 30379 21695 30385
rect 21637 30345 21649 30379
rect 21683 30376 21695 30379
rect 21910 30376 21916 30388
rect 21683 30348 21916 30376
rect 21683 30345 21695 30348
rect 21637 30339 21695 30345
rect 21910 30336 21916 30348
rect 21968 30376 21974 30388
rect 21968 30348 22094 30376
rect 21968 30336 21974 30348
rect 17420 30280 20300 30308
rect 17310 30200 17316 30252
rect 17368 30240 17374 30252
rect 17420 30249 17448 30280
rect 17405 30243 17463 30249
rect 17405 30240 17417 30243
rect 17368 30212 17417 30240
rect 17368 30200 17374 30212
rect 17405 30209 17417 30212
rect 17451 30209 17463 30243
rect 17405 30203 17463 30209
rect 17672 30243 17730 30249
rect 17672 30209 17684 30243
rect 17718 30240 17730 30243
rect 18690 30240 18696 30252
rect 17718 30212 18696 30240
rect 17718 30209 17730 30212
rect 17672 30203 17730 30209
rect 18690 30200 18696 30212
rect 18748 30200 18754 30252
rect 19334 30200 19340 30252
rect 19392 30240 19398 30252
rect 19429 30243 19487 30249
rect 19429 30240 19441 30243
rect 19392 30212 19441 30240
rect 19392 30200 19398 30212
rect 19429 30209 19441 30212
rect 19475 30209 19487 30243
rect 19429 30203 19487 30209
rect 18785 30107 18843 30113
rect 18785 30073 18797 30107
rect 18831 30104 18843 30107
rect 19352 30104 19380 30200
rect 20272 30181 20300 30280
rect 20530 30249 20536 30252
rect 20524 30203 20536 30249
rect 20530 30200 20536 30203
rect 20588 30200 20594 30252
rect 22066 30240 22094 30348
rect 22373 30243 22431 30249
rect 22373 30240 22385 30243
rect 22066 30212 22385 30240
rect 22373 30209 22385 30212
rect 22419 30209 22431 30243
rect 22373 30203 22431 30209
rect 22741 30243 22799 30249
rect 22741 30209 22753 30243
rect 22787 30240 22799 30243
rect 26142 30240 26148 30252
rect 22787 30212 26148 30240
rect 22787 30209 22799 30212
rect 22741 30203 22799 30209
rect 26142 30200 26148 30212
rect 26200 30200 26206 30252
rect 20257 30175 20315 30181
rect 20257 30141 20269 30175
rect 20303 30141 20315 30175
rect 20257 30135 20315 30141
rect 18831 30076 19380 30104
rect 18831 30073 18843 30076
rect 18785 30067 18843 30073
rect 934 29996 940 30048
rect 992 30036 998 30048
rect 10686 30036 10692 30048
rect 992 30008 10692 30036
rect 992 29996 998 30008
rect 10686 29996 10692 30008
rect 10744 29996 10750 30048
rect 18874 29996 18880 30048
rect 18932 29996 18938 30048
rect 20272 30036 20300 30135
rect 21821 30107 21879 30113
rect 21821 30104 21833 30107
rect 21192 30076 21833 30104
rect 20622 30036 20628 30048
rect 20272 30008 20628 30036
rect 20622 29996 20628 30008
rect 20680 29996 20686 30048
rect 20898 29996 20904 30048
rect 20956 30036 20962 30048
rect 21192 30036 21220 30076
rect 21821 30073 21833 30076
rect 21867 30073 21879 30107
rect 21821 30067 21879 30073
rect 20956 30008 21220 30036
rect 20956 29996 20962 30008
rect 22186 29996 22192 30048
rect 22244 30036 22250 30048
rect 22557 30039 22615 30045
rect 22557 30036 22569 30039
rect 22244 30008 22569 30036
rect 22244 29996 22250 30008
rect 22557 30005 22569 30008
rect 22603 30005 22615 30039
rect 22557 29999 22615 30005
rect 1104 29946 32844 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 32844 29946
rect 1104 29872 32844 29894
rect 1210 29792 1216 29844
rect 1268 29832 1274 29844
rect 8846 29832 8852 29844
rect 1268 29804 8852 29832
rect 1268 29792 1274 29804
rect 8846 29792 8852 29804
rect 8904 29832 8910 29844
rect 9125 29835 9183 29841
rect 9125 29832 9137 29835
rect 8904 29804 9137 29832
rect 8904 29792 8910 29804
rect 9125 29801 9137 29804
rect 9171 29801 9183 29835
rect 9125 29795 9183 29801
rect 9858 29792 9864 29844
rect 9916 29832 9922 29844
rect 10321 29835 10379 29841
rect 10321 29832 10333 29835
rect 9916 29804 10333 29832
rect 9916 29792 9922 29804
rect 10321 29801 10333 29804
rect 10367 29801 10379 29835
rect 10321 29795 10379 29801
rect 15933 29835 15991 29841
rect 15933 29801 15945 29835
rect 15979 29832 15991 29835
rect 17126 29832 17132 29844
rect 15979 29804 17132 29832
rect 15979 29801 15991 29804
rect 15933 29795 15991 29801
rect 17126 29792 17132 29804
rect 17184 29832 17190 29844
rect 17184 29804 18000 29832
rect 17184 29792 17190 29804
rect 1026 29724 1032 29776
rect 1084 29764 1090 29776
rect 7190 29764 7196 29776
rect 1084 29736 7196 29764
rect 1084 29724 1090 29736
rect 7190 29724 7196 29736
rect 7248 29724 7254 29776
rect 9398 29724 9404 29776
rect 9456 29764 9462 29776
rect 9493 29767 9551 29773
rect 9493 29764 9505 29767
rect 9456 29736 9505 29764
rect 9456 29724 9462 29736
rect 9493 29733 9505 29736
rect 9539 29733 9551 29767
rect 9493 29727 9551 29733
rect 10229 29767 10287 29773
rect 10229 29733 10241 29767
rect 10275 29764 10287 29767
rect 11698 29764 11704 29776
rect 10275 29736 11704 29764
rect 10275 29733 10287 29736
rect 10229 29727 10287 29733
rect 11698 29724 11704 29736
rect 11756 29724 11762 29776
rect 5626 29656 5632 29708
rect 5684 29696 5690 29708
rect 5684 29668 10548 29696
rect 5684 29656 5690 29668
rect 3145 29631 3203 29637
rect 3145 29597 3157 29631
rect 3191 29597 3203 29631
rect 3145 29591 3203 29597
rect 3160 29560 3188 29591
rect 3234 29588 3240 29640
rect 3292 29588 3298 29640
rect 7006 29588 7012 29640
rect 7064 29628 7070 29640
rect 10520 29637 10548 29668
rect 17310 29656 17316 29708
rect 17368 29656 17374 29708
rect 17972 29705 18000 29804
rect 18690 29792 18696 29844
rect 18748 29792 18754 29844
rect 20530 29792 20536 29844
rect 20588 29832 20594 29844
rect 20717 29835 20775 29841
rect 20717 29832 20729 29835
rect 20588 29804 20729 29832
rect 20588 29792 20594 29804
rect 20717 29801 20729 29804
rect 20763 29801 20775 29835
rect 20717 29795 20775 29801
rect 23385 29835 23443 29841
rect 23385 29801 23397 29835
rect 23431 29832 23443 29835
rect 23658 29832 23664 29844
rect 23431 29804 23664 29832
rect 23431 29801 23443 29804
rect 23385 29795 23443 29801
rect 23658 29792 23664 29804
rect 23716 29792 23722 29844
rect 17957 29699 18015 29705
rect 17957 29665 17969 29699
rect 18003 29665 18015 29699
rect 17957 29659 18015 29665
rect 20622 29656 20628 29708
rect 20680 29696 20686 29708
rect 22005 29699 22063 29705
rect 22005 29696 22017 29699
rect 20680 29668 22017 29696
rect 20680 29656 20686 29668
rect 22005 29665 22017 29668
rect 22051 29665 22063 29699
rect 23676 29696 23704 29792
rect 24029 29699 24087 29705
rect 24029 29696 24041 29699
rect 23676 29668 24041 29696
rect 22005 29659 22063 29665
rect 24029 29665 24041 29668
rect 24075 29665 24087 29699
rect 24029 29659 24087 29665
rect 9309 29631 9367 29637
rect 9309 29628 9321 29631
rect 7064 29600 9321 29628
rect 7064 29588 7070 29600
rect 9309 29597 9321 29600
rect 9355 29597 9367 29631
rect 9309 29591 9367 29597
rect 9677 29631 9735 29637
rect 9677 29597 9689 29631
rect 9723 29597 9735 29631
rect 9677 29591 9735 29597
rect 10045 29631 10103 29637
rect 10045 29597 10057 29631
rect 10091 29597 10103 29631
rect 10045 29591 10103 29597
rect 10505 29631 10563 29637
rect 10505 29597 10517 29631
rect 10551 29597 10563 29631
rect 10505 29591 10563 29597
rect 10597 29631 10655 29637
rect 10597 29597 10609 29631
rect 10643 29597 10655 29631
rect 10597 29591 10655 29597
rect 3160 29532 3464 29560
rect 3436 29504 3464 29532
rect 9122 29520 9128 29572
rect 9180 29560 9186 29572
rect 9692 29560 9720 29591
rect 9180 29532 9720 29560
rect 9180 29520 9186 29532
rect 2961 29495 3019 29501
rect 2961 29461 2973 29495
rect 3007 29492 3019 29495
rect 3326 29492 3332 29504
rect 3007 29464 3332 29492
rect 3007 29461 3019 29464
rect 2961 29455 3019 29461
rect 3326 29452 3332 29464
rect 3384 29452 3390 29504
rect 3418 29452 3424 29504
rect 3476 29452 3482 29504
rect 5258 29452 5264 29504
rect 5316 29492 5322 29504
rect 10060 29492 10088 29591
rect 10226 29520 10232 29572
rect 10284 29560 10290 29572
rect 10612 29560 10640 29591
rect 10686 29588 10692 29640
rect 10744 29628 10750 29640
rect 16574 29628 16580 29640
rect 10744 29600 16580 29628
rect 10744 29588 10750 29600
rect 16574 29588 16580 29600
rect 16632 29588 16638 29640
rect 17494 29588 17500 29640
rect 17552 29628 17558 29640
rect 18141 29631 18199 29637
rect 18141 29628 18153 29631
rect 17552 29600 18153 29628
rect 17552 29588 17558 29600
rect 18141 29597 18153 29600
rect 18187 29597 18199 29631
rect 18141 29591 18199 29597
rect 18509 29631 18567 29637
rect 18509 29597 18521 29631
rect 18555 29628 18567 29631
rect 18874 29628 18880 29640
rect 18555 29600 18880 29628
rect 18555 29597 18567 29600
rect 18509 29591 18567 29597
rect 18874 29588 18880 29600
rect 18932 29588 18938 29640
rect 20898 29588 20904 29640
rect 20956 29588 20962 29640
rect 21008 29600 21220 29628
rect 10284 29532 10640 29560
rect 17068 29563 17126 29569
rect 10284 29520 10290 29532
rect 17068 29529 17080 29563
rect 17114 29560 17126 29563
rect 17218 29560 17224 29572
rect 17114 29532 17224 29560
rect 17114 29529 17126 29532
rect 17068 29523 17126 29529
rect 17218 29520 17224 29532
rect 17276 29520 17282 29572
rect 18325 29563 18383 29569
rect 18325 29560 18337 29563
rect 17328 29532 18337 29560
rect 5316 29464 10088 29492
rect 5316 29452 5322 29464
rect 10502 29452 10508 29504
rect 10560 29492 10566 29504
rect 10781 29495 10839 29501
rect 10781 29492 10793 29495
rect 10560 29464 10793 29492
rect 10560 29452 10566 29464
rect 10781 29461 10793 29464
rect 10827 29461 10839 29495
rect 10781 29455 10839 29461
rect 16850 29452 16856 29504
rect 16908 29492 16914 29504
rect 17328 29492 17356 29532
rect 18325 29529 18337 29532
rect 18371 29529 18383 29563
rect 18325 29523 18383 29529
rect 16908 29464 17356 29492
rect 16908 29452 16914 29464
rect 17402 29452 17408 29504
rect 17460 29452 17466 29504
rect 18340 29492 18368 29523
rect 18414 29520 18420 29572
rect 18472 29560 18478 29572
rect 21008 29569 21036 29600
rect 20993 29563 21051 29569
rect 20993 29560 21005 29563
rect 18472 29532 21005 29560
rect 18472 29520 18478 29532
rect 20993 29529 21005 29532
rect 21039 29529 21051 29563
rect 20993 29523 21051 29529
rect 21085 29563 21143 29569
rect 21085 29529 21097 29563
rect 21131 29529 21143 29563
rect 21192 29560 21220 29600
rect 21266 29588 21272 29640
rect 21324 29588 21330 29640
rect 21913 29631 21971 29637
rect 21913 29597 21925 29631
rect 21959 29628 21971 29631
rect 21959 29600 25728 29628
rect 21959 29597 21971 29600
rect 21913 29591 21971 29597
rect 22272 29563 22330 29569
rect 21192 29532 22232 29560
rect 21085 29523 21143 29529
rect 21100 29492 21128 29523
rect 22204 29504 22232 29532
rect 22272 29529 22284 29563
rect 22318 29560 22330 29563
rect 22462 29560 22468 29572
rect 22318 29532 22468 29560
rect 22318 29529 22330 29532
rect 22272 29523 22330 29529
rect 22462 29520 22468 29532
rect 22520 29520 22526 29572
rect 24486 29520 24492 29572
rect 24544 29560 24550 29572
rect 25510 29563 25568 29569
rect 25510 29560 25522 29563
rect 24544 29532 25522 29560
rect 24544 29520 24550 29532
rect 25510 29529 25522 29532
rect 25556 29529 25568 29563
rect 25700 29560 25728 29600
rect 25774 29588 25780 29640
rect 25832 29588 25838 29640
rect 28994 29560 29000 29572
rect 25700 29532 29000 29560
rect 25510 29523 25568 29529
rect 28994 29520 29000 29532
rect 29052 29520 29058 29572
rect 21729 29495 21787 29501
rect 21729 29492 21741 29495
rect 18340 29464 21741 29492
rect 21729 29461 21741 29464
rect 21775 29492 21787 29495
rect 22094 29492 22100 29504
rect 21775 29464 22100 29492
rect 21775 29461 21787 29464
rect 21729 29455 21787 29461
rect 22094 29452 22100 29464
rect 22152 29452 22158 29504
rect 22186 29452 22192 29504
rect 22244 29452 22250 29504
rect 22370 29452 22376 29504
rect 22428 29492 22434 29504
rect 23477 29495 23535 29501
rect 23477 29492 23489 29495
rect 22428 29464 23489 29492
rect 22428 29452 22434 29464
rect 23477 29461 23489 29464
rect 23523 29461 23535 29495
rect 23477 29455 23535 29461
rect 24397 29495 24455 29501
rect 24397 29461 24409 29495
rect 24443 29492 24455 29495
rect 25314 29492 25320 29504
rect 24443 29464 25320 29492
rect 24443 29461 24455 29464
rect 24397 29455 24455 29461
rect 25314 29452 25320 29464
rect 25372 29452 25378 29504
rect 1104 29402 32844 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 32844 29402
rect 1104 29328 32844 29350
rect 3510 29288 3516 29300
rect 2516 29260 3516 29288
rect 1394 29112 1400 29164
rect 1452 29112 1458 29164
rect 2516 29161 2544 29260
rect 3510 29248 3516 29260
rect 3568 29248 3574 29300
rect 3697 29291 3755 29297
rect 3697 29257 3709 29291
rect 3743 29288 3755 29291
rect 3743 29260 8984 29288
rect 3743 29257 3755 29260
rect 3697 29251 3755 29257
rect 2774 29180 2780 29232
rect 2832 29220 2838 29232
rect 2832 29192 3188 29220
rect 2832 29180 2838 29192
rect 2501 29155 2559 29161
rect 2501 29121 2513 29155
rect 2547 29121 2559 29155
rect 2501 29115 2559 29121
rect 2961 29155 3019 29161
rect 2961 29121 2973 29155
rect 3007 29152 3019 29155
rect 3050 29152 3056 29164
rect 3007 29124 3056 29152
rect 3007 29121 3019 29124
rect 2961 29115 3019 29121
rect 3050 29112 3056 29124
rect 3108 29112 3114 29164
rect 3160 29161 3188 29192
rect 3418 29180 3424 29232
rect 3476 29220 3482 29232
rect 3476 29192 5304 29220
rect 3476 29180 3482 29192
rect 3988 29161 4016 29192
rect 3145 29155 3203 29161
rect 3145 29121 3157 29155
rect 3191 29121 3203 29155
rect 3145 29115 3203 29121
rect 3513 29155 3571 29161
rect 3513 29121 3525 29155
rect 3559 29121 3571 29155
rect 3513 29115 3571 29121
rect 3973 29155 4031 29161
rect 3973 29121 3985 29155
rect 4019 29121 4031 29155
rect 3973 29115 4031 29121
rect 4249 29155 4307 29161
rect 4249 29121 4261 29155
rect 4295 29121 4307 29155
rect 4249 29115 4307 29121
rect 2222 29044 2228 29096
rect 2280 29084 2286 29096
rect 3528 29084 3556 29115
rect 2280 29056 3556 29084
rect 4264 29084 4292 29115
rect 4338 29112 4344 29164
rect 4396 29152 4402 29164
rect 4433 29155 4491 29161
rect 4433 29152 4445 29155
rect 4396 29124 4445 29152
rect 4396 29112 4402 29124
rect 4433 29121 4445 29124
rect 4479 29121 4491 29155
rect 4433 29115 4491 29121
rect 4706 29112 4712 29164
rect 4764 29112 4770 29164
rect 5276 29161 5304 29192
rect 7208 29192 7880 29220
rect 7208 29164 7236 29192
rect 5169 29155 5227 29161
rect 5169 29121 5181 29155
rect 5215 29121 5227 29155
rect 5169 29115 5227 29121
rect 5261 29155 5319 29161
rect 5261 29121 5273 29155
rect 5307 29121 5319 29155
rect 5261 29115 5319 29121
rect 4614 29084 4620 29096
rect 4264 29056 4620 29084
rect 2280 29044 2286 29056
rect 4614 29044 4620 29056
rect 4672 29044 4678 29096
rect 2685 29019 2743 29025
rect 2685 28985 2697 29019
rect 2731 29016 2743 29019
rect 2866 29016 2872 29028
rect 2731 28988 2872 29016
rect 2731 28985 2743 28988
rect 2685 28979 2743 28985
rect 2866 28976 2872 28988
rect 2924 28976 2930 29028
rect 5184 29016 5212 29115
rect 7190 29112 7196 29164
rect 7248 29112 7254 29164
rect 7466 29112 7472 29164
rect 7524 29112 7530 29164
rect 7558 29112 7564 29164
rect 7616 29152 7622 29164
rect 7745 29155 7803 29161
rect 7745 29152 7757 29155
rect 7616 29124 7757 29152
rect 7616 29112 7622 29124
rect 7745 29121 7757 29124
rect 7791 29121 7803 29155
rect 7745 29115 7803 29121
rect 3988 28988 5580 29016
rect 1581 28951 1639 28957
rect 1581 28917 1593 28951
rect 1627 28948 1639 28951
rect 1670 28948 1676 28960
rect 1627 28920 1676 28948
rect 1627 28917 1639 28920
rect 1581 28911 1639 28917
rect 1670 28908 1676 28920
rect 1728 28908 1734 28960
rect 2777 28951 2835 28957
rect 2777 28917 2789 28951
rect 2823 28948 2835 28951
rect 2958 28948 2964 28960
rect 2823 28920 2964 28948
rect 2823 28917 2835 28920
rect 2777 28911 2835 28917
rect 2958 28908 2964 28920
rect 3016 28908 3022 28960
rect 3142 28908 3148 28960
rect 3200 28948 3206 28960
rect 3329 28951 3387 28957
rect 3329 28948 3341 28951
rect 3200 28920 3341 28948
rect 3200 28908 3206 28920
rect 3329 28917 3341 28920
rect 3375 28917 3387 28951
rect 3329 28911 3387 28917
rect 3786 28908 3792 28960
rect 3844 28908 3850 28960
rect 3878 28908 3884 28960
rect 3936 28948 3942 28960
rect 3988 28948 4016 28988
rect 3936 28920 4016 28948
rect 4065 28951 4123 28957
rect 3936 28908 3942 28920
rect 4065 28917 4077 28951
rect 4111 28948 4123 28951
rect 4246 28948 4252 28960
rect 4111 28920 4252 28948
rect 4111 28917 4123 28920
rect 4065 28911 4123 28917
rect 4246 28908 4252 28920
rect 4304 28908 4310 28960
rect 4632 28957 4660 28988
rect 4617 28951 4675 28957
rect 4617 28917 4629 28951
rect 4663 28948 4675 28951
rect 4663 28920 4697 28948
rect 4663 28917 4675 28920
rect 4617 28911 4675 28917
rect 4890 28908 4896 28960
rect 4948 28908 4954 28960
rect 4982 28908 4988 28960
rect 5040 28908 5046 28960
rect 5442 28908 5448 28960
rect 5500 28908 5506 28960
rect 5552 28948 5580 28988
rect 6730 28976 6736 29028
rect 6788 29016 6794 29028
rect 7009 29019 7067 29025
rect 7009 29016 7021 29019
rect 6788 28988 7021 29016
rect 6788 28976 6794 28988
rect 7009 28985 7021 28988
rect 7055 28985 7067 29019
rect 7484 29016 7512 29112
rect 7852 29025 7880 29192
rect 8018 29112 8024 29164
rect 8076 29112 8082 29164
rect 8846 29112 8852 29164
rect 8904 29112 8910 29164
rect 8956 29161 8984 29260
rect 9122 29248 9128 29300
rect 9180 29248 9186 29300
rect 9674 29248 9680 29300
rect 9732 29248 9738 29300
rect 9766 29248 9772 29300
rect 9824 29288 9830 29300
rect 10505 29291 10563 29297
rect 10505 29288 10517 29291
rect 9824 29260 10517 29288
rect 9824 29248 9830 29260
rect 10505 29257 10517 29260
rect 10551 29257 10563 29291
rect 12805 29291 12863 29297
rect 12805 29288 12817 29291
rect 10505 29251 10563 29257
rect 12406 29260 12817 29288
rect 9030 29180 9036 29232
rect 9088 29220 9094 29232
rect 9088 29192 9996 29220
rect 9088 29180 9094 29192
rect 8941 29155 8999 29161
rect 8941 29121 8953 29155
rect 8987 29121 8999 29155
rect 8941 29115 8999 29121
rect 9398 29112 9404 29164
rect 9456 29112 9462 29164
rect 9766 29152 9772 29164
rect 9508 29124 9772 29152
rect 8662 29044 8668 29096
rect 8720 29084 8726 29096
rect 9508 29084 9536 29124
rect 9766 29112 9772 29124
rect 9824 29112 9830 29164
rect 9858 29112 9864 29164
rect 9916 29112 9922 29164
rect 9968 29161 9996 29192
rect 10042 29180 10048 29232
rect 10100 29220 10106 29232
rect 10100 29192 11744 29220
rect 10100 29180 10106 29192
rect 9953 29155 10011 29161
rect 9953 29121 9965 29155
rect 9999 29121 10011 29155
rect 9953 29115 10011 29121
rect 10413 29155 10471 29161
rect 10413 29121 10425 29155
rect 10459 29152 10471 29155
rect 10594 29152 10600 29164
rect 10459 29124 10600 29152
rect 10459 29121 10471 29124
rect 10413 29115 10471 29121
rect 10594 29112 10600 29124
rect 10652 29112 10658 29164
rect 10689 29155 10747 29161
rect 10689 29121 10701 29155
rect 10735 29121 10747 29155
rect 10689 29115 10747 29121
rect 10781 29155 10839 29161
rect 10781 29121 10793 29155
rect 10827 29152 10839 29155
rect 10962 29152 10968 29164
rect 10827 29124 10968 29152
rect 10827 29121 10839 29124
rect 10781 29115 10839 29121
rect 8720 29056 9536 29084
rect 8720 29044 8726 29056
rect 9674 29044 9680 29096
rect 9732 29084 9738 29096
rect 10704 29084 10732 29115
rect 10962 29112 10968 29124
rect 11020 29112 11026 29164
rect 11716 29161 11744 29192
rect 11057 29155 11115 29161
rect 11057 29121 11069 29155
rect 11103 29121 11115 29155
rect 11057 29115 11115 29121
rect 11701 29155 11759 29161
rect 11701 29121 11713 29155
rect 11747 29121 11759 29155
rect 11701 29115 11759 29121
rect 12161 29155 12219 29161
rect 12161 29121 12173 29155
rect 12207 29152 12219 29155
rect 12253 29155 12311 29161
rect 12253 29152 12265 29155
rect 12207 29124 12265 29152
rect 12207 29121 12219 29124
rect 12161 29115 12219 29121
rect 12253 29121 12265 29124
rect 12299 29152 12311 29155
rect 12406 29152 12434 29260
rect 12805 29257 12817 29260
rect 12851 29257 12863 29291
rect 12805 29251 12863 29257
rect 15930 29248 15936 29300
rect 15988 29248 15994 29300
rect 16301 29291 16359 29297
rect 16301 29257 16313 29291
rect 16347 29288 16359 29291
rect 16390 29288 16396 29300
rect 16347 29260 16396 29288
rect 16347 29257 16359 29260
rect 16301 29251 16359 29257
rect 16390 29248 16396 29260
rect 16448 29288 16454 29300
rect 16448 29260 18552 29288
rect 16448 29248 16454 29260
rect 12299 29124 12434 29152
rect 12299 29121 12311 29124
rect 12253 29115 12311 29121
rect 9732 29056 10732 29084
rect 9732 29044 9738 29056
rect 7561 29019 7619 29025
rect 7561 29016 7573 29019
rect 7484 28988 7573 29016
rect 7009 28979 7067 28985
rect 7561 28985 7573 28988
rect 7607 28985 7619 29019
rect 7561 28979 7619 28985
rect 7837 29019 7895 29025
rect 7837 28985 7849 29019
rect 7883 28985 7895 29019
rect 7837 28979 7895 28985
rect 8386 28976 8392 29028
rect 8444 29016 8450 29028
rect 11072 29016 11100 29115
rect 12710 29112 12716 29164
rect 12768 29112 12774 29164
rect 12989 29155 13047 29161
rect 12989 29121 13001 29155
rect 13035 29152 13047 29155
rect 13262 29152 13268 29164
rect 13035 29124 13268 29152
rect 13035 29121 13047 29124
rect 12989 29115 13047 29121
rect 13262 29112 13268 29124
rect 13320 29112 13326 29164
rect 15948 29152 15976 29248
rect 16850 29180 16856 29232
rect 16908 29180 16914 29232
rect 16945 29223 17003 29229
rect 16945 29189 16957 29223
rect 16991 29220 17003 29223
rect 18414 29220 18420 29232
rect 16991 29192 18420 29220
rect 16991 29189 17003 29192
rect 16945 29183 17003 29189
rect 18414 29180 18420 29192
rect 18472 29180 18478 29232
rect 18524 29220 18552 29260
rect 22462 29248 22468 29300
rect 22520 29248 22526 29300
rect 24486 29248 24492 29300
rect 24544 29248 24550 29300
rect 18524 29192 19334 29220
rect 16117 29155 16175 29161
rect 16117 29152 16129 29155
rect 15948 29124 16129 29152
rect 16117 29121 16129 29124
rect 16163 29121 16175 29155
rect 16117 29115 16175 29121
rect 16298 29112 16304 29164
rect 16356 29152 16362 29164
rect 16669 29155 16727 29161
rect 16669 29152 16681 29155
rect 16356 29124 16681 29152
rect 16356 29112 16362 29124
rect 16669 29121 16681 29124
rect 16715 29121 16727 29155
rect 16669 29115 16727 29121
rect 17037 29155 17095 29161
rect 17037 29121 17049 29155
rect 17083 29152 17095 29155
rect 17402 29152 17408 29164
rect 17083 29124 17408 29152
rect 17083 29121 17095 29124
rect 17037 29115 17095 29121
rect 17402 29112 17408 29124
rect 17460 29112 17466 29164
rect 17957 29155 18015 29161
rect 17957 29121 17969 29155
rect 18003 29121 18015 29155
rect 18233 29155 18291 29161
rect 18233 29152 18245 29155
rect 17957 29115 18015 29121
rect 18156 29124 18245 29152
rect 11146 29044 11152 29096
rect 11204 29084 11210 29096
rect 17972 29084 18000 29115
rect 11204 29056 18000 29084
rect 11204 29044 11210 29056
rect 18156 29028 18184 29124
rect 18233 29121 18245 29124
rect 18279 29121 18291 29155
rect 18233 29115 18291 29121
rect 19306 29084 19334 29192
rect 22094 29180 22100 29232
rect 22152 29180 22158 29232
rect 24121 29223 24179 29229
rect 24121 29220 24133 29223
rect 23860 29192 24133 29220
rect 20162 29112 20168 29164
rect 20220 29112 20226 29164
rect 21910 29112 21916 29164
rect 21968 29112 21974 29164
rect 22186 29112 22192 29164
rect 22244 29112 22250 29164
rect 22281 29155 22339 29161
rect 22281 29121 22293 29155
rect 22327 29152 22339 29155
rect 22370 29152 22376 29164
rect 22327 29124 22376 29152
rect 22327 29121 22339 29124
rect 22281 29115 22339 29121
rect 22370 29112 22376 29124
rect 22428 29112 22434 29164
rect 23477 29155 23535 29161
rect 23477 29121 23489 29155
rect 23523 29121 23535 29155
rect 23477 29115 23535 29121
rect 23492 29084 23520 29115
rect 23750 29084 23756 29096
rect 19306 29056 22048 29084
rect 8444 28988 11100 29016
rect 8444 28976 8450 28988
rect 11238 28976 11244 29028
rect 11296 29016 11302 29028
rect 12066 29016 12072 29028
rect 11296 28988 12072 29016
rect 11296 28976 11302 28988
rect 12066 28976 12072 28988
rect 12124 28976 12130 29028
rect 12437 29019 12495 29025
rect 12437 28985 12449 29019
rect 12483 29016 12495 29019
rect 12894 29016 12900 29028
rect 12483 28988 12900 29016
rect 12483 28985 12495 28988
rect 12437 28979 12495 28985
rect 12894 28976 12900 28988
rect 12952 28976 12958 29028
rect 17218 28976 17224 29028
rect 17276 28976 17282 29028
rect 18138 28976 18144 29028
rect 18196 28976 18202 29028
rect 22020 29016 22048 29056
rect 23492 29056 23756 29084
rect 23492 29016 23520 29056
rect 23750 29044 23756 29056
rect 23808 29044 23814 29096
rect 18340 28988 18552 29016
rect 22020 28988 23520 29016
rect 23860 29016 23888 29192
rect 24121 29189 24133 29192
rect 24167 29189 24179 29223
rect 24121 29183 24179 29189
rect 24213 29223 24271 29229
rect 24213 29189 24225 29223
rect 24259 29220 24271 29223
rect 29914 29220 29920 29232
rect 24259 29192 29920 29220
rect 24259 29189 24271 29192
rect 24213 29183 24271 29189
rect 29914 29180 29920 29192
rect 29972 29180 29978 29232
rect 23937 29155 23995 29161
rect 23937 29121 23949 29155
rect 23983 29121 23995 29155
rect 23937 29115 23995 29121
rect 24305 29155 24363 29161
rect 24305 29121 24317 29155
rect 24351 29152 24363 29155
rect 24581 29155 24639 29161
rect 24581 29152 24593 29155
rect 24351 29124 24593 29152
rect 24351 29121 24363 29124
rect 24305 29115 24363 29121
rect 24581 29121 24593 29124
rect 24627 29121 24639 29155
rect 24581 29115 24639 29121
rect 25225 29155 25283 29161
rect 25225 29121 25237 29155
rect 25271 29152 25283 29155
rect 25314 29152 25320 29164
rect 25271 29124 25320 29152
rect 25271 29121 25283 29124
rect 25225 29115 25283 29121
rect 23952 29084 23980 29115
rect 25314 29112 25320 29124
rect 25372 29112 25378 29164
rect 24394 29084 24400 29096
rect 23952 29056 24400 29084
rect 24394 29044 24400 29056
rect 24452 29044 24458 29096
rect 30374 29016 30380 29028
rect 23860 28988 30380 29016
rect 5902 28948 5908 28960
rect 5552 28920 5908 28948
rect 5902 28908 5908 28920
rect 5960 28908 5966 28960
rect 7098 28908 7104 28960
rect 7156 28948 7162 28960
rect 7285 28951 7343 28957
rect 7285 28948 7297 28951
rect 7156 28920 7297 28948
rect 7156 28908 7162 28920
rect 7285 28917 7297 28920
rect 7331 28917 7343 28951
rect 7285 28911 7343 28917
rect 8202 28908 8208 28960
rect 8260 28948 8266 28960
rect 8665 28951 8723 28957
rect 8665 28948 8677 28951
rect 8260 28920 8677 28948
rect 8260 28908 8266 28920
rect 8665 28917 8677 28920
rect 8711 28917 8723 28951
rect 8665 28911 8723 28917
rect 9214 28908 9220 28960
rect 9272 28908 9278 28960
rect 9858 28908 9864 28960
rect 9916 28948 9922 28960
rect 10137 28951 10195 28957
rect 10137 28948 10149 28951
rect 9916 28920 10149 28948
rect 9916 28908 9922 28920
rect 10137 28917 10149 28920
rect 10183 28917 10195 28951
rect 10137 28911 10195 28917
rect 10229 28951 10287 28957
rect 10229 28917 10241 28951
rect 10275 28948 10287 28951
rect 10686 28948 10692 28960
rect 10275 28920 10692 28948
rect 10275 28917 10287 28920
rect 10229 28911 10287 28917
rect 10686 28908 10692 28920
rect 10744 28908 10750 28960
rect 10778 28908 10784 28960
rect 10836 28948 10842 28960
rect 10965 28951 11023 28957
rect 10965 28948 10977 28951
rect 10836 28920 10977 28948
rect 10836 28908 10842 28920
rect 10965 28917 10977 28920
rect 11011 28917 11023 28951
rect 10965 28911 11023 28917
rect 11514 28908 11520 28960
rect 11572 28908 11578 28960
rect 11974 28908 11980 28960
rect 12032 28908 12038 28960
rect 12529 28951 12587 28957
rect 12529 28917 12541 28951
rect 12575 28948 12587 28951
rect 12802 28948 12808 28960
rect 12575 28920 12808 28948
rect 12575 28917 12587 28920
rect 12529 28911 12587 28917
rect 12802 28908 12808 28920
rect 12860 28908 12866 28960
rect 15838 28908 15844 28960
rect 15896 28948 15902 28960
rect 18340 28948 18368 28988
rect 15896 28920 18368 28948
rect 15896 28908 15902 28920
rect 18414 28908 18420 28960
rect 18472 28908 18478 28960
rect 18524 28948 18552 28988
rect 30374 28976 30380 28988
rect 30432 28976 30438 29028
rect 19610 28948 19616 28960
rect 18524 28920 19616 28948
rect 19610 28908 19616 28920
rect 19668 28908 19674 28960
rect 19886 28908 19892 28960
rect 19944 28948 19950 28960
rect 20349 28951 20407 28957
rect 20349 28948 20361 28951
rect 19944 28920 20361 28948
rect 19944 28908 19950 28920
rect 20349 28917 20361 28920
rect 20395 28917 20407 28951
rect 20349 28911 20407 28917
rect 23661 28951 23719 28957
rect 23661 28917 23673 28951
rect 23707 28948 23719 28951
rect 23750 28948 23756 28960
rect 23707 28920 23756 28948
rect 23707 28917 23719 28920
rect 23661 28911 23719 28917
rect 23750 28908 23756 28920
rect 23808 28908 23814 28960
rect 1104 28858 32844 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 32844 28858
rect 1104 28784 32844 28806
rect 2866 28704 2872 28756
rect 2924 28744 2930 28756
rect 2961 28747 3019 28753
rect 2961 28744 2973 28747
rect 2924 28716 2973 28744
rect 2924 28704 2930 28716
rect 2961 28713 2973 28716
rect 3007 28713 3019 28747
rect 2961 28707 3019 28713
rect 3973 28747 4031 28753
rect 3973 28713 3985 28747
rect 4019 28744 4031 28747
rect 4062 28744 4068 28756
rect 4019 28716 4068 28744
rect 4019 28713 4031 28716
rect 3973 28707 4031 28713
rect 4062 28704 4068 28716
rect 4120 28704 4126 28756
rect 4338 28704 4344 28756
rect 4396 28744 4402 28756
rect 4890 28744 4896 28756
rect 4396 28716 4896 28744
rect 4396 28704 4402 28716
rect 4890 28704 4896 28716
rect 4948 28744 4954 28756
rect 5810 28744 5816 28756
rect 4948 28716 5816 28744
rect 4948 28704 4954 28716
rect 5810 28704 5816 28716
rect 5868 28704 5874 28756
rect 6089 28747 6147 28753
rect 6089 28713 6101 28747
rect 6135 28744 6147 28747
rect 8018 28744 8024 28756
rect 6135 28716 8024 28744
rect 6135 28713 6147 28716
rect 6089 28707 6147 28713
rect 8018 28704 8024 28716
rect 8076 28704 8082 28756
rect 10410 28744 10416 28756
rect 8128 28716 10416 28744
rect 2777 28679 2835 28685
rect 2777 28645 2789 28679
rect 2823 28676 2835 28679
rect 4614 28676 4620 28688
rect 2823 28648 4620 28676
rect 2823 28645 2835 28648
rect 2777 28639 2835 28645
rect 4614 28636 4620 28648
rect 4672 28636 4678 28688
rect 5350 28636 5356 28688
rect 5408 28636 5414 28688
rect 3142 28568 3148 28620
rect 3200 28568 3206 28620
rect 4798 28568 4804 28620
rect 4856 28608 4862 28620
rect 4893 28611 4951 28617
rect 4893 28608 4905 28611
rect 4856 28580 4905 28608
rect 4856 28568 4862 28580
rect 4893 28577 4905 28580
rect 4939 28608 4951 28611
rect 4982 28608 4988 28620
rect 4939 28580 4988 28608
rect 4939 28577 4951 28580
rect 4893 28571 4951 28577
rect 4982 28568 4988 28580
rect 5040 28568 5046 28620
rect 5721 28611 5779 28617
rect 5721 28577 5733 28611
rect 5767 28577 5779 28611
rect 5721 28571 5779 28577
rect 1394 28500 1400 28552
rect 1452 28500 1458 28552
rect 1670 28549 1676 28552
rect 1664 28540 1676 28549
rect 1631 28512 1676 28540
rect 1664 28503 1676 28512
rect 1670 28500 1676 28503
rect 1728 28500 1734 28552
rect 2498 28500 2504 28552
rect 2556 28540 2562 28552
rect 3326 28540 3332 28552
rect 2556 28512 3332 28540
rect 2556 28500 2562 28512
rect 3326 28500 3332 28512
rect 3384 28500 3390 28552
rect 3789 28543 3847 28549
rect 3789 28509 3801 28543
rect 3835 28509 3847 28543
rect 3789 28503 3847 28509
rect 2869 28475 2927 28481
rect 2869 28441 2881 28475
rect 2915 28472 2927 28475
rect 2958 28472 2964 28484
rect 2915 28444 2964 28472
rect 2915 28441 2927 28444
rect 2869 28435 2927 28441
rect 2958 28432 2964 28444
rect 3016 28432 3022 28484
rect 3694 28472 3700 28484
rect 3252 28444 3700 28472
rect 2314 28364 2320 28416
rect 2372 28404 2378 28416
rect 2682 28404 2688 28416
rect 2372 28376 2688 28404
rect 2372 28364 2378 28376
rect 2682 28364 2688 28376
rect 2740 28404 2746 28416
rect 3252 28404 3280 28444
rect 3694 28432 3700 28444
rect 3752 28472 3758 28484
rect 3804 28472 3832 28503
rect 4246 28500 4252 28552
rect 4304 28500 4310 28552
rect 4338 28500 4344 28552
rect 4396 28500 4402 28552
rect 5629 28543 5687 28549
rect 5629 28540 5641 28543
rect 4448 28512 5641 28540
rect 3752 28444 3832 28472
rect 3752 28432 3758 28444
rect 2740 28376 3280 28404
rect 2740 28364 2746 28376
rect 3326 28364 3332 28416
rect 3384 28404 3390 28416
rect 3513 28407 3571 28413
rect 3513 28404 3525 28407
rect 3384 28376 3525 28404
rect 3384 28364 3390 28376
rect 3513 28373 3525 28376
rect 3559 28373 3571 28407
rect 3513 28367 3571 28373
rect 4062 28364 4068 28416
rect 4120 28404 4126 28416
rect 4448 28404 4476 28512
rect 5629 28509 5641 28512
rect 5675 28509 5687 28543
rect 5736 28540 5764 28571
rect 5810 28568 5816 28620
rect 5868 28568 5874 28620
rect 5902 28568 5908 28620
rect 5960 28568 5966 28620
rect 6638 28568 6644 28620
rect 6696 28608 6702 28620
rect 8128 28608 8156 28716
rect 10410 28704 10416 28716
rect 10468 28704 10474 28756
rect 10778 28704 10784 28756
rect 10836 28744 10842 28756
rect 12434 28744 12440 28756
rect 10836 28716 12440 28744
rect 10836 28704 10842 28716
rect 12434 28704 12440 28716
rect 12492 28704 12498 28756
rect 12526 28704 12532 28756
rect 12584 28704 12590 28756
rect 12710 28704 12716 28756
rect 12768 28744 12774 28756
rect 13541 28747 13599 28753
rect 13541 28744 13553 28747
rect 12768 28716 13553 28744
rect 12768 28704 12774 28716
rect 8481 28679 8539 28685
rect 8481 28645 8493 28679
rect 8527 28676 8539 28679
rect 8570 28676 8576 28688
rect 8527 28648 8576 28676
rect 8527 28645 8539 28648
rect 8481 28639 8539 28645
rect 8570 28636 8576 28648
rect 8628 28676 8634 28688
rect 9493 28679 9551 28685
rect 8628 28648 9352 28676
rect 8628 28636 8634 28648
rect 9214 28608 9220 28620
rect 6696 28580 8156 28608
rect 8588 28580 9220 28608
rect 6696 28568 6702 28580
rect 5994 28540 6000 28552
rect 5736 28512 6000 28540
rect 5629 28503 5687 28509
rect 5353 28475 5411 28481
rect 5353 28472 5365 28475
rect 4540 28444 5365 28472
rect 4540 28416 4568 28444
rect 5353 28441 5365 28444
rect 5399 28441 5411 28475
rect 5353 28435 5411 28441
rect 4120 28376 4476 28404
rect 4120 28364 4126 28376
rect 4522 28364 4528 28416
rect 4580 28364 4586 28416
rect 4614 28364 4620 28416
rect 4672 28364 4678 28416
rect 4801 28407 4859 28413
rect 4801 28373 4813 28407
rect 4847 28404 4859 28407
rect 5644 28404 5672 28503
rect 5994 28500 6000 28512
rect 6052 28500 6058 28552
rect 6730 28500 6736 28552
rect 6788 28540 6794 28552
rect 6825 28543 6883 28549
rect 6825 28540 6837 28543
rect 6788 28512 6837 28540
rect 6788 28500 6794 28512
rect 6825 28509 6837 28512
rect 6871 28509 6883 28543
rect 6825 28503 6883 28509
rect 6917 28543 6975 28549
rect 6917 28509 6929 28543
rect 6963 28540 6975 28543
rect 7098 28540 7104 28552
rect 6963 28512 7104 28540
rect 6963 28509 6975 28512
rect 6917 28503 6975 28509
rect 7098 28500 7104 28512
rect 7156 28500 7162 28552
rect 7190 28500 7196 28552
rect 7248 28500 7254 28552
rect 7653 28543 7711 28549
rect 7653 28540 7665 28543
rect 7300 28512 7665 28540
rect 5718 28432 5724 28484
rect 5776 28472 5782 28484
rect 7300 28472 7328 28512
rect 7653 28509 7665 28512
rect 7699 28509 7711 28543
rect 7653 28503 7711 28509
rect 8021 28543 8079 28549
rect 8021 28509 8033 28543
rect 8067 28540 8079 28543
rect 8202 28540 8208 28552
rect 8067 28512 8208 28540
rect 8067 28509 8079 28512
rect 8021 28503 8079 28509
rect 8202 28500 8208 28512
rect 8260 28500 8266 28552
rect 8294 28500 8300 28552
rect 8352 28500 8358 28552
rect 8588 28549 8616 28580
rect 9214 28568 9220 28580
rect 9272 28568 9278 28620
rect 8573 28543 8631 28549
rect 8573 28509 8585 28543
rect 8619 28509 8631 28543
rect 8573 28503 8631 28509
rect 8754 28500 8760 28552
rect 8812 28540 8818 28552
rect 9324 28549 9352 28648
rect 9493 28645 9505 28679
rect 9539 28676 9551 28679
rect 11146 28676 11152 28688
rect 9539 28648 11152 28676
rect 9539 28645 9551 28648
rect 9493 28639 9551 28645
rect 11146 28636 11152 28648
rect 11204 28636 11210 28688
rect 11882 28636 11888 28688
rect 11940 28636 11946 28688
rect 12066 28636 12072 28688
rect 12124 28676 12130 28688
rect 12124 28648 12848 28676
rect 12124 28636 12130 28648
rect 12710 28608 12716 28620
rect 10244 28580 11560 28608
rect 8941 28543 8999 28549
rect 8941 28540 8953 28543
rect 8812 28512 8953 28540
rect 8812 28500 8818 28512
rect 8941 28509 8953 28512
rect 8987 28509 8999 28543
rect 9324 28543 9391 28549
rect 9324 28512 9345 28543
rect 8941 28503 8999 28509
rect 9333 28509 9345 28512
rect 9379 28509 9391 28543
rect 9333 28503 9391 28509
rect 9766 28500 9772 28552
rect 9824 28500 9830 28552
rect 10244 28549 10272 28580
rect 11532 28552 11560 28580
rect 11716 28580 12388 28608
rect 10229 28543 10287 28549
rect 10229 28509 10241 28543
rect 10275 28509 10287 28543
rect 10229 28503 10287 28509
rect 10502 28500 10508 28552
rect 10560 28500 10566 28552
rect 10778 28500 10784 28552
rect 10836 28500 10842 28552
rect 10870 28500 10876 28552
rect 10928 28500 10934 28552
rect 11333 28543 11391 28549
rect 11333 28509 11345 28543
rect 11379 28540 11391 28543
rect 11422 28540 11428 28552
rect 11379 28512 11428 28540
rect 11379 28509 11391 28512
rect 11333 28503 11391 28509
rect 11422 28500 11428 28512
rect 11480 28500 11486 28552
rect 11514 28500 11520 28552
rect 11572 28500 11578 28552
rect 11716 28549 11744 28580
rect 12360 28552 12388 28580
rect 12636 28580 12716 28608
rect 11701 28543 11759 28549
rect 11701 28509 11713 28543
rect 11747 28509 11759 28543
rect 11701 28503 11759 28509
rect 11974 28500 11980 28552
rect 12032 28500 12038 28552
rect 12342 28500 12348 28552
rect 12400 28500 12406 28552
rect 12636 28549 12664 28580
rect 12710 28568 12716 28580
rect 12768 28568 12774 28620
rect 12820 28549 12848 28648
rect 13170 28636 13176 28688
rect 13228 28676 13234 28688
rect 13265 28679 13323 28685
rect 13265 28676 13277 28679
rect 13228 28648 13277 28676
rect 13228 28636 13234 28648
rect 13265 28645 13277 28648
rect 13311 28645 13323 28679
rect 13265 28639 13323 28645
rect 12621 28543 12679 28549
rect 12621 28509 12633 28543
rect 12667 28509 12679 28543
rect 12621 28503 12679 28509
rect 12805 28543 12863 28549
rect 12805 28509 12817 28543
rect 12851 28509 12863 28543
rect 12805 28503 12863 28509
rect 12894 28500 12900 28552
rect 12952 28500 12958 28552
rect 12986 28500 12992 28552
rect 13044 28500 13050 28552
rect 13464 28549 13492 28716
rect 13541 28713 13553 28716
rect 13587 28713 13599 28747
rect 13541 28707 13599 28713
rect 16022 28704 16028 28756
rect 16080 28744 16086 28756
rect 16485 28747 16543 28753
rect 16485 28744 16497 28747
rect 16080 28716 16497 28744
rect 16080 28704 16086 28716
rect 16485 28713 16497 28716
rect 16531 28744 16543 28747
rect 17310 28744 17316 28756
rect 16531 28716 17316 28744
rect 16531 28713 16543 28716
rect 16485 28707 16543 28713
rect 17310 28704 17316 28716
rect 17368 28744 17374 28756
rect 19426 28744 19432 28756
rect 17368 28716 19432 28744
rect 17368 28704 17374 28716
rect 19426 28704 19432 28716
rect 19484 28704 19490 28756
rect 19886 28704 19892 28756
rect 19944 28704 19950 28756
rect 19978 28704 19984 28756
rect 20036 28744 20042 28756
rect 23201 28747 23259 28753
rect 23201 28744 23213 28747
rect 20036 28716 23213 28744
rect 20036 28704 20042 28716
rect 23201 28713 23213 28716
rect 23247 28713 23259 28747
rect 23201 28707 23259 28713
rect 23753 28747 23811 28753
rect 23753 28713 23765 28747
rect 23799 28713 23811 28747
rect 23753 28707 23811 28713
rect 13906 28636 13912 28688
rect 13964 28676 13970 28688
rect 14369 28679 14427 28685
rect 14369 28676 14381 28679
rect 13964 28648 14381 28676
rect 13964 28636 13970 28648
rect 14369 28645 14381 28648
rect 14415 28645 14427 28679
rect 14369 28639 14427 28645
rect 17954 28636 17960 28688
rect 18012 28676 18018 28688
rect 18012 28648 18368 28676
rect 18012 28636 18018 28648
rect 13538 28568 13544 28620
rect 13596 28608 13602 28620
rect 18230 28608 18236 28620
rect 13596 28580 18236 28608
rect 13596 28568 13602 28580
rect 18230 28568 18236 28580
rect 18288 28568 18294 28620
rect 13449 28543 13507 28549
rect 13449 28509 13461 28543
rect 13495 28509 13507 28543
rect 13449 28503 13507 28509
rect 13725 28543 13783 28549
rect 13725 28509 13737 28543
rect 13771 28509 13783 28543
rect 14274 28540 14280 28552
rect 13725 28503 13783 28509
rect 14200 28512 14280 28540
rect 5776 28444 7328 28472
rect 9125 28475 9183 28481
rect 5776 28432 5782 28444
rect 9125 28441 9137 28475
rect 9171 28441 9183 28475
rect 9125 28435 9183 28441
rect 9217 28475 9275 28481
rect 9217 28441 9229 28475
rect 9263 28472 9275 28475
rect 9263 28444 9444 28472
rect 9263 28441 9275 28444
rect 9217 28435 9275 28441
rect 4847 28376 5672 28404
rect 4847 28373 4859 28376
rect 4801 28367 4859 28373
rect 6638 28364 6644 28416
rect 6696 28364 6702 28416
rect 7101 28407 7159 28413
rect 7101 28373 7113 28407
rect 7147 28404 7159 28407
rect 7190 28404 7196 28416
rect 7147 28376 7196 28404
rect 7147 28373 7159 28376
rect 7101 28367 7159 28373
rect 7190 28364 7196 28376
rect 7248 28364 7254 28416
rect 7377 28407 7435 28413
rect 7377 28373 7389 28407
rect 7423 28404 7435 28407
rect 7466 28404 7472 28416
rect 7423 28376 7472 28404
rect 7423 28373 7435 28376
rect 7377 28367 7435 28373
rect 7466 28364 7472 28376
rect 7524 28364 7530 28416
rect 7742 28364 7748 28416
rect 7800 28404 7806 28416
rect 7837 28407 7895 28413
rect 7837 28404 7849 28407
rect 7800 28376 7849 28404
rect 7800 28364 7806 28376
rect 7837 28373 7849 28376
rect 7883 28373 7895 28407
rect 7837 28367 7895 28373
rect 8205 28407 8263 28413
rect 8205 28373 8217 28407
rect 8251 28404 8263 28407
rect 8294 28404 8300 28416
rect 8251 28376 8300 28404
rect 8251 28373 8263 28376
rect 8205 28367 8263 28373
rect 8294 28364 8300 28376
rect 8352 28364 8358 28416
rect 8757 28407 8815 28413
rect 8757 28373 8769 28407
rect 8803 28404 8815 28407
rect 9030 28404 9036 28416
rect 8803 28376 9036 28404
rect 8803 28373 8815 28376
rect 8757 28367 8815 28373
rect 9030 28364 9036 28376
rect 9088 28404 9094 28416
rect 9140 28404 9168 28435
rect 9416 28416 9444 28444
rect 9582 28432 9588 28484
rect 9640 28472 9646 28484
rect 10134 28472 10140 28484
rect 9640 28444 10140 28472
rect 9640 28432 9646 28444
rect 10134 28432 10140 28444
rect 10192 28432 10198 28484
rect 10689 28475 10747 28481
rect 10689 28441 10701 28475
rect 10735 28472 10747 28475
rect 10735 28444 11560 28472
rect 10735 28441 10747 28444
rect 10689 28435 10747 28441
rect 9088 28376 9168 28404
rect 9088 28364 9094 28376
rect 9398 28364 9404 28416
rect 9456 28364 9462 28416
rect 9950 28364 9956 28416
rect 10008 28364 10014 28416
rect 10413 28407 10471 28413
rect 10413 28373 10425 28407
rect 10459 28404 10471 28407
rect 10704 28404 10732 28435
rect 10459 28376 10732 28404
rect 10459 28373 10471 28376
rect 10413 28367 10471 28373
rect 11054 28364 11060 28416
rect 11112 28364 11118 28416
rect 11532 28404 11560 28444
rect 11606 28432 11612 28484
rect 11664 28472 11670 28484
rect 11992 28472 12020 28500
rect 11664 28444 12020 28472
rect 12161 28475 12219 28481
rect 11664 28432 11670 28444
rect 12161 28441 12173 28475
rect 12207 28441 12219 28475
rect 12161 28435 12219 28441
rect 12253 28475 12311 28481
rect 12253 28441 12265 28475
rect 12299 28472 12311 28475
rect 12526 28472 12532 28484
rect 12299 28444 12532 28472
rect 12299 28441 12311 28444
rect 12253 28435 12311 28441
rect 11974 28404 11980 28416
rect 11532 28376 11980 28404
rect 11974 28364 11980 28376
rect 12032 28404 12038 28416
rect 12176 28404 12204 28435
rect 12526 28432 12532 28444
rect 12584 28432 12590 28484
rect 13740 28472 13768 28503
rect 14200 28472 14228 28512
rect 14274 28500 14280 28512
rect 14332 28500 14338 28552
rect 14550 28500 14556 28552
rect 14608 28540 14614 28552
rect 15286 28540 15292 28552
rect 14608 28512 15292 28540
rect 14608 28500 14614 28512
rect 15286 28500 15292 28512
rect 15344 28500 15350 28552
rect 16301 28543 16359 28549
rect 15764 28512 16252 28540
rect 15764 28472 15792 28512
rect 12820 28444 13768 28472
rect 14016 28444 14228 28472
rect 14292 28444 15792 28472
rect 12032 28376 12204 28404
rect 12032 28364 12038 28376
rect 12434 28364 12440 28416
rect 12492 28404 12498 28416
rect 12820 28404 12848 28444
rect 12492 28376 12848 28404
rect 13173 28407 13231 28413
rect 12492 28364 12498 28376
rect 13173 28373 13185 28407
rect 13219 28404 13231 28407
rect 14016 28404 14044 28444
rect 13219 28376 14044 28404
rect 13219 28373 13231 28376
rect 13173 28367 13231 28373
rect 14090 28364 14096 28416
rect 14148 28404 14154 28416
rect 14292 28404 14320 28444
rect 15838 28432 15844 28484
rect 15896 28432 15902 28484
rect 16022 28432 16028 28484
rect 16080 28432 16086 28484
rect 16224 28472 16252 28512
rect 16301 28509 16313 28543
rect 16347 28540 16359 28543
rect 16390 28540 16396 28552
rect 16347 28512 16396 28540
rect 16347 28509 16359 28512
rect 16301 28503 16359 28509
rect 16390 28500 16396 28512
rect 16448 28500 16454 28552
rect 17957 28543 18015 28549
rect 16592 28512 17908 28540
rect 16592 28472 16620 28512
rect 16224 28444 16620 28472
rect 17310 28432 17316 28484
rect 17368 28432 17374 28484
rect 17497 28475 17555 28481
rect 17497 28441 17509 28475
rect 17543 28472 17555 28475
rect 17880 28472 17908 28512
rect 17957 28509 17969 28543
rect 18003 28540 18015 28543
rect 18046 28540 18052 28552
rect 18003 28512 18052 28540
rect 18003 28509 18015 28512
rect 17957 28503 18015 28509
rect 18046 28500 18052 28512
rect 18104 28500 18110 28552
rect 18340 28549 18368 28648
rect 18414 28636 18420 28688
rect 18472 28676 18478 28688
rect 19334 28676 19340 28688
rect 18472 28648 19340 28676
rect 18472 28636 18478 28648
rect 19334 28636 19340 28648
rect 19392 28636 19398 28688
rect 19720 28648 20300 28676
rect 18325 28543 18383 28549
rect 18325 28509 18337 28543
rect 18371 28509 18383 28543
rect 18325 28503 18383 28509
rect 18414 28500 18420 28552
rect 18472 28540 18478 28552
rect 19720 28540 19748 28648
rect 19889 28611 19947 28617
rect 19889 28577 19901 28611
rect 19935 28608 19947 28611
rect 20162 28608 20168 28620
rect 19935 28580 20168 28608
rect 19935 28577 19947 28580
rect 19889 28571 19947 28577
rect 20162 28568 20168 28580
rect 20220 28568 20226 28620
rect 20272 28617 20300 28648
rect 20346 28636 20352 28688
rect 20404 28676 20410 28688
rect 23768 28676 23796 28707
rect 20404 28648 23796 28676
rect 20404 28636 20410 28648
rect 20257 28611 20315 28617
rect 20257 28577 20269 28611
rect 20303 28577 20315 28611
rect 20257 28571 20315 28577
rect 21726 28568 21732 28620
rect 21784 28608 21790 28620
rect 21784 28580 23980 28608
rect 21784 28568 21790 28580
rect 18472 28512 19748 28540
rect 19997 28543 20055 28549
rect 18472 28500 18478 28512
rect 19997 28509 20009 28543
rect 20043 28540 20055 28543
rect 20530 28540 20536 28552
rect 20043 28512 20536 28540
rect 20043 28509 20055 28512
rect 19997 28503 20055 28509
rect 20530 28500 20536 28512
rect 20588 28500 20594 28552
rect 23198 28500 23204 28552
rect 23256 28500 23262 28552
rect 23382 28500 23388 28552
rect 23440 28500 23446 28552
rect 23750 28500 23756 28552
rect 23808 28500 23814 28552
rect 23952 28549 23980 28580
rect 23937 28543 23995 28549
rect 23937 28509 23949 28543
rect 23983 28540 23995 28543
rect 24486 28540 24492 28552
rect 23983 28512 24492 28540
rect 23983 28509 23995 28512
rect 23937 28503 23995 28509
rect 24486 28500 24492 28512
rect 24544 28500 24550 28552
rect 18141 28475 18199 28481
rect 18141 28472 18153 28475
rect 17543 28444 17816 28472
rect 17880 28444 18153 28472
rect 17543 28441 17555 28444
rect 17497 28435 17555 28441
rect 14148 28376 14320 28404
rect 14148 28364 14154 28376
rect 14458 28364 14464 28416
rect 14516 28404 14522 28416
rect 15010 28404 15016 28416
rect 14516 28376 15016 28404
rect 14516 28364 14522 28376
rect 15010 28364 15016 28376
rect 15068 28364 15074 28416
rect 16206 28364 16212 28416
rect 16264 28364 16270 28416
rect 17678 28364 17684 28416
rect 17736 28364 17742 28416
rect 17788 28413 17816 28444
rect 18141 28441 18153 28444
rect 18187 28472 18199 28475
rect 18230 28472 18236 28484
rect 18187 28444 18236 28472
rect 18187 28441 18199 28444
rect 18141 28435 18199 28441
rect 18230 28432 18236 28444
rect 18288 28432 18294 28484
rect 19705 28475 19763 28481
rect 19705 28472 19717 28475
rect 18432 28444 19717 28472
rect 17773 28407 17831 28413
rect 17773 28373 17785 28407
rect 17819 28404 17831 28407
rect 18432 28404 18460 28444
rect 19705 28441 19717 28444
rect 19751 28472 19763 28475
rect 23400 28472 23428 28500
rect 19751 28444 23428 28472
rect 19751 28441 19763 28444
rect 19705 28435 19763 28441
rect 23474 28432 23480 28484
rect 23532 28472 23538 28484
rect 29086 28472 29092 28484
rect 23532 28444 29092 28472
rect 23532 28432 23538 28444
rect 29086 28432 29092 28444
rect 29144 28432 29150 28484
rect 17819 28376 18460 28404
rect 18509 28407 18567 28413
rect 17819 28373 17831 28376
rect 17773 28367 17831 28373
rect 18509 28373 18521 28407
rect 18555 28404 18567 28407
rect 18966 28404 18972 28416
rect 18555 28376 18972 28404
rect 18555 28373 18567 28376
rect 18509 28367 18567 28373
rect 18966 28364 18972 28376
rect 19024 28364 19030 28416
rect 19426 28364 19432 28416
rect 19484 28404 19490 28416
rect 19978 28404 19984 28416
rect 19484 28376 19984 28404
rect 19484 28364 19490 28376
rect 19978 28364 19984 28376
rect 20036 28364 20042 28416
rect 20162 28364 20168 28416
rect 20220 28364 20226 28416
rect 23566 28364 23572 28416
rect 23624 28364 23630 28416
rect 23934 28364 23940 28416
rect 23992 28404 23998 28416
rect 24121 28407 24179 28413
rect 24121 28404 24133 28407
rect 23992 28376 24133 28404
rect 23992 28364 23998 28376
rect 24121 28373 24133 28376
rect 24167 28373 24179 28407
rect 24121 28367 24179 28373
rect 1104 28314 32844 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 32844 28314
rect 1104 28240 32844 28262
rect 2777 28203 2835 28209
rect 2777 28169 2789 28203
rect 2823 28200 2835 28203
rect 3234 28200 3240 28212
rect 2823 28172 3240 28200
rect 2823 28169 2835 28172
rect 2777 28163 2835 28169
rect 3234 28160 3240 28172
rect 3292 28160 3298 28212
rect 5350 28160 5356 28212
rect 5408 28200 5414 28212
rect 5997 28203 6055 28209
rect 5997 28200 6009 28203
rect 5408 28172 6009 28200
rect 5408 28160 5414 28172
rect 3326 28092 3332 28144
rect 3384 28132 3390 28144
rect 3786 28132 3792 28144
rect 3384 28104 3792 28132
rect 3384 28092 3390 28104
rect 3786 28092 3792 28104
rect 3844 28092 3850 28144
rect 3973 28135 4031 28141
rect 3973 28101 3985 28135
rect 4019 28132 4031 28135
rect 4338 28132 4344 28144
rect 4019 28104 4344 28132
rect 4019 28101 4031 28104
rect 3973 28095 4031 28101
rect 4338 28092 4344 28104
rect 4396 28092 4402 28144
rect 4433 28135 4491 28141
rect 4433 28101 4445 28135
rect 4479 28132 4491 28135
rect 4798 28132 4804 28144
rect 4479 28104 4804 28132
rect 4479 28101 4491 28104
rect 4433 28095 4491 28101
rect 4798 28092 4804 28104
rect 4856 28132 4862 28144
rect 4893 28135 4951 28141
rect 4893 28132 4905 28135
rect 4856 28104 4905 28132
rect 4856 28092 4862 28104
rect 4893 28101 4905 28104
rect 4939 28101 4951 28135
rect 4893 28095 4951 28101
rect 1670 28073 1676 28076
rect 1664 28027 1676 28073
rect 1670 28024 1676 28027
rect 1728 28024 1734 28076
rect 3142 28024 3148 28076
rect 3200 28064 3206 28076
rect 3538 28067 3596 28073
rect 3538 28064 3550 28067
rect 3200 28036 3550 28064
rect 3200 28024 3206 28036
rect 3538 28033 3550 28036
rect 3584 28033 3596 28067
rect 3538 28027 3596 28033
rect 4246 28024 4252 28076
rect 4304 28064 4310 28076
rect 5442 28064 5448 28076
rect 4304 28036 5448 28064
rect 4304 28024 4310 28036
rect 5442 28024 5448 28036
rect 5500 28024 5506 28076
rect 5736 28073 5764 28172
rect 5997 28169 6009 28172
rect 6043 28169 6055 28203
rect 5997 28163 6055 28169
rect 6638 28160 6644 28212
rect 6696 28160 6702 28212
rect 7190 28200 7196 28212
rect 6748 28172 7196 28200
rect 6656 28132 6684 28160
rect 6564 28104 6684 28132
rect 5721 28067 5779 28073
rect 5721 28033 5733 28067
rect 5767 28033 5779 28067
rect 5721 28027 5779 28033
rect 6178 28024 6184 28076
rect 6236 28024 6242 28076
rect 6365 28067 6423 28073
rect 6365 28033 6377 28067
rect 6411 28064 6423 28067
rect 6454 28064 6460 28076
rect 6411 28036 6460 28064
rect 6411 28033 6423 28036
rect 6365 28027 6423 28033
rect 6454 28024 6460 28036
rect 6512 28024 6518 28076
rect 6564 28073 6592 28104
rect 6549 28067 6607 28073
rect 6549 28033 6561 28067
rect 6595 28033 6607 28067
rect 6549 28027 6607 28033
rect 6638 28024 6644 28076
rect 6696 28024 6702 28076
rect 6748 28073 6776 28172
rect 7190 28160 7196 28172
rect 7248 28160 7254 28212
rect 8205 28203 8263 28209
rect 8205 28169 8217 28203
rect 8251 28200 8263 28203
rect 8386 28200 8392 28212
rect 8251 28172 8392 28200
rect 8251 28169 8263 28172
rect 8205 28163 8263 28169
rect 8386 28160 8392 28172
rect 8444 28160 8450 28212
rect 8481 28203 8539 28209
rect 8481 28169 8493 28203
rect 8527 28200 8539 28203
rect 9766 28200 9772 28212
rect 8527 28172 9772 28200
rect 8527 28169 8539 28172
rect 8481 28163 8539 28169
rect 9766 28160 9772 28172
rect 9824 28160 9830 28212
rect 9858 28160 9864 28212
rect 9916 28200 9922 28212
rect 11054 28200 11060 28212
rect 9916 28172 11060 28200
rect 9916 28160 9922 28172
rect 11054 28160 11060 28172
rect 11112 28160 11118 28212
rect 11333 28203 11391 28209
rect 11333 28169 11345 28203
rect 11379 28169 11391 28203
rect 11333 28163 11391 28169
rect 7558 28132 7564 28144
rect 6840 28104 7564 28132
rect 6733 28067 6791 28073
rect 6733 28033 6745 28067
rect 6779 28033 6791 28067
rect 6733 28027 6791 28033
rect 1394 27956 1400 28008
rect 1452 27956 1458 28008
rect 2958 27956 2964 28008
rect 3016 27996 3022 28008
rect 3053 27999 3111 28005
rect 3053 27996 3065 27999
rect 3016 27968 3065 27996
rect 3016 27956 3022 27968
rect 3053 27965 3065 27968
rect 3099 27965 3111 27999
rect 3053 27959 3111 27965
rect 3234 27956 3240 28008
rect 3292 27996 3298 28008
rect 3421 27999 3479 28005
rect 3421 27996 3433 27999
rect 3292 27968 3433 27996
rect 3292 27956 3298 27968
rect 3421 27965 3433 27968
rect 3467 27965 3479 27999
rect 3421 27959 3479 27965
rect 4525 27999 4583 28005
rect 4525 27965 4537 27999
rect 4571 27996 4583 27999
rect 5629 27999 5687 28005
rect 4571 27968 5028 27996
rect 4571 27965 4583 27968
rect 4525 27959 4583 27965
rect 5000 27940 5028 27968
rect 5629 27965 5641 27999
rect 5675 27996 5687 27999
rect 6840 27996 6868 28104
rect 7558 28092 7564 28104
rect 7616 28092 7622 28144
rect 8662 28132 8668 28144
rect 8312 28104 8668 28132
rect 7009 28067 7067 28073
rect 7009 28033 7021 28067
rect 7055 28033 7067 28067
rect 7009 28027 7067 28033
rect 5675 27968 6224 27996
rect 5675 27965 5687 27968
rect 5629 27959 5687 27965
rect 3973 27931 4031 27937
rect 3973 27897 3985 27931
rect 4019 27928 4031 27931
rect 4062 27928 4068 27940
rect 4019 27900 4068 27928
rect 4019 27897 4031 27900
rect 3973 27891 4031 27897
rect 4062 27888 4068 27900
rect 4120 27888 4126 27940
rect 4614 27888 4620 27940
rect 4672 27928 4678 27940
rect 4893 27931 4951 27937
rect 4893 27928 4905 27931
rect 4672 27900 4905 27928
rect 4672 27888 4678 27900
rect 4893 27897 4905 27900
rect 4939 27897 4951 27931
rect 4893 27891 4951 27897
rect 4982 27888 4988 27940
rect 5040 27928 5046 27940
rect 5905 27931 5963 27937
rect 5905 27928 5917 27931
rect 5040 27900 5917 27928
rect 5040 27888 5046 27900
rect 5905 27897 5917 27900
rect 5951 27928 5963 27931
rect 5994 27928 6000 27940
rect 5951 27900 6000 27928
rect 5951 27897 5963 27900
rect 5905 27891 5963 27897
rect 5994 27888 6000 27900
rect 6052 27888 6058 27940
rect 6196 27928 6224 27968
rect 6656 27968 6868 27996
rect 6656 27928 6684 27968
rect 6196 27900 6684 27928
rect 7024 27928 7052 28027
rect 7190 28024 7196 28076
rect 7248 28024 7254 28076
rect 7466 28024 7472 28076
rect 7524 28024 7530 28076
rect 7742 28024 7748 28076
rect 7800 28024 7806 28076
rect 8018 28024 8024 28076
rect 8076 28024 8082 28076
rect 8312 28073 8340 28104
rect 8662 28092 8668 28104
rect 8720 28092 8726 28144
rect 8754 28092 8760 28144
rect 8812 28092 8818 28144
rect 8849 28135 8907 28141
rect 8849 28101 8861 28135
rect 8895 28132 8907 28135
rect 9398 28132 9404 28144
rect 8895 28104 9404 28132
rect 8895 28101 8907 28104
rect 8849 28095 8907 28101
rect 9398 28092 9404 28104
rect 9456 28092 9462 28144
rect 9582 28092 9588 28144
rect 9640 28132 9646 28144
rect 11238 28132 11244 28144
rect 9640 28104 10180 28132
rect 9640 28092 9646 28104
rect 8297 28067 8355 28073
rect 8297 28033 8309 28067
rect 8343 28033 8355 28067
rect 8297 28027 8355 28033
rect 8570 28024 8576 28076
rect 8628 28024 8634 28076
rect 8941 28067 8999 28073
rect 8941 28033 8953 28067
rect 8987 28064 8999 28067
rect 9030 28064 9036 28076
rect 8987 28036 9036 28064
rect 8987 28033 8999 28036
rect 8941 28027 8999 28033
rect 9030 28024 9036 28036
rect 9088 28024 9094 28076
rect 9490 28024 9496 28076
rect 9548 28024 9554 28076
rect 9769 28067 9827 28073
rect 9769 28033 9781 28067
rect 9815 28064 9827 28067
rect 9858 28064 9864 28076
rect 9815 28036 9864 28064
rect 9815 28033 9827 28036
rect 9769 28027 9827 28033
rect 9858 28024 9864 28036
rect 9916 28024 9922 28076
rect 10042 28024 10048 28076
rect 10100 28024 10106 28076
rect 10152 28073 10180 28104
rect 10428 28104 11244 28132
rect 10137 28067 10195 28073
rect 10137 28033 10149 28067
rect 10183 28033 10195 28067
rect 10137 28027 10195 28033
rect 10321 28068 10379 28073
rect 10428 28068 10456 28104
rect 11238 28092 11244 28104
rect 11296 28092 11302 28144
rect 10321 28067 10456 28068
rect 10321 28033 10333 28067
rect 10367 28040 10456 28067
rect 10597 28057 10655 28063
rect 10597 28054 10609 28057
rect 10367 28033 10379 28040
rect 10321 28027 10379 28033
rect 10520 28026 10609 28054
rect 7098 27956 7104 28008
rect 7156 27996 7162 28008
rect 7558 27996 7564 28008
rect 7156 27968 7564 27996
rect 7156 27956 7162 27968
rect 7558 27956 7564 27968
rect 7616 27956 7622 28008
rect 7653 27999 7711 28005
rect 7653 27965 7665 27999
rect 7699 27996 7711 27999
rect 10226 27996 10232 28008
rect 7699 27968 10232 27996
rect 7699 27965 7711 27968
rect 7653 27959 7711 27965
rect 10226 27956 10232 27968
rect 10284 27956 10290 28008
rect 8662 27928 8668 27940
rect 7024 27900 8668 27928
rect 8662 27888 8668 27900
rect 8720 27888 8726 27940
rect 9122 27888 9128 27940
rect 9180 27888 9186 27940
rect 9674 27928 9680 27940
rect 9232 27900 9680 27928
rect 3602 27820 3608 27872
rect 3660 27860 3666 27872
rect 3697 27863 3755 27869
rect 3697 27860 3709 27863
rect 3660 27832 3709 27860
rect 3660 27820 3666 27832
rect 3697 27829 3709 27832
rect 3743 27829 3755 27863
rect 3697 27823 3755 27829
rect 4709 27863 4767 27869
rect 4709 27829 4721 27863
rect 4755 27860 4767 27863
rect 5810 27860 5816 27872
rect 4755 27832 5816 27860
rect 4755 27829 4767 27832
rect 4709 27823 4767 27829
rect 5810 27820 5816 27832
rect 5868 27820 5874 27872
rect 6914 27820 6920 27872
rect 6972 27820 6978 27872
rect 7834 27820 7840 27872
rect 7892 27860 7898 27872
rect 7929 27863 7987 27869
rect 7929 27860 7941 27863
rect 7892 27832 7941 27860
rect 7892 27820 7898 27832
rect 7929 27829 7941 27832
rect 7975 27829 7987 27863
rect 7929 27823 7987 27829
rect 8754 27820 8760 27872
rect 8812 27860 8818 27872
rect 9232 27860 9260 27900
rect 9674 27888 9680 27900
rect 9732 27928 9738 27940
rect 9861 27931 9919 27937
rect 9861 27928 9873 27931
rect 9732 27900 9873 27928
rect 9732 27888 9738 27900
rect 9861 27897 9873 27900
rect 9907 27897 9919 27931
rect 9861 27891 9919 27897
rect 10134 27888 10140 27940
rect 10192 27928 10198 27940
rect 10520 27928 10548 28026
rect 10597 28023 10609 28026
rect 10643 28023 10655 28057
rect 10778 28024 10784 28076
rect 10836 28024 10842 28076
rect 10873 28067 10931 28073
rect 10873 28033 10885 28067
rect 10919 28033 10931 28067
rect 10873 28027 10931 28033
rect 10597 28017 10655 28023
rect 10888 27996 10916 28027
rect 11146 28024 11152 28076
rect 11204 28024 11210 28076
rect 11348 28064 11376 28163
rect 11422 28160 11428 28212
rect 11480 28200 11486 28212
rect 12526 28200 12532 28212
rect 11480 28172 12532 28200
rect 11480 28160 11486 28172
rect 12526 28160 12532 28172
rect 12584 28160 12590 28212
rect 12713 28203 12771 28209
rect 12713 28169 12725 28203
rect 12759 28200 12771 28203
rect 12986 28200 12992 28212
rect 12759 28172 12992 28200
rect 12759 28169 12771 28172
rect 12713 28163 12771 28169
rect 11885 28135 11943 28141
rect 11885 28101 11897 28135
rect 11931 28101 11943 28135
rect 12728 28132 12756 28163
rect 12986 28160 12992 28172
rect 13044 28160 13050 28212
rect 13354 28160 13360 28212
rect 13412 28200 13418 28212
rect 13412 28172 13768 28200
rect 13412 28160 13418 28172
rect 13740 28141 13768 28172
rect 14550 28160 14556 28212
rect 14608 28200 14614 28212
rect 15381 28203 15439 28209
rect 15381 28200 15393 28203
rect 14608 28172 15393 28200
rect 14608 28160 14614 28172
rect 15381 28169 15393 28172
rect 15427 28200 15439 28203
rect 22370 28200 22376 28212
rect 15427 28172 22376 28200
rect 15427 28169 15439 28172
rect 15381 28163 15439 28169
rect 22370 28160 22376 28172
rect 22428 28160 22434 28212
rect 11885 28095 11943 28101
rect 11992 28104 12756 28132
rect 13725 28135 13783 28141
rect 11514 28064 11520 28076
rect 11348 28036 11520 28064
rect 11514 28024 11520 28036
rect 11572 28064 11578 28076
rect 11609 28067 11667 28073
rect 11609 28064 11621 28067
rect 11572 28036 11621 28064
rect 11572 28024 11578 28036
rect 11609 28033 11621 28036
rect 11655 28033 11667 28067
rect 11609 28027 11667 28033
rect 11793 28067 11851 28073
rect 11793 28033 11805 28067
rect 11839 28033 11851 28067
rect 11793 28027 11851 28033
rect 10192 27900 10548 27928
rect 10796 27968 10916 27996
rect 10192 27888 10198 27900
rect 8812 27832 9260 27860
rect 8812 27820 8818 27832
rect 9306 27820 9312 27872
rect 9364 27820 9370 27872
rect 9582 27820 9588 27872
rect 9640 27820 9646 27872
rect 10410 27820 10416 27872
rect 10468 27860 10474 27872
rect 10796 27860 10824 27968
rect 11238 27956 11244 28008
rect 11296 27996 11302 28008
rect 11808 27996 11836 28027
rect 11296 27968 11836 27996
rect 11900 27996 11928 28095
rect 11992 28073 12020 28104
rect 13725 28101 13737 28135
rect 13771 28101 13783 28135
rect 13725 28095 13783 28101
rect 14274 28092 14280 28144
rect 14332 28132 14338 28144
rect 14332 28104 18276 28132
rect 14332 28092 14338 28104
rect 11977 28067 12035 28073
rect 11977 28033 11989 28067
rect 12023 28033 12035 28067
rect 11977 28027 12035 28033
rect 12437 28067 12495 28073
rect 12437 28033 12449 28067
rect 12483 28033 12495 28067
rect 12437 28027 12495 28033
rect 12452 27996 12480 28027
rect 12526 28024 12532 28076
rect 12584 28024 12590 28076
rect 12710 28024 12716 28076
rect 12768 28064 12774 28076
rect 12989 28067 13047 28073
rect 12989 28064 13001 28067
rect 12768 28036 13001 28064
rect 12768 28024 12774 28036
rect 12989 28033 13001 28036
rect 13035 28033 13047 28067
rect 12989 28027 13047 28033
rect 14001 28067 14059 28073
rect 14001 28033 14013 28067
rect 14047 28064 14059 28067
rect 14090 28064 14096 28076
rect 14047 28036 14096 28064
rect 14047 28033 14059 28036
rect 14001 28027 14059 28033
rect 14090 28024 14096 28036
rect 14148 28024 14154 28076
rect 14645 28067 14703 28073
rect 14645 28033 14657 28067
rect 14691 28033 14703 28067
rect 14645 28027 14703 28033
rect 12802 27996 12808 28008
rect 11900 27968 12808 27996
rect 11296 27956 11302 27968
rect 12802 27956 12808 27968
rect 12860 27956 12866 28008
rect 13722 27956 13728 28008
rect 13780 27996 13786 28008
rect 13817 27999 13875 28005
rect 13817 27996 13829 27999
rect 13780 27968 13829 27996
rect 13780 27956 13786 27968
rect 13817 27965 13829 27968
rect 13863 27965 13875 27999
rect 14660 27996 14688 28027
rect 14826 28024 14832 28076
rect 14884 28024 14890 28076
rect 15010 28024 15016 28076
rect 15068 28024 15074 28076
rect 15102 28024 15108 28076
rect 15160 28064 15166 28076
rect 15197 28067 15255 28073
rect 15197 28064 15209 28067
rect 15160 28036 15209 28064
rect 15160 28024 15166 28036
rect 15197 28033 15209 28036
rect 15243 28033 15255 28067
rect 15197 28027 15255 28033
rect 16574 28024 16580 28076
rect 16632 28064 16638 28076
rect 18248 28073 18276 28104
rect 18322 28092 18328 28144
rect 18380 28132 18386 28144
rect 18380 28104 20208 28132
rect 18380 28092 18386 28104
rect 17865 28067 17923 28073
rect 17865 28064 17877 28067
rect 16632 28036 17877 28064
rect 16632 28024 16638 28036
rect 17865 28033 17877 28036
rect 17911 28033 17923 28067
rect 17865 28027 17923 28033
rect 18233 28067 18291 28073
rect 18233 28033 18245 28067
rect 18279 28033 18291 28067
rect 18233 28027 18291 28033
rect 19150 28024 19156 28076
rect 19208 28064 19214 28076
rect 19521 28067 19579 28073
rect 19521 28064 19533 28067
rect 19208 28036 19533 28064
rect 19208 28024 19214 28036
rect 19521 28033 19533 28036
rect 19567 28033 19579 28067
rect 19521 28027 19579 28033
rect 19610 28024 19616 28076
rect 19668 28064 19674 28076
rect 20180 28073 20208 28104
rect 20254 28092 20260 28144
rect 20312 28132 20318 28144
rect 20312 28104 22692 28132
rect 20312 28092 20318 28104
rect 19797 28067 19855 28073
rect 19797 28064 19809 28067
rect 19668 28036 19809 28064
rect 19668 28024 19674 28036
rect 19797 28033 19809 28036
rect 19843 28033 19855 28067
rect 19797 28027 19855 28033
rect 20165 28067 20223 28073
rect 20165 28033 20177 28067
rect 20211 28033 20223 28067
rect 20165 28027 20223 28033
rect 20530 28024 20536 28076
rect 20588 28064 20594 28076
rect 22005 28067 22063 28073
rect 22005 28064 22017 28067
rect 20588 28036 22017 28064
rect 20588 28024 20594 28036
rect 22005 28033 22017 28036
rect 22051 28033 22063 28067
rect 22005 28027 22063 28033
rect 22278 28024 22284 28076
rect 22336 28024 22342 28076
rect 22554 28024 22560 28076
rect 22612 28024 22618 28076
rect 22664 28064 22692 28104
rect 23290 28092 23296 28144
rect 23348 28092 23354 28144
rect 25590 28092 25596 28144
rect 25648 28092 25654 28144
rect 23569 28067 23627 28073
rect 23569 28064 23581 28067
rect 22664 28036 23581 28064
rect 23569 28033 23581 28036
rect 23615 28033 23627 28067
rect 23569 28027 23627 28033
rect 23750 28024 23756 28076
rect 23808 28024 23814 28076
rect 24854 28024 24860 28076
rect 24912 28024 24918 28076
rect 25133 28067 25191 28073
rect 25133 28033 25145 28067
rect 25179 28064 25191 28067
rect 25498 28064 25504 28076
rect 25179 28036 25504 28064
rect 25179 28033 25191 28036
rect 25133 28027 25191 28033
rect 25498 28024 25504 28036
rect 25556 28024 25562 28076
rect 15120 27996 15148 28024
rect 14660 27968 15148 27996
rect 13817 27959 13875 27965
rect 15286 27956 15292 28008
rect 15344 27996 15350 28008
rect 16666 27996 16672 28008
rect 15344 27968 16672 27996
rect 15344 27956 15350 27968
rect 16666 27956 16672 27968
rect 16724 27956 16730 28008
rect 16945 27999 17003 28005
rect 16945 27965 16957 27999
rect 16991 27965 17003 27999
rect 16945 27959 17003 27965
rect 17221 27999 17279 28005
rect 17221 27965 17233 27999
rect 17267 27965 17279 27999
rect 17221 27959 17279 27965
rect 11422 27888 11428 27940
rect 11480 27928 11486 27940
rect 16960 27928 16988 27959
rect 11480 27900 16988 27928
rect 11480 27888 11486 27900
rect 10468 27832 10824 27860
rect 10468 27820 10474 27832
rect 10870 27820 10876 27872
rect 10928 27860 10934 27872
rect 11057 27863 11115 27869
rect 11057 27860 11069 27863
rect 10928 27832 11069 27860
rect 10928 27820 10934 27832
rect 11057 27829 11069 27832
rect 11103 27829 11115 27863
rect 11057 27823 11115 27829
rect 12158 27820 12164 27872
rect 12216 27820 12222 27872
rect 12250 27820 12256 27872
rect 12308 27820 12314 27872
rect 12802 27820 12808 27872
rect 12860 27820 12866 27872
rect 12986 27820 12992 27872
rect 13044 27860 13050 27872
rect 13538 27860 13544 27872
rect 13044 27832 13544 27860
rect 13044 27820 13050 27832
rect 13538 27820 13544 27832
rect 13596 27820 13602 27872
rect 13906 27820 13912 27872
rect 13964 27820 13970 27872
rect 14185 27863 14243 27869
rect 14185 27829 14197 27863
rect 14231 27860 14243 27863
rect 14366 27860 14372 27872
rect 14231 27832 14372 27860
rect 14231 27829 14243 27832
rect 14185 27823 14243 27829
rect 14366 27820 14372 27832
rect 14424 27820 14430 27872
rect 14458 27820 14464 27872
rect 14516 27860 14522 27872
rect 14553 27863 14611 27869
rect 14553 27860 14565 27863
rect 14516 27832 14565 27860
rect 14516 27820 14522 27832
rect 14553 27829 14565 27832
rect 14599 27860 14611 27863
rect 14642 27860 14648 27872
rect 14599 27832 14648 27860
rect 14599 27829 14611 27832
rect 14553 27823 14611 27829
rect 14642 27820 14648 27832
rect 14700 27820 14706 27872
rect 16850 27820 16856 27872
rect 16908 27860 16914 27872
rect 17236 27860 17264 27959
rect 18138 27956 18144 28008
rect 18196 27996 18202 28008
rect 18325 27999 18383 28005
rect 18325 27996 18337 27999
rect 18196 27968 18337 27996
rect 18196 27956 18202 27968
rect 18325 27965 18337 27968
rect 18371 27996 18383 27999
rect 19242 27996 19248 28008
rect 18371 27968 19248 27996
rect 18371 27965 18383 27968
rect 18325 27959 18383 27965
rect 19242 27956 19248 27968
rect 19300 27956 19306 28008
rect 19705 27999 19763 28005
rect 19705 27965 19717 27999
rect 19751 27996 19763 27999
rect 20346 27996 20352 28008
rect 19751 27968 20352 27996
rect 19751 27965 19763 27968
rect 19705 27959 19763 27965
rect 20346 27956 20352 27968
rect 20404 27996 20410 28008
rect 20441 27999 20499 28005
rect 20441 27996 20453 27999
rect 20404 27968 20453 27996
rect 20404 27956 20410 27968
rect 20441 27965 20453 27968
rect 20487 27965 20499 27999
rect 20441 27959 20499 27965
rect 22094 27956 22100 28008
rect 22152 27956 22158 28008
rect 23477 27999 23535 28005
rect 23477 27965 23489 27999
rect 23523 27996 23535 27999
rect 23768 27996 23796 28024
rect 23523 27968 23796 27996
rect 23523 27965 23535 27968
rect 23477 27959 23535 27965
rect 24762 27956 24768 28008
rect 24820 27996 24826 28008
rect 24949 27999 25007 28005
rect 24949 27996 24961 27999
rect 24820 27968 24961 27996
rect 24820 27956 24826 27968
rect 24949 27965 24961 27968
rect 24995 27965 25007 27999
rect 24949 27959 25007 27965
rect 17770 27888 17776 27940
rect 17828 27928 17834 27940
rect 18049 27931 18107 27937
rect 18049 27928 18061 27931
rect 17828 27900 18061 27928
rect 17828 27888 17834 27900
rect 18049 27897 18061 27900
rect 18095 27928 18107 27931
rect 21726 27928 21732 27940
rect 18095 27900 21732 27928
rect 18095 27897 18107 27900
rect 18049 27891 18107 27897
rect 21726 27888 21732 27900
rect 21784 27888 21790 27940
rect 21818 27888 21824 27940
rect 21876 27888 21882 27940
rect 22373 27931 22431 27937
rect 22373 27928 22385 27931
rect 22296 27900 22385 27928
rect 16908 27832 17264 27860
rect 16908 27820 16914 27832
rect 17954 27820 17960 27872
rect 18012 27860 18018 27872
rect 18233 27863 18291 27869
rect 18233 27860 18245 27863
rect 18012 27832 18245 27860
rect 18012 27820 18018 27832
rect 18233 27829 18245 27832
rect 18279 27829 18291 27863
rect 18233 27823 18291 27829
rect 18598 27820 18604 27872
rect 18656 27820 18662 27872
rect 19797 27863 19855 27869
rect 19797 27829 19809 27863
rect 19843 27860 19855 27863
rect 19886 27860 19892 27872
rect 19843 27832 19892 27860
rect 19843 27829 19855 27832
rect 19797 27823 19855 27829
rect 19886 27820 19892 27832
rect 19944 27820 19950 27872
rect 19981 27863 20039 27869
rect 19981 27829 19993 27863
rect 20027 27860 20039 27863
rect 20438 27860 20444 27872
rect 20027 27832 20444 27860
rect 20027 27829 20039 27832
rect 19981 27823 20039 27829
rect 20438 27820 20444 27832
rect 20496 27820 20502 27872
rect 22296 27869 22324 27900
rect 22373 27897 22385 27900
rect 22419 27928 22431 27931
rect 23753 27931 23811 27937
rect 22419 27900 23704 27928
rect 22419 27897 22431 27900
rect 22373 27891 22431 27897
rect 22281 27863 22339 27869
rect 22281 27829 22293 27863
rect 22327 27829 22339 27863
rect 22281 27823 22339 27829
rect 23382 27820 23388 27872
rect 23440 27820 23446 27872
rect 23676 27860 23704 27900
rect 23753 27897 23765 27931
rect 23799 27928 23811 27931
rect 25590 27928 25596 27940
rect 23799 27900 25596 27928
rect 23799 27897 23811 27900
rect 23753 27891 23811 27897
rect 25590 27888 25596 27900
rect 25648 27888 25654 27940
rect 24762 27860 24768 27872
rect 23676 27832 24768 27860
rect 24762 27820 24768 27832
rect 24820 27820 24826 27872
rect 25130 27820 25136 27872
rect 25188 27820 25194 27872
rect 25314 27820 25320 27872
rect 25372 27820 25378 27872
rect 25498 27820 25504 27872
rect 25556 27820 25562 27872
rect 1104 27770 32844 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 32844 27770
rect 1104 27696 32844 27718
rect 1581 27659 1639 27665
rect 1581 27625 1593 27659
rect 1627 27656 1639 27659
rect 1670 27656 1676 27668
rect 1627 27628 1676 27656
rect 1627 27625 1639 27628
rect 1581 27619 1639 27625
rect 1670 27616 1676 27628
rect 1728 27616 1734 27668
rect 4798 27616 4804 27668
rect 4856 27656 4862 27668
rect 5166 27656 5172 27668
rect 4856 27628 5172 27656
rect 4856 27616 4862 27628
rect 5166 27616 5172 27628
rect 5224 27616 5230 27668
rect 7282 27616 7288 27668
rect 7340 27616 7346 27668
rect 7374 27616 7380 27668
rect 7432 27616 7438 27668
rect 7834 27616 7840 27668
rect 7892 27656 7898 27668
rect 9677 27659 9735 27665
rect 7892 27628 8340 27656
rect 7892 27616 7898 27628
rect 2222 27548 2228 27600
rect 2280 27548 2286 27600
rect 2958 27588 2964 27600
rect 2608 27560 2964 27588
rect 2498 27480 2504 27532
rect 2556 27480 2562 27532
rect 2608 27529 2636 27560
rect 2958 27548 2964 27560
rect 3016 27588 3022 27600
rect 3513 27591 3571 27597
rect 3016 27560 3280 27588
rect 3016 27548 3022 27560
rect 2593 27523 2651 27529
rect 2593 27489 2605 27523
rect 2639 27489 2651 27523
rect 2593 27483 2651 27489
rect 2866 27480 2872 27532
rect 2924 27480 2930 27532
rect 3252 27529 3280 27560
rect 3513 27557 3525 27591
rect 3559 27588 3571 27591
rect 3694 27588 3700 27600
rect 3559 27560 3700 27588
rect 3559 27557 3571 27560
rect 3513 27551 3571 27557
rect 3694 27548 3700 27560
rect 3752 27548 3758 27600
rect 3973 27591 4031 27597
rect 3973 27557 3985 27591
rect 4019 27588 4031 27591
rect 4062 27588 4068 27600
rect 4019 27560 4068 27588
rect 4019 27557 4031 27560
rect 3973 27551 4031 27557
rect 4062 27548 4068 27560
rect 4120 27548 4126 27600
rect 4893 27591 4951 27597
rect 4893 27588 4905 27591
rect 4356 27560 4905 27588
rect 3237 27523 3295 27529
rect 3237 27489 3249 27523
rect 3283 27489 3295 27523
rect 3237 27483 3295 27489
rect 3326 27480 3332 27532
rect 3384 27529 3390 27532
rect 3384 27523 3412 27529
rect 3400 27489 3412 27523
rect 3384 27483 3412 27489
rect 3384 27480 3390 27483
rect 1397 27455 1455 27461
rect 1397 27421 1409 27455
rect 1443 27452 1455 27455
rect 1486 27452 1492 27464
rect 1443 27424 1492 27452
rect 1443 27421 1455 27424
rect 1397 27415 1455 27421
rect 1486 27412 1492 27424
rect 1544 27412 1550 27464
rect 2409 27455 2467 27461
rect 2409 27421 2421 27455
rect 2455 27421 2467 27455
rect 2409 27415 2467 27421
rect 2685 27455 2743 27461
rect 2685 27421 2697 27455
rect 2731 27421 2743 27455
rect 2685 27415 2743 27421
rect 2424 27316 2452 27415
rect 2700 27384 2728 27415
rect 3050 27412 3056 27464
rect 3108 27452 3114 27464
rect 4246 27452 4252 27464
rect 3108 27424 4252 27452
rect 3108 27412 3114 27424
rect 4246 27412 4252 27424
rect 4304 27412 4310 27464
rect 4356 27452 4384 27560
rect 4893 27557 4905 27560
rect 4939 27588 4951 27591
rect 4982 27588 4988 27600
rect 4939 27560 4988 27588
rect 4939 27557 4951 27560
rect 4893 27551 4951 27557
rect 4982 27548 4988 27560
rect 5040 27548 5046 27600
rect 5626 27548 5632 27600
rect 5684 27548 5690 27600
rect 6365 27591 6423 27597
rect 6365 27557 6377 27591
rect 6411 27557 6423 27591
rect 6365 27551 6423 27557
rect 4433 27523 4491 27529
rect 4433 27489 4445 27523
rect 4479 27520 4491 27523
rect 4614 27520 4620 27532
rect 4479 27492 4620 27520
rect 4479 27489 4491 27492
rect 4433 27483 4491 27489
rect 4614 27480 4620 27492
rect 4672 27520 4678 27532
rect 5353 27523 5411 27529
rect 5353 27520 5365 27523
rect 4672 27492 5365 27520
rect 4672 27480 4678 27492
rect 5353 27489 5365 27492
rect 5399 27489 5411 27523
rect 6380 27520 6408 27551
rect 6546 27548 6552 27600
rect 6604 27588 6610 27600
rect 7466 27588 7472 27600
rect 6604 27560 7472 27588
rect 6604 27548 6610 27560
rect 7466 27548 7472 27560
rect 7524 27548 7530 27600
rect 7653 27591 7711 27597
rect 7653 27557 7665 27591
rect 7699 27588 7711 27591
rect 8018 27588 8024 27600
rect 7699 27560 8024 27588
rect 7699 27557 7711 27560
rect 7653 27551 7711 27557
rect 5353 27483 5411 27489
rect 5920 27492 6408 27520
rect 6932 27492 7512 27520
rect 4525 27455 4583 27461
rect 4525 27452 4537 27455
rect 4356 27424 4537 27452
rect 4525 27421 4537 27424
rect 4571 27421 4583 27455
rect 5920 27452 5948 27492
rect 6104 27461 6132 27492
rect 6932 27464 6960 27492
rect 4525 27415 4583 27421
rect 4632 27424 5948 27452
rect 5997 27455 6055 27461
rect 3142 27384 3148 27396
rect 2700 27356 3148 27384
rect 3142 27344 3148 27356
rect 3200 27344 3206 27396
rect 3878 27344 3884 27396
rect 3936 27384 3942 27396
rect 3973 27387 4031 27393
rect 3973 27384 3985 27387
rect 3936 27356 3985 27384
rect 3936 27344 3942 27356
rect 3973 27353 3985 27356
rect 4019 27353 4031 27387
rect 3973 27347 4031 27353
rect 3234 27316 3240 27328
rect 2424 27288 3240 27316
rect 3234 27276 3240 27288
rect 3292 27276 3298 27328
rect 3418 27276 3424 27328
rect 3476 27316 3482 27328
rect 4632 27316 4660 27424
rect 5997 27421 6009 27455
rect 6043 27421 6055 27455
rect 5997 27415 6055 27421
rect 6089 27455 6147 27461
rect 6089 27421 6101 27455
rect 6135 27421 6147 27455
rect 6089 27415 6147 27421
rect 4893 27387 4951 27393
rect 4893 27353 4905 27387
rect 4939 27384 4951 27387
rect 4982 27384 4988 27396
rect 4939 27356 4988 27384
rect 4939 27353 4951 27356
rect 4893 27347 4951 27353
rect 4982 27344 4988 27356
rect 5040 27344 5046 27396
rect 5445 27387 5503 27393
rect 5445 27353 5457 27387
rect 5491 27384 5503 27387
rect 5534 27384 5540 27396
rect 5491 27356 5540 27384
rect 5491 27353 5503 27356
rect 5445 27347 5503 27353
rect 5534 27344 5540 27356
rect 5592 27344 5598 27396
rect 6012 27384 6040 27415
rect 6362 27412 6368 27464
rect 6420 27452 6426 27464
rect 6549 27455 6607 27461
rect 6549 27452 6561 27455
rect 6420 27424 6561 27452
rect 6420 27412 6426 27424
rect 6549 27421 6561 27424
rect 6595 27421 6607 27455
rect 6549 27415 6607 27421
rect 6825 27455 6883 27461
rect 6825 27421 6837 27455
rect 6871 27452 6883 27455
rect 6914 27452 6920 27464
rect 6871 27424 6920 27452
rect 6871 27421 6883 27424
rect 6825 27415 6883 27421
rect 6914 27412 6920 27424
rect 6972 27412 6978 27464
rect 7101 27455 7159 27461
rect 7101 27421 7113 27455
rect 7147 27452 7159 27455
rect 7374 27452 7380 27464
rect 7147 27424 7380 27452
rect 7147 27421 7159 27424
rect 7101 27415 7159 27421
rect 7374 27412 7380 27424
rect 7432 27412 7438 27464
rect 6012 27356 6316 27384
rect 6288 27328 6316 27356
rect 6454 27344 6460 27396
rect 6512 27384 6518 27396
rect 7484 27384 7512 27492
rect 7561 27455 7619 27461
rect 7561 27421 7573 27455
rect 7607 27452 7619 27455
rect 7668 27452 7696 27551
rect 8018 27548 8024 27560
rect 8076 27548 8082 27600
rect 8205 27591 8263 27597
rect 8205 27557 8217 27591
rect 8251 27557 8263 27591
rect 8205 27551 8263 27557
rect 8220 27520 8248 27551
rect 7607 27424 7696 27452
rect 7760 27492 8248 27520
rect 7607 27421 7619 27424
rect 7561 27415 7619 27421
rect 7760 27384 7788 27492
rect 7837 27455 7895 27461
rect 7837 27421 7849 27455
rect 7883 27452 7895 27455
rect 7926 27452 7932 27464
rect 7883 27424 7932 27452
rect 7883 27421 7895 27424
rect 7837 27415 7895 27421
rect 7926 27412 7932 27424
rect 7984 27412 7990 27464
rect 8113 27455 8171 27461
rect 8113 27421 8125 27455
rect 8159 27421 8171 27455
rect 8312 27452 8340 27628
rect 9677 27625 9689 27659
rect 9723 27656 9735 27659
rect 9723 27628 10916 27656
rect 9723 27625 9735 27628
rect 9677 27619 9735 27625
rect 9582 27548 9588 27600
rect 9640 27588 9646 27600
rect 9640 27560 10732 27588
rect 9640 27548 9646 27560
rect 9306 27480 9312 27532
rect 9364 27480 9370 27532
rect 9950 27520 9956 27532
rect 9416 27492 9956 27520
rect 8389 27455 8447 27461
rect 8389 27452 8401 27455
rect 8312 27424 8401 27452
rect 8113 27415 8171 27421
rect 8389 27421 8401 27424
rect 8435 27421 8447 27455
rect 8389 27415 8447 27421
rect 8128 27384 8156 27415
rect 8478 27412 8484 27464
rect 8536 27452 8542 27464
rect 8573 27455 8631 27461
rect 8573 27452 8585 27455
rect 8536 27424 8585 27452
rect 8536 27412 8542 27424
rect 8573 27421 8585 27424
rect 8619 27421 8631 27455
rect 8573 27415 8631 27421
rect 9125 27455 9183 27461
rect 9125 27421 9137 27455
rect 9171 27452 9183 27455
rect 9324 27452 9352 27480
rect 9416 27461 9444 27492
rect 9950 27480 9956 27492
rect 10008 27480 10014 27532
rect 9171 27424 9352 27452
rect 9401 27455 9459 27461
rect 9171 27421 9183 27424
rect 9125 27415 9183 27421
rect 9401 27421 9413 27455
rect 9447 27421 9459 27455
rect 9401 27415 9459 27421
rect 9493 27455 9551 27461
rect 9493 27421 9505 27455
rect 9539 27452 9551 27455
rect 9582 27452 9588 27464
rect 9539 27424 9588 27452
rect 9539 27421 9551 27424
rect 9493 27415 9551 27421
rect 9582 27412 9588 27424
rect 9640 27412 9646 27464
rect 9674 27412 9680 27464
rect 9732 27452 9738 27464
rect 9769 27455 9827 27461
rect 9769 27452 9781 27455
rect 9732 27424 9781 27452
rect 9732 27412 9738 27424
rect 9769 27421 9781 27424
rect 9815 27421 9827 27455
rect 9769 27415 9827 27421
rect 10134 27412 10140 27464
rect 10192 27412 10198 27464
rect 10226 27412 10232 27464
rect 10284 27452 10290 27464
rect 10284 27424 10548 27452
rect 10284 27412 10290 27424
rect 6512 27356 7328 27384
rect 7484 27356 7788 27384
rect 7852 27356 8156 27384
rect 9309 27387 9367 27393
rect 6512 27344 6518 27356
rect 3476 27288 4660 27316
rect 4709 27319 4767 27325
rect 3476 27276 3482 27288
rect 4709 27285 4721 27319
rect 4755 27316 4767 27319
rect 5074 27316 5080 27328
rect 4755 27288 5080 27316
rect 4755 27285 4767 27288
rect 4709 27279 4767 27285
rect 5074 27276 5080 27288
rect 5132 27276 5138 27328
rect 5626 27276 5632 27328
rect 5684 27316 5690 27328
rect 5813 27319 5871 27325
rect 5813 27316 5825 27319
rect 5684 27288 5825 27316
rect 5684 27276 5690 27288
rect 5813 27285 5825 27288
rect 5859 27285 5871 27319
rect 5813 27279 5871 27285
rect 6270 27276 6276 27328
rect 6328 27276 6334 27328
rect 7009 27319 7067 27325
rect 7009 27285 7021 27319
rect 7055 27316 7067 27319
rect 7190 27316 7196 27328
rect 7055 27288 7196 27316
rect 7055 27285 7067 27288
rect 7009 27279 7067 27285
rect 7190 27276 7196 27288
rect 7248 27276 7254 27328
rect 7300 27316 7328 27356
rect 7852 27316 7880 27356
rect 9309 27353 9321 27387
rect 9355 27353 9367 27387
rect 9309 27347 9367 27353
rect 7300 27288 7880 27316
rect 7926 27276 7932 27328
rect 7984 27276 7990 27328
rect 8757 27319 8815 27325
rect 8757 27285 8769 27319
rect 8803 27316 8815 27319
rect 9122 27316 9128 27328
rect 8803 27288 9128 27316
rect 8803 27285 8815 27288
rect 8757 27279 8815 27285
rect 9122 27276 9128 27288
rect 9180 27316 9186 27328
rect 9324 27316 9352 27347
rect 9858 27344 9864 27396
rect 9916 27384 9922 27396
rect 9953 27387 10011 27393
rect 9953 27384 9965 27387
rect 9916 27356 9965 27384
rect 9916 27344 9922 27356
rect 9953 27353 9965 27356
rect 9999 27353 10011 27387
rect 9953 27347 10011 27353
rect 10045 27387 10103 27393
rect 10045 27353 10057 27387
rect 10091 27384 10103 27387
rect 10410 27384 10416 27396
rect 10091 27356 10416 27384
rect 10091 27353 10103 27356
rect 10045 27347 10103 27353
rect 9180 27288 9352 27316
rect 9180 27276 9186 27288
rect 9398 27276 9404 27328
rect 9456 27316 9462 27328
rect 10060 27316 10088 27347
rect 10410 27344 10416 27356
rect 10468 27344 10474 27396
rect 10520 27384 10548 27424
rect 10594 27412 10600 27464
rect 10652 27412 10658 27464
rect 10704 27452 10732 27560
rect 10888 27520 10916 27628
rect 11054 27616 11060 27668
rect 11112 27656 11118 27668
rect 12526 27656 12532 27668
rect 11112 27628 12532 27656
rect 11112 27616 11118 27628
rect 12526 27616 12532 27628
rect 12584 27616 12590 27668
rect 14550 27616 14556 27668
rect 14608 27616 14614 27668
rect 15010 27616 15016 27668
rect 15068 27616 15074 27668
rect 15194 27616 15200 27668
rect 15252 27616 15258 27668
rect 16022 27616 16028 27668
rect 16080 27616 16086 27668
rect 16390 27616 16396 27668
rect 16448 27656 16454 27668
rect 16761 27659 16819 27665
rect 16761 27656 16773 27659
rect 16448 27628 16773 27656
rect 16448 27616 16454 27628
rect 16761 27625 16773 27628
rect 16807 27625 16819 27659
rect 17586 27656 17592 27668
rect 16761 27619 16819 27625
rect 16868 27628 17592 27656
rect 10962 27548 10968 27600
rect 11020 27588 11026 27600
rect 11241 27591 11299 27597
rect 11241 27588 11253 27591
rect 11020 27560 11253 27588
rect 11020 27548 11026 27560
rect 11241 27557 11253 27560
rect 11287 27557 11299 27591
rect 11241 27551 11299 27557
rect 11330 27548 11336 27600
rect 11388 27548 11394 27600
rect 12250 27548 12256 27600
rect 12308 27588 12314 27600
rect 12345 27591 12403 27597
rect 12345 27588 12357 27591
rect 12308 27560 12357 27588
rect 12308 27548 12314 27560
rect 12345 27557 12357 27560
rect 12391 27557 12403 27591
rect 12345 27551 12403 27557
rect 12618 27548 12624 27600
rect 12676 27588 12682 27600
rect 12676 27560 12756 27588
rect 12676 27548 12682 27560
rect 11348 27520 11376 27548
rect 12728 27520 12756 27560
rect 12986 27548 12992 27600
rect 13044 27548 13050 27600
rect 14918 27520 14924 27532
rect 10888 27492 11376 27520
rect 11992 27492 12664 27520
rect 12728 27492 13308 27520
rect 11992 27464 12020 27492
rect 10965 27455 11023 27461
rect 10965 27452 10977 27455
rect 10704 27424 10977 27452
rect 10965 27421 10977 27424
rect 11011 27421 11023 27455
rect 10965 27415 11023 27421
rect 11330 27412 11336 27464
rect 11388 27452 11394 27464
rect 11425 27455 11483 27461
rect 11425 27452 11437 27455
rect 11388 27424 11437 27452
rect 11388 27412 11394 27424
rect 11425 27421 11437 27424
rect 11471 27421 11483 27455
rect 11425 27415 11483 27421
rect 11514 27412 11520 27464
rect 11572 27412 11578 27464
rect 11793 27455 11851 27461
rect 11793 27452 11805 27455
rect 11716 27424 11805 27452
rect 10781 27387 10839 27393
rect 10781 27384 10793 27387
rect 10520 27356 10793 27384
rect 10781 27353 10793 27356
rect 10827 27353 10839 27387
rect 10781 27347 10839 27353
rect 10870 27344 10876 27396
rect 10928 27344 10934 27396
rect 9456 27288 10088 27316
rect 10321 27319 10379 27325
rect 9456 27276 9462 27288
rect 10321 27285 10333 27319
rect 10367 27316 10379 27319
rect 11054 27316 11060 27328
rect 10367 27288 11060 27316
rect 10367 27285 10379 27288
rect 10321 27279 10379 27285
rect 11054 27276 11060 27288
rect 11112 27276 11118 27328
rect 11146 27276 11152 27328
rect 11204 27276 11210 27328
rect 11422 27276 11428 27328
rect 11480 27316 11486 27328
rect 11716 27325 11744 27424
rect 11793 27421 11805 27424
rect 11839 27421 11851 27455
rect 11793 27415 11851 27421
rect 11974 27412 11980 27464
rect 12032 27412 12038 27464
rect 12161 27455 12219 27461
rect 12161 27421 12173 27455
rect 12207 27448 12219 27455
rect 12342 27448 12348 27464
rect 12207 27421 12348 27448
rect 12161 27420 12348 27421
rect 12161 27415 12219 27420
rect 12342 27412 12348 27420
rect 12400 27412 12406 27464
rect 12437 27455 12495 27461
rect 12437 27421 12449 27455
rect 12483 27452 12495 27455
rect 12526 27452 12532 27464
rect 12483 27424 12532 27452
rect 12483 27421 12495 27424
rect 12437 27415 12495 27421
rect 12526 27412 12532 27424
rect 12584 27412 12590 27464
rect 12636 27461 12664 27492
rect 12621 27455 12679 27461
rect 12621 27421 12633 27455
rect 12667 27421 12679 27455
rect 12621 27415 12679 27421
rect 12802 27412 12808 27464
rect 12860 27412 12866 27464
rect 13280 27461 13308 27492
rect 14108 27492 14924 27520
rect 13265 27455 13323 27461
rect 13265 27421 13277 27455
rect 13311 27421 13323 27455
rect 13265 27415 13323 27421
rect 11882 27344 11888 27396
rect 11940 27384 11946 27396
rect 12069 27387 12127 27393
rect 12069 27384 12081 27387
rect 11940 27356 12081 27384
rect 11940 27344 11946 27356
rect 12069 27353 12081 27356
rect 12115 27353 12127 27387
rect 12069 27347 12127 27353
rect 12713 27387 12771 27393
rect 12713 27353 12725 27387
rect 12759 27353 12771 27387
rect 12713 27347 12771 27353
rect 11701 27319 11759 27325
rect 11701 27316 11713 27319
rect 11480 27288 11713 27316
rect 11480 27276 11486 27288
rect 11701 27285 11713 27288
rect 11747 27316 11759 27319
rect 12728 27316 12756 27347
rect 11747 27288 12756 27316
rect 12820 27316 12848 27412
rect 13081 27319 13139 27325
rect 13081 27316 13093 27319
rect 12820 27288 13093 27316
rect 11747 27285 11759 27288
rect 11701 27279 11759 27285
rect 13081 27285 13093 27288
rect 13127 27285 13139 27319
rect 13081 27279 13139 27285
rect 13354 27276 13360 27328
rect 13412 27316 13418 27328
rect 14108 27325 14136 27492
rect 14384 27461 14412 27492
rect 14918 27480 14924 27492
rect 14976 27480 14982 27532
rect 15028 27461 15056 27616
rect 15565 27591 15623 27597
rect 15565 27557 15577 27591
rect 15611 27588 15623 27591
rect 15611 27560 16068 27588
rect 15611 27557 15623 27560
rect 15565 27551 15623 27557
rect 16040 27529 16068 27560
rect 16298 27548 16304 27600
rect 16356 27548 16362 27600
rect 16868 27529 16896 27628
rect 17586 27616 17592 27628
rect 17644 27616 17650 27668
rect 17954 27616 17960 27668
rect 18012 27656 18018 27668
rect 18874 27656 18880 27668
rect 18012 27628 18880 27656
rect 18012 27616 18018 27628
rect 18874 27616 18880 27628
rect 18932 27616 18938 27668
rect 19334 27616 19340 27668
rect 19392 27656 19398 27668
rect 20254 27656 20260 27668
rect 19392 27628 20260 27656
rect 19392 27616 19398 27628
rect 20254 27616 20260 27628
rect 20312 27616 20318 27668
rect 20438 27616 20444 27668
rect 20496 27616 20502 27668
rect 22462 27616 22468 27668
rect 22520 27616 22526 27668
rect 23661 27659 23719 27665
rect 22664 27628 22876 27656
rect 22664 27588 22692 27628
rect 16960 27560 18920 27588
rect 16025 27523 16083 27529
rect 16025 27489 16037 27523
rect 16071 27489 16083 27523
rect 16025 27483 16083 27489
rect 16853 27523 16911 27529
rect 16853 27489 16865 27523
rect 16899 27489 16911 27523
rect 16853 27483 16911 27489
rect 14277 27455 14335 27461
rect 14277 27421 14289 27455
rect 14323 27421 14335 27455
rect 14277 27415 14335 27421
rect 14369 27455 14427 27461
rect 14369 27421 14381 27455
rect 14415 27421 14427 27455
rect 14369 27415 14427 27421
rect 14553 27455 14611 27461
rect 14553 27421 14565 27455
rect 14599 27452 14611 27455
rect 15013 27455 15071 27461
rect 14599 27424 14872 27452
rect 14599 27421 14611 27424
rect 14553 27415 14611 27421
rect 14292 27384 14320 27415
rect 14292 27356 14596 27384
rect 14568 27328 14596 27356
rect 14093 27319 14151 27325
rect 14093 27316 14105 27319
rect 13412 27288 14105 27316
rect 13412 27276 13418 27288
rect 14093 27285 14105 27288
rect 14139 27285 14151 27319
rect 14093 27279 14151 27285
rect 14550 27276 14556 27328
rect 14608 27276 14614 27328
rect 14642 27276 14648 27328
rect 14700 27316 14706 27328
rect 14844 27325 14872 27424
rect 15013 27421 15025 27455
rect 15059 27421 15071 27455
rect 15013 27415 15071 27421
rect 15194 27412 15200 27464
rect 15252 27452 15258 27464
rect 15289 27455 15347 27461
rect 15289 27452 15301 27455
rect 15252 27424 15301 27452
rect 15252 27412 15258 27424
rect 15289 27421 15301 27424
rect 15335 27421 15347 27455
rect 15289 27415 15347 27421
rect 15378 27412 15384 27464
rect 15436 27412 15442 27464
rect 15933 27455 15991 27461
rect 15933 27421 15945 27455
rect 15979 27421 15991 27455
rect 15933 27415 15991 27421
rect 14918 27344 14924 27396
rect 14976 27384 14982 27396
rect 15105 27387 15163 27393
rect 15105 27384 15117 27387
rect 14976 27356 15117 27384
rect 14976 27344 14982 27356
rect 15105 27353 15117 27356
rect 15151 27353 15163 27387
rect 15948 27384 15976 27415
rect 16482 27412 16488 27464
rect 16540 27412 16546 27464
rect 16960 27452 16988 27560
rect 18414 27480 18420 27532
rect 18472 27520 18478 27532
rect 18785 27523 18843 27529
rect 18785 27520 18797 27523
rect 18472 27492 18797 27520
rect 18472 27480 18478 27492
rect 18785 27489 18797 27492
rect 18831 27489 18843 27523
rect 18892 27520 18920 27560
rect 19076 27560 19472 27588
rect 19076 27520 19104 27560
rect 18892 27492 19104 27520
rect 18785 27483 18843 27489
rect 19242 27480 19248 27532
rect 19300 27480 19306 27532
rect 16592 27424 16988 27452
rect 17037 27455 17095 27461
rect 16592 27384 16620 27424
rect 17037 27421 17049 27455
rect 17083 27421 17095 27455
rect 17037 27415 17095 27421
rect 16761 27387 16819 27393
rect 16761 27384 16773 27387
rect 15948 27356 16620 27384
rect 16684 27356 16773 27384
rect 15105 27347 15163 27353
rect 14737 27319 14795 27325
rect 14737 27316 14749 27319
rect 14700 27288 14749 27316
rect 14700 27276 14706 27288
rect 14737 27285 14749 27288
rect 14783 27285 14795 27319
rect 14737 27279 14795 27285
rect 14829 27319 14887 27325
rect 14829 27285 14841 27319
rect 14875 27316 14887 27319
rect 16298 27316 16304 27328
rect 14875 27288 16304 27316
rect 14875 27285 14887 27288
rect 14829 27279 14887 27285
rect 16298 27276 16304 27288
rect 16356 27276 16362 27328
rect 16684 27325 16712 27356
rect 16761 27353 16773 27356
rect 16807 27384 16819 27387
rect 16942 27384 16948 27396
rect 16807 27356 16948 27384
rect 16807 27353 16819 27356
rect 16761 27347 16819 27353
rect 16942 27344 16948 27356
rect 17000 27344 17006 27396
rect 17052 27384 17080 27415
rect 17218 27412 17224 27464
rect 17276 27452 17282 27464
rect 17313 27455 17371 27461
rect 17313 27452 17325 27455
rect 17276 27424 17325 27452
rect 17276 27412 17282 27424
rect 17313 27421 17325 27424
rect 17359 27421 17371 27455
rect 17313 27415 17371 27421
rect 17770 27412 17776 27464
rect 17828 27412 17834 27464
rect 18690 27412 18696 27464
rect 18748 27412 18754 27464
rect 19444 27452 19472 27560
rect 19812 27560 22692 27588
rect 22741 27591 22799 27597
rect 19518 27480 19524 27532
rect 19576 27480 19582 27532
rect 19812 27452 19840 27560
rect 22741 27557 22753 27591
rect 22787 27557 22799 27591
rect 22848 27588 22876 27628
rect 23661 27625 23673 27659
rect 23707 27656 23719 27659
rect 24210 27656 24216 27668
rect 23707 27628 24216 27656
rect 23707 27625 23719 27628
rect 23661 27619 23719 27625
rect 24210 27616 24216 27628
rect 24268 27616 24274 27668
rect 25590 27616 25596 27668
rect 25648 27616 25654 27668
rect 26142 27616 26148 27668
rect 26200 27656 26206 27668
rect 29730 27656 29736 27668
rect 26200 27628 29736 27656
rect 26200 27616 26206 27628
rect 29730 27616 29736 27628
rect 29788 27616 29794 27668
rect 23753 27591 23811 27597
rect 23753 27588 23765 27591
rect 22848 27560 23765 27588
rect 22741 27551 22799 27557
rect 23753 27557 23765 27560
rect 23799 27557 23811 27591
rect 23753 27551 23811 27557
rect 20254 27480 20260 27532
rect 20312 27520 20318 27532
rect 20312 27492 20576 27520
rect 20312 27480 20318 27492
rect 19444 27424 19840 27452
rect 19978 27412 19984 27464
rect 20036 27452 20042 27464
rect 20349 27455 20407 27461
rect 20349 27452 20361 27455
rect 20036 27424 20361 27452
rect 20036 27412 20042 27424
rect 20349 27421 20361 27424
rect 20395 27421 20407 27455
rect 20349 27415 20407 27421
rect 20441 27455 20499 27461
rect 20441 27421 20453 27455
rect 20487 27421 20499 27455
rect 20548 27452 20576 27492
rect 22370 27480 22376 27532
rect 22428 27480 22434 27532
rect 22756 27520 22784 27551
rect 25314 27548 25320 27600
rect 25372 27588 25378 27600
rect 25372 27560 25820 27588
rect 25372 27548 25378 27560
rect 25792 27529 25820 27560
rect 25777 27523 25835 27529
rect 22756 27492 25636 27520
rect 22557 27455 22615 27461
rect 22557 27452 22569 27455
rect 20548 27424 22569 27452
rect 20441 27415 20499 27421
rect 22557 27421 22569 27424
rect 22603 27452 22615 27455
rect 23566 27452 23572 27464
rect 22603 27424 23572 27452
rect 22603 27421 22615 27424
rect 22557 27415 22615 27421
rect 17862 27384 17868 27396
rect 17052 27356 17868 27384
rect 16669 27319 16727 27325
rect 16669 27285 16681 27319
rect 16715 27285 16727 27319
rect 16669 27279 16727 27285
rect 17221 27319 17279 27325
rect 17221 27285 17233 27319
rect 17267 27316 17279 27319
rect 17310 27316 17316 27328
rect 17267 27288 17316 27316
rect 17267 27285 17279 27288
rect 17221 27279 17279 27285
rect 17310 27276 17316 27288
rect 17368 27276 17374 27328
rect 17512 27325 17540 27356
rect 17862 27344 17868 27356
rect 17920 27344 17926 27396
rect 19426 27384 19432 27396
rect 18984 27356 19432 27384
rect 17497 27319 17555 27325
rect 17497 27285 17509 27319
rect 17543 27285 17555 27319
rect 17497 27279 17555 27285
rect 17586 27276 17592 27328
rect 17644 27316 17650 27328
rect 18984 27316 19012 27356
rect 19426 27344 19432 27356
rect 19484 27344 19490 27396
rect 20165 27387 20223 27393
rect 20165 27384 20177 27387
rect 19628 27356 20177 27384
rect 19628 27328 19656 27356
rect 20165 27353 20177 27356
rect 20211 27353 20223 27387
rect 20456 27384 20484 27415
rect 23566 27412 23572 27424
rect 23624 27412 23630 27464
rect 23934 27412 23940 27464
rect 23992 27412 23998 27464
rect 25608 27461 25636 27492
rect 25777 27489 25789 27523
rect 25823 27520 25835 27523
rect 26510 27520 26516 27532
rect 25823 27492 26516 27520
rect 25823 27489 25835 27492
rect 25777 27483 25835 27489
rect 26510 27480 26516 27492
rect 26568 27480 26574 27532
rect 24029 27455 24087 27461
rect 24029 27421 24041 27455
rect 24075 27421 24087 27455
rect 24029 27415 24087 27421
rect 25593 27455 25651 27461
rect 25593 27421 25605 27455
rect 25639 27421 25651 27455
rect 25593 27415 25651 27421
rect 25869 27455 25927 27461
rect 25869 27421 25881 27455
rect 25915 27452 25927 27455
rect 25958 27452 25964 27464
rect 25915 27424 25964 27452
rect 25915 27421 25927 27424
rect 25869 27415 25927 27421
rect 20456 27356 22140 27384
rect 20165 27347 20223 27353
rect 17644 27288 19012 27316
rect 19061 27319 19119 27325
rect 17644 27276 17650 27288
rect 19061 27285 19073 27319
rect 19107 27316 19119 27319
rect 19242 27316 19248 27328
rect 19107 27288 19248 27316
rect 19107 27285 19119 27288
rect 19061 27279 19119 27285
rect 19242 27276 19248 27288
rect 19300 27276 19306 27328
rect 19610 27276 19616 27328
rect 19668 27276 19674 27328
rect 19702 27276 19708 27328
rect 19760 27316 19766 27328
rect 19978 27316 19984 27328
rect 19760 27288 19984 27316
rect 19760 27276 19766 27288
rect 19978 27276 19984 27288
rect 20036 27276 20042 27328
rect 20625 27319 20683 27325
rect 20625 27285 20637 27319
rect 20671 27316 20683 27319
rect 22002 27316 22008 27328
rect 20671 27288 22008 27316
rect 20671 27285 20683 27288
rect 20625 27279 20683 27285
rect 22002 27276 22008 27288
rect 22060 27276 22066 27328
rect 22112 27316 22140 27356
rect 22278 27344 22284 27396
rect 22336 27344 22342 27396
rect 23842 27344 23848 27396
rect 23900 27384 23906 27396
rect 24044 27384 24072 27415
rect 25958 27412 25964 27424
rect 26016 27412 26022 27464
rect 23900 27356 24072 27384
rect 23900 27344 23906 27356
rect 24118 27344 24124 27396
rect 24176 27384 24182 27396
rect 24213 27387 24271 27393
rect 24213 27384 24225 27387
rect 24176 27356 24225 27384
rect 24176 27344 24182 27356
rect 24213 27353 24225 27356
rect 24259 27353 24271 27387
rect 26605 27387 26663 27393
rect 26605 27384 26617 27387
rect 24213 27347 24271 27353
rect 24320 27356 26617 27384
rect 22922 27316 22928 27328
rect 22112 27288 22928 27316
rect 22922 27276 22928 27288
rect 22980 27276 22986 27328
rect 23934 27276 23940 27328
rect 23992 27316 23998 27328
rect 24320 27316 24348 27356
rect 26605 27353 26617 27356
rect 26651 27353 26663 27387
rect 26605 27347 26663 27353
rect 26786 27344 26792 27396
rect 26844 27344 26850 27396
rect 23992 27288 24348 27316
rect 26053 27319 26111 27325
rect 23992 27276 23998 27288
rect 26053 27285 26065 27319
rect 26099 27316 26111 27319
rect 26878 27316 26884 27328
rect 26099 27288 26884 27316
rect 26099 27285 26111 27288
rect 26053 27279 26111 27285
rect 26878 27276 26884 27288
rect 26936 27276 26942 27328
rect 26973 27319 27031 27325
rect 26973 27285 26985 27319
rect 27019 27316 27031 27319
rect 27338 27316 27344 27328
rect 27019 27288 27344 27316
rect 27019 27285 27031 27288
rect 26973 27279 27031 27285
rect 27338 27276 27344 27288
rect 27396 27276 27402 27328
rect 1104 27226 32844 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 32844 27226
rect 1104 27152 32844 27174
rect 3050 27112 3056 27124
rect 2056 27084 3056 27112
rect 2056 26985 2084 27084
rect 3050 27072 3056 27084
rect 3108 27072 3114 27124
rect 3510 27072 3516 27124
rect 3568 27112 3574 27124
rect 3973 27115 4031 27121
rect 3973 27112 3985 27115
rect 3568 27084 3985 27112
rect 3568 27072 3574 27084
rect 3973 27081 3985 27084
rect 4019 27081 4031 27115
rect 3973 27075 4031 27081
rect 4617 27115 4675 27121
rect 4617 27081 4629 27115
rect 4663 27112 4675 27115
rect 4706 27112 4712 27124
rect 4663 27084 4712 27112
rect 4663 27081 4675 27084
rect 4617 27075 4675 27081
rect 2774 27044 2780 27056
rect 2240 27016 2780 27044
rect 2041 26979 2099 26985
rect 2041 26945 2053 26979
rect 2087 26945 2099 26979
rect 2041 26939 2099 26945
rect 2240 26849 2268 27016
rect 2774 27004 2780 27016
rect 2832 27044 2838 27056
rect 3988 27044 4016 27075
rect 4706 27072 4712 27084
rect 4764 27112 4770 27124
rect 4985 27115 5043 27121
rect 4985 27112 4997 27115
rect 4764 27084 4997 27112
rect 4764 27072 4770 27084
rect 4985 27081 4997 27084
rect 5031 27081 5043 27115
rect 4985 27075 5043 27081
rect 5074 27072 5080 27124
rect 5132 27112 5138 27124
rect 6454 27112 6460 27124
rect 5132 27084 6460 27112
rect 5132 27072 5138 27084
rect 6454 27072 6460 27084
rect 6512 27072 6518 27124
rect 6549 27115 6607 27121
rect 6549 27081 6561 27115
rect 6595 27112 6607 27115
rect 6638 27112 6644 27124
rect 6595 27084 6644 27112
rect 6595 27081 6607 27084
rect 6549 27075 6607 27081
rect 6638 27072 6644 27084
rect 6696 27112 6702 27124
rect 6696 27084 6776 27112
rect 6696 27072 6702 27084
rect 6178 27044 6184 27056
rect 2832 27016 3004 27044
rect 3988 27016 4476 27044
rect 2832 27004 2838 27016
rect 2314 26936 2320 26988
rect 2372 26936 2378 26988
rect 2866 26936 2872 26988
rect 2924 26936 2930 26988
rect 2976 26985 3004 27016
rect 2961 26979 3019 26985
rect 2961 26945 2973 26979
rect 3007 26945 3019 26979
rect 2961 26939 3019 26945
rect 3234 26936 3240 26988
rect 3292 26936 3298 26988
rect 3510 26936 3516 26988
rect 3568 26936 3574 26988
rect 3786 26936 3792 26988
rect 3844 26936 3850 26988
rect 3878 26936 3884 26988
rect 3936 26976 3942 26988
rect 4448 26985 4476 27016
rect 5368 27016 6184 27044
rect 4065 26979 4123 26985
rect 4065 26976 4077 26979
rect 3936 26948 4077 26976
rect 3936 26936 3942 26948
rect 4065 26945 4077 26948
rect 4111 26945 4123 26979
rect 4065 26939 4123 26945
rect 4433 26979 4491 26985
rect 4433 26945 4445 26979
rect 4479 26945 4491 26979
rect 4433 26939 4491 26945
rect 4706 26936 4712 26988
rect 4764 26936 4770 26988
rect 4890 26936 4896 26988
rect 4948 26976 4954 26988
rect 5194 26979 5252 26985
rect 5194 26976 5206 26979
rect 4948 26948 5206 26976
rect 4948 26936 4954 26948
rect 5194 26945 5206 26948
rect 5240 26976 5252 26979
rect 5368 26976 5396 27016
rect 6178 27004 6184 27016
rect 6236 27004 6242 27056
rect 5537 26979 5595 26985
rect 5537 26976 5549 26979
rect 5240 26948 5396 26976
rect 5460 26948 5549 26976
rect 5240 26945 5252 26948
rect 5194 26939 5252 26945
rect 2590 26868 2596 26920
rect 2648 26868 2654 26920
rect 2777 26911 2835 26917
rect 2777 26877 2789 26911
rect 2823 26908 2835 26911
rect 2823 26880 2857 26908
rect 2823 26877 2835 26880
rect 2777 26871 2835 26877
rect 2225 26843 2283 26849
rect 2225 26809 2237 26843
rect 2271 26809 2283 26843
rect 2225 26803 2283 26809
rect 2501 26843 2559 26849
rect 2501 26809 2513 26843
rect 2547 26840 2559 26843
rect 2792 26840 2820 26871
rect 3050 26868 3056 26920
rect 3108 26868 3114 26920
rect 3252 26908 3280 26936
rect 3252 26880 3740 26908
rect 2958 26840 2964 26852
rect 2547 26812 2964 26840
rect 2547 26809 2559 26812
rect 2501 26803 2559 26809
rect 2958 26800 2964 26812
rect 3016 26800 3022 26852
rect 3712 26849 3740 26880
rect 3970 26868 3976 26920
rect 4028 26908 4034 26920
rect 4614 26908 4620 26920
rect 4028 26880 4620 26908
rect 4028 26868 4034 26880
rect 4614 26868 4620 26880
rect 4672 26908 4678 26920
rect 5077 26911 5135 26917
rect 5077 26908 5089 26911
rect 4672 26880 5089 26908
rect 4672 26868 4678 26880
rect 5077 26877 5089 26880
rect 5123 26877 5135 26911
rect 5077 26871 5135 26877
rect 3697 26843 3755 26849
rect 3697 26809 3709 26843
rect 3743 26840 3755 26843
rect 4062 26840 4068 26852
rect 3743 26812 4068 26840
rect 3743 26809 3755 26812
rect 3697 26803 3755 26809
rect 4062 26800 4068 26812
rect 4120 26800 4126 26852
rect 5460 26840 5488 26948
rect 5537 26945 5549 26948
rect 5583 26945 5595 26979
rect 5537 26939 5595 26945
rect 5626 26936 5632 26988
rect 5684 26976 5690 26988
rect 5813 26979 5871 26985
rect 5813 26976 5825 26979
rect 5684 26948 5825 26976
rect 5684 26936 5690 26948
rect 5813 26945 5825 26948
rect 5859 26945 5871 26979
rect 5813 26939 5871 26945
rect 6365 26979 6423 26985
rect 6365 26945 6377 26979
rect 6411 26945 6423 26979
rect 6365 26939 6423 26945
rect 6380 26908 6408 26939
rect 6546 26936 6552 26988
rect 6604 26976 6610 26988
rect 6641 26979 6699 26985
rect 6641 26976 6653 26979
rect 6604 26948 6653 26976
rect 6604 26936 6610 26948
rect 6641 26945 6653 26948
rect 6687 26945 6699 26979
rect 6748 26976 6776 27084
rect 7006 27072 7012 27124
rect 7064 27112 7070 27124
rect 7193 27115 7251 27121
rect 7193 27112 7205 27115
rect 7064 27084 7205 27112
rect 7064 27072 7070 27084
rect 7193 27081 7205 27084
rect 7239 27081 7251 27115
rect 7193 27075 7251 27081
rect 7282 27072 7288 27124
rect 7340 27072 7346 27124
rect 7466 27072 7472 27124
rect 7524 27112 7530 27124
rect 7524 27084 7696 27112
rect 7524 27072 7530 27084
rect 6825 27047 6883 27053
rect 6825 27013 6837 27047
rect 6871 27044 6883 27047
rect 7098 27044 7104 27056
rect 6871 27016 7104 27044
rect 6871 27013 6883 27016
rect 6825 27007 6883 27013
rect 7098 27004 7104 27016
rect 7156 27004 7162 27056
rect 7300 27044 7328 27072
rect 7561 27047 7619 27053
rect 7561 27044 7573 27047
rect 7300 27016 7573 27044
rect 7561 27013 7573 27016
rect 7607 27013 7619 27047
rect 7668 27044 7696 27084
rect 9490 27072 9496 27124
rect 9548 27112 9554 27124
rect 9548 27084 10088 27112
rect 9548 27072 9554 27084
rect 7668 27016 8064 27044
rect 7561 27007 7619 27013
rect 6917 26979 6975 26985
rect 6917 26976 6929 26979
rect 6748 26948 6929 26976
rect 6641 26939 6699 26945
rect 6917 26945 6929 26948
rect 6963 26945 6975 26979
rect 6917 26939 6975 26945
rect 6822 26908 6828 26920
rect 6380 26880 6828 26908
rect 6380 26840 6408 26880
rect 6822 26868 6828 26880
rect 6880 26868 6886 26920
rect 4172 26812 5488 26840
rect 5920 26812 6408 26840
rect 6932 26840 6960 26939
rect 7006 26936 7012 26988
rect 7064 26936 7070 26988
rect 7190 26936 7196 26988
rect 7248 26976 7254 26988
rect 7285 26979 7343 26985
rect 7285 26976 7297 26979
rect 7248 26948 7297 26976
rect 7248 26936 7254 26948
rect 7285 26945 7297 26948
rect 7331 26945 7343 26979
rect 7285 26939 7343 26945
rect 7300 26908 7328 26939
rect 7466 26936 7472 26988
rect 7524 26936 7530 26988
rect 7650 26936 7656 26988
rect 7708 26936 7714 26988
rect 7834 26936 7840 26988
rect 7892 26976 7898 26988
rect 7929 26979 7987 26985
rect 7929 26976 7941 26979
rect 7892 26948 7941 26976
rect 7892 26936 7898 26948
rect 7929 26945 7941 26948
rect 7975 26945 7987 26979
rect 8036 26976 8064 27016
rect 8754 27004 8760 27056
rect 8812 27044 8818 27056
rect 8941 27047 8999 27053
rect 8941 27044 8953 27047
rect 8812 27016 8953 27044
rect 8812 27004 8818 27016
rect 8941 27013 8953 27016
rect 8987 27013 8999 27047
rect 9766 27044 9772 27056
rect 8941 27007 8999 27013
rect 9508 27016 9772 27044
rect 8113 26979 8171 26985
rect 8113 26976 8125 26979
rect 8036 26948 8125 26976
rect 7929 26939 7987 26945
rect 8113 26945 8125 26948
rect 8159 26945 8171 26979
rect 8113 26939 8171 26945
rect 8205 26979 8263 26985
rect 8205 26945 8217 26979
rect 8251 26945 8263 26979
rect 8205 26939 8263 26945
rect 8297 26979 8355 26985
rect 8297 26945 8309 26979
rect 8343 26945 8355 26979
rect 8297 26939 8355 26945
rect 7742 26908 7748 26920
rect 7300 26880 7748 26908
rect 7742 26868 7748 26880
rect 7800 26868 7806 26920
rect 8220 26908 8248 26939
rect 7852 26880 8248 26908
rect 7852 26840 7880 26880
rect 6932 26812 7880 26840
rect 3142 26732 3148 26784
rect 3200 26772 3206 26784
rect 3421 26775 3479 26781
rect 3421 26772 3433 26775
rect 3200 26744 3433 26772
rect 3200 26732 3206 26744
rect 3421 26741 3433 26744
rect 3467 26741 3479 26775
rect 3421 26735 3479 26741
rect 3510 26732 3516 26784
rect 3568 26772 3574 26784
rect 4172 26772 4200 26812
rect 5920 26784 5948 26812
rect 8110 26800 8116 26852
rect 8168 26840 8174 26852
rect 8312 26840 8340 26939
rect 8386 26936 8392 26988
rect 8444 26976 8450 26988
rect 8849 26979 8907 26985
rect 8849 26976 8861 26979
rect 8444 26948 8861 26976
rect 8444 26936 8450 26948
rect 8849 26945 8861 26948
rect 8895 26945 8907 26979
rect 8849 26939 8907 26945
rect 9030 26936 9036 26988
rect 9088 26936 9094 26988
rect 9122 26936 9128 26988
rect 9180 26976 9186 26988
rect 9217 26979 9275 26985
rect 9217 26976 9229 26979
rect 9180 26948 9229 26976
rect 9180 26936 9186 26948
rect 9217 26945 9229 26948
rect 9263 26945 9275 26979
rect 9217 26939 9275 26945
rect 9306 26936 9312 26988
rect 9364 26936 9370 26988
rect 9508 26985 9536 27016
rect 9766 27004 9772 27016
rect 9824 27004 9830 27056
rect 9493 26979 9551 26985
rect 9493 26945 9505 26979
rect 9539 26945 9551 26979
rect 9493 26939 9551 26945
rect 9585 26979 9643 26985
rect 9585 26945 9597 26979
rect 9631 26945 9643 26979
rect 9585 26939 9643 26945
rect 9677 26979 9735 26985
rect 9677 26945 9689 26979
rect 9723 26976 9735 26979
rect 9950 26976 9956 26988
rect 9723 26948 9956 26976
rect 9723 26945 9735 26948
rect 9677 26939 9735 26945
rect 9398 26868 9404 26920
rect 9456 26908 9462 26920
rect 9600 26908 9628 26939
rect 9950 26936 9956 26948
rect 10008 26936 10014 26988
rect 10060 26976 10088 27084
rect 10226 27072 10232 27124
rect 10284 27072 10290 27124
rect 10410 27072 10416 27124
rect 10468 27112 10474 27124
rect 10597 27115 10655 27121
rect 10597 27112 10609 27115
rect 10468 27084 10609 27112
rect 10468 27072 10474 27084
rect 10597 27081 10609 27084
rect 10643 27081 10655 27115
rect 11698 27112 11704 27124
rect 10597 27075 10655 27081
rect 11348 27084 11704 27112
rect 10137 27047 10195 27053
rect 10137 27013 10149 27047
rect 10183 27044 10195 27047
rect 10244 27044 10272 27072
rect 11238 27044 11244 27056
rect 10183 27016 11244 27044
rect 10183 27013 10195 27016
rect 10137 27007 10195 27013
rect 11238 27004 11244 27016
rect 11296 27004 11302 27056
rect 10229 26979 10287 26985
rect 10229 26976 10241 26979
rect 10060 26948 10241 26976
rect 10229 26945 10241 26948
rect 10275 26945 10287 26979
rect 10229 26939 10287 26945
rect 10321 26979 10379 26985
rect 10321 26945 10333 26979
rect 10367 26945 10379 26979
rect 10321 26939 10379 26945
rect 10781 26979 10839 26985
rect 10781 26945 10793 26979
rect 10827 26976 10839 26979
rect 10962 26976 10968 26988
rect 10827 26948 10968 26976
rect 10827 26945 10839 26948
rect 10781 26939 10839 26945
rect 9456 26880 9628 26908
rect 9456 26868 9462 26880
rect 9766 26868 9772 26920
rect 9824 26908 9830 26920
rect 10336 26908 10364 26939
rect 10962 26936 10968 26948
rect 11020 26936 11026 26988
rect 11054 26936 11060 26988
rect 11112 26976 11118 26988
rect 11348 26976 11376 27084
rect 11698 27072 11704 27084
rect 11756 27072 11762 27124
rect 11790 27072 11796 27124
rect 11848 27112 11854 27124
rect 12526 27112 12532 27124
rect 11848 27084 12532 27112
rect 11848 27072 11854 27084
rect 12526 27072 12532 27084
rect 12584 27072 12590 27124
rect 13722 27072 13728 27124
rect 13780 27112 13786 27124
rect 14369 27115 14427 27121
rect 14369 27112 14381 27115
rect 13780 27084 14381 27112
rect 13780 27072 13786 27084
rect 14369 27081 14381 27084
rect 14415 27112 14427 27115
rect 14415 27084 14780 27112
rect 14415 27081 14427 27084
rect 14369 27075 14427 27081
rect 13354 27044 13360 27056
rect 11112 26948 11376 26976
rect 12360 27016 13360 27044
rect 11112 26936 11118 26948
rect 9824 26880 10364 26908
rect 9824 26868 9830 26880
rect 10410 26868 10416 26920
rect 10468 26908 10474 26920
rect 12360 26908 12388 27016
rect 13354 27004 13360 27016
rect 13412 27004 13418 27056
rect 13630 27044 13636 27056
rect 13464 27016 13636 27044
rect 12434 26936 12440 26988
rect 12492 26976 12498 26988
rect 13081 26979 13139 26985
rect 13081 26976 13093 26979
rect 12492 26948 13093 26976
rect 12492 26936 12498 26948
rect 13081 26945 13093 26948
rect 13127 26976 13139 26979
rect 13170 26976 13176 26988
rect 13127 26948 13176 26976
rect 13127 26945 13139 26948
rect 13081 26939 13139 26945
rect 13170 26936 13176 26948
rect 13228 26936 13234 26988
rect 13464 26985 13492 27016
rect 13630 27004 13636 27016
rect 13688 27004 13694 27056
rect 14458 27004 14464 27056
rect 14516 27004 14522 27056
rect 13272 26979 13330 26985
rect 13272 26945 13284 26979
rect 13318 26945 13330 26979
rect 13272 26939 13330 26945
rect 13449 26979 13507 26985
rect 13449 26945 13461 26979
rect 13495 26945 13507 26979
rect 13449 26939 13507 26945
rect 13541 26979 13599 26985
rect 13541 26945 13553 26979
rect 13587 26976 13599 26979
rect 13722 26976 13728 26988
rect 13587 26948 13728 26976
rect 13587 26945 13599 26948
rect 13541 26939 13599 26945
rect 10468 26880 12388 26908
rect 10468 26868 10474 26880
rect 12986 26868 12992 26920
rect 13044 26908 13050 26920
rect 13280 26908 13308 26939
rect 13722 26936 13728 26948
rect 13780 26936 13786 26988
rect 13998 26936 14004 26988
rect 14056 26936 14062 26988
rect 14182 26936 14188 26988
rect 14240 26936 14246 26988
rect 14752 26985 14780 27084
rect 14918 27072 14924 27124
rect 14976 27072 14982 27124
rect 15010 27072 15016 27124
rect 15068 27112 15074 27124
rect 22278 27112 22284 27124
rect 15068 27084 22284 27112
rect 15068 27072 15074 27084
rect 22278 27072 22284 27084
rect 22336 27072 22342 27124
rect 22554 27072 22560 27124
rect 22612 27112 22618 27124
rect 22612 27084 25176 27112
rect 22612 27072 22618 27084
rect 14826 27004 14832 27056
rect 14884 27044 14890 27056
rect 14884 27016 17172 27044
rect 14884 27004 14890 27016
rect 14737 26979 14795 26985
rect 14292 26948 14688 26976
rect 13044 26880 13308 26908
rect 13044 26868 13050 26880
rect 13354 26868 13360 26920
rect 13412 26908 13418 26920
rect 13817 26911 13875 26917
rect 13817 26908 13829 26911
rect 13412 26880 13829 26908
rect 13412 26868 13418 26880
rect 13817 26877 13829 26880
rect 13863 26908 13875 26911
rect 14292 26908 14320 26948
rect 13863 26880 14320 26908
rect 14553 26911 14611 26917
rect 13863 26877 13875 26880
rect 13817 26871 13875 26877
rect 14553 26877 14565 26911
rect 14599 26877 14611 26911
rect 14660 26908 14688 26948
rect 14737 26945 14749 26979
rect 14783 26945 14795 26979
rect 14737 26939 14795 26945
rect 15930 26936 15936 26988
rect 15988 26976 15994 26988
rect 16393 26979 16451 26985
rect 16393 26976 16405 26979
rect 15988 26948 16405 26976
rect 15988 26936 15994 26948
rect 16393 26945 16405 26948
rect 16439 26945 16451 26979
rect 16393 26939 16451 26945
rect 16850 26936 16856 26988
rect 16908 26936 16914 26988
rect 17144 26976 17172 27016
rect 17310 27004 17316 27056
rect 17368 27004 17374 27056
rect 18506 27004 18512 27056
rect 18564 27004 18570 27056
rect 18598 27004 18604 27056
rect 18656 27044 18662 27056
rect 19518 27044 19524 27056
rect 18656 27016 19524 27044
rect 18656 27004 18662 27016
rect 17589 26979 17647 26985
rect 17589 26976 17601 26979
rect 17144 26948 17601 26976
rect 17589 26945 17601 26948
rect 17635 26945 17647 26979
rect 17589 26939 17647 26945
rect 18230 26936 18236 26988
rect 18288 26976 18294 26988
rect 18800 26985 18828 27016
rect 19518 27004 19524 27016
rect 19576 27004 19582 27056
rect 20714 27004 20720 27056
rect 20772 27044 20778 27056
rect 23477 27047 23535 27053
rect 20772 27016 23428 27044
rect 20772 27004 20778 27016
rect 18325 26979 18383 26985
rect 18325 26976 18337 26979
rect 18288 26948 18337 26976
rect 18288 26936 18294 26948
rect 18325 26945 18337 26948
rect 18371 26945 18383 26979
rect 18325 26939 18383 26945
rect 18785 26979 18843 26985
rect 18785 26945 18797 26979
rect 18831 26945 18843 26979
rect 18785 26939 18843 26945
rect 19242 26936 19248 26988
rect 19300 26976 19306 26988
rect 19610 26976 19616 26994
rect 19300 26948 19616 26976
rect 19300 26936 19306 26948
rect 19610 26942 19616 26948
rect 19668 26942 19674 26994
rect 19705 26979 19763 26985
rect 19705 26945 19717 26979
rect 19751 26976 19763 26979
rect 19978 26976 19984 26988
rect 19751 26948 19984 26976
rect 19751 26945 19763 26948
rect 19613 26939 19671 26942
rect 19705 26939 19763 26945
rect 19978 26936 19984 26948
rect 20036 26936 20042 26988
rect 20438 26936 20444 26988
rect 20496 26976 20502 26988
rect 20496 26948 21404 26976
rect 20496 26936 20502 26948
rect 15562 26908 15568 26920
rect 14660 26880 15568 26908
rect 14553 26871 14611 26877
rect 13906 26840 13912 26852
rect 8168 26812 8340 26840
rect 8404 26812 13912 26840
rect 8168 26800 8174 26812
rect 3568 26744 4200 26772
rect 3568 26732 3574 26744
rect 4246 26732 4252 26784
rect 4304 26772 4310 26784
rect 4706 26772 4712 26784
rect 4304 26744 4712 26772
rect 4304 26732 4310 26744
rect 4706 26732 4712 26744
rect 4764 26732 4770 26784
rect 4798 26732 4804 26784
rect 4856 26772 4862 26784
rect 5353 26775 5411 26781
rect 5353 26772 5365 26775
rect 4856 26744 5365 26772
rect 4856 26732 4862 26744
rect 5353 26741 5365 26744
rect 5399 26741 5411 26775
rect 5353 26735 5411 26741
rect 5721 26775 5779 26781
rect 5721 26741 5733 26775
rect 5767 26772 5779 26775
rect 5902 26772 5908 26784
rect 5767 26744 5908 26772
rect 5767 26741 5779 26744
rect 5721 26735 5779 26741
rect 5902 26732 5908 26744
rect 5960 26732 5966 26784
rect 5994 26732 6000 26784
rect 6052 26732 6058 26784
rect 6822 26732 6828 26784
rect 6880 26772 6886 26784
rect 7650 26772 7656 26784
rect 6880 26744 7656 26772
rect 6880 26732 6886 26744
rect 7650 26732 7656 26744
rect 7708 26732 7714 26784
rect 7837 26775 7895 26781
rect 7837 26741 7849 26775
rect 7883 26772 7895 26775
rect 8404 26772 8432 26812
rect 13906 26800 13912 26812
rect 13964 26800 13970 26852
rect 13998 26800 14004 26852
rect 14056 26840 14062 26852
rect 14568 26840 14596 26871
rect 15562 26868 15568 26880
rect 15620 26868 15626 26920
rect 17126 26868 17132 26920
rect 17184 26908 17190 26920
rect 17405 26911 17463 26917
rect 17405 26908 17417 26911
rect 17184 26880 17417 26908
rect 17184 26868 17190 26880
rect 17405 26877 17417 26880
rect 17451 26877 17463 26911
rect 17405 26871 17463 26877
rect 18693 26911 18751 26917
rect 18693 26877 18705 26911
rect 18739 26908 18751 26911
rect 19521 26911 19579 26917
rect 19521 26908 19533 26911
rect 18739 26880 19533 26908
rect 18739 26877 18751 26880
rect 18693 26871 18751 26877
rect 19521 26877 19533 26880
rect 19567 26908 19579 26911
rect 19886 26908 19892 26920
rect 19567 26880 19892 26908
rect 19567 26877 19579 26880
rect 19521 26871 19579 26877
rect 19886 26868 19892 26880
rect 19944 26868 19950 26920
rect 20806 26908 20812 26920
rect 20640 26880 20812 26908
rect 14734 26840 14740 26852
rect 14056 26812 14504 26840
rect 14568 26812 14740 26840
rect 14056 26800 14062 26812
rect 7883 26744 8432 26772
rect 7883 26741 7895 26744
rect 7837 26735 7895 26741
rect 8478 26732 8484 26784
rect 8536 26732 8542 26784
rect 8570 26732 8576 26784
rect 8628 26772 8634 26784
rect 8665 26775 8723 26781
rect 8665 26772 8677 26775
rect 8628 26744 8677 26772
rect 8628 26732 8634 26744
rect 8665 26741 8677 26744
rect 8711 26741 8723 26775
rect 8665 26735 8723 26741
rect 9858 26732 9864 26784
rect 9916 26732 9922 26784
rect 10226 26732 10232 26784
rect 10284 26772 10290 26784
rect 10505 26775 10563 26781
rect 10505 26772 10517 26775
rect 10284 26744 10517 26772
rect 10284 26732 10290 26744
rect 10505 26741 10517 26744
rect 10551 26741 10563 26775
rect 10505 26735 10563 26741
rect 10778 26732 10784 26784
rect 10836 26772 10842 26784
rect 10873 26775 10931 26781
rect 10873 26772 10885 26775
rect 10836 26744 10885 26772
rect 10836 26732 10842 26744
rect 10873 26741 10885 26744
rect 10919 26741 10931 26775
rect 10873 26735 10931 26741
rect 12986 26732 12992 26784
rect 13044 26732 13050 26784
rect 13538 26732 13544 26784
rect 13596 26732 13602 26784
rect 13725 26775 13783 26781
rect 13725 26741 13737 26775
rect 13771 26772 13783 26775
rect 13814 26772 13820 26784
rect 13771 26744 13820 26772
rect 13771 26741 13783 26744
rect 13725 26735 13783 26741
rect 13814 26732 13820 26744
rect 13872 26732 13878 26784
rect 14476 26781 14504 26812
rect 14734 26800 14740 26812
rect 14792 26800 14798 26852
rect 16482 26800 16488 26852
rect 16540 26840 16546 26852
rect 17037 26843 17095 26849
rect 17037 26840 17049 26843
rect 16540 26812 17049 26840
rect 16540 26800 16546 26812
rect 17037 26809 17049 26812
rect 17083 26840 17095 26843
rect 17083 26812 17908 26840
rect 17083 26809 17095 26812
rect 17037 26803 17095 26809
rect 14461 26775 14519 26781
rect 14461 26741 14473 26775
rect 14507 26741 14519 26775
rect 14461 26735 14519 26741
rect 16022 26732 16028 26784
rect 16080 26772 16086 26784
rect 16209 26775 16267 26781
rect 16209 26772 16221 26775
rect 16080 26744 16221 26772
rect 16080 26732 16086 26744
rect 16209 26741 16221 26744
rect 16255 26741 16267 26775
rect 16209 26735 16267 26741
rect 17402 26732 17408 26784
rect 17460 26732 17466 26784
rect 17770 26732 17776 26784
rect 17828 26732 17834 26784
rect 17880 26772 17908 26812
rect 18782 26800 18788 26852
rect 18840 26840 18846 26852
rect 18969 26843 19027 26849
rect 18969 26840 18981 26843
rect 18840 26812 18981 26840
rect 18840 26800 18846 26812
rect 18969 26809 18981 26812
rect 19015 26809 19027 26843
rect 18969 26803 19027 26809
rect 19242 26800 19248 26852
rect 19300 26800 19306 26852
rect 20640 26840 20668 26880
rect 20806 26868 20812 26880
rect 20864 26868 20870 26920
rect 19904 26812 20668 26840
rect 21376 26840 21404 26948
rect 21450 26936 21456 26988
rect 21508 26976 21514 26988
rect 22465 26979 22523 26985
rect 22465 26976 22477 26979
rect 21508 26948 22477 26976
rect 21508 26936 21514 26948
rect 22465 26945 22477 26948
rect 22511 26945 22523 26979
rect 22465 26939 22523 26945
rect 22554 26936 22560 26988
rect 22612 26976 22618 26988
rect 22649 26979 22707 26985
rect 22649 26976 22661 26979
rect 22612 26948 22661 26976
rect 22612 26936 22618 26948
rect 22649 26945 22661 26948
rect 22695 26945 22707 26979
rect 22649 26939 22707 26945
rect 23290 26936 23296 26988
rect 23348 26936 23354 26988
rect 23400 26976 23428 27016
rect 23477 27013 23489 27047
rect 23523 27044 23535 27047
rect 23750 27044 23756 27056
rect 23523 27016 23756 27044
rect 23523 27013 23535 27016
rect 23477 27007 23535 27013
rect 23750 27004 23756 27016
rect 23808 27004 23814 27056
rect 25148 26985 25176 27084
rect 28258 27072 28264 27124
rect 28316 27072 28322 27124
rect 23569 26979 23627 26985
rect 23569 26976 23581 26979
rect 23400 26948 23581 26976
rect 23569 26945 23581 26948
rect 23615 26945 23627 26979
rect 23569 26939 23627 26945
rect 24949 26979 25007 26985
rect 24949 26945 24961 26979
rect 24995 26945 25007 26979
rect 24949 26939 25007 26945
rect 25133 26979 25191 26985
rect 25133 26945 25145 26979
rect 25179 26945 25191 26979
rect 25133 26939 25191 26945
rect 25225 26979 25283 26985
rect 25225 26945 25237 26979
rect 25271 26976 25283 26979
rect 25406 26976 25412 26988
rect 25271 26948 25412 26976
rect 25271 26945 25283 26948
rect 25225 26939 25283 26945
rect 22002 26840 22008 26852
rect 21376 26812 22008 26840
rect 19904 26784 19932 26812
rect 22002 26800 22008 26812
rect 22060 26840 22066 26852
rect 24964 26840 24992 26939
rect 25406 26936 25412 26948
rect 25464 26936 25470 26988
rect 25590 26936 25596 26988
rect 25648 26936 25654 26988
rect 25869 26979 25927 26985
rect 25869 26945 25881 26979
rect 25915 26976 25927 26979
rect 25958 26976 25964 26988
rect 25915 26948 25964 26976
rect 25915 26945 25927 26948
rect 25869 26939 25927 26945
rect 25958 26936 25964 26948
rect 26016 26936 26022 26988
rect 26970 26936 26976 26988
rect 27028 26936 27034 26988
rect 27246 26936 27252 26988
rect 27304 26936 27310 26988
rect 28276 26976 28304 27072
rect 29914 27004 29920 27056
rect 29972 27044 29978 27056
rect 31205 27047 31263 27053
rect 31205 27044 31217 27047
rect 29972 27016 31217 27044
rect 29972 27004 29978 27016
rect 31205 27013 31217 27016
rect 31251 27013 31263 27047
rect 31205 27007 31263 27013
rect 28629 26979 28687 26985
rect 28629 26976 28641 26979
rect 28276 26948 28641 26976
rect 28629 26945 28641 26948
rect 28675 26945 28687 26979
rect 28629 26939 28687 26945
rect 30926 26936 30932 26988
rect 30984 26936 30990 26988
rect 31113 26979 31171 26985
rect 31113 26945 31125 26979
rect 31159 26945 31171 26979
rect 31113 26939 31171 26945
rect 25685 26911 25743 26917
rect 25685 26877 25697 26911
rect 25731 26877 25743 26911
rect 25685 26871 25743 26877
rect 22060 26812 24992 26840
rect 25409 26843 25467 26849
rect 22060 26800 22066 26812
rect 25409 26809 25421 26843
rect 25455 26840 25467 26843
rect 25700 26840 25728 26871
rect 30374 26868 30380 26920
rect 30432 26908 30438 26920
rect 31128 26908 31156 26939
rect 31294 26936 31300 26988
rect 31352 26936 31358 26988
rect 32490 26936 32496 26988
rect 32548 26936 32554 26988
rect 30432 26880 31156 26908
rect 30432 26868 30438 26880
rect 25455 26812 25728 26840
rect 25455 26809 25467 26812
rect 25409 26803 25467 26809
rect 27062 26800 27068 26852
rect 27120 26840 27126 26852
rect 29822 26840 29828 26852
rect 27120 26812 29828 26840
rect 27120 26800 27126 26812
rect 29822 26800 29828 26812
rect 29880 26800 29886 26852
rect 19150 26772 19156 26784
rect 17880 26744 19156 26772
rect 19150 26732 19156 26744
rect 19208 26732 19214 26784
rect 19518 26732 19524 26784
rect 19576 26732 19582 26784
rect 19610 26732 19616 26784
rect 19668 26772 19674 26784
rect 19794 26772 19800 26784
rect 19668 26744 19800 26772
rect 19668 26732 19674 26744
rect 19794 26732 19800 26744
rect 19852 26732 19858 26784
rect 19886 26732 19892 26784
rect 19944 26732 19950 26784
rect 20162 26732 20168 26784
rect 20220 26772 20226 26784
rect 22462 26772 22468 26784
rect 20220 26744 22468 26772
rect 20220 26732 20226 26744
rect 22462 26732 22468 26744
rect 22520 26732 22526 26784
rect 22830 26732 22836 26784
rect 22888 26732 22894 26784
rect 23109 26775 23167 26781
rect 23109 26741 23121 26775
rect 23155 26772 23167 26775
rect 23198 26772 23204 26784
rect 23155 26744 23204 26772
rect 23155 26741 23167 26744
rect 23109 26735 23167 26741
rect 23198 26732 23204 26744
rect 23256 26732 23262 26784
rect 23750 26732 23756 26784
rect 23808 26732 23814 26784
rect 25222 26732 25228 26784
rect 25280 26732 25286 26784
rect 25682 26732 25688 26784
rect 25740 26732 25746 26784
rect 26050 26732 26056 26784
rect 26108 26732 26114 26784
rect 27154 26732 27160 26784
rect 27212 26732 27218 26784
rect 27430 26732 27436 26784
rect 27488 26732 27494 26784
rect 28350 26732 28356 26784
rect 28408 26772 28414 26784
rect 28445 26775 28503 26781
rect 28445 26772 28457 26775
rect 28408 26744 28457 26772
rect 28408 26732 28414 26744
rect 28445 26741 28457 26744
rect 28491 26741 28503 26775
rect 28445 26735 28503 26741
rect 31386 26732 31392 26784
rect 31444 26772 31450 26784
rect 31481 26775 31539 26781
rect 31481 26772 31493 26775
rect 31444 26744 31493 26772
rect 31444 26732 31450 26744
rect 31481 26741 31493 26744
rect 31527 26741 31539 26775
rect 31481 26735 31539 26741
rect 31662 26732 31668 26784
rect 31720 26772 31726 26784
rect 32309 26775 32367 26781
rect 32309 26772 32321 26775
rect 31720 26744 32321 26772
rect 31720 26732 31726 26744
rect 32309 26741 32321 26744
rect 32355 26741 32367 26775
rect 32309 26735 32367 26741
rect 1104 26682 32844 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 32844 26682
rect 1104 26608 32844 26630
rect 2777 26571 2835 26577
rect 2777 26537 2789 26571
rect 2823 26568 2835 26571
rect 3786 26568 3792 26580
rect 2823 26540 3792 26568
rect 2823 26537 2835 26540
rect 2777 26531 2835 26537
rect 3786 26528 3792 26540
rect 3844 26528 3850 26580
rect 4154 26528 4160 26580
rect 4212 26568 4218 26580
rect 4890 26568 4896 26580
rect 4212 26540 4896 26568
rect 4212 26528 4218 26540
rect 4890 26528 4896 26540
rect 4948 26528 4954 26580
rect 5445 26571 5503 26577
rect 5445 26537 5457 26571
rect 5491 26568 5503 26571
rect 5534 26568 5540 26580
rect 5491 26540 5540 26568
rect 5491 26537 5503 26540
rect 5445 26531 5503 26537
rect 5534 26528 5540 26540
rect 5592 26528 5598 26580
rect 6730 26568 6736 26580
rect 5828 26540 6736 26568
rect 3694 26460 3700 26512
rect 3752 26500 3758 26512
rect 3881 26503 3939 26509
rect 3881 26500 3893 26503
rect 3752 26472 3893 26500
rect 3752 26460 3758 26472
rect 3881 26469 3893 26472
rect 3927 26469 3939 26503
rect 3881 26463 3939 26469
rect 3970 26460 3976 26512
rect 4028 26500 4034 26512
rect 5074 26500 5080 26512
rect 4028 26472 5080 26500
rect 4028 26460 4034 26472
rect 5074 26460 5080 26472
rect 5132 26460 5138 26512
rect 5169 26503 5227 26509
rect 5169 26469 5181 26503
rect 5215 26500 5227 26503
rect 5828 26500 5856 26540
rect 6730 26528 6736 26540
rect 6788 26528 6794 26580
rect 7006 26528 7012 26580
rect 7064 26568 7070 26580
rect 7834 26568 7840 26580
rect 7064 26540 7840 26568
rect 7064 26528 7070 26540
rect 7834 26528 7840 26540
rect 7892 26528 7898 26580
rect 8110 26528 8116 26580
rect 8168 26528 8174 26580
rect 8938 26528 8944 26580
rect 8996 26568 9002 26580
rect 9398 26568 9404 26580
rect 8996 26540 9404 26568
rect 8996 26528 9002 26540
rect 9398 26528 9404 26540
rect 9456 26528 9462 26580
rect 9858 26528 9864 26580
rect 9916 26568 9922 26580
rect 9916 26540 13584 26568
rect 9916 26528 9922 26540
rect 5215 26472 5580 26500
rect 5215 26469 5227 26472
rect 5169 26463 5227 26469
rect 2866 26392 2872 26444
rect 2924 26432 2930 26444
rect 3329 26435 3387 26441
rect 3329 26432 3341 26435
rect 2924 26404 3341 26432
rect 2924 26392 2930 26404
rect 3329 26401 3341 26404
rect 3375 26401 3387 26435
rect 3329 26395 3387 26401
rect 1394 26324 1400 26376
rect 1452 26324 1458 26376
rect 2958 26324 2964 26376
rect 3016 26324 3022 26376
rect 3344 26364 3372 26395
rect 4062 26392 4068 26444
rect 4120 26432 4126 26444
rect 4341 26435 4399 26441
rect 4341 26432 4353 26435
rect 4120 26404 4353 26432
rect 4120 26392 4126 26404
rect 4341 26401 4353 26404
rect 4387 26401 4399 26435
rect 4341 26395 4399 26401
rect 4522 26392 4528 26444
rect 4580 26432 4586 26444
rect 5350 26432 5356 26444
rect 4580 26404 5356 26432
rect 4580 26392 4586 26404
rect 4433 26367 4491 26373
rect 3344 26336 3924 26364
rect 1670 26305 1676 26308
rect 1664 26259 1676 26305
rect 1670 26256 1676 26259
rect 1728 26256 1734 26308
rect 2774 26256 2780 26308
rect 2832 26296 2838 26308
rect 3446 26299 3504 26305
rect 3446 26296 3458 26299
rect 2832 26268 3458 26296
rect 2832 26256 2838 26268
rect 3446 26265 3458 26268
rect 3492 26296 3504 26299
rect 3694 26296 3700 26308
rect 3492 26268 3700 26296
rect 3492 26265 3504 26268
rect 3446 26259 3504 26265
rect 3694 26256 3700 26268
rect 3752 26256 3758 26308
rect 3896 26305 3924 26336
rect 4433 26333 4445 26367
rect 4479 26364 4491 26367
rect 4614 26364 4620 26376
rect 4479 26336 4620 26364
rect 4479 26333 4491 26336
rect 4433 26327 4491 26333
rect 4614 26324 4620 26336
rect 4672 26324 4678 26376
rect 4706 26324 4712 26376
rect 4764 26324 4770 26376
rect 5000 26373 5028 26404
rect 5350 26392 5356 26404
rect 5408 26392 5414 26444
rect 5552 26376 5580 26472
rect 5736 26472 5856 26500
rect 6089 26503 6147 26509
rect 4985 26367 5043 26373
rect 4985 26333 4997 26367
rect 5031 26333 5043 26367
rect 4985 26327 5043 26333
rect 5258 26324 5264 26376
rect 5316 26324 5322 26376
rect 5534 26324 5540 26376
rect 5592 26324 5598 26376
rect 5736 26373 5764 26472
rect 6089 26469 6101 26503
rect 6135 26500 6147 26503
rect 6178 26500 6184 26512
rect 6135 26472 6184 26500
rect 6135 26469 6147 26472
rect 6089 26463 6147 26469
rect 6178 26460 6184 26472
rect 6236 26460 6242 26512
rect 6362 26460 6368 26512
rect 6420 26500 6426 26512
rect 6641 26503 6699 26509
rect 6641 26500 6653 26503
rect 6420 26472 6653 26500
rect 6420 26460 6426 26472
rect 6641 26469 6653 26472
rect 6687 26469 6699 26503
rect 6641 26463 6699 26469
rect 6380 26432 6408 26460
rect 5828 26404 6408 26432
rect 5828 26373 5856 26404
rect 5721 26367 5779 26373
rect 5721 26333 5733 26367
rect 5767 26333 5779 26367
rect 5721 26327 5779 26333
rect 5813 26367 5871 26373
rect 5813 26333 5825 26367
rect 5859 26333 5871 26367
rect 5813 26327 5871 26333
rect 5905 26367 5963 26373
rect 5905 26333 5917 26367
rect 5951 26364 5963 26367
rect 6178 26364 6184 26376
rect 5951 26336 6184 26364
rect 5951 26333 5963 26336
rect 5905 26327 5963 26333
rect 6178 26324 6184 26336
rect 6236 26324 6242 26376
rect 6365 26367 6423 26373
rect 6365 26333 6377 26367
rect 6411 26333 6423 26367
rect 6365 26327 6423 26333
rect 3881 26299 3939 26305
rect 3881 26265 3893 26299
rect 3927 26265 3939 26299
rect 6380 26296 6408 26327
rect 6454 26324 6460 26376
rect 6512 26364 6518 26376
rect 7024 26373 7052 26528
rect 7561 26503 7619 26509
rect 7561 26469 7573 26503
rect 7607 26500 7619 26503
rect 7607 26472 11008 26500
rect 7607 26469 7619 26472
rect 7561 26463 7619 26469
rect 7282 26392 7288 26444
rect 7340 26432 7346 26444
rect 7340 26404 7696 26432
rect 7340 26392 7346 26404
rect 7668 26373 7696 26404
rect 9306 26392 9312 26444
rect 9364 26432 9370 26444
rect 10134 26432 10140 26444
rect 9364 26404 10140 26432
rect 9364 26392 9370 26404
rect 10134 26392 10140 26404
rect 10192 26392 10198 26444
rect 10980 26432 11008 26472
rect 11054 26460 11060 26512
rect 11112 26500 11118 26512
rect 11149 26503 11207 26509
rect 11149 26500 11161 26503
rect 11112 26472 11161 26500
rect 11112 26460 11118 26472
rect 11149 26469 11161 26472
rect 11195 26469 11207 26503
rect 12250 26500 12256 26512
rect 11149 26463 11207 26469
rect 11716 26472 12256 26500
rect 11716 26432 11744 26472
rect 12250 26460 12256 26472
rect 12308 26460 12314 26512
rect 13078 26500 13084 26512
rect 12406 26472 13084 26500
rect 12406 26432 12434 26472
rect 13078 26460 13084 26472
rect 13136 26460 13142 26512
rect 10980 26404 11744 26432
rect 11808 26404 12434 26432
rect 13556 26432 13584 26540
rect 13630 26528 13636 26580
rect 13688 26568 13694 26580
rect 14826 26568 14832 26580
rect 13688 26540 14832 26568
rect 13688 26528 13694 26540
rect 14826 26528 14832 26540
rect 14884 26528 14890 26580
rect 15010 26528 15016 26580
rect 15068 26528 15074 26580
rect 15194 26528 15200 26580
rect 15252 26528 15258 26580
rect 16022 26528 16028 26580
rect 16080 26528 16086 26580
rect 18141 26571 18199 26577
rect 16224 26540 17954 26568
rect 13909 26503 13967 26509
rect 13909 26469 13921 26503
rect 13955 26500 13967 26503
rect 14182 26500 14188 26512
rect 13955 26472 14188 26500
rect 13955 26469 13967 26472
rect 13909 26463 13967 26469
rect 14182 26460 14188 26472
rect 14240 26500 14246 26512
rect 14458 26500 14464 26512
rect 14240 26472 14464 26500
rect 14240 26460 14246 26472
rect 14458 26460 14464 26472
rect 14516 26460 14522 26512
rect 16224 26500 16252 26540
rect 14752 26472 16252 26500
rect 16485 26503 16543 26509
rect 14752 26432 14780 26472
rect 16485 26469 16497 26503
rect 16531 26500 16543 26503
rect 17402 26500 17408 26512
rect 16531 26472 17408 26500
rect 16531 26469 16543 26472
rect 16485 26463 16543 26469
rect 17402 26460 17408 26472
rect 17460 26460 17466 26512
rect 17926 26500 17954 26540
rect 18141 26537 18153 26571
rect 18187 26568 18199 26571
rect 18414 26568 18420 26580
rect 18187 26540 18420 26568
rect 18187 26537 18199 26540
rect 18141 26531 18199 26537
rect 18414 26528 18420 26540
rect 18472 26568 18478 26580
rect 19518 26568 19524 26580
rect 18472 26540 19524 26568
rect 18472 26528 18478 26540
rect 19518 26528 19524 26540
rect 19576 26568 19582 26580
rect 19576 26540 20300 26568
rect 19576 26528 19582 26540
rect 18690 26500 18696 26512
rect 17926 26472 18696 26500
rect 13556 26404 14780 26432
rect 6825 26367 6883 26373
rect 6825 26364 6837 26367
rect 6512 26336 6837 26364
rect 6512 26324 6518 26336
rect 6825 26333 6837 26336
rect 6871 26333 6883 26367
rect 6825 26327 6883 26333
rect 7009 26367 7067 26373
rect 7009 26333 7021 26367
rect 7055 26333 7067 26367
rect 7377 26367 7435 26373
rect 7377 26364 7389 26367
rect 7009 26327 7067 26333
rect 7116 26336 7389 26364
rect 6914 26296 6920 26308
rect 3881 26259 3939 26265
rect 5736 26268 6408 26296
rect 6472 26268 6920 26296
rect 5736 26240 5764 26268
rect 3142 26188 3148 26240
rect 3200 26228 3206 26240
rect 3237 26231 3295 26237
rect 3237 26228 3249 26231
rect 3200 26200 3249 26228
rect 3200 26188 3206 26200
rect 3237 26197 3249 26200
rect 3283 26197 3295 26231
rect 3237 26191 3295 26197
rect 3605 26231 3663 26237
rect 3605 26197 3617 26231
rect 3651 26228 3663 26231
rect 3970 26228 3976 26240
rect 3651 26200 3976 26228
rect 3651 26197 3663 26200
rect 3605 26191 3663 26197
rect 3970 26188 3976 26200
rect 4028 26188 4034 26240
rect 4617 26231 4675 26237
rect 4617 26197 4629 26231
rect 4663 26228 4675 26231
rect 5626 26228 5632 26240
rect 4663 26200 5632 26228
rect 4663 26197 4675 26200
rect 4617 26191 4675 26197
rect 5626 26188 5632 26200
rect 5684 26188 5690 26240
rect 5718 26188 5724 26240
rect 5776 26188 5782 26240
rect 6178 26188 6184 26240
rect 6236 26228 6242 26240
rect 6472 26228 6500 26268
rect 6914 26256 6920 26268
rect 6972 26296 6978 26308
rect 7116 26296 7144 26336
rect 7377 26333 7389 26336
rect 7423 26333 7435 26367
rect 7377 26327 7435 26333
rect 7653 26367 7711 26373
rect 7653 26333 7665 26367
rect 7699 26333 7711 26367
rect 7653 26327 7711 26333
rect 7742 26324 7748 26376
rect 7800 26364 7806 26376
rect 7929 26367 7987 26373
rect 7929 26364 7941 26367
rect 7800 26336 7941 26364
rect 7800 26324 7806 26336
rect 7929 26333 7941 26336
rect 7975 26333 7987 26367
rect 7929 26327 7987 26333
rect 8294 26324 8300 26376
rect 8352 26364 8358 26376
rect 8941 26367 8999 26373
rect 8941 26364 8953 26367
rect 8352 26336 8953 26364
rect 8352 26324 8358 26336
rect 8941 26333 8953 26336
rect 8987 26333 8999 26367
rect 8941 26327 8999 26333
rect 9214 26324 9220 26376
rect 9272 26324 9278 26376
rect 9861 26367 9919 26373
rect 9861 26364 9873 26367
rect 9324 26336 9873 26364
rect 6972 26268 7144 26296
rect 7193 26299 7251 26305
rect 6972 26256 6978 26268
rect 7193 26265 7205 26299
rect 7239 26265 7251 26299
rect 7193 26259 7251 26265
rect 6236 26200 6500 26228
rect 6549 26231 6607 26237
rect 6236 26188 6242 26200
rect 6549 26197 6561 26231
rect 6595 26228 6607 26231
rect 6638 26228 6644 26240
rect 6595 26200 6644 26228
rect 6595 26197 6607 26200
rect 6549 26191 6607 26197
rect 6638 26188 6644 26200
rect 6696 26188 6702 26240
rect 6730 26188 6736 26240
rect 6788 26228 6794 26240
rect 7208 26228 7236 26259
rect 7282 26256 7288 26308
rect 7340 26296 7346 26308
rect 8110 26296 8116 26308
rect 7340 26268 8116 26296
rect 7340 26256 7346 26268
rect 8110 26256 8116 26268
rect 8168 26256 8174 26308
rect 9324 26296 9352 26336
rect 9861 26333 9873 26336
rect 9907 26333 9919 26367
rect 9861 26327 9919 26333
rect 10321 26367 10379 26373
rect 10321 26333 10333 26367
rect 10367 26364 10379 26367
rect 10686 26364 10692 26376
rect 10367 26336 10692 26364
rect 10367 26333 10379 26336
rect 10321 26327 10379 26333
rect 10686 26324 10692 26336
rect 10744 26324 10750 26376
rect 10778 26324 10784 26376
rect 10836 26364 10842 26376
rect 11238 26364 11244 26376
rect 10836 26336 11244 26364
rect 10836 26324 10842 26336
rect 11238 26324 11244 26336
rect 11296 26324 11302 26376
rect 11333 26367 11391 26373
rect 11333 26333 11345 26367
rect 11379 26333 11391 26367
rect 11333 26327 11391 26333
rect 8312 26268 9352 26296
rect 8312 26240 8340 26268
rect 9490 26256 9496 26308
rect 9548 26296 9554 26308
rect 9548 26268 10180 26296
rect 9548 26256 9554 26268
rect 7466 26228 7472 26240
rect 6788 26200 7472 26228
rect 6788 26188 6794 26200
rect 7466 26188 7472 26200
rect 7524 26188 7530 26240
rect 8294 26188 8300 26240
rect 8352 26188 8358 26240
rect 8754 26188 8760 26240
rect 8812 26228 8818 26240
rect 9125 26231 9183 26237
rect 9125 26228 9137 26231
rect 8812 26200 9137 26228
rect 8812 26188 8818 26200
rect 9125 26197 9137 26200
rect 9171 26197 9183 26231
rect 9125 26191 9183 26197
rect 9214 26188 9220 26240
rect 9272 26228 9278 26240
rect 9401 26231 9459 26237
rect 9401 26228 9413 26231
rect 9272 26200 9413 26228
rect 9272 26188 9278 26200
rect 9401 26197 9413 26200
rect 9447 26197 9459 26231
rect 9401 26191 9459 26197
rect 10042 26188 10048 26240
rect 10100 26188 10106 26240
rect 10152 26237 10180 26268
rect 11348 26240 11376 26327
rect 11698 26324 11704 26376
rect 11756 26324 11762 26376
rect 11808 26373 11836 26404
rect 14826 26392 14832 26444
rect 14884 26392 14890 26444
rect 18049 26435 18107 26441
rect 18049 26401 18061 26435
rect 18095 26432 18107 26435
rect 18417 26435 18475 26441
rect 18417 26432 18429 26435
rect 18095 26404 18429 26432
rect 18095 26401 18107 26404
rect 18049 26395 18107 26401
rect 18417 26401 18429 26404
rect 18463 26432 18475 26435
rect 18463 26404 18552 26432
rect 18463 26401 18475 26404
rect 18417 26395 18475 26401
rect 11793 26367 11851 26373
rect 11793 26333 11805 26367
rect 11839 26333 11851 26367
rect 11793 26327 11851 26333
rect 11882 26324 11888 26376
rect 11940 26364 11946 26376
rect 12161 26367 12219 26373
rect 12161 26364 12173 26367
rect 11940 26336 12173 26364
rect 11940 26324 11946 26336
rect 12161 26333 12173 26336
rect 12207 26333 12219 26367
rect 12161 26327 12219 26333
rect 12710 26324 12716 26376
rect 12768 26364 12774 26376
rect 12768 26336 12940 26364
rect 12768 26324 12774 26336
rect 11422 26256 11428 26308
rect 11480 26256 11486 26308
rect 11514 26256 11520 26308
rect 11572 26296 11578 26308
rect 11977 26299 12035 26305
rect 11977 26296 11989 26299
rect 11572 26268 11989 26296
rect 11572 26256 11578 26268
rect 11977 26265 11989 26268
rect 12023 26265 12035 26299
rect 11977 26259 12035 26265
rect 12069 26299 12127 26305
rect 12069 26265 12081 26299
rect 12115 26296 12127 26299
rect 12802 26296 12808 26308
rect 12115 26268 12808 26296
rect 12115 26265 12127 26268
rect 12069 26259 12127 26265
rect 12802 26256 12808 26268
rect 12860 26256 12866 26308
rect 12912 26296 12940 26336
rect 13354 26324 13360 26376
rect 13412 26364 13418 26376
rect 13449 26367 13507 26373
rect 13449 26364 13461 26367
rect 13412 26336 13461 26364
rect 13412 26324 13418 26336
rect 13449 26333 13461 26336
rect 13495 26333 13507 26367
rect 13449 26327 13507 26333
rect 13722 26324 13728 26376
rect 13780 26324 13786 26376
rect 15010 26324 15016 26376
rect 15068 26324 15074 26376
rect 15286 26324 15292 26376
rect 15344 26364 15350 26376
rect 16209 26367 16267 26373
rect 16209 26364 16221 26367
rect 15344 26336 16221 26364
rect 15344 26324 15350 26336
rect 16209 26333 16221 26336
rect 16255 26333 16267 26367
rect 16209 26327 16267 26333
rect 14737 26299 14795 26305
rect 12912 26268 14688 26296
rect 10137 26231 10195 26237
rect 10137 26197 10149 26231
rect 10183 26197 10195 26231
rect 10137 26191 10195 26197
rect 11330 26188 11336 26240
rect 11388 26228 11394 26240
rect 11882 26228 11888 26240
rect 11388 26200 11888 26228
rect 11388 26188 11394 26200
rect 11882 26188 11888 26200
rect 11940 26188 11946 26240
rect 12345 26231 12403 26237
rect 12345 26197 12357 26231
rect 12391 26228 12403 26231
rect 13170 26228 13176 26240
rect 12391 26200 13176 26228
rect 12391 26197 12403 26200
rect 12345 26191 12403 26197
rect 13170 26188 13176 26200
rect 13228 26188 13234 26240
rect 14660 26228 14688 26268
rect 14737 26265 14749 26299
rect 14783 26296 14795 26299
rect 14826 26296 14832 26308
rect 14783 26268 14832 26296
rect 14783 26265 14795 26268
rect 14737 26259 14795 26265
rect 14826 26256 14832 26268
rect 14884 26256 14890 26308
rect 16025 26299 16083 26305
rect 14936 26268 15976 26296
rect 14936 26228 14964 26268
rect 14660 26200 14964 26228
rect 15948 26228 15976 26268
rect 16025 26265 16037 26299
rect 16071 26296 16083 26299
rect 16114 26296 16120 26308
rect 16071 26268 16120 26296
rect 16071 26265 16083 26268
rect 16025 26259 16083 26265
rect 16114 26256 16120 26268
rect 16172 26256 16178 26308
rect 16224 26296 16252 26327
rect 16298 26324 16304 26376
rect 16356 26324 16362 26376
rect 18141 26367 18199 26373
rect 18141 26333 18153 26367
rect 18187 26364 18199 26367
rect 18230 26364 18236 26376
rect 18187 26336 18236 26364
rect 18187 26333 18199 26336
rect 18141 26327 18199 26333
rect 18230 26324 18236 26336
rect 18288 26324 18294 26376
rect 16482 26296 16488 26308
rect 16224 26268 16488 26296
rect 16482 26256 16488 26268
rect 16540 26256 16546 26308
rect 17218 26296 17224 26308
rect 16592 26268 17224 26296
rect 16592 26228 16620 26268
rect 17218 26256 17224 26268
rect 17276 26256 17282 26308
rect 17586 26256 17592 26308
rect 17644 26296 17650 26308
rect 17865 26299 17923 26305
rect 17865 26296 17877 26299
rect 17644 26268 17877 26296
rect 17644 26256 17650 26268
rect 17865 26265 17877 26268
rect 17911 26265 17923 26299
rect 18524 26296 18552 26404
rect 18616 26373 18644 26472
rect 18690 26460 18696 26472
rect 18748 26500 18754 26512
rect 20162 26500 20168 26512
rect 18748 26472 20168 26500
rect 18748 26460 18754 26472
rect 20162 26460 20168 26472
rect 20220 26460 20226 26512
rect 20272 26500 20300 26540
rect 22830 26528 22836 26580
rect 22888 26568 22894 26580
rect 23109 26571 23167 26577
rect 23109 26568 23121 26571
rect 22888 26540 23121 26568
rect 22888 26528 22894 26540
rect 23109 26537 23121 26540
rect 23155 26537 23167 26571
rect 24854 26568 24860 26580
rect 23109 26531 23167 26537
rect 23216 26540 24860 26568
rect 21358 26500 21364 26512
rect 20272 26472 21364 26500
rect 21358 26460 21364 26472
rect 21416 26460 21422 26512
rect 21637 26503 21695 26509
rect 21637 26469 21649 26503
rect 21683 26500 21695 26503
rect 21726 26500 21732 26512
rect 21683 26472 21732 26500
rect 21683 26469 21695 26472
rect 21637 26463 21695 26469
rect 21726 26460 21732 26472
rect 21784 26500 21790 26512
rect 23216 26500 23244 26540
rect 24854 26528 24860 26540
rect 24912 26528 24918 26580
rect 25590 26528 25596 26580
rect 25648 26568 25654 26580
rect 26605 26571 26663 26577
rect 26605 26568 26617 26571
rect 25648 26540 26617 26568
rect 25648 26528 25654 26540
rect 26605 26537 26617 26540
rect 26651 26537 26663 26571
rect 26605 26531 26663 26537
rect 26970 26528 26976 26580
rect 27028 26528 27034 26580
rect 27430 26528 27436 26580
rect 27488 26568 27494 26580
rect 27617 26571 27675 26577
rect 27617 26568 27629 26571
rect 27488 26540 27629 26568
rect 27488 26528 27494 26540
rect 27617 26537 27629 26540
rect 27663 26537 27675 26571
rect 27617 26531 27675 26537
rect 21784 26472 23244 26500
rect 21784 26460 21790 26472
rect 23474 26460 23480 26512
rect 23532 26500 23538 26512
rect 23569 26503 23627 26509
rect 23569 26500 23581 26503
rect 23532 26472 23581 26500
rect 23532 26460 23538 26472
rect 23569 26469 23581 26472
rect 23615 26469 23627 26503
rect 23569 26463 23627 26469
rect 25682 26460 25688 26512
rect 25740 26500 25746 26512
rect 25958 26500 25964 26512
rect 25740 26472 25964 26500
rect 25740 26460 25746 26472
rect 25958 26460 25964 26472
rect 26016 26460 26022 26512
rect 27632 26500 27660 26531
rect 27890 26528 27896 26580
rect 27948 26528 27954 26580
rect 28350 26528 28356 26580
rect 28408 26528 28414 26580
rect 31294 26528 31300 26580
rect 31352 26568 31358 26580
rect 31849 26571 31907 26577
rect 31849 26568 31861 26571
rect 31352 26540 31861 26568
rect 31352 26528 31358 26540
rect 31849 26537 31861 26540
rect 31895 26537 31907 26571
rect 31849 26531 31907 26537
rect 27632 26472 28396 26500
rect 19886 26432 19892 26444
rect 18708 26404 19892 26432
rect 18708 26376 18736 26404
rect 19886 26392 19892 26404
rect 19944 26392 19950 26444
rect 19978 26392 19984 26444
rect 20036 26432 20042 26444
rect 21910 26432 21916 26444
rect 20036 26404 21916 26432
rect 20036 26392 20042 26404
rect 21910 26392 21916 26404
rect 21968 26392 21974 26444
rect 22738 26392 22744 26444
rect 22796 26432 22802 26444
rect 23017 26435 23075 26441
rect 23017 26432 23029 26435
rect 22796 26404 23029 26432
rect 22796 26392 22802 26404
rect 23017 26401 23029 26404
rect 23063 26401 23075 26435
rect 23017 26395 23075 26401
rect 18601 26367 18659 26373
rect 18601 26333 18613 26367
rect 18647 26333 18659 26367
rect 18601 26327 18659 26333
rect 18690 26324 18696 26376
rect 18748 26324 18754 26376
rect 18782 26324 18788 26376
rect 18840 26324 18846 26376
rect 18874 26324 18880 26376
rect 18932 26364 18938 26376
rect 20438 26364 20444 26376
rect 18932 26336 20444 26364
rect 18932 26324 18938 26336
rect 20438 26324 20444 26336
rect 20496 26324 20502 26376
rect 21361 26367 21419 26373
rect 20824 26336 21312 26364
rect 20824 26296 20852 26336
rect 18524 26268 20852 26296
rect 17865 26259 17923 26265
rect 21174 26256 21180 26308
rect 21232 26256 21238 26308
rect 21284 26296 21312 26336
rect 21361 26333 21373 26367
rect 21407 26364 21419 26367
rect 21726 26364 21732 26376
rect 21407 26336 21732 26364
rect 21407 26333 21419 26336
rect 21361 26327 21419 26333
rect 21726 26324 21732 26336
rect 21784 26324 21790 26376
rect 21818 26324 21824 26376
rect 21876 26324 21882 26376
rect 23032 26360 23060 26395
rect 23198 26392 23204 26444
rect 23256 26392 23262 26444
rect 23750 26392 23756 26444
rect 23808 26432 23814 26444
rect 26881 26435 26939 26441
rect 26881 26432 26893 26435
rect 23808 26404 26893 26432
rect 23808 26392 23814 26404
rect 26881 26401 26893 26404
rect 26927 26401 26939 26435
rect 26881 26395 26939 26401
rect 26970 26392 26976 26444
rect 27028 26432 27034 26444
rect 27890 26432 27896 26444
rect 27028 26404 27896 26432
rect 27028 26392 27034 26404
rect 23109 26367 23167 26373
rect 23109 26360 23121 26367
rect 23032 26333 23121 26360
rect 23155 26333 23167 26367
rect 23032 26332 23167 26333
rect 23109 26327 23167 26332
rect 23385 26367 23443 26373
rect 23385 26333 23397 26367
rect 23431 26364 23443 26367
rect 24302 26364 24308 26376
rect 23431 26336 24308 26364
rect 23431 26333 23443 26336
rect 23385 26327 23443 26333
rect 24302 26324 24308 26336
rect 24360 26324 24366 26376
rect 26789 26367 26847 26373
rect 26789 26333 26801 26367
rect 26835 26364 26847 26367
rect 27154 26364 27160 26376
rect 26835 26336 27160 26364
rect 26835 26333 26847 26336
rect 26789 26327 26847 26333
rect 27154 26324 27160 26336
rect 27212 26364 27218 26376
rect 27632 26373 27660 26404
rect 27890 26392 27896 26404
rect 27948 26432 27954 26444
rect 28368 26441 28396 26472
rect 28442 26460 28448 26512
rect 28500 26500 28506 26512
rect 28721 26503 28779 26509
rect 28721 26500 28733 26503
rect 28500 26472 28733 26500
rect 28500 26460 28506 26472
rect 28721 26469 28733 26472
rect 28767 26469 28779 26503
rect 28721 26463 28779 26469
rect 28353 26435 28411 26441
rect 27948 26404 28304 26432
rect 27948 26392 27954 26404
rect 27525 26367 27583 26373
rect 27525 26364 27537 26367
rect 27212 26336 27537 26364
rect 27212 26324 27218 26336
rect 27525 26333 27537 26336
rect 27571 26333 27583 26367
rect 27525 26327 27583 26333
rect 27617 26367 27675 26373
rect 27617 26333 27629 26367
rect 27663 26333 27675 26367
rect 27617 26327 27675 26333
rect 21542 26296 21548 26308
rect 21284 26268 21548 26296
rect 21542 26256 21548 26268
rect 21600 26256 21606 26308
rect 23290 26256 23296 26308
rect 23348 26296 23354 26308
rect 25314 26296 25320 26308
rect 23348 26268 25320 26296
rect 23348 26256 23354 26268
rect 25314 26256 25320 26268
rect 25372 26256 25378 26308
rect 27062 26256 27068 26308
rect 27120 26256 27126 26308
rect 27540 26296 27568 26327
rect 27706 26324 27712 26376
rect 27764 26324 27770 26376
rect 28276 26373 28304 26404
rect 28353 26401 28365 26435
rect 28399 26401 28411 26435
rect 28353 26395 28411 26401
rect 28261 26367 28319 26373
rect 28261 26333 28273 26367
rect 28307 26333 28319 26367
rect 28537 26367 28595 26373
rect 28537 26364 28549 26367
rect 28261 26327 28319 26333
rect 28368 26336 28549 26364
rect 27540 26268 27844 26296
rect 15948 26200 16620 26228
rect 18322 26188 18328 26240
rect 18380 26188 18386 26240
rect 18506 26188 18512 26240
rect 18564 26228 18570 26240
rect 22830 26228 22836 26240
rect 18564 26200 22836 26228
rect 18564 26188 18570 26200
rect 22830 26188 22836 26200
rect 22888 26188 22894 26240
rect 27246 26188 27252 26240
rect 27304 26188 27310 26240
rect 27816 26228 27844 26268
rect 28368 26228 28396 26336
rect 28537 26333 28549 26336
rect 28583 26364 28595 26367
rect 29270 26364 29276 26376
rect 28583 26336 29276 26364
rect 28583 26333 28595 26336
rect 28537 26327 28595 26333
rect 29270 26324 29276 26336
rect 29328 26324 29334 26376
rect 31573 26367 31631 26373
rect 31573 26333 31585 26367
rect 31619 26364 31631 26367
rect 31754 26364 31760 26376
rect 31619 26336 31760 26364
rect 31619 26333 31631 26336
rect 31573 26327 31631 26333
rect 31754 26324 31760 26336
rect 31812 26324 31818 26376
rect 32490 26324 32496 26376
rect 32548 26324 32554 26376
rect 27816 26200 28396 26228
rect 30926 26188 30932 26240
rect 30984 26188 30990 26240
rect 1104 26138 32844 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 32844 26138
rect 1104 26064 32844 26086
rect 1581 26027 1639 26033
rect 1581 25993 1593 26027
rect 1627 26024 1639 26027
rect 1670 26024 1676 26036
rect 1627 25996 1676 26024
rect 1627 25993 1639 25996
rect 1581 25987 1639 25993
rect 1670 25984 1676 25996
rect 1728 25984 1734 26036
rect 2866 25984 2872 26036
rect 2924 26024 2930 26036
rect 3053 26027 3111 26033
rect 3053 26024 3065 26027
rect 2924 25996 3065 26024
rect 2924 25984 2930 25996
rect 3053 25993 3065 25996
rect 3099 26024 3111 26027
rect 3513 26027 3571 26033
rect 3513 26024 3525 26027
rect 3099 25996 3525 26024
rect 3099 25993 3111 25996
rect 3053 25987 3111 25993
rect 3513 25993 3525 25996
rect 3559 25993 3571 26027
rect 3513 25987 3571 25993
rect 4709 26027 4767 26033
rect 4709 25993 4721 26027
rect 4755 25993 4767 26027
rect 5626 26024 5632 26036
rect 4709 25987 4767 25993
rect 5276 25996 5632 26024
rect 2958 25916 2964 25968
rect 3016 25956 3022 25968
rect 3237 25959 3295 25965
rect 3237 25956 3249 25959
rect 3016 25928 3249 25956
rect 3016 25916 3022 25928
rect 3237 25925 3249 25928
rect 3283 25956 3295 25959
rect 3789 25959 3847 25965
rect 3789 25956 3801 25959
rect 3283 25928 3801 25956
rect 3283 25925 3295 25928
rect 3237 25919 3295 25925
rect 3789 25925 3801 25928
rect 3835 25925 3847 25959
rect 4724 25956 4752 25987
rect 5276 25965 5304 25996
rect 5626 25984 5632 25996
rect 5684 25984 5690 26036
rect 5905 26027 5963 26033
rect 5905 25993 5917 26027
rect 5951 26024 5963 26027
rect 6546 26024 6552 26036
rect 5951 25996 6552 26024
rect 5951 25993 5963 25996
rect 5905 25987 5963 25993
rect 6546 25984 6552 25996
rect 6604 25984 6610 26036
rect 6638 25984 6644 26036
rect 6696 26024 6702 26036
rect 7009 26027 7067 26033
rect 7009 26024 7021 26027
rect 6696 25996 7021 26024
rect 6696 25984 6702 25996
rect 7009 25993 7021 25996
rect 7055 26024 7067 26027
rect 8386 26024 8392 26036
rect 7055 25996 8392 26024
rect 7055 25993 7067 25996
rect 7009 25987 7067 25993
rect 8386 25984 8392 25996
rect 8444 25984 8450 26036
rect 8665 26027 8723 26033
rect 8665 25993 8677 26027
rect 8711 26024 8723 26027
rect 9030 26024 9036 26036
rect 8711 25996 9036 26024
rect 8711 25993 8723 25996
rect 8665 25987 8723 25993
rect 9030 25984 9036 25996
rect 9088 25984 9094 26036
rect 9401 26027 9459 26033
rect 9401 25993 9413 26027
rect 9447 26024 9459 26027
rect 9490 26024 9496 26036
rect 9447 25996 9496 26024
rect 9447 25993 9459 25996
rect 9401 25987 9459 25993
rect 9490 25984 9496 25996
rect 9548 25984 9554 26036
rect 9861 26027 9919 26033
rect 9861 25993 9873 26027
rect 9907 25993 9919 26027
rect 9861 25987 9919 25993
rect 5261 25959 5319 25965
rect 5261 25956 5273 25959
rect 4724 25928 5273 25956
rect 3789 25919 3847 25925
rect 5261 25925 5273 25928
rect 5307 25925 5319 25959
rect 5261 25919 5319 25925
rect 5534 25916 5540 25968
rect 5592 25956 5598 25968
rect 5592 25928 6776 25956
rect 5592 25916 5598 25928
rect 842 25848 848 25900
rect 900 25888 906 25900
rect 1397 25891 1455 25897
rect 1397 25888 1409 25891
rect 900 25860 1409 25888
rect 900 25848 906 25860
rect 1397 25857 1409 25860
rect 1443 25857 1455 25891
rect 1397 25851 1455 25857
rect 2774 25848 2780 25900
rect 2832 25888 2838 25900
rect 2869 25891 2927 25897
rect 2869 25888 2881 25891
rect 2832 25860 2881 25888
rect 2832 25848 2838 25860
rect 2869 25857 2881 25860
rect 2915 25857 2927 25891
rect 2869 25851 2927 25857
rect 3142 25848 3148 25900
rect 3200 25848 3206 25900
rect 3326 25848 3332 25900
rect 3384 25888 3390 25900
rect 3694 25888 3700 25900
rect 3384 25860 3700 25888
rect 3384 25848 3390 25860
rect 3694 25848 3700 25860
rect 3752 25848 3758 25900
rect 4065 25891 4123 25897
rect 4065 25857 4077 25891
rect 4111 25888 4123 25891
rect 4154 25888 4160 25900
rect 4111 25860 4160 25888
rect 4111 25857 4123 25860
rect 4065 25851 4123 25857
rect 4154 25848 4160 25860
rect 4212 25848 4218 25900
rect 4522 25848 4528 25900
rect 4580 25848 4586 25900
rect 4801 25891 4859 25897
rect 4801 25857 4813 25891
rect 4847 25888 4859 25891
rect 4982 25888 4988 25900
rect 4847 25860 4988 25888
rect 4847 25857 4859 25860
rect 4801 25851 4859 25857
rect 4982 25848 4988 25860
rect 5040 25848 5046 25900
rect 5074 25848 5080 25900
rect 5132 25848 5138 25900
rect 5166 25848 5172 25900
rect 5224 25888 5230 25900
rect 5353 25891 5411 25897
rect 5353 25888 5365 25891
rect 5224 25860 5365 25888
rect 5224 25848 5230 25860
rect 5353 25857 5365 25860
rect 5399 25857 5411 25891
rect 5353 25851 5411 25857
rect 5445 25892 5503 25897
rect 5445 25891 5512 25892
rect 5445 25857 5457 25891
rect 5491 25857 5512 25891
rect 5445 25851 5512 25857
rect 5721 25891 5779 25897
rect 5721 25857 5733 25891
rect 5767 25888 5779 25891
rect 5902 25888 5908 25900
rect 5767 25860 5908 25888
rect 5767 25857 5779 25860
rect 5721 25851 5779 25857
rect 3160 25820 3188 25848
rect 3881 25823 3939 25829
rect 3881 25820 3893 25823
rect 3160 25792 3893 25820
rect 3881 25789 3893 25792
rect 3927 25789 3939 25823
rect 5484 25820 5512 25851
rect 5902 25848 5908 25860
rect 5960 25848 5966 25900
rect 5997 25891 6055 25897
rect 5997 25857 6009 25891
rect 6043 25888 6055 25891
rect 6086 25888 6092 25900
rect 6043 25860 6092 25888
rect 6043 25857 6055 25860
rect 5997 25851 6055 25857
rect 6086 25848 6092 25860
rect 6144 25848 6150 25900
rect 6362 25848 6368 25900
rect 6420 25848 6426 25900
rect 6546 25848 6552 25900
rect 6604 25848 6610 25900
rect 6748 25897 6776 25928
rect 7650 25916 7656 25968
rect 7708 25956 7714 25968
rect 8294 25956 8300 25968
rect 7708 25928 8300 25956
rect 7708 25916 7714 25928
rect 8294 25916 8300 25928
rect 8352 25916 8358 25968
rect 8941 25959 8999 25965
rect 8941 25925 8953 25959
rect 8987 25956 8999 25959
rect 9876 25956 9904 25987
rect 11422 25984 11428 26036
rect 11480 26024 11486 26036
rect 11790 26024 11796 26036
rect 11480 25996 11796 26024
rect 11480 25984 11486 25996
rect 11790 25984 11796 25996
rect 11848 25984 11854 26036
rect 12526 25984 12532 26036
rect 12584 26024 12590 26036
rect 13722 26024 13728 26036
rect 12584 25996 13728 26024
rect 12584 25984 12590 25996
rect 13722 25984 13728 25996
rect 13780 26024 13786 26036
rect 19794 26024 19800 26036
rect 13780 25996 19800 26024
rect 13780 25984 13786 25996
rect 19794 25984 19800 25996
rect 19852 25984 19858 26036
rect 20165 26027 20223 26033
rect 20165 25993 20177 26027
rect 20211 25993 20223 26027
rect 20165 25987 20223 25993
rect 10597 25959 10655 25965
rect 10597 25956 10609 25959
rect 8987 25928 10609 25956
rect 8987 25925 8999 25928
rect 8941 25919 8999 25925
rect 10597 25925 10609 25928
rect 10643 25956 10655 25959
rect 11514 25956 11520 25968
rect 10643 25928 11520 25956
rect 10643 25925 10655 25928
rect 10597 25919 10655 25925
rect 11514 25916 11520 25928
rect 11572 25916 11578 25968
rect 13188 25928 15884 25956
rect 6641 25891 6699 25897
rect 6641 25857 6653 25891
rect 6687 25857 6699 25891
rect 6641 25851 6699 25857
rect 6733 25891 6791 25897
rect 6733 25857 6745 25891
rect 6779 25857 6791 25891
rect 6733 25851 6791 25857
rect 5810 25820 5816 25832
rect 5484 25792 5816 25820
rect 3881 25783 3939 25789
rect 5810 25780 5816 25792
rect 5868 25780 5874 25832
rect 6656 25820 6684 25851
rect 6914 25848 6920 25900
rect 6972 25848 6978 25900
rect 7190 25848 7196 25900
rect 7248 25848 7254 25900
rect 7285 25891 7343 25897
rect 7285 25857 7297 25891
rect 7331 25857 7343 25891
rect 7285 25851 7343 25857
rect 6932 25820 6960 25848
rect 5920 25792 6960 25820
rect 3421 25755 3479 25761
rect 3421 25721 3433 25755
rect 3467 25752 3479 25755
rect 5258 25752 5264 25764
rect 3467 25724 5264 25752
rect 3467 25721 3479 25724
rect 3421 25715 3479 25721
rect 5258 25712 5264 25724
rect 5316 25712 5322 25764
rect 5920 25752 5948 25792
rect 7098 25780 7104 25832
rect 7156 25820 7162 25832
rect 7300 25820 7328 25851
rect 8110 25848 8116 25900
rect 8168 25888 8174 25900
rect 8205 25891 8263 25897
rect 8205 25888 8217 25891
rect 8168 25860 8217 25888
rect 8168 25848 8174 25860
rect 8205 25857 8217 25860
rect 8251 25857 8263 25891
rect 8205 25851 8263 25857
rect 8386 25848 8392 25900
rect 8444 25888 8450 25900
rect 8481 25891 8539 25897
rect 8481 25888 8493 25891
rect 8444 25860 8493 25888
rect 8444 25848 8450 25860
rect 8481 25857 8493 25860
rect 8527 25857 8539 25891
rect 8481 25851 8539 25857
rect 8754 25848 8760 25900
rect 8812 25848 8818 25900
rect 9033 25891 9091 25897
rect 9033 25857 9045 25891
rect 9079 25857 9091 25891
rect 9033 25851 9091 25857
rect 9125 25891 9183 25897
rect 9125 25857 9137 25891
rect 9171 25857 9183 25891
rect 9125 25851 9183 25857
rect 7156 25792 7328 25820
rect 7156 25780 7162 25792
rect 8294 25780 8300 25832
rect 8352 25820 8358 25832
rect 8938 25820 8944 25832
rect 8352 25792 8944 25820
rect 8352 25780 8358 25792
rect 8938 25780 8944 25792
rect 8996 25780 9002 25832
rect 5552 25724 5948 25752
rect 6181 25755 6239 25761
rect 3694 25644 3700 25696
rect 3752 25684 3758 25696
rect 3789 25687 3847 25693
rect 3789 25684 3801 25687
rect 3752 25656 3801 25684
rect 3752 25644 3758 25656
rect 3789 25653 3801 25656
rect 3835 25653 3847 25687
rect 3789 25647 3847 25653
rect 4062 25644 4068 25696
rect 4120 25684 4126 25696
rect 4249 25687 4307 25693
rect 4249 25684 4261 25687
rect 4120 25656 4261 25684
rect 4120 25644 4126 25656
rect 4249 25653 4261 25656
rect 4295 25653 4307 25687
rect 4249 25647 4307 25653
rect 4985 25687 5043 25693
rect 4985 25653 4997 25687
rect 5031 25684 5043 25687
rect 5166 25684 5172 25696
rect 5031 25656 5172 25684
rect 5031 25653 5043 25656
rect 4985 25647 5043 25653
rect 5166 25644 5172 25656
rect 5224 25684 5230 25696
rect 5552 25684 5580 25724
rect 6181 25721 6193 25755
rect 6227 25752 6239 25755
rect 6822 25752 6828 25764
rect 6227 25724 6828 25752
rect 6227 25721 6239 25724
rect 6181 25715 6239 25721
rect 6822 25712 6828 25724
rect 6880 25712 6886 25764
rect 6917 25755 6975 25761
rect 6917 25721 6929 25755
rect 6963 25752 6975 25755
rect 9048 25752 9076 25851
rect 9140 25820 9168 25851
rect 9398 25848 9404 25900
rect 9456 25888 9462 25900
rect 9585 25891 9643 25897
rect 9585 25888 9597 25891
rect 9456 25860 9597 25888
rect 9456 25848 9462 25860
rect 9585 25857 9597 25860
rect 9631 25857 9643 25891
rect 9585 25851 9643 25857
rect 9674 25848 9680 25900
rect 9732 25848 9738 25900
rect 10318 25848 10324 25900
rect 10376 25888 10382 25900
rect 10413 25891 10471 25897
rect 10413 25888 10425 25891
rect 10376 25860 10425 25888
rect 10376 25848 10382 25860
rect 10413 25857 10425 25860
rect 10459 25857 10471 25891
rect 10413 25851 10471 25857
rect 10502 25848 10508 25900
rect 10560 25888 10566 25900
rect 10689 25891 10747 25897
rect 10689 25888 10701 25891
rect 10560 25860 10701 25888
rect 10560 25848 10566 25860
rect 10689 25857 10701 25860
rect 10735 25857 10747 25891
rect 10689 25851 10747 25857
rect 10781 25891 10839 25897
rect 10781 25857 10793 25891
rect 10827 25888 10839 25891
rect 11330 25888 11336 25900
rect 10827 25860 11336 25888
rect 10827 25857 10839 25860
rect 10781 25851 10839 25857
rect 9490 25820 9496 25832
rect 9140 25792 9496 25820
rect 9490 25780 9496 25792
rect 9548 25820 9554 25832
rect 10796 25820 10824 25851
rect 11330 25848 11336 25860
rect 11388 25848 11394 25900
rect 11422 25848 11428 25900
rect 11480 25888 11486 25900
rect 13188 25897 13216 25928
rect 13173 25891 13231 25897
rect 13173 25888 13185 25891
rect 11480 25860 13185 25888
rect 11480 25848 11486 25860
rect 13173 25857 13185 25860
rect 13219 25857 13231 25891
rect 13173 25851 13231 25857
rect 13449 25891 13507 25897
rect 13449 25857 13461 25891
rect 13495 25888 13507 25891
rect 14274 25888 14280 25900
rect 13495 25860 14280 25888
rect 13495 25857 13507 25860
rect 13449 25851 13507 25857
rect 9548 25792 10824 25820
rect 9548 25780 9554 25792
rect 11514 25780 11520 25832
rect 11572 25820 11578 25832
rect 11698 25820 11704 25832
rect 11572 25792 11704 25820
rect 11572 25780 11578 25792
rect 11698 25780 11704 25792
rect 11756 25780 11762 25832
rect 12618 25780 12624 25832
rect 12676 25820 12682 25832
rect 13464 25820 13492 25851
rect 14274 25848 14280 25860
rect 14332 25848 14338 25900
rect 12676 25792 13492 25820
rect 15856 25820 15884 25928
rect 16666 25916 16672 25968
rect 16724 25956 16730 25968
rect 16724 25928 17080 25956
rect 16724 25916 16730 25928
rect 16758 25848 16764 25900
rect 16816 25848 16822 25900
rect 16942 25848 16948 25900
rect 17000 25848 17006 25900
rect 17052 25888 17080 25928
rect 17402 25916 17408 25968
rect 17460 25956 17466 25968
rect 20180 25956 20208 25987
rect 20806 25984 20812 26036
rect 20864 26024 20870 26036
rect 21910 26024 21916 26036
rect 20864 25996 21916 26024
rect 20864 25984 20870 25996
rect 21910 25984 21916 25996
rect 21968 25984 21974 26036
rect 22830 25984 22836 26036
rect 22888 26024 22894 26036
rect 25406 26024 25412 26036
rect 22888 25996 25412 26024
rect 22888 25984 22894 25996
rect 25406 25984 25412 25996
rect 25464 25984 25470 26036
rect 30098 26024 30104 26036
rect 29840 25996 30104 26024
rect 29840 25965 29868 25996
rect 30098 25984 30104 25996
rect 30156 25984 30162 26036
rect 30193 26027 30251 26033
rect 30193 25993 30205 26027
rect 30239 25993 30251 26027
rect 30193 25987 30251 25993
rect 29825 25959 29883 25965
rect 17460 25928 20024 25956
rect 20180 25928 23704 25956
rect 17460 25916 17466 25928
rect 18141 25891 18199 25897
rect 18141 25888 18153 25891
rect 17052 25860 18153 25888
rect 18141 25857 18153 25860
rect 18187 25857 18199 25891
rect 18141 25851 18199 25857
rect 18325 25891 18383 25897
rect 18325 25857 18337 25891
rect 18371 25888 18383 25891
rect 18414 25888 18420 25900
rect 18371 25860 18420 25888
rect 18371 25857 18383 25860
rect 18325 25851 18383 25857
rect 18414 25848 18420 25860
rect 18472 25848 18478 25900
rect 19334 25848 19340 25900
rect 19392 25888 19398 25900
rect 19429 25891 19487 25897
rect 19429 25888 19441 25891
rect 19392 25860 19441 25888
rect 19392 25848 19398 25860
rect 19429 25857 19441 25860
rect 19475 25857 19487 25891
rect 19429 25851 19487 25857
rect 19610 25848 19616 25900
rect 19668 25888 19674 25900
rect 19705 25891 19763 25897
rect 19705 25888 19717 25891
rect 19668 25860 19717 25888
rect 19668 25848 19674 25860
rect 19705 25857 19717 25860
rect 19751 25857 19763 25891
rect 19705 25851 19763 25857
rect 19886 25848 19892 25900
rect 19944 25848 19950 25900
rect 19996 25897 20024 25928
rect 19981 25891 20039 25897
rect 19981 25857 19993 25891
rect 20027 25857 20039 25891
rect 19981 25851 20039 25857
rect 20254 25848 20260 25900
rect 20312 25848 20318 25900
rect 20438 25848 20444 25900
rect 20496 25848 20502 25900
rect 20990 25848 20996 25900
rect 21048 25848 21054 25900
rect 21174 25848 21180 25900
rect 21232 25888 21238 25900
rect 21269 25891 21327 25897
rect 21269 25888 21281 25891
rect 21232 25860 21281 25888
rect 21232 25848 21238 25860
rect 21269 25857 21281 25860
rect 21315 25857 21327 25891
rect 21269 25851 21327 25857
rect 21821 25891 21879 25897
rect 21821 25857 21833 25891
rect 21867 25857 21879 25891
rect 21821 25851 21879 25857
rect 18690 25820 18696 25832
rect 15856 25792 18696 25820
rect 12676 25780 12682 25792
rect 18690 25780 18696 25792
rect 18748 25780 18754 25832
rect 20714 25820 20720 25832
rect 19260 25792 20720 25820
rect 9122 25752 9128 25764
rect 6963 25724 8708 25752
rect 9048 25724 9128 25752
rect 6963 25721 6975 25724
rect 6917 25715 6975 25721
rect 5224 25656 5580 25684
rect 5629 25687 5687 25693
rect 5224 25644 5230 25656
rect 5629 25653 5641 25687
rect 5675 25684 5687 25687
rect 7098 25684 7104 25696
rect 5675 25656 7104 25684
rect 5675 25653 5687 25656
rect 5629 25647 5687 25653
rect 7098 25644 7104 25656
rect 7156 25644 7162 25696
rect 7190 25644 7196 25696
rect 7248 25684 7254 25696
rect 7469 25687 7527 25693
rect 7469 25684 7481 25687
rect 7248 25656 7481 25684
rect 7248 25644 7254 25656
rect 7469 25653 7481 25656
rect 7515 25684 7527 25687
rect 8294 25684 8300 25696
rect 7515 25656 8300 25684
rect 7515 25653 7527 25656
rect 7469 25647 7527 25653
rect 8294 25644 8300 25656
rect 8352 25644 8358 25696
rect 8389 25687 8447 25693
rect 8389 25653 8401 25687
rect 8435 25684 8447 25687
rect 8570 25684 8576 25696
rect 8435 25656 8576 25684
rect 8435 25653 8447 25656
rect 8389 25647 8447 25653
rect 8570 25644 8576 25656
rect 8628 25644 8634 25696
rect 8680 25684 8708 25724
rect 9122 25712 9128 25724
rect 9180 25712 9186 25764
rect 9309 25755 9367 25761
rect 9309 25721 9321 25755
rect 9355 25752 9367 25755
rect 15746 25752 15752 25764
rect 9355 25724 15752 25752
rect 9355 25721 9367 25724
rect 9309 25715 9367 25721
rect 15746 25712 15752 25724
rect 15804 25712 15810 25764
rect 17218 25712 17224 25764
rect 17276 25752 17282 25764
rect 17494 25752 17500 25764
rect 17276 25724 17500 25752
rect 17276 25712 17282 25724
rect 17494 25712 17500 25724
rect 17552 25712 17558 25764
rect 10778 25684 10784 25696
rect 8680 25656 10784 25684
rect 10778 25644 10784 25656
rect 10836 25644 10842 25696
rect 10962 25644 10968 25696
rect 11020 25644 11026 25696
rect 12986 25644 12992 25696
rect 13044 25644 13050 25696
rect 13078 25644 13084 25696
rect 13136 25684 13142 25696
rect 13265 25687 13323 25693
rect 13265 25684 13277 25687
rect 13136 25656 13277 25684
rect 13136 25644 13142 25656
rect 13265 25653 13277 25656
rect 13311 25653 13323 25687
rect 13265 25647 13323 25653
rect 13906 25644 13912 25696
rect 13964 25684 13970 25696
rect 19260 25684 19288 25792
rect 20714 25780 20720 25792
rect 20772 25780 20778 25832
rect 20806 25780 20812 25832
rect 20864 25820 20870 25832
rect 21836 25820 21864 25851
rect 21910 25848 21916 25900
rect 21968 25888 21974 25900
rect 22005 25891 22063 25897
rect 22005 25888 22017 25891
rect 21968 25860 22017 25888
rect 21968 25848 21974 25860
rect 22005 25857 22017 25860
rect 22051 25888 22063 25891
rect 22646 25888 22652 25900
rect 22051 25860 22652 25888
rect 22051 25857 22063 25860
rect 22005 25851 22063 25857
rect 22646 25848 22652 25860
rect 22704 25848 22710 25900
rect 23106 25848 23112 25900
rect 23164 25888 23170 25900
rect 23385 25891 23443 25897
rect 23385 25888 23397 25891
rect 23164 25860 23397 25888
rect 23164 25848 23170 25860
rect 23385 25857 23397 25860
rect 23431 25857 23443 25891
rect 23385 25851 23443 25857
rect 23474 25848 23480 25900
rect 23532 25888 23538 25900
rect 23676 25897 23704 25928
rect 29825 25925 29837 25959
rect 29871 25925 29883 25959
rect 29825 25919 29883 25925
rect 29914 25916 29920 25968
rect 29972 25916 29978 25968
rect 30208 25956 30236 25987
rect 30530 25959 30588 25965
rect 30530 25956 30542 25959
rect 30208 25928 30542 25956
rect 30530 25925 30542 25928
rect 30576 25925 30588 25959
rect 30530 25919 30588 25925
rect 23569 25891 23627 25897
rect 23569 25888 23581 25891
rect 23532 25860 23581 25888
rect 23532 25848 23538 25860
rect 23569 25857 23581 25860
rect 23615 25857 23627 25891
rect 23569 25851 23627 25857
rect 23661 25891 23719 25897
rect 23661 25857 23673 25891
rect 23707 25857 23719 25891
rect 23661 25851 23719 25857
rect 24029 25891 24087 25897
rect 24029 25857 24041 25891
rect 24075 25888 24087 25891
rect 24578 25888 24584 25900
rect 24075 25860 24584 25888
rect 24075 25857 24087 25860
rect 24029 25851 24087 25857
rect 24578 25848 24584 25860
rect 24636 25848 24642 25900
rect 29638 25848 29644 25900
rect 29696 25848 29702 25900
rect 30009 25891 30067 25897
rect 30009 25857 30021 25891
rect 30055 25888 30067 25891
rect 30926 25888 30932 25900
rect 30055 25860 30932 25888
rect 30055 25857 30067 25860
rect 30009 25851 30067 25857
rect 30926 25848 30932 25860
rect 30984 25848 30990 25900
rect 32122 25848 32128 25900
rect 32180 25888 32186 25900
rect 32217 25891 32275 25897
rect 32217 25888 32229 25891
rect 32180 25860 32229 25888
rect 32180 25848 32186 25860
rect 32217 25857 32229 25860
rect 32263 25857 32275 25891
rect 32217 25851 32275 25857
rect 25498 25820 25504 25832
rect 20864 25792 21864 25820
rect 21928 25792 25504 25820
rect 20864 25780 20870 25792
rect 19518 25712 19524 25764
rect 19576 25752 19582 25764
rect 19613 25755 19671 25761
rect 19613 25752 19625 25755
rect 19576 25724 19625 25752
rect 19576 25712 19582 25724
rect 19613 25721 19625 25724
rect 19659 25721 19671 25755
rect 20625 25755 20683 25761
rect 20625 25752 20637 25755
rect 19613 25715 19671 25721
rect 20180 25724 20637 25752
rect 13964 25656 19288 25684
rect 13964 25644 13970 25656
rect 19334 25644 19340 25696
rect 19392 25644 19398 25696
rect 19978 25644 19984 25696
rect 20036 25684 20042 25696
rect 20180 25684 20208 25724
rect 20625 25721 20637 25724
rect 20671 25721 20683 25755
rect 21928 25752 21956 25792
rect 25498 25780 25504 25792
rect 25556 25780 25562 25832
rect 25774 25780 25780 25832
rect 25832 25820 25838 25832
rect 30285 25823 30343 25829
rect 30285 25820 30297 25823
rect 25832 25792 30297 25820
rect 25832 25780 25838 25792
rect 30285 25789 30297 25792
rect 30331 25789 30343 25823
rect 30285 25783 30343 25789
rect 20625 25715 20683 25721
rect 20732 25724 21956 25752
rect 22189 25755 22247 25761
rect 20036 25656 20208 25684
rect 20036 25644 20042 25656
rect 20254 25644 20260 25696
rect 20312 25644 20318 25696
rect 20438 25644 20444 25696
rect 20496 25684 20502 25696
rect 20732 25684 20760 25724
rect 22189 25721 22201 25755
rect 22235 25752 22247 25755
rect 23842 25752 23848 25764
rect 22235 25724 23848 25752
rect 22235 25721 22247 25724
rect 22189 25715 22247 25721
rect 23842 25712 23848 25724
rect 23900 25712 23906 25764
rect 23937 25755 23995 25761
rect 23937 25721 23949 25755
rect 23983 25752 23995 25755
rect 29454 25752 29460 25764
rect 23983 25724 29460 25752
rect 23983 25721 23995 25724
rect 23937 25715 23995 25721
rect 29454 25712 29460 25724
rect 29512 25712 29518 25764
rect 20496 25656 20760 25684
rect 20496 25644 20502 25656
rect 20990 25644 20996 25696
rect 21048 25684 21054 25696
rect 21177 25687 21235 25693
rect 21177 25684 21189 25687
rect 21048 25656 21189 25684
rect 21048 25644 21054 25656
rect 21177 25653 21189 25656
rect 21223 25684 21235 25687
rect 21358 25684 21364 25696
rect 21223 25656 21364 25684
rect 21223 25653 21235 25656
rect 21177 25647 21235 25653
rect 21358 25644 21364 25656
rect 21416 25644 21422 25696
rect 21450 25644 21456 25696
rect 21508 25644 21514 25696
rect 21542 25644 21548 25696
rect 21600 25684 21606 25696
rect 21821 25687 21879 25693
rect 21821 25684 21833 25687
rect 21600 25656 21833 25684
rect 21600 25644 21606 25656
rect 21821 25653 21833 25656
rect 21867 25653 21879 25687
rect 21821 25647 21879 25653
rect 22922 25644 22928 25696
rect 22980 25684 22986 25696
rect 23201 25687 23259 25693
rect 23201 25684 23213 25687
rect 22980 25656 23213 25684
rect 22980 25644 22986 25656
rect 23201 25653 23213 25656
rect 23247 25653 23259 25687
rect 23201 25647 23259 25653
rect 23658 25644 23664 25696
rect 23716 25644 23722 25696
rect 24210 25644 24216 25696
rect 24268 25644 24274 25696
rect 24946 25644 24952 25696
rect 25004 25684 25010 25696
rect 25958 25684 25964 25696
rect 25004 25656 25964 25684
rect 25004 25644 25010 25656
rect 25958 25644 25964 25656
rect 26016 25644 26022 25696
rect 30300 25684 30328 25783
rect 31754 25780 31760 25832
rect 31812 25780 31818 25832
rect 31665 25755 31723 25761
rect 31665 25721 31677 25755
rect 31711 25752 31723 25755
rect 31772 25752 31800 25780
rect 32214 25752 32220 25764
rect 31711 25724 32220 25752
rect 31711 25721 31723 25724
rect 31665 25715 31723 25721
rect 32214 25712 32220 25724
rect 32272 25712 32278 25764
rect 30926 25684 30932 25696
rect 30300 25656 30932 25684
rect 30926 25644 30932 25656
rect 30984 25644 30990 25696
rect 31754 25644 31760 25696
rect 31812 25684 31818 25696
rect 32401 25687 32459 25693
rect 32401 25684 32413 25687
rect 31812 25656 32413 25684
rect 31812 25644 31818 25656
rect 32401 25653 32413 25656
rect 32447 25653 32459 25687
rect 32401 25647 32459 25653
rect 1104 25594 32844 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 32844 25594
rect 1104 25520 32844 25542
rect 2777 25483 2835 25489
rect 2777 25449 2789 25483
rect 2823 25480 2835 25483
rect 3878 25480 3884 25492
rect 2823 25452 3884 25480
rect 2823 25449 2835 25452
rect 2777 25443 2835 25449
rect 3878 25440 3884 25452
rect 3936 25440 3942 25492
rect 6178 25440 6184 25492
rect 6236 25480 6242 25492
rect 6457 25483 6515 25489
rect 6457 25480 6469 25483
rect 6236 25452 6469 25480
rect 6236 25440 6242 25452
rect 6457 25449 6469 25452
rect 6503 25449 6515 25483
rect 6457 25443 6515 25449
rect 6546 25440 6552 25492
rect 6604 25480 6610 25492
rect 6730 25480 6736 25492
rect 6604 25452 6736 25480
rect 6604 25440 6610 25452
rect 6730 25440 6736 25452
rect 6788 25440 6794 25492
rect 6914 25440 6920 25492
rect 6972 25480 6978 25492
rect 8478 25480 8484 25492
rect 6972 25452 8484 25480
rect 6972 25440 6978 25452
rect 8478 25440 8484 25452
rect 8536 25440 8542 25492
rect 8754 25440 8760 25492
rect 8812 25480 8818 25492
rect 9306 25480 9312 25492
rect 8812 25452 9312 25480
rect 8812 25440 8818 25452
rect 9306 25440 9312 25452
rect 9364 25440 9370 25492
rect 9674 25480 9680 25492
rect 9416 25452 9680 25480
rect 4065 25415 4123 25421
rect 4065 25381 4077 25415
rect 4111 25412 4123 25415
rect 4614 25412 4620 25424
rect 4111 25384 4620 25412
rect 4111 25381 4123 25384
rect 4065 25375 4123 25381
rect 4614 25372 4620 25384
rect 4672 25372 4678 25424
rect 5445 25415 5503 25421
rect 5445 25381 5457 25415
rect 5491 25381 5503 25415
rect 5445 25375 5503 25381
rect 4338 25344 4344 25356
rect 3896 25316 4344 25344
rect 1394 25236 1400 25288
rect 1452 25236 1458 25288
rect 3050 25236 3056 25288
rect 3108 25236 3114 25288
rect 3142 25236 3148 25288
rect 3200 25236 3206 25288
rect 3602 25236 3608 25288
rect 3660 25236 3666 25288
rect 3896 25285 3924 25316
rect 4338 25304 4344 25316
rect 4396 25304 4402 25356
rect 5460 25344 5488 25375
rect 6086 25372 6092 25424
rect 6144 25412 6150 25424
rect 9416 25412 9444 25452
rect 9674 25440 9680 25452
rect 9732 25440 9738 25492
rect 10321 25483 10379 25489
rect 10321 25449 10333 25483
rect 10367 25480 10379 25483
rect 11422 25480 11428 25492
rect 10367 25452 11428 25480
rect 10367 25449 10379 25452
rect 10321 25443 10379 25449
rect 11422 25440 11428 25452
rect 11480 25440 11486 25492
rect 12802 25440 12808 25492
rect 12860 25480 12866 25492
rect 13078 25480 13084 25492
rect 12860 25452 13084 25480
rect 12860 25440 12866 25452
rect 13078 25440 13084 25452
rect 13136 25440 13142 25492
rect 13633 25483 13691 25489
rect 13633 25449 13645 25483
rect 13679 25480 13691 25483
rect 13722 25480 13728 25492
rect 13679 25452 13728 25480
rect 13679 25449 13691 25452
rect 13633 25443 13691 25449
rect 13722 25440 13728 25452
rect 13780 25440 13786 25492
rect 16761 25483 16819 25489
rect 16761 25449 16773 25483
rect 16807 25480 16819 25483
rect 17037 25483 17095 25489
rect 17037 25480 17049 25483
rect 16807 25452 17049 25480
rect 16807 25449 16819 25452
rect 16761 25443 16819 25449
rect 17037 25449 17049 25452
rect 17083 25449 17095 25483
rect 17037 25443 17095 25449
rect 17405 25483 17463 25489
rect 17405 25449 17417 25483
rect 17451 25480 17463 25483
rect 17494 25480 17500 25492
rect 17451 25452 17500 25480
rect 17451 25449 17463 25452
rect 17405 25443 17463 25449
rect 17494 25440 17500 25452
rect 17552 25440 17558 25492
rect 19613 25483 19671 25489
rect 19613 25449 19625 25483
rect 19659 25480 19671 25483
rect 19702 25480 19708 25492
rect 19659 25452 19708 25480
rect 19659 25449 19671 25452
rect 19613 25443 19671 25449
rect 19702 25440 19708 25452
rect 19760 25440 19766 25492
rect 20162 25440 20168 25492
rect 20220 25480 20226 25492
rect 20438 25480 20444 25492
rect 20220 25452 20444 25480
rect 20220 25440 20226 25452
rect 20438 25440 20444 25452
rect 20496 25440 20502 25492
rect 20533 25483 20591 25489
rect 20533 25449 20545 25483
rect 20579 25480 20591 25483
rect 20806 25480 20812 25492
rect 20579 25452 20812 25480
rect 20579 25449 20591 25452
rect 20533 25443 20591 25449
rect 20806 25440 20812 25452
rect 20864 25440 20870 25492
rect 21358 25440 21364 25492
rect 21416 25440 21422 25492
rect 22738 25440 22744 25492
rect 22796 25440 22802 25492
rect 23658 25440 23664 25492
rect 23716 25440 23722 25492
rect 24210 25440 24216 25492
rect 24268 25480 24274 25492
rect 24268 25452 24532 25480
rect 24268 25440 24274 25452
rect 6144 25384 9444 25412
rect 6144 25372 6150 25384
rect 9582 25372 9588 25424
rect 9640 25372 9646 25424
rect 11238 25412 11244 25424
rect 9692 25384 11244 25412
rect 6454 25344 6460 25356
rect 5460 25316 6460 25344
rect 3881 25279 3939 25285
rect 3881 25245 3893 25279
rect 3927 25245 3939 25279
rect 3881 25239 3939 25245
rect 4154 25236 4160 25288
rect 4212 25236 4218 25288
rect 4433 25279 4491 25285
rect 4433 25245 4445 25279
rect 4479 25245 4491 25279
rect 4433 25239 4491 25245
rect 1670 25217 1676 25220
rect 1664 25171 1676 25217
rect 1670 25168 1676 25171
rect 1728 25168 1734 25220
rect 4448 25208 4476 25239
rect 5258 25236 5264 25288
rect 5316 25236 5322 25288
rect 5736 25285 5764 25316
rect 6454 25304 6460 25316
rect 6512 25304 6518 25356
rect 8570 25304 8576 25356
rect 8628 25344 8634 25356
rect 8628 25316 9444 25344
rect 8628 25304 8634 25316
rect 5721 25279 5779 25285
rect 5721 25245 5733 25279
rect 5767 25245 5779 25279
rect 5721 25239 5779 25245
rect 5810 25236 5816 25288
rect 5868 25236 5874 25288
rect 6089 25279 6147 25285
rect 6089 25276 6101 25279
rect 5920 25248 6101 25276
rect 4706 25208 4712 25220
rect 3344 25180 4476 25208
rect 4540 25180 4712 25208
rect 3344 25152 3372 25180
rect 2866 25100 2872 25152
rect 2924 25100 2930 25152
rect 3326 25100 3332 25152
rect 3384 25100 3390 25152
rect 3418 25100 3424 25152
rect 3476 25100 3482 25152
rect 4341 25143 4399 25149
rect 4341 25109 4353 25143
rect 4387 25140 4399 25143
rect 4540 25140 4568 25180
rect 4706 25168 4712 25180
rect 4764 25168 4770 25220
rect 5626 25168 5632 25220
rect 5684 25208 5690 25220
rect 5920 25208 5948 25248
rect 6089 25245 6101 25248
rect 6135 25245 6147 25279
rect 6089 25239 6147 25245
rect 6178 25236 6184 25288
rect 6236 25236 6242 25288
rect 6546 25276 6552 25288
rect 6288 25248 6552 25276
rect 5684 25180 5948 25208
rect 5997 25211 6055 25217
rect 5684 25168 5690 25180
rect 5997 25177 6009 25211
rect 6043 25208 6055 25211
rect 6288 25208 6316 25248
rect 6546 25236 6552 25248
rect 6604 25236 6610 25288
rect 6638 25236 6644 25288
rect 6696 25236 6702 25288
rect 6822 25236 6828 25288
rect 6880 25276 6886 25288
rect 6917 25279 6975 25285
rect 6917 25276 6929 25279
rect 6880 25248 6929 25276
rect 6880 25236 6886 25248
rect 6917 25245 6929 25248
rect 6963 25276 6975 25279
rect 8386 25276 8392 25288
rect 6963 25248 8392 25276
rect 6963 25245 6975 25248
rect 6917 25239 6975 25245
rect 8386 25236 8392 25248
rect 8444 25236 8450 25288
rect 8938 25236 8944 25288
rect 8996 25236 9002 25288
rect 9030 25236 9036 25288
rect 9088 25276 9094 25288
rect 9416 25285 9444 25316
rect 9125 25279 9183 25285
rect 9125 25276 9137 25279
rect 9088 25248 9137 25276
rect 9088 25236 9094 25248
rect 9125 25245 9137 25248
rect 9171 25245 9183 25279
rect 9125 25239 9183 25245
rect 9401 25279 9459 25285
rect 9401 25245 9413 25279
rect 9447 25245 9459 25279
rect 9401 25239 9459 25245
rect 9490 25236 9496 25288
rect 9548 25276 9554 25288
rect 9692 25285 9720 25384
rect 11238 25372 11244 25384
rect 11296 25372 11302 25424
rect 11698 25372 11704 25424
rect 11756 25412 11762 25424
rect 11756 25384 12480 25412
rect 11756 25372 11762 25384
rect 9950 25344 9956 25356
rect 9876 25316 9956 25344
rect 9876 25285 9904 25316
rect 9950 25304 9956 25316
rect 10008 25304 10014 25356
rect 11146 25344 11152 25356
rect 10796 25316 11152 25344
rect 9677 25279 9735 25285
rect 9677 25276 9689 25279
rect 9548 25248 9689 25276
rect 9548 25236 9554 25248
rect 9677 25245 9689 25248
rect 9723 25245 9735 25279
rect 9677 25239 9735 25245
rect 9861 25279 9919 25285
rect 9861 25245 9873 25279
rect 9907 25245 9919 25279
rect 9861 25239 9919 25245
rect 10045 25279 10103 25285
rect 10045 25245 10057 25279
rect 10091 25276 10103 25279
rect 10134 25276 10140 25288
rect 10091 25248 10140 25276
rect 10091 25245 10103 25248
rect 10045 25239 10103 25245
rect 10134 25236 10140 25248
rect 10192 25236 10198 25288
rect 10502 25236 10508 25288
rect 10560 25236 10566 25288
rect 10796 25285 10824 25316
rect 11146 25304 11152 25316
rect 11204 25344 11210 25356
rect 11204 25316 11744 25344
rect 11204 25304 11210 25316
rect 10781 25279 10839 25285
rect 10781 25245 10793 25279
rect 10827 25245 10839 25279
rect 10781 25239 10839 25245
rect 10965 25279 11023 25285
rect 10965 25245 10977 25279
rect 11011 25245 11023 25279
rect 10965 25239 11023 25245
rect 11057 25279 11115 25285
rect 11057 25245 11069 25279
rect 11103 25276 11115 25279
rect 11238 25276 11244 25288
rect 11103 25248 11244 25276
rect 11103 25245 11115 25248
rect 11057 25239 11115 25245
rect 6043 25180 6316 25208
rect 6380 25180 9444 25208
rect 6043 25177 6055 25180
rect 5997 25171 6055 25177
rect 4387 25112 4568 25140
rect 4617 25143 4675 25149
rect 4387 25109 4399 25112
rect 4341 25103 4399 25109
rect 4617 25109 4629 25143
rect 4663 25140 4675 25143
rect 4798 25140 4804 25152
rect 4663 25112 4804 25140
rect 4663 25109 4675 25112
rect 4617 25103 4675 25109
rect 4798 25100 4804 25112
rect 4856 25100 4862 25152
rect 5537 25143 5595 25149
rect 5537 25109 5549 25143
rect 5583 25140 5595 25143
rect 5810 25140 5816 25152
rect 5583 25112 5816 25140
rect 5583 25109 5595 25112
rect 5537 25103 5595 25109
rect 5810 25100 5816 25112
rect 5868 25100 5874 25152
rect 6380 25149 6408 25180
rect 6365 25143 6423 25149
rect 6365 25109 6377 25143
rect 6411 25109 6423 25143
rect 6365 25103 6423 25109
rect 6454 25100 6460 25152
rect 6512 25140 6518 25152
rect 7926 25140 7932 25152
rect 6512 25112 7932 25140
rect 6512 25100 6518 25112
rect 7926 25100 7932 25112
rect 7984 25100 7990 25152
rect 9416 25140 9444 25180
rect 9950 25168 9956 25220
rect 10008 25168 10014 25220
rect 10134 25140 10140 25152
rect 9416 25112 10140 25140
rect 10134 25100 10140 25112
rect 10192 25100 10198 25152
rect 10229 25143 10287 25149
rect 10229 25109 10241 25143
rect 10275 25140 10287 25143
rect 10410 25140 10416 25152
rect 10275 25112 10416 25140
rect 10275 25109 10287 25112
rect 10229 25103 10287 25109
rect 10410 25100 10416 25112
rect 10468 25100 10474 25152
rect 10980 25140 11008 25239
rect 11238 25236 11244 25248
rect 11296 25236 11302 25288
rect 11422 25236 11428 25288
rect 11480 25236 11486 25288
rect 11514 25236 11520 25288
rect 11572 25276 11578 25288
rect 11716 25285 11744 25316
rect 11609 25279 11667 25285
rect 11609 25276 11621 25279
rect 11572 25248 11621 25276
rect 11572 25236 11578 25248
rect 11609 25245 11621 25248
rect 11655 25245 11667 25279
rect 11609 25239 11667 25245
rect 11701 25279 11759 25285
rect 11701 25245 11713 25279
rect 11747 25245 11759 25279
rect 11701 25239 11759 25245
rect 11790 25236 11796 25288
rect 11848 25236 11854 25288
rect 12069 25279 12127 25285
rect 12069 25245 12081 25279
rect 12115 25245 12127 25279
rect 12069 25239 12127 25245
rect 12084 25208 12112 25239
rect 12342 25236 12348 25288
rect 12400 25236 12406 25288
rect 12452 25285 12480 25384
rect 12618 25372 12624 25424
rect 12676 25372 12682 25424
rect 13265 25415 13323 25421
rect 13265 25381 13277 25415
rect 13311 25412 13323 25415
rect 13311 25384 13492 25412
rect 13311 25381 13323 25384
rect 13265 25375 13323 25381
rect 13464 25353 13492 25384
rect 15286 25372 15292 25424
rect 15344 25412 15350 25424
rect 16114 25412 16120 25424
rect 15344 25384 16120 25412
rect 15344 25372 15350 25384
rect 16114 25372 16120 25384
rect 16172 25372 16178 25424
rect 16945 25415 17003 25421
rect 16945 25381 16957 25415
rect 16991 25412 17003 25415
rect 17218 25412 17224 25424
rect 16991 25384 17224 25412
rect 16991 25381 17003 25384
rect 16945 25375 17003 25381
rect 17218 25372 17224 25384
rect 17276 25372 17282 25424
rect 19245 25415 19303 25421
rect 19245 25381 19257 25415
rect 19291 25381 19303 25415
rect 19245 25375 19303 25381
rect 13449 25347 13507 25353
rect 13449 25313 13461 25347
rect 13495 25313 13507 25347
rect 13449 25307 13507 25313
rect 13722 25304 13728 25356
rect 13780 25344 13786 25356
rect 17034 25344 17040 25356
rect 13780 25316 17040 25344
rect 13780 25304 13786 25316
rect 17034 25304 17040 25316
rect 17092 25304 17098 25356
rect 18414 25344 18420 25356
rect 17328 25316 18420 25344
rect 12437 25279 12495 25285
rect 12437 25245 12449 25279
rect 12483 25245 12495 25279
rect 12437 25239 12495 25245
rect 12618 25236 12624 25288
rect 12676 25276 12682 25288
rect 12986 25276 12992 25288
rect 12676 25248 12992 25276
rect 12676 25236 12682 25248
rect 12986 25236 12992 25248
rect 13044 25236 13050 25288
rect 13078 25236 13084 25288
rect 13136 25236 13142 25288
rect 13633 25279 13691 25285
rect 13633 25245 13645 25279
rect 13679 25276 13691 25279
rect 14366 25276 14372 25288
rect 13679 25248 14372 25276
rect 13679 25245 13691 25248
rect 13633 25239 13691 25245
rect 14366 25236 14372 25248
rect 14424 25236 14430 25288
rect 14461 25279 14519 25285
rect 14461 25245 14473 25279
rect 14507 25276 14519 25279
rect 14550 25276 14556 25288
rect 14507 25248 14556 25276
rect 14507 25245 14519 25248
rect 14461 25239 14519 25245
rect 14550 25236 14556 25248
rect 14608 25276 14614 25288
rect 15194 25276 15200 25288
rect 14608 25248 15200 25276
rect 14608 25236 14614 25248
rect 15194 25236 15200 25248
rect 15252 25236 15258 25288
rect 15933 25279 15991 25285
rect 15933 25245 15945 25279
rect 15979 25276 15991 25279
rect 16022 25276 16028 25288
rect 15979 25248 16028 25276
rect 15979 25245 15991 25248
rect 15933 25239 15991 25245
rect 16022 25236 16028 25248
rect 16080 25236 16086 25288
rect 16390 25236 16396 25288
rect 16448 25276 16454 25288
rect 16577 25279 16635 25285
rect 16577 25276 16589 25279
rect 16448 25248 16589 25276
rect 16448 25236 16454 25248
rect 16577 25245 16589 25248
rect 16623 25245 16635 25279
rect 16577 25239 16635 25245
rect 16666 25236 16672 25288
rect 16724 25236 16730 25288
rect 17218 25236 17224 25288
rect 17276 25236 17282 25288
rect 11808 25180 12112 25208
rect 11808 25152 11836 25180
rect 12250 25168 12256 25220
rect 12308 25168 12314 25220
rect 12805 25211 12863 25217
rect 12805 25177 12817 25211
rect 12851 25177 12863 25211
rect 12805 25171 12863 25177
rect 11241 25143 11299 25149
rect 11241 25140 11253 25143
rect 10980 25112 11253 25140
rect 11241 25109 11253 25112
rect 11287 25140 11299 25143
rect 11790 25140 11796 25152
rect 11287 25112 11796 25140
rect 11287 25109 11299 25112
rect 11241 25103 11299 25109
rect 11790 25100 11796 25112
rect 11848 25100 11854 25152
rect 11977 25143 12035 25149
rect 11977 25109 11989 25143
rect 12023 25140 12035 25143
rect 12526 25140 12532 25152
rect 12023 25112 12532 25140
rect 12023 25109 12035 25112
rect 11977 25103 12035 25109
rect 12526 25100 12532 25112
rect 12584 25100 12590 25152
rect 12820 25140 12848 25171
rect 13354 25168 13360 25220
rect 13412 25168 13418 25220
rect 16114 25168 16120 25220
rect 16172 25168 16178 25220
rect 16301 25211 16359 25217
rect 16301 25177 16313 25211
rect 16347 25208 16359 25211
rect 17328 25208 17356 25316
rect 18414 25304 18420 25316
rect 18472 25304 18478 25356
rect 19150 25304 19156 25356
rect 19208 25344 19214 25356
rect 19260 25344 19288 25375
rect 19886 25372 19892 25424
rect 19944 25412 19950 25424
rect 19944 25384 20576 25412
rect 19944 25372 19950 25384
rect 20349 25347 20407 25353
rect 20349 25344 20361 25347
rect 19208 25316 20361 25344
rect 19208 25304 19214 25316
rect 20349 25313 20361 25316
rect 20395 25313 20407 25347
rect 20548 25344 20576 25384
rect 20714 25372 20720 25424
rect 20772 25372 20778 25424
rect 20993 25415 21051 25421
rect 20993 25381 21005 25415
rect 21039 25412 21051 25415
rect 21082 25412 21088 25424
rect 21039 25384 21088 25412
rect 21039 25381 21051 25384
rect 20993 25375 21051 25381
rect 21082 25372 21088 25384
rect 21140 25372 21146 25424
rect 21174 25372 21180 25424
rect 21232 25372 21238 25424
rect 21637 25415 21695 25421
rect 21637 25381 21649 25415
rect 21683 25412 21695 25415
rect 21683 25384 22600 25412
rect 21683 25381 21695 25384
rect 21637 25375 21695 25381
rect 21192 25344 21220 25372
rect 21450 25344 21456 25356
rect 20548 25316 21220 25344
rect 21284 25316 21456 25344
rect 20349 25307 20407 25313
rect 17402 25236 17408 25288
rect 17460 25236 17466 25288
rect 17494 25236 17500 25288
rect 17552 25236 17558 25288
rect 17681 25279 17739 25285
rect 17681 25245 17693 25279
rect 17727 25245 17739 25279
rect 17681 25239 17739 25245
rect 16347 25180 17356 25208
rect 17512 25208 17540 25236
rect 17696 25208 17724 25239
rect 17770 25236 17776 25288
rect 17828 25236 17834 25288
rect 18049 25279 18107 25285
rect 18049 25245 18061 25279
rect 18095 25276 18107 25279
rect 18506 25276 18512 25288
rect 18095 25248 18512 25276
rect 18095 25245 18107 25248
rect 18049 25239 18107 25245
rect 18506 25236 18512 25248
rect 18564 25236 18570 25288
rect 19426 25236 19432 25288
rect 19484 25236 19490 25288
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25276 19671 25279
rect 19702 25276 19708 25288
rect 19659 25248 19708 25276
rect 19659 25245 19671 25248
rect 19613 25239 19671 25245
rect 19702 25236 19708 25248
rect 19760 25236 19766 25288
rect 19978 25236 19984 25288
rect 20036 25276 20042 25288
rect 20257 25279 20315 25285
rect 20257 25276 20269 25279
rect 20036 25248 20269 25276
rect 20036 25236 20042 25248
rect 20257 25245 20269 25248
rect 20303 25245 20315 25279
rect 20257 25239 20315 25245
rect 20530 25236 20536 25288
rect 20588 25236 20594 25288
rect 20809 25279 20867 25285
rect 20809 25245 20821 25279
rect 20855 25276 20867 25279
rect 21174 25276 21180 25288
rect 20855 25248 21180 25276
rect 20855 25245 20867 25248
rect 20809 25239 20867 25245
rect 21174 25236 21180 25248
rect 21232 25236 21238 25288
rect 21284 25285 21312 25316
rect 21450 25304 21456 25316
rect 21508 25304 21514 25356
rect 22572 25344 22600 25384
rect 22646 25372 22652 25424
rect 22704 25412 22710 25424
rect 23474 25412 23480 25424
rect 22704 25384 23480 25412
rect 22704 25372 22710 25384
rect 23474 25372 23480 25384
rect 23532 25372 23538 25424
rect 24504 25412 24532 25452
rect 24854 25440 24860 25492
rect 24912 25480 24918 25492
rect 25041 25483 25099 25489
rect 25041 25480 25053 25483
rect 24912 25452 25053 25480
rect 24912 25440 24918 25452
rect 25041 25449 25053 25452
rect 25087 25449 25099 25483
rect 25041 25443 25099 25449
rect 25501 25483 25559 25489
rect 25501 25449 25513 25483
rect 25547 25480 25559 25483
rect 25774 25480 25780 25492
rect 25547 25452 25780 25480
rect 25547 25449 25559 25452
rect 25501 25443 25559 25449
rect 25774 25440 25780 25452
rect 25832 25440 25838 25492
rect 25958 25440 25964 25492
rect 26016 25440 26022 25492
rect 26329 25483 26387 25489
rect 26329 25449 26341 25483
rect 26375 25449 26387 25483
rect 26329 25443 26387 25449
rect 26344 25412 26372 25443
rect 29546 25440 29552 25492
rect 29604 25440 29610 25492
rect 29638 25440 29644 25492
rect 29696 25480 29702 25492
rect 29917 25483 29975 25489
rect 29917 25480 29929 25483
rect 29696 25452 29929 25480
rect 29696 25440 29702 25452
rect 29917 25449 29929 25452
rect 29963 25449 29975 25483
rect 29917 25443 29975 25449
rect 32490 25440 32496 25492
rect 32548 25440 32554 25492
rect 24504 25384 25360 25412
rect 21652 25316 22048 25344
rect 22572 25316 24164 25344
rect 21269 25279 21327 25285
rect 21269 25245 21281 25279
rect 21315 25245 21327 25279
rect 21269 25239 21327 25245
rect 21361 25279 21419 25285
rect 21361 25245 21373 25279
rect 21407 25276 21419 25279
rect 21542 25276 21548 25288
rect 21407 25248 21548 25276
rect 21407 25245 21419 25248
rect 21361 25239 21419 25245
rect 21542 25236 21548 25248
rect 21600 25236 21606 25288
rect 21652 25208 21680 25316
rect 21910 25236 21916 25288
rect 21968 25236 21974 25288
rect 22020 25276 22048 25316
rect 22646 25276 22652 25288
rect 22020 25248 22652 25276
rect 22646 25236 22652 25248
rect 22704 25236 22710 25288
rect 22738 25236 22744 25288
rect 22796 25276 22802 25288
rect 22925 25279 22983 25285
rect 22925 25276 22937 25279
rect 22796 25248 22937 25276
rect 22796 25236 22802 25248
rect 22925 25245 22937 25248
rect 22971 25245 22983 25279
rect 22925 25239 22983 25245
rect 23106 25236 23112 25288
rect 23164 25276 23170 25288
rect 23952 25285 23980 25316
rect 23201 25279 23259 25285
rect 23201 25276 23213 25279
rect 23164 25248 23213 25276
rect 23164 25236 23170 25248
rect 23201 25245 23213 25248
rect 23247 25245 23259 25279
rect 23201 25239 23259 25245
rect 23937 25279 23995 25285
rect 23937 25245 23949 25279
rect 23983 25245 23995 25279
rect 23937 25239 23995 25245
rect 24029 25279 24087 25285
rect 24029 25245 24041 25279
rect 24075 25245 24087 25279
rect 24136 25276 24164 25316
rect 24946 25304 24952 25356
rect 25004 25344 25010 25356
rect 25133 25347 25191 25353
rect 25133 25344 25145 25347
rect 25004 25316 25145 25344
rect 25004 25304 25010 25316
rect 25133 25313 25145 25316
rect 25179 25313 25191 25347
rect 25133 25307 25191 25313
rect 25332 25285 25360 25384
rect 25424 25384 26372 25412
rect 25317 25279 25375 25285
rect 24136 25248 25176 25276
rect 24029 25239 24087 25245
rect 24044 25208 24072 25239
rect 17512 25180 17724 25208
rect 17880 25180 21680 25208
rect 21744 25180 24072 25208
rect 16347 25177 16359 25180
rect 16301 25171 16359 25177
rect 12986 25140 12992 25152
rect 12820 25112 12992 25140
rect 12986 25100 12992 25112
rect 13044 25100 13050 25152
rect 13817 25143 13875 25149
rect 13817 25109 13829 25143
rect 13863 25140 13875 25143
rect 14182 25140 14188 25152
rect 13863 25112 14188 25140
rect 13863 25109 13875 25112
rect 13817 25103 13875 25109
rect 14182 25100 14188 25112
rect 14240 25100 14246 25152
rect 14277 25143 14335 25149
rect 14277 25109 14289 25143
rect 14323 25140 14335 25143
rect 14366 25140 14372 25152
rect 14323 25112 14372 25140
rect 14323 25109 14335 25112
rect 14277 25103 14335 25109
rect 14366 25100 14372 25112
rect 14424 25140 14430 25152
rect 16132 25140 16160 25168
rect 16592 25152 16620 25180
rect 14424 25112 16160 25140
rect 14424 25100 14430 25112
rect 16390 25100 16396 25152
rect 16448 25100 16454 25152
rect 16574 25100 16580 25152
rect 16632 25100 16638 25152
rect 16850 25100 16856 25152
rect 16908 25140 16914 25152
rect 17497 25143 17555 25149
rect 17497 25140 17509 25143
rect 16908 25112 17509 25140
rect 16908 25100 16914 25112
rect 17497 25109 17509 25112
rect 17543 25140 17555 25143
rect 17880 25140 17908 25180
rect 17543 25112 17908 25140
rect 17957 25143 18015 25149
rect 17543 25109 17555 25112
rect 17497 25103 17555 25109
rect 17957 25109 17969 25143
rect 18003 25140 18015 25143
rect 18046 25140 18052 25152
rect 18003 25112 18052 25140
rect 18003 25109 18015 25112
rect 17957 25103 18015 25109
rect 18046 25100 18052 25112
rect 18104 25100 18110 25152
rect 18230 25100 18236 25152
rect 18288 25100 18294 25152
rect 18414 25100 18420 25152
rect 18472 25140 18478 25152
rect 21744 25140 21772 25180
rect 24210 25168 24216 25220
rect 24268 25168 24274 25220
rect 25038 25168 25044 25220
rect 25096 25168 25102 25220
rect 25148 25208 25176 25248
rect 25317 25245 25329 25279
rect 25363 25245 25375 25279
rect 25317 25239 25375 25245
rect 25424 25208 25452 25384
rect 25590 25304 25596 25356
rect 25648 25344 25654 25356
rect 25777 25347 25835 25353
rect 25777 25344 25789 25347
rect 25648 25316 25789 25344
rect 25648 25304 25654 25316
rect 25777 25313 25789 25316
rect 25823 25313 25835 25347
rect 25777 25307 25835 25313
rect 26510 25304 26516 25356
rect 26568 25344 26574 25356
rect 27430 25344 27436 25356
rect 26568 25316 27436 25344
rect 26568 25304 26574 25316
rect 27430 25304 27436 25316
rect 27488 25304 27494 25356
rect 30926 25304 30932 25356
rect 30984 25344 30990 25356
rect 31113 25347 31171 25353
rect 31113 25344 31125 25347
rect 30984 25316 31125 25344
rect 30984 25304 30990 25316
rect 31113 25313 31125 25316
rect 31159 25313 31171 25347
rect 31113 25307 31171 25313
rect 25498 25236 25504 25288
rect 25556 25276 25562 25288
rect 25961 25279 26019 25285
rect 25961 25276 25973 25279
rect 25556 25248 25973 25276
rect 25556 25236 25562 25248
rect 25961 25245 25973 25248
rect 26007 25245 26019 25279
rect 25961 25239 26019 25245
rect 26602 25236 26608 25288
rect 26660 25236 26666 25288
rect 29454 25236 29460 25288
rect 29512 25276 29518 25288
rect 29549 25279 29607 25285
rect 29549 25276 29561 25279
rect 29512 25248 29561 25276
rect 29512 25236 29518 25248
rect 29549 25245 29561 25248
rect 29595 25245 29607 25279
rect 29549 25239 29607 25245
rect 29638 25236 29644 25288
rect 29696 25236 29702 25288
rect 31386 25285 31392 25288
rect 31021 25279 31079 25285
rect 31021 25245 31033 25279
rect 31067 25245 31079 25279
rect 31380 25276 31392 25285
rect 31347 25248 31392 25276
rect 31021 25239 31079 25245
rect 31380 25239 31392 25248
rect 25148 25180 25452 25208
rect 25685 25211 25743 25217
rect 25685 25177 25697 25211
rect 25731 25177 25743 25211
rect 25685 25171 25743 25177
rect 18472 25112 21772 25140
rect 18472 25100 18478 25112
rect 22094 25100 22100 25152
rect 22152 25100 22158 25152
rect 23109 25143 23167 25149
rect 23109 25109 23121 25143
rect 23155 25140 23167 25143
rect 23198 25140 23204 25152
rect 23155 25112 23204 25140
rect 23155 25109 23167 25112
rect 23109 25103 23167 25109
rect 23198 25100 23204 25112
rect 23256 25100 23262 25152
rect 23382 25100 23388 25152
rect 23440 25100 23446 25152
rect 23753 25143 23811 25149
rect 23753 25109 23765 25143
rect 23799 25140 23811 25143
rect 24118 25140 24124 25152
rect 23799 25112 24124 25140
rect 23799 25109 23811 25112
rect 23753 25103 23811 25109
rect 24118 25100 24124 25112
rect 24176 25100 24182 25152
rect 24762 25100 24768 25152
rect 24820 25140 24826 25152
rect 25700 25140 25728 25171
rect 26234 25168 26240 25220
rect 26292 25208 26298 25220
rect 26329 25211 26387 25217
rect 26329 25208 26341 25211
rect 26292 25180 26341 25208
rect 26292 25168 26298 25180
rect 26329 25177 26341 25180
rect 26375 25208 26387 25211
rect 26510 25208 26516 25220
rect 26375 25180 26516 25208
rect 26375 25177 26387 25180
rect 26329 25171 26387 25177
rect 26510 25168 26516 25180
rect 26568 25168 26574 25220
rect 31036 25208 31064 25239
rect 31386 25236 31392 25239
rect 31444 25236 31450 25288
rect 31846 25208 31852 25220
rect 31036 25180 31852 25208
rect 31846 25168 31852 25180
rect 31904 25168 31910 25220
rect 24820 25112 25728 25140
rect 24820 25100 24826 25112
rect 26142 25100 26148 25152
rect 26200 25100 26206 25152
rect 26786 25100 26792 25152
rect 26844 25100 26850 25152
rect 30834 25100 30840 25152
rect 30892 25100 30898 25152
rect 1104 25050 32844 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 32844 25050
rect 1104 24976 32844 24998
rect 2041 24939 2099 24945
rect 2041 24905 2053 24939
rect 2087 24936 2099 24939
rect 2087 24908 2728 24936
rect 2087 24905 2099 24908
rect 2041 24899 2099 24905
rect 2700 24880 2728 24908
rect 3510 24896 3516 24948
rect 3568 24896 3574 24948
rect 3970 24896 3976 24948
rect 4028 24896 4034 24948
rect 5258 24896 5264 24948
rect 5316 24936 5322 24948
rect 5994 24936 6000 24948
rect 5316 24908 6000 24936
rect 5316 24896 5322 24908
rect 5994 24896 6000 24908
rect 6052 24936 6058 24948
rect 6638 24936 6644 24948
rect 6052 24908 6644 24936
rect 6052 24896 6058 24908
rect 6638 24896 6644 24908
rect 6696 24896 6702 24948
rect 9030 24936 9036 24948
rect 6794 24908 9036 24936
rect 2682 24828 2688 24880
rect 2740 24868 2746 24880
rect 2777 24871 2835 24877
rect 2777 24868 2789 24871
rect 2740 24840 2789 24868
rect 2740 24828 2746 24840
rect 2777 24837 2789 24840
rect 2823 24837 2835 24871
rect 2777 24831 2835 24837
rect 2866 24828 2872 24880
rect 2924 24868 2930 24880
rect 3329 24871 3387 24877
rect 3329 24868 3341 24871
rect 2924 24840 3341 24868
rect 2924 24828 2930 24840
rect 3329 24837 3341 24840
rect 3375 24868 3387 24871
rect 3375 24840 5212 24868
rect 3375 24837 3387 24840
rect 3329 24831 3387 24837
rect 1857 24803 1915 24809
rect 1857 24769 1869 24803
rect 1903 24800 1915 24803
rect 2038 24800 2044 24812
rect 1903 24772 2044 24800
rect 1903 24769 1915 24772
rect 1857 24763 1915 24769
rect 2038 24760 2044 24772
rect 2096 24760 2102 24812
rect 2133 24803 2191 24809
rect 2133 24769 2145 24803
rect 2179 24800 2191 24803
rect 2314 24800 2320 24812
rect 2179 24772 2320 24800
rect 2179 24769 2191 24772
rect 2133 24763 2191 24769
rect 2314 24760 2320 24772
rect 2372 24760 2378 24812
rect 2406 24760 2412 24812
rect 2464 24760 2470 24812
rect 3786 24760 3792 24812
rect 3844 24760 3850 24812
rect 4062 24760 4068 24812
rect 4120 24760 4126 24812
rect 5184 24809 5212 24840
rect 5534 24828 5540 24880
rect 5592 24828 5598 24880
rect 5169 24803 5227 24809
rect 5169 24769 5181 24803
rect 5215 24769 5227 24803
rect 5169 24763 5227 24769
rect 5353 24803 5411 24809
rect 5353 24769 5365 24803
rect 5399 24769 5411 24803
rect 5353 24763 5411 24769
rect 3237 24735 3295 24741
rect 3237 24701 3249 24735
rect 3283 24732 3295 24735
rect 4154 24732 4160 24744
rect 3283 24704 4160 24732
rect 3283 24701 3295 24704
rect 3237 24695 3295 24701
rect 2317 24667 2375 24673
rect 2317 24633 2329 24667
rect 2363 24664 2375 24667
rect 2777 24667 2835 24673
rect 2777 24664 2789 24667
rect 2363 24636 2789 24664
rect 2363 24633 2375 24636
rect 2317 24627 2375 24633
rect 2777 24633 2789 24636
rect 2823 24664 2835 24667
rect 3142 24664 3148 24676
rect 2823 24636 3148 24664
rect 2823 24633 2835 24636
rect 2777 24627 2835 24633
rect 3142 24624 3148 24636
rect 3200 24624 3206 24676
rect 2590 24556 2596 24608
rect 2648 24596 2654 24608
rect 3252 24596 3280 24695
rect 4154 24692 4160 24704
rect 4212 24692 4218 24744
rect 4338 24692 4344 24744
rect 4396 24692 4402 24744
rect 5368 24732 5396 24763
rect 5626 24760 5632 24812
rect 5684 24760 5690 24812
rect 5721 24803 5779 24809
rect 5721 24769 5733 24803
rect 5767 24800 5779 24803
rect 5810 24800 5816 24812
rect 5767 24772 5816 24800
rect 5767 24769 5779 24772
rect 5721 24763 5779 24769
rect 5810 24760 5816 24772
rect 5868 24800 5874 24812
rect 6086 24800 6092 24812
rect 5868 24772 6092 24800
rect 5868 24760 5874 24772
rect 6086 24760 6092 24772
rect 6144 24760 6150 24812
rect 6178 24760 6184 24812
rect 6236 24800 6242 24812
rect 6794 24800 6822 24908
rect 9030 24896 9036 24908
rect 9088 24896 9094 24948
rect 9950 24936 9956 24948
rect 9140 24908 9956 24936
rect 7190 24828 7196 24880
rect 7248 24828 7254 24880
rect 8662 24868 8668 24880
rect 7944 24840 8668 24868
rect 6236 24772 6822 24800
rect 7009 24803 7067 24809
rect 6236 24760 6242 24772
rect 7009 24769 7021 24803
rect 7055 24769 7067 24803
rect 7009 24763 7067 24769
rect 7285 24803 7343 24809
rect 7285 24769 7297 24803
rect 7331 24769 7343 24803
rect 7285 24763 7343 24769
rect 7377 24803 7435 24809
rect 7377 24769 7389 24803
rect 7423 24800 7435 24803
rect 7834 24800 7840 24812
rect 7423 24772 7840 24800
rect 7423 24769 7435 24772
rect 7377 24763 7435 24769
rect 7024 24732 7052 24763
rect 5368 24704 7052 24732
rect 6012 24676 6040 24704
rect 3602 24624 3608 24676
rect 3660 24664 3666 24676
rect 4062 24664 4068 24676
rect 3660 24636 4068 24664
rect 3660 24624 3666 24636
rect 4062 24624 4068 24636
rect 4120 24664 4126 24676
rect 4985 24667 5043 24673
rect 4985 24664 4997 24667
rect 4120 24636 4997 24664
rect 4120 24624 4126 24636
rect 4985 24633 4997 24636
rect 5031 24633 5043 24667
rect 4985 24627 5043 24633
rect 5902 24624 5908 24676
rect 5960 24624 5966 24676
rect 5994 24624 6000 24676
rect 6052 24624 6058 24676
rect 6914 24624 6920 24676
rect 6972 24664 6978 24676
rect 7300 24664 7328 24763
rect 7834 24760 7840 24772
rect 7892 24760 7898 24812
rect 7944 24664 7972 24840
rect 8662 24828 8668 24840
rect 8720 24828 8726 24880
rect 9140 24824 9168 24908
rect 9950 24896 9956 24908
rect 10008 24896 10014 24948
rect 11514 24896 11520 24948
rect 11572 24936 11578 24948
rect 12250 24936 12256 24948
rect 11572 24908 12256 24936
rect 11572 24896 11578 24908
rect 12250 24896 12256 24908
rect 12308 24896 12314 24948
rect 16390 24936 16396 24948
rect 12406 24908 16396 24936
rect 9217 24827 9275 24833
rect 10042 24828 10048 24880
rect 10100 24868 10106 24880
rect 12406 24868 12434 24908
rect 16390 24896 16396 24908
rect 16448 24896 16454 24948
rect 16666 24896 16672 24948
rect 16724 24896 16730 24948
rect 17862 24896 17868 24948
rect 17920 24936 17926 24948
rect 19886 24936 19892 24948
rect 17920 24908 19892 24936
rect 17920 24896 17926 24908
rect 19886 24896 19892 24908
rect 19944 24896 19950 24948
rect 20162 24896 20168 24948
rect 20220 24896 20226 24948
rect 21361 24939 21419 24945
rect 21361 24936 21373 24939
rect 20456 24908 21373 24936
rect 10100 24840 12434 24868
rect 12636 24840 13308 24868
rect 10100 24828 10106 24840
rect 9217 24824 9229 24827
rect 8297 24803 8355 24809
rect 8297 24769 8309 24803
rect 8343 24769 8355 24803
rect 8297 24763 8355 24769
rect 6972 24636 7328 24664
rect 7392 24636 7972 24664
rect 8312 24664 8340 24763
rect 8478 24760 8484 24812
rect 8536 24760 8542 24812
rect 8570 24760 8576 24812
rect 8628 24800 8634 24812
rect 8757 24803 8815 24809
rect 8757 24800 8769 24803
rect 8628 24772 8769 24800
rect 8628 24760 8634 24772
rect 8757 24769 8769 24772
rect 8803 24769 8815 24803
rect 9140 24796 9229 24824
rect 9217 24793 9229 24796
rect 9263 24793 9275 24827
rect 9217 24787 9275 24793
rect 9309 24806 9367 24809
rect 9309 24803 9444 24806
rect 8757 24763 8815 24769
rect 9309 24769 9321 24803
rect 9355 24778 9444 24803
rect 9355 24769 9367 24778
rect 9309 24763 9367 24769
rect 9416 24732 9444 24778
rect 9585 24803 9643 24809
rect 9585 24769 9597 24803
rect 9631 24790 9643 24803
rect 9674 24790 9680 24812
rect 9631 24769 9680 24790
rect 9585 24763 9680 24769
rect 9600 24762 9680 24763
rect 9674 24760 9680 24762
rect 9732 24760 9738 24812
rect 11514 24760 11520 24812
rect 11572 24760 11578 24812
rect 11698 24760 11704 24812
rect 11756 24760 11762 24812
rect 11790 24760 11796 24812
rect 11848 24760 11854 24812
rect 11885 24803 11943 24809
rect 11885 24769 11897 24803
rect 11931 24800 11943 24803
rect 12342 24800 12348 24812
rect 11931 24772 12348 24800
rect 11931 24769 11943 24772
rect 11885 24763 11943 24769
rect 12342 24760 12348 24772
rect 12400 24760 12406 24812
rect 9766 24732 9772 24744
rect 9416 24704 9772 24732
rect 9766 24692 9772 24704
rect 9824 24692 9830 24744
rect 12250 24692 12256 24744
rect 12308 24732 12314 24744
rect 12636 24732 12664 24840
rect 13280 24812 13308 24840
rect 13906 24828 13912 24880
rect 13964 24868 13970 24880
rect 14182 24868 14188 24880
rect 13964 24840 14188 24868
rect 13964 24828 13970 24840
rect 14182 24828 14188 24840
rect 14240 24828 14246 24880
rect 16114 24828 16120 24880
rect 16172 24868 16178 24880
rect 17957 24871 18015 24877
rect 16172 24840 17264 24868
rect 16172 24828 16178 24840
rect 12805 24803 12863 24809
rect 12805 24769 12817 24803
rect 12851 24769 12863 24803
rect 12805 24763 12863 24769
rect 12308 24704 12664 24732
rect 12308 24692 12314 24704
rect 8478 24664 8484 24676
rect 8312 24636 8484 24664
rect 6972 24624 6978 24636
rect 2648 24568 3280 24596
rect 2648 24556 2654 24568
rect 3694 24556 3700 24608
rect 3752 24596 3758 24608
rect 6546 24596 6552 24608
rect 3752 24568 6552 24596
rect 3752 24556 3758 24568
rect 6546 24556 6552 24568
rect 6604 24596 6610 24608
rect 7392 24596 7420 24636
rect 8478 24624 8484 24636
rect 8536 24664 8542 24676
rect 9033 24667 9091 24673
rect 9033 24664 9045 24667
rect 8536 24636 9045 24664
rect 8536 24624 8542 24636
rect 9033 24633 9045 24636
rect 9079 24633 9091 24667
rect 11514 24664 11520 24676
rect 9033 24627 9091 24633
rect 9416 24636 11520 24664
rect 6604 24568 7420 24596
rect 7561 24599 7619 24605
rect 6604 24556 6610 24568
rect 7561 24565 7573 24599
rect 7607 24596 7619 24599
rect 7742 24596 7748 24608
rect 7607 24568 7748 24596
rect 7607 24565 7619 24568
rect 7561 24559 7619 24565
rect 7742 24556 7748 24568
rect 7800 24556 7806 24608
rect 8941 24599 8999 24605
rect 8941 24565 8953 24599
rect 8987 24596 8999 24599
rect 9416 24596 9444 24636
rect 11514 24624 11520 24636
rect 11572 24624 11578 24676
rect 12820 24664 12848 24763
rect 13262 24760 13268 24812
rect 13320 24760 13326 24812
rect 13446 24760 13452 24812
rect 13504 24760 13510 24812
rect 13814 24760 13820 24812
rect 13872 24800 13878 24812
rect 14093 24803 14151 24809
rect 14093 24800 14105 24803
rect 13872 24772 14105 24800
rect 13872 24760 13878 24772
rect 14093 24769 14105 24772
rect 14139 24769 14151 24803
rect 14093 24763 14151 24769
rect 14369 24803 14427 24809
rect 14369 24769 14381 24803
rect 14415 24800 14427 24803
rect 14642 24800 14648 24812
rect 14415 24772 14648 24800
rect 14415 24769 14427 24772
rect 14369 24763 14427 24769
rect 14642 24760 14648 24772
rect 14700 24760 14706 24812
rect 14826 24760 14832 24812
rect 14884 24760 14890 24812
rect 15013 24803 15071 24809
rect 15013 24769 15025 24803
rect 15059 24800 15071 24803
rect 15102 24800 15108 24812
rect 15059 24772 15108 24800
rect 15059 24769 15071 24772
rect 15013 24763 15071 24769
rect 15102 24760 15108 24772
rect 15160 24760 15166 24812
rect 16298 24760 16304 24812
rect 16356 24800 16362 24812
rect 16666 24800 16672 24812
rect 16356 24772 16672 24800
rect 16356 24760 16362 24772
rect 16666 24760 16672 24772
rect 16724 24760 16730 24812
rect 16850 24760 16856 24812
rect 16908 24760 16914 24812
rect 16942 24760 16948 24812
rect 17000 24760 17006 24812
rect 17129 24803 17187 24809
rect 17129 24769 17141 24803
rect 17175 24769 17187 24803
rect 17129 24763 17187 24769
rect 13906 24732 13912 24744
rect 13648 24704 13912 24732
rect 13078 24664 13084 24676
rect 11992 24636 12848 24664
rect 12912 24636 13084 24664
rect 8987 24568 9444 24596
rect 8987 24565 8999 24568
rect 8941 24559 8999 24565
rect 9490 24556 9496 24608
rect 9548 24556 9554 24608
rect 9769 24599 9827 24605
rect 9769 24565 9781 24599
rect 9815 24596 9827 24599
rect 9950 24596 9956 24608
rect 9815 24568 9956 24596
rect 9815 24565 9827 24568
rect 9769 24559 9827 24565
rect 9950 24556 9956 24568
rect 10008 24596 10014 24608
rect 10686 24596 10692 24608
rect 10008 24568 10692 24596
rect 10008 24556 10014 24568
rect 10686 24556 10692 24568
rect 10744 24556 10750 24608
rect 11330 24556 11336 24608
rect 11388 24596 11394 24608
rect 11992 24596 12020 24636
rect 11388 24568 12020 24596
rect 12069 24599 12127 24605
rect 11388 24556 11394 24568
rect 12069 24565 12081 24599
rect 12115 24596 12127 24599
rect 12250 24596 12256 24608
rect 12115 24568 12256 24596
rect 12115 24565 12127 24568
rect 12069 24559 12127 24565
rect 12250 24556 12256 24568
rect 12308 24556 12314 24608
rect 12434 24556 12440 24608
rect 12492 24596 12498 24608
rect 12912 24596 12940 24636
rect 13078 24624 13084 24636
rect 13136 24624 13142 24676
rect 13648 24673 13676 24704
rect 13906 24692 13912 24704
rect 13964 24692 13970 24744
rect 14277 24735 14335 24741
rect 14277 24701 14289 24735
rect 14323 24732 14335 24735
rect 14918 24732 14924 24744
rect 14323 24704 14924 24732
rect 14323 24701 14335 24704
rect 14277 24695 14335 24701
rect 14918 24692 14924 24704
rect 14976 24692 14982 24744
rect 13633 24667 13691 24673
rect 13633 24633 13645 24667
rect 13679 24633 13691 24667
rect 13633 24627 13691 24633
rect 15930 24624 15936 24676
rect 15988 24664 15994 24676
rect 17144 24664 17172 24763
rect 17236 24732 17264 24840
rect 17957 24837 17969 24871
rect 18003 24868 18015 24871
rect 18230 24868 18236 24880
rect 18003 24840 18236 24868
rect 18003 24837 18015 24840
rect 17957 24831 18015 24837
rect 18230 24828 18236 24840
rect 18288 24828 18294 24880
rect 20180 24868 20208 24896
rect 18340 24840 20208 24868
rect 17586 24760 17592 24812
rect 17644 24760 17650 24812
rect 17773 24803 17831 24809
rect 17773 24769 17785 24803
rect 17819 24800 17831 24803
rect 18046 24800 18052 24812
rect 17819 24772 18052 24800
rect 17819 24769 17831 24772
rect 17773 24763 17831 24769
rect 18046 24760 18052 24772
rect 18104 24760 18110 24812
rect 18138 24760 18144 24812
rect 18196 24760 18202 24812
rect 18340 24809 18368 24840
rect 20254 24828 20260 24880
rect 20312 24868 20318 24880
rect 20312 24840 20392 24868
rect 20312 24828 20318 24840
rect 18325 24803 18383 24809
rect 18325 24769 18337 24803
rect 18371 24769 18383 24803
rect 18325 24763 18383 24769
rect 18340 24732 18368 24763
rect 18414 24760 18420 24812
rect 18472 24760 18478 24812
rect 18969 24803 19027 24809
rect 18969 24800 18981 24803
rect 18616 24772 18981 24800
rect 17236 24704 18368 24732
rect 15988 24636 17172 24664
rect 15988 24624 15994 24636
rect 18046 24624 18052 24676
rect 18104 24664 18110 24676
rect 18616 24673 18644 24772
rect 18969 24769 18981 24772
rect 19015 24769 19027 24803
rect 18969 24763 19027 24769
rect 19150 24760 19156 24812
rect 19208 24760 19214 24812
rect 19245 24803 19303 24809
rect 19245 24769 19257 24803
rect 19291 24800 19303 24803
rect 19334 24800 19340 24812
rect 19291 24772 19340 24800
rect 19291 24769 19303 24772
rect 19245 24763 19303 24769
rect 19334 24760 19340 24772
rect 19392 24760 19398 24812
rect 19610 24760 19616 24812
rect 19668 24800 19674 24812
rect 19668 24772 19840 24800
rect 19668 24760 19674 24772
rect 19812 24732 19840 24772
rect 19886 24760 19892 24812
rect 19944 24760 19950 24812
rect 19978 24760 19984 24812
rect 20036 24800 20042 24812
rect 20165 24803 20223 24809
rect 20165 24800 20177 24803
rect 20036 24772 20177 24800
rect 20036 24760 20042 24772
rect 20165 24769 20177 24772
rect 20211 24769 20223 24803
rect 20165 24763 20223 24769
rect 20257 24735 20315 24741
rect 20257 24732 20269 24735
rect 19812 24704 20269 24732
rect 20257 24701 20269 24704
rect 20303 24701 20315 24735
rect 20364 24732 20392 24840
rect 20456 24809 20484 24908
rect 21361 24905 21373 24908
rect 21407 24936 21419 24939
rect 22554 24936 22560 24948
rect 21407 24908 22560 24936
rect 21407 24905 21419 24908
rect 21361 24899 21419 24905
rect 22554 24896 22560 24908
rect 22612 24896 22618 24948
rect 22738 24896 22744 24948
rect 22796 24896 22802 24948
rect 22848 24908 23704 24936
rect 22005 24871 22063 24877
rect 22005 24837 22017 24871
rect 22051 24868 22063 24871
rect 22094 24868 22100 24880
rect 22051 24840 22100 24868
rect 22051 24837 22063 24840
rect 20441 24803 20499 24809
rect 20441 24769 20453 24803
rect 20487 24769 20499 24803
rect 20441 24763 20499 24769
rect 20717 24803 20775 24809
rect 20717 24769 20729 24803
rect 20763 24769 20775 24803
rect 20717 24763 20775 24769
rect 21177 24803 21235 24809
rect 21177 24769 21189 24803
rect 21223 24800 21235 24803
rect 21358 24800 21364 24812
rect 21223 24772 21364 24800
rect 21223 24769 21235 24772
rect 21177 24763 21235 24769
rect 20732 24732 20760 24763
rect 21358 24760 21364 24772
rect 21416 24760 21422 24812
rect 21450 24784 21456 24836
rect 21508 24784 21514 24836
rect 22005 24831 22063 24837
rect 22094 24828 22100 24840
rect 22152 24868 22158 24880
rect 22848 24868 22876 24908
rect 22152 24840 22876 24868
rect 22152 24828 22158 24840
rect 22922 24828 22928 24880
rect 22980 24868 22986 24880
rect 23676 24868 23704 24908
rect 23750 24896 23756 24948
rect 23808 24896 23814 24948
rect 24854 24936 24860 24948
rect 23860 24908 24860 24936
rect 23860 24868 23888 24908
rect 24854 24896 24860 24908
rect 24912 24896 24918 24948
rect 27985 24939 28043 24945
rect 27985 24905 27997 24939
rect 28031 24905 28043 24939
rect 27985 24899 28043 24905
rect 22980 24840 23612 24868
rect 23676 24840 23888 24868
rect 22980 24828 22986 24840
rect 22186 24760 22192 24812
rect 22244 24760 22250 24812
rect 22462 24760 22468 24812
rect 22520 24760 22526 24812
rect 22554 24760 22560 24812
rect 22612 24760 22618 24812
rect 23106 24760 23112 24812
rect 23164 24800 23170 24812
rect 23293 24803 23351 24809
rect 23293 24800 23305 24803
rect 23164 24772 23305 24800
rect 23164 24760 23170 24772
rect 23293 24769 23305 24772
rect 23339 24769 23351 24803
rect 23293 24763 23351 24769
rect 23385 24803 23443 24809
rect 23385 24769 23397 24803
rect 23431 24769 23443 24803
rect 23385 24763 23443 24769
rect 20364 24704 20760 24732
rect 20809 24735 20867 24741
rect 20257 24695 20315 24701
rect 20809 24701 20821 24735
rect 20855 24732 20867 24735
rect 21450 24732 21456 24744
rect 20855 24704 21456 24732
rect 20855 24701 20867 24704
rect 20809 24695 20867 24701
rect 21450 24692 21456 24704
rect 21508 24692 21514 24744
rect 21560 24704 23060 24732
rect 18601 24667 18659 24673
rect 18104 24636 18368 24664
rect 18104 24624 18110 24636
rect 12492 24568 12940 24596
rect 12492 24556 12498 24568
rect 12986 24556 12992 24608
rect 13044 24556 13050 24608
rect 14366 24556 14372 24608
rect 14424 24556 14430 24608
rect 14550 24556 14556 24608
rect 14608 24556 14614 24608
rect 14642 24556 14648 24608
rect 14700 24556 14706 24608
rect 17129 24599 17187 24605
rect 17129 24565 17141 24599
rect 17175 24596 17187 24599
rect 17402 24596 17408 24608
rect 17175 24568 17408 24596
rect 17175 24565 17187 24568
rect 17129 24559 17187 24565
rect 17402 24556 17408 24568
rect 17460 24556 17466 24608
rect 18230 24556 18236 24608
rect 18288 24556 18294 24608
rect 18340 24596 18368 24636
rect 18601 24633 18613 24667
rect 18647 24633 18659 24667
rect 21085 24667 21143 24673
rect 18601 24627 18659 24633
rect 18708 24636 21036 24664
rect 18708 24596 18736 24636
rect 18340 24568 18736 24596
rect 19242 24556 19248 24608
rect 19300 24556 19306 24608
rect 19426 24556 19432 24608
rect 19484 24556 19490 24608
rect 19886 24556 19892 24608
rect 19944 24596 19950 24608
rect 20073 24599 20131 24605
rect 20073 24596 20085 24599
rect 19944 24568 20085 24596
rect 19944 24556 19950 24568
rect 20073 24565 20085 24568
rect 20119 24565 20131 24599
rect 20073 24559 20131 24565
rect 20162 24556 20168 24608
rect 20220 24556 20226 24608
rect 20530 24556 20536 24608
rect 20588 24596 20594 24608
rect 20625 24599 20683 24605
rect 20625 24596 20637 24599
rect 20588 24568 20637 24596
rect 20588 24556 20594 24568
rect 20625 24565 20637 24568
rect 20671 24565 20683 24599
rect 20625 24559 20683 24565
rect 20714 24556 20720 24608
rect 20772 24556 20778 24608
rect 21008 24596 21036 24636
rect 21085 24633 21097 24667
rect 21131 24664 21143 24667
rect 21266 24664 21272 24676
rect 21131 24636 21272 24664
rect 21131 24633 21143 24636
rect 21085 24627 21143 24633
rect 21266 24624 21272 24636
rect 21324 24624 21330 24676
rect 21560 24596 21588 24704
rect 21818 24624 21824 24676
rect 21876 24624 21882 24676
rect 22094 24624 22100 24676
rect 22152 24664 22158 24676
rect 22281 24667 22339 24673
rect 22281 24664 22293 24667
rect 22152 24636 22293 24664
rect 22152 24624 22158 24636
rect 22281 24633 22293 24636
rect 22327 24633 22339 24667
rect 22281 24627 22339 24633
rect 22738 24624 22744 24676
rect 22796 24664 22802 24676
rect 22925 24667 22983 24673
rect 22925 24664 22937 24667
rect 22796 24636 22937 24664
rect 22796 24624 22802 24636
rect 22925 24633 22937 24636
rect 22971 24633 22983 24667
rect 23032 24664 23060 24704
rect 23198 24692 23204 24744
rect 23256 24692 23262 24744
rect 23400 24664 23428 24763
rect 23474 24760 23480 24812
rect 23532 24760 23538 24812
rect 23584 24800 23612 24840
rect 24210 24828 24216 24880
rect 24268 24868 24274 24880
rect 26694 24868 26700 24880
rect 24268 24840 26700 24868
rect 24268 24828 24274 24840
rect 26694 24828 26700 24840
rect 26752 24828 26758 24880
rect 23845 24803 23903 24809
rect 23845 24800 23857 24803
rect 23584 24772 23857 24800
rect 23845 24769 23857 24772
rect 23891 24769 23903 24803
rect 23845 24763 23903 24769
rect 23934 24760 23940 24812
rect 23992 24800 23998 24812
rect 24029 24803 24087 24809
rect 24029 24800 24041 24803
rect 23992 24772 24041 24800
rect 23992 24760 23998 24772
rect 24029 24769 24041 24772
rect 24075 24769 24087 24803
rect 24029 24763 24087 24769
rect 26786 24760 26792 24812
rect 26844 24800 26850 24812
rect 27525 24803 27583 24809
rect 27525 24800 27537 24803
rect 26844 24772 27537 24800
rect 26844 24760 26850 24772
rect 27525 24769 27537 24772
rect 27571 24769 27583 24803
rect 27525 24763 27583 24769
rect 27801 24803 27859 24809
rect 27801 24769 27813 24803
rect 27847 24769 27859 24803
rect 28000 24800 28028 24899
rect 28074 24800 28080 24812
rect 28000 24772 28080 24800
rect 27801 24763 27859 24769
rect 24213 24735 24271 24741
rect 24213 24701 24225 24735
rect 24259 24732 24271 24735
rect 24302 24732 24308 24744
rect 24259 24704 24308 24732
rect 24259 24701 24271 24704
rect 24213 24695 24271 24701
rect 24302 24692 24308 24704
rect 24360 24692 24366 24744
rect 23032 24636 23428 24664
rect 22925 24627 22983 24633
rect 23842 24624 23848 24676
rect 23900 24664 23906 24676
rect 25958 24664 25964 24676
rect 23900 24636 25964 24664
rect 23900 24624 23906 24636
rect 25958 24624 25964 24636
rect 26016 24624 26022 24676
rect 27709 24667 27767 24673
rect 27709 24633 27721 24667
rect 27755 24664 27767 24667
rect 27816 24664 27844 24763
rect 28074 24760 28080 24772
rect 28132 24760 28138 24812
rect 28166 24760 28172 24812
rect 28224 24760 28230 24812
rect 28258 24760 28264 24812
rect 28316 24800 28322 24812
rect 28445 24803 28503 24809
rect 28445 24800 28457 24803
rect 28316 24772 28457 24800
rect 28316 24760 28322 24772
rect 28445 24769 28457 24772
rect 28491 24769 28503 24803
rect 28445 24763 28503 24769
rect 29362 24760 29368 24812
rect 29420 24800 29426 24812
rect 30193 24803 30251 24809
rect 30193 24800 30205 24803
rect 29420 24772 30205 24800
rect 29420 24760 29426 24772
rect 30193 24769 30205 24772
rect 30239 24800 30251 24803
rect 31570 24800 31576 24812
rect 30239 24772 31576 24800
rect 30239 24769 30251 24772
rect 30193 24763 30251 24769
rect 31570 24760 31576 24772
rect 31628 24760 31634 24812
rect 31846 24760 31852 24812
rect 31904 24760 31910 24812
rect 32214 24760 32220 24812
rect 32272 24760 32278 24812
rect 28353 24735 28411 24741
rect 28353 24701 28365 24735
rect 28399 24732 28411 24735
rect 28534 24732 28540 24744
rect 28399 24704 28540 24732
rect 28399 24701 28411 24704
rect 28353 24695 28411 24701
rect 28534 24692 28540 24704
rect 28592 24692 28598 24744
rect 30466 24692 30472 24744
rect 30524 24692 30530 24744
rect 28258 24664 28264 24676
rect 27755 24636 28264 24664
rect 27755 24633 27767 24636
rect 27709 24627 27767 24633
rect 28258 24624 28264 24636
rect 28316 24624 28322 24676
rect 28629 24667 28687 24673
rect 28629 24633 28641 24667
rect 28675 24664 28687 24667
rect 29638 24664 29644 24676
rect 28675 24636 29644 24664
rect 28675 24633 28687 24636
rect 28629 24627 28687 24633
rect 29638 24624 29644 24636
rect 29696 24624 29702 24676
rect 21008 24568 21588 24596
rect 21634 24556 21640 24608
rect 21692 24596 21698 24608
rect 22830 24596 22836 24608
rect 21692 24568 22836 24596
rect 21692 24556 21698 24568
rect 22830 24556 22836 24568
rect 22888 24556 22894 24608
rect 23290 24556 23296 24608
rect 23348 24556 23354 24608
rect 23382 24556 23388 24608
rect 23440 24556 23446 24608
rect 24302 24556 24308 24608
rect 24360 24596 24366 24608
rect 24486 24596 24492 24608
rect 24360 24568 24492 24596
rect 24360 24556 24366 24568
rect 24486 24556 24492 24568
rect 24544 24556 24550 24608
rect 25130 24556 25136 24608
rect 25188 24596 25194 24608
rect 28169 24599 28227 24605
rect 28169 24596 28181 24599
rect 25188 24568 28181 24596
rect 25188 24556 25194 24568
rect 28169 24565 28181 24568
rect 28215 24565 28227 24599
rect 28169 24559 28227 24565
rect 29178 24556 29184 24608
rect 29236 24596 29242 24608
rect 31297 24599 31355 24605
rect 31297 24596 31309 24599
rect 29236 24568 31309 24596
rect 29236 24556 29242 24568
rect 31297 24565 31309 24568
rect 31343 24565 31355 24599
rect 31297 24559 31355 24565
rect 32401 24599 32459 24605
rect 32401 24565 32413 24599
rect 32447 24596 32459 24599
rect 32490 24596 32496 24608
rect 32447 24568 32496 24596
rect 32447 24565 32459 24568
rect 32401 24559 32459 24565
rect 32490 24556 32496 24568
rect 32548 24556 32554 24608
rect 1104 24506 32844 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 32844 24506
rect 1104 24432 32844 24454
rect 1581 24395 1639 24401
rect 1581 24361 1593 24395
rect 1627 24392 1639 24395
rect 1670 24392 1676 24404
rect 1627 24364 1676 24392
rect 1627 24361 1639 24364
rect 1581 24355 1639 24361
rect 1670 24352 1676 24364
rect 1728 24352 1734 24404
rect 2130 24352 2136 24404
rect 2188 24352 2194 24404
rect 3418 24392 3424 24404
rect 2884 24364 3424 24392
rect 2682 24324 2688 24336
rect 2332 24296 2688 24324
rect 2332 24265 2360 24296
rect 2682 24284 2688 24296
rect 2740 24284 2746 24336
rect 2884 24333 2912 24364
rect 3418 24352 3424 24364
rect 3476 24352 3482 24404
rect 3605 24395 3663 24401
rect 3605 24361 3617 24395
rect 3651 24392 3663 24395
rect 3694 24392 3700 24404
rect 3651 24364 3700 24392
rect 3651 24361 3663 24364
rect 3605 24355 3663 24361
rect 3694 24352 3700 24364
rect 3752 24352 3758 24404
rect 4338 24352 4344 24404
rect 4396 24392 4402 24404
rect 4706 24392 4712 24404
rect 4396 24364 4712 24392
rect 4396 24352 4402 24364
rect 4706 24352 4712 24364
rect 4764 24352 4770 24404
rect 5350 24352 5356 24404
rect 5408 24352 5414 24404
rect 6178 24392 6184 24404
rect 5552 24364 6184 24392
rect 2869 24327 2927 24333
rect 2869 24293 2881 24327
rect 2915 24293 2927 24327
rect 2869 24287 2927 24293
rect 3881 24327 3939 24333
rect 3881 24293 3893 24327
rect 3927 24324 3939 24327
rect 4154 24324 4160 24336
rect 3927 24296 4160 24324
rect 3927 24293 3939 24296
rect 3881 24287 3939 24293
rect 4154 24284 4160 24296
rect 4212 24284 4218 24336
rect 4617 24327 4675 24333
rect 4617 24293 4629 24327
rect 4663 24324 4675 24327
rect 5552 24324 5580 24364
rect 6178 24352 6184 24364
rect 6236 24352 6242 24404
rect 6365 24395 6423 24401
rect 6365 24361 6377 24395
rect 6411 24392 6423 24395
rect 6914 24392 6920 24404
rect 6411 24364 6920 24392
rect 6411 24361 6423 24364
rect 6365 24355 6423 24361
rect 4663 24296 5580 24324
rect 4663 24293 4675 24296
rect 4617 24287 4675 24293
rect 5626 24284 5632 24336
rect 5684 24324 5690 24336
rect 6380 24324 6408 24355
rect 6914 24352 6920 24364
rect 6972 24352 6978 24404
rect 8757 24395 8815 24401
rect 8757 24361 8769 24395
rect 8803 24392 8815 24395
rect 8938 24392 8944 24404
rect 8803 24364 8944 24392
rect 8803 24361 8815 24364
rect 8757 24355 8815 24361
rect 8938 24352 8944 24364
rect 8996 24352 9002 24404
rect 9306 24352 9312 24404
rect 9364 24392 9370 24404
rect 11057 24395 11115 24401
rect 11057 24392 11069 24395
rect 9364 24364 9996 24392
rect 9364 24352 9370 24364
rect 5684 24296 6408 24324
rect 5684 24284 5690 24296
rect 2317 24259 2375 24265
rect 2317 24225 2329 24259
rect 2363 24225 2375 24259
rect 2317 24219 2375 24225
rect 2409 24259 2467 24265
rect 2409 24225 2421 24259
rect 2455 24256 2467 24259
rect 3142 24256 3148 24268
rect 2455 24228 3148 24256
rect 2455 24225 2467 24228
rect 2409 24219 2467 24225
rect 3142 24216 3148 24228
rect 3200 24216 3206 24268
rect 3326 24216 3332 24268
rect 3384 24256 3390 24268
rect 3421 24259 3479 24265
rect 3421 24256 3433 24259
rect 3384 24228 3433 24256
rect 3384 24216 3390 24228
rect 3421 24225 3433 24228
rect 3467 24225 3479 24259
rect 3421 24219 3479 24225
rect 3970 24216 3976 24268
rect 4028 24256 4034 24268
rect 4341 24259 4399 24265
rect 4341 24256 4353 24259
rect 4028 24228 4353 24256
rect 4028 24216 4034 24228
rect 4341 24225 4353 24228
rect 4387 24225 4399 24259
rect 4341 24219 4399 24225
rect 4448 24228 5028 24256
rect 842 24148 848 24200
rect 900 24188 906 24200
rect 1397 24191 1455 24197
rect 1397 24188 1409 24191
rect 900 24160 1409 24188
rect 900 24148 906 24160
rect 1397 24157 1409 24160
rect 1443 24157 1455 24191
rect 1397 24151 1455 24157
rect 1854 24148 1860 24200
rect 1912 24148 1918 24200
rect 2501 24191 2559 24197
rect 2501 24157 2513 24191
rect 2547 24157 2559 24191
rect 2501 24151 2559 24157
rect 2516 24120 2544 24151
rect 2590 24148 2596 24200
rect 2648 24148 2654 24200
rect 2682 24148 2688 24200
rect 2740 24188 2746 24200
rect 4448 24188 4476 24228
rect 5000 24197 5028 24228
rect 2740 24160 4476 24188
rect 4709 24191 4767 24197
rect 2740 24148 2746 24160
rect 2774 24120 2780 24132
rect 2516 24092 2780 24120
rect 2774 24080 2780 24092
rect 2832 24080 2838 24132
rect 2884 24129 2912 24160
rect 4709 24157 4721 24191
rect 4755 24157 4767 24191
rect 4709 24151 4767 24157
rect 4985 24191 5043 24197
rect 4985 24157 4997 24191
rect 5031 24157 5043 24191
rect 4985 24151 5043 24157
rect 2869 24123 2927 24129
rect 2869 24089 2881 24123
rect 2915 24089 2927 24123
rect 3881 24123 3939 24129
rect 3881 24120 3893 24123
rect 2869 24083 2927 24089
rect 3344 24092 3893 24120
rect 3344 24064 3372 24092
rect 3881 24089 3893 24092
rect 3927 24120 3939 24123
rect 4715 24120 4743 24151
rect 5442 24148 5448 24200
rect 5500 24148 5506 24200
rect 5721 24191 5779 24197
rect 5721 24157 5733 24191
rect 5767 24188 5779 24191
rect 5920 24188 5948 24296
rect 6730 24284 6736 24336
rect 6788 24324 6794 24336
rect 7650 24324 7656 24336
rect 6788 24296 7656 24324
rect 6788 24284 6794 24296
rect 7650 24284 7656 24296
rect 7708 24284 7714 24336
rect 9493 24327 9551 24333
rect 9493 24293 9505 24327
rect 9539 24324 9551 24327
rect 9674 24324 9680 24336
rect 9539 24296 9680 24324
rect 9539 24293 9551 24296
rect 9493 24287 9551 24293
rect 9674 24284 9680 24296
rect 9732 24284 9738 24336
rect 6012 24228 7236 24256
rect 6012 24200 6040 24228
rect 5767 24160 5948 24188
rect 5767 24157 5779 24160
rect 5721 24151 5779 24157
rect 5994 24148 6000 24200
rect 6052 24148 6058 24200
rect 6086 24148 6092 24200
rect 6144 24148 6150 24200
rect 6546 24148 6552 24200
rect 6604 24148 6610 24200
rect 6914 24148 6920 24200
rect 6972 24148 6978 24200
rect 7006 24148 7012 24200
rect 7064 24188 7070 24200
rect 7208 24197 7236 24228
rect 8956 24228 9904 24256
rect 8956 24200 8984 24228
rect 7101 24191 7159 24197
rect 7101 24188 7113 24191
rect 7064 24160 7113 24188
rect 7064 24148 7070 24160
rect 7101 24157 7113 24160
rect 7147 24157 7159 24191
rect 7101 24151 7159 24157
rect 7193 24191 7251 24197
rect 7193 24157 7205 24191
rect 7239 24157 7251 24191
rect 7193 24151 7251 24157
rect 7285 24191 7343 24197
rect 7285 24157 7297 24191
rect 7331 24188 7343 24191
rect 7374 24188 7380 24200
rect 7331 24160 7380 24188
rect 7331 24157 7343 24160
rect 7285 24151 7343 24157
rect 7374 24148 7380 24160
rect 7432 24148 7438 24200
rect 8573 24191 8631 24197
rect 8573 24157 8585 24191
rect 8619 24188 8631 24191
rect 8662 24188 8668 24200
rect 8619 24160 8668 24188
rect 8619 24157 8631 24160
rect 8573 24151 8631 24157
rect 8662 24148 8668 24160
rect 8720 24148 8726 24200
rect 8938 24148 8944 24200
rect 8996 24148 9002 24200
rect 9217 24191 9275 24197
rect 9217 24188 9229 24191
rect 9048 24160 9229 24188
rect 3927 24092 4743 24120
rect 3927 24089 3939 24092
rect 3881 24083 3939 24089
rect 4798 24080 4804 24132
rect 4856 24120 4862 24132
rect 5077 24123 5135 24129
rect 5077 24120 5089 24123
rect 4856 24092 5089 24120
rect 4856 24080 4862 24092
rect 5077 24089 5089 24092
rect 5123 24089 5135 24123
rect 5077 24083 5135 24089
rect 5194 24123 5252 24129
rect 5194 24089 5206 24123
rect 5240 24089 5252 24123
rect 5194 24083 5252 24089
rect 2041 24055 2099 24061
rect 2041 24021 2053 24055
rect 2087 24052 2099 24055
rect 3326 24052 3332 24064
rect 2087 24024 3332 24052
rect 2087 24021 2099 24024
rect 2041 24015 2099 24021
rect 3326 24012 3332 24024
rect 3384 24012 3390 24064
rect 3418 24012 3424 24064
rect 3476 24052 3482 24064
rect 4433 24055 4491 24061
rect 4433 24052 4445 24055
rect 3476 24024 4445 24052
rect 3476 24012 3482 24024
rect 4433 24021 4445 24024
rect 4479 24052 4491 24055
rect 5209 24052 5237 24083
rect 5534 24080 5540 24132
rect 5592 24120 5598 24132
rect 5905 24123 5963 24129
rect 5905 24120 5917 24123
rect 5592 24092 5917 24120
rect 5592 24080 5598 24092
rect 5905 24089 5917 24092
rect 5951 24089 5963 24123
rect 6730 24120 6736 24132
rect 5905 24083 5963 24089
rect 6196 24092 6736 24120
rect 6196 24064 6224 24092
rect 6730 24080 6736 24092
rect 6788 24080 6794 24132
rect 8846 24120 8852 24132
rect 7392 24092 8852 24120
rect 4479 24024 5237 24052
rect 5629 24055 5687 24061
rect 4479 24021 4491 24024
rect 4433 24015 4491 24021
rect 5629 24021 5641 24055
rect 5675 24052 5687 24055
rect 6178 24052 6184 24064
rect 5675 24024 6184 24052
rect 5675 24021 5687 24024
rect 5629 24015 5687 24021
rect 6178 24012 6184 24024
rect 6236 24012 6242 24064
rect 6273 24055 6331 24061
rect 6273 24021 6285 24055
rect 6319 24052 6331 24055
rect 7392 24052 7420 24092
rect 8846 24080 8852 24092
rect 8904 24080 8910 24132
rect 9048 24120 9076 24160
rect 9217 24157 9229 24160
rect 9263 24157 9275 24191
rect 9217 24151 9275 24157
rect 8956 24092 9076 24120
rect 6319 24024 7420 24052
rect 6319 24021 6331 24024
rect 6273 24015 6331 24021
rect 7466 24012 7472 24064
rect 7524 24012 7530 24064
rect 8478 24012 8484 24064
rect 8536 24052 8542 24064
rect 8956 24052 8984 24092
rect 9122 24080 9128 24132
rect 9180 24080 9186 24132
rect 9232 24120 9260 24151
rect 9306 24148 9312 24200
rect 9364 24148 9370 24200
rect 9876 24197 9904 24228
rect 9968 24197 9996 24364
rect 10520 24364 11069 24392
rect 10134 24216 10140 24268
rect 10192 24256 10198 24268
rect 10192 24228 10456 24256
rect 10192 24216 10198 24228
rect 10428 24197 10456 24228
rect 10520 24200 10548 24364
rect 11057 24361 11069 24364
rect 11103 24392 11115 24395
rect 11146 24392 11152 24404
rect 11103 24364 11152 24392
rect 11103 24361 11115 24364
rect 11057 24355 11115 24361
rect 11146 24352 11152 24364
rect 11204 24352 11210 24404
rect 11333 24395 11391 24401
rect 11333 24361 11345 24395
rect 11379 24392 11391 24395
rect 11422 24392 11428 24404
rect 11379 24364 11428 24392
rect 11379 24361 11391 24364
rect 11333 24355 11391 24361
rect 11422 24352 11428 24364
rect 11480 24352 11486 24404
rect 12986 24352 12992 24404
rect 13044 24392 13050 24404
rect 16298 24392 16304 24404
rect 13044 24364 16304 24392
rect 13044 24352 13050 24364
rect 16298 24352 16304 24364
rect 16356 24352 16362 24404
rect 16390 24352 16396 24404
rect 16448 24392 16454 24404
rect 18138 24392 18144 24404
rect 16448 24364 18144 24392
rect 16448 24352 16454 24364
rect 18138 24352 18144 24364
rect 18196 24352 18202 24404
rect 19334 24352 19340 24404
rect 19392 24392 19398 24404
rect 20530 24392 20536 24404
rect 19392 24364 20536 24392
rect 19392 24352 19398 24364
rect 20530 24352 20536 24364
rect 20588 24352 20594 24404
rect 20717 24395 20775 24401
rect 20717 24361 20729 24395
rect 20763 24392 20775 24395
rect 20806 24392 20812 24404
rect 20763 24364 20812 24392
rect 20763 24361 20775 24364
rect 20717 24355 20775 24361
rect 20806 24352 20812 24364
rect 20864 24352 20870 24404
rect 21085 24395 21143 24401
rect 21085 24361 21097 24395
rect 21131 24361 21143 24395
rect 21085 24355 21143 24361
rect 10781 24327 10839 24333
rect 10781 24293 10793 24327
rect 10827 24293 10839 24327
rect 10781 24287 10839 24293
rect 10796 24256 10824 24287
rect 11514 24284 11520 24336
rect 11572 24324 11578 24336
rect 14458 24324 14464 24336
rect 11572 24296 14464 24324
rect 11572 24284 11578 24296
rect 14458 24284 14464 24296
rect 14516 24284 14522 24336
rect 15102 24284 15108 24336
rect 15160 24324 15166 24336
rect 19610 24324 19616 24336
rect 15160 24296 19616 24324
rect 15160 24284 15166 24296
rect 19610 24284 19616 24296
rect 19668 24284 19674 24336
rect 21100 24324 21128 24355
rect 21542 24352 21548 24404
rect 21600 24392 21606 24404
rect 22186 24392 22192 24404
rect 21600 24364 22192 24392
rect 21600 24352 21606 24364
rect 22186 24352 22192 24364
rect 22244 24392 22250 24404
rect 22646 24392 22652 24404
rect 22244 24364 22652 24392
rect 22244 24352 22250 24364
rect 22646 24352 22652 24364
rect 22704 24352 22710 24404
rect 23845 24395 23903 24401
rect 23845 24361 23857 24395
rect 23891 24392 23903 24395
rect 24854 24392 24860 24404
rect 23891 24364 24860 24392
rect 23891 24361 23903 24364
rect 23845 24355 23903 24361
rect 24854 24352 24860 24364
rect 24912 24352 24918 24404
rect 25222 24352 25228 24404
rect 25280 24392 25286 24404
rect 25317 24395 25375 24401
rect 25317 24392 25329 24395
rect 25280 24364 25329 24392
rect 25280 24352 25286 24364
rect 25317 24361 25329 24364
rect 25363 24361 25375 24395
rect 25317 24355 25375 24361
rect 25685 24395 25743 24401
rect 25685 24361 25697 24395
rect 25731 24392 25743 24395
rect 27890 24392 27896 24404
rect 25731 24364 27896 24392
rect 25731 24361 25743 24364
rect 25685 24355 25743 24361
rect 27890 24352 27896 24364
rect 27948 24352 27954 24404
rect 28074 24352 28080 24404
rect 28132 24352 28138 24404
rect 28169 24395 28227 24401
rect 28169 24361 28181 24395
rect 28215 24361 28227 24395
rect 28169 24355 28227 24361
rect 21174 24324 21180 24336
rect 21100 24296 21180 24324
rect 21174 24284 21180 24296
rect 21232 24324 21238 24336
rect 28184 24324 28212 24355
rect 21232 24296 28212 24324
rect 21232 24284 21238 24296
rect 10796 24228 12940 24256
rect 9585 24191 9643 24197
rect 9585 24157 9597 24191
rect 9631 24157 9643 24191
rect 9585 24151 9643 24157
rect 9861 24191 9919 24197
rect 9861 24157 9873 24191
rect 9907 24157 9919 24191
rect 9861 24151 9919 24157
rect 9953 24191 10011 24197
rect 9953 24157 9965 24191
rect 9999 24157 10011 24191
rect 9953 24151 10011 24157
rect 10229 24191 10287 24197
rect 10229 24157 10241 24191
rect 10275 24188 10287 24191
rect 10413 24191 10471 24197
rect 10275 24160 10364 24188
rect 10275 24157 10287 24160
rect 10229 24151 10287 24157
rect 9600 24120 9628 24151
rect 9232 24092 9628 24120
rect 9769 24123 9827 24129
rect 9769 24089 9781 24123
rect 9815 24089 9827 24123
rect 9769 24083 9827 24089
rect 8536 24024 8984 24052
rect 9140 24052 9168 24080
rect 9784 24052 9812 24083
rect 9140 24024 9812 24052
rect 8536 24012 8542 24024
rect 9950 24012 9956 24064
rect 10008 24052 10014 24064
rect 10137 24055 10195 24061
rect 10137 24052 10149 24055
rect 10008 24024 10149 24052
rect 10008 24012 10014 24024
rect 10137 24021 10149 24024
rect 10183 24021 10195 24055
rect 10336 24052 10364 24160
rect 10413 24157 10425 24191
rect 10459 24157 10471 24191
rect 10413 24151 10471 24157
rect 10428 24120 10456 24151
rect 10502 24148 10508 24200
rect 10560 24148 10566 24200
rect 10594 24148 10600 24200
rect 10652 24148 10658 24200
rect 10686 24148 10692 24200
rect 10744 24188 10750 24200
rect 10873 24191 10931 24197
rect 10873 24188 10885 24191
rect 10744 24160 10885 24188
rect 10744 24148 10750 24160
rect 10873 24157 10885 24160
rect 10919 24157 10931 24191
rect 10873 24151 10931 24157
rect 11149 24191 11207 24197
rect 11149 24157 11161 24191
rect 11195 24188 11207 24191
rect 11238 24188 11244 24200
rect 11195 24160 11244 24188
rect 11195 24157 11207 24160
rect 11149 24151 11207 24157
rect 10778 24120 10784 24132
rect 10428 24092 10784 24120
rect 10778 24080 10784 24092
rect 10836 24080 10842 24132
rect 10888 24120 10916 24151
rect 11238 24148 11244 24160
rect 11296 24148 11302 24200
rect 12912 24188 12940 24228
rect 13170 24216 13176 24268
rect 13228 24256 13234 24268
rect 20162 24256 20168 24268
rect 13228 24228 20168 24256
rect 13228 24216 13234 24228
rect 20162 24216 20168 24228
rect 20220 24216 20226 24268
rect 20993 24259 21051 24265
rect 20993 24225 21005 24259
rect 21039 24256 21051 24259
rect 21634 24256 21640 24268
rect 21039 24228 21640 24256
rect 21039 24225 21051 24228
rect 20993 24219 21051 24225
rect 21634 24216 21640 24228
rect 21692 24216 21698 24268
rect 24210 24216 24216 24268
rect 24268 24256 24274 24268
rect 27985 24259 28043 24265
rect 24268 24228 27844 24256
rect 24268 24216 24274 24228
rect 14090 24188 14096 24200
rect 12912 24160 14096 24188
rect 14090 24148 14096 24160
rect 14148 24148 14154 24200
rect 14182 24148 14188 24200
rect 14240 24188 14246 24200
rect 20806 24188 20812 24200
rect 14240 24160 20812 24188
rect 14240 24148 14246 24160
rect 20806 24148 20812 24160
rect 20864 24188 20870 24200
rect 21085 24191 21143 24197
rect 21085 24188 21097 24191
rect 20864 24160 21097 24188
rect 20864 24148 20870 24160
rect 21085 24157 21097 24160
rect 21131 24157 21143 24191
rect 21085 24151 21143 24157
rect 21174 24148 21180 24200
rect 21232 24188 21238 24200
rect 21453 24191 21511 24197
rect 21453 24188 21465 24191
rect 21232 24160 21465 24188
rect 21232 24148 21238 24160
rect 21453 24157 21465 24160
rect 21499 24157 21511 24191
rect 21729 24191 21787 24197
rect 21729 24188 21741 24191
rect 21453 24151 21511 24157
rect 21560 24160 21741 24188
rect 11882 24120 11888 24132
rect 10888 24092 11888 24120
rect 11882 24080 11888 24092
rect 11940 24080 11946 24132
rect 11977 24123 12035 24129
rect 11977 24089 11989 24123
rect 12023 24089 12035 24123
rect 11977 24083 12035 24089
rect 12161 24123 12219 24129
rect 12161 24089 12173 24123
rect 12207 24120 12219 24123
rect 12618 24120 12624 24132
rect 12207 24092 12624 24120
rect 12207 24089 12219 24092
rect 12161 24083 12219 24089
rect 11422 24052 11428 24064
rect 10336 24024 11428 24052
rect 10137 24015 10195 24021
rect 11422 24012 11428 24024
rect 11480 24012 11486 24064
rect 11790 24012 11796 24064
rect 11848 24012 11854 24064
rect 11992 24052 12020 24083
rect 12618 24080 12624 24092
rect 12676 24120 12682 24132
rect 13078 24120 13084 24132
rect 12676 24092 13084 24120
rect 12676 24080 12682 24092
rect 13078 24080 13084 24092
rect 13136 24080 13142 24132
rect 14274 24080 14280 24132
rect 14332 24120 14338 24132
rect 21560 24120 21588 24160
rect 21729 24157 21741 24160
rect 21775 24157 21787 24191
rect 21729 24151 21787 24157
rect 22833 24191 22891 24197
rect 22833 24157 22845 24191
rect 22879 24188 22891 24191
rect 23014 24188 23020 24200
rect 22879 24160 23020 24188
rect 22879 24157 22891 24160
rect 22833 24151 22891 24157
rect 23014 24148 23020 24160
rect 23072 24148 23078 24200
rect 23658 24148 23664 24200
rect 23716 24188 23722 24200
rect 25317 24191 25375 24197
rect 25317 24188 25329 24191
rect 23716 24160 25329 24188
rect 23716 24148 23722 24160
rect 25317 24157 25329 24160
rect 25363 24157 25375 24191
rect 25317 24151 25375 24157
rect 25406 24148 25412 24200
rect 25464 24148 25470 24200
rect 27816 24197 27844 24228
rect 27985 24225 27997 24259
rect 28031 24256 28043 24259
rect 28184 24256 28212 24296
rect 29825 24327 29883 24333
rect 29825 24293 29837 24327
rect 29871 24324 29883 24327
rect 29914 24324 29920 24336
rect 29871 24296 29920 24324
rect 29871 24293 29883 24296
rect 29825 24287 29883 24293
rect 29914 24284 29920 24296
rect 29972 24284 29978 24336
rect 31481 24327 31539 24333
rect 31481 24293 31493 24327
rect 31527 24324 31539 24327
rect 31527 24296 31754 24324
rect 31527 24293 31539 24296
rect 31481 24287 31539 24293
rect 28031 24228 28212 24256
rect 28031 24225 28043 24228
rect 27985 24219 28043 24225
rect 28258 24216 28264 24268
rect 28316 24216 28322 24268
rect 29362 24256 29368 24268
rect 29012 24228 29368 24256
rect 27801 24191 27859 24197
rect 27801 24157 27813 24191
rect 27847 24157 27859 24191
rect 27801 24151 27859 24157
rect 28169 24191 28227 24197
rect 28169 24157 28181 24191
rect 28215 24157 28227 24191
rect 28169 24151 28227 24157
rect 14332 24092 21588 24120
rect 21637 24123 21695 24129
rect 14332 24080 14338 24092
rect 21637 24089 21649 24123
rect 21683 24089 21695 24123
rect 21637 24083 21695 24089
rect 12802 24052 12808 24064
rect 11992 24024 12808 24052
rect 12802 24012 12808 24024
rect 12860 24052 12866 24064
rect 13722 24052 13728 24064
rect 12860 24024 13728 24052
rect 12860 24012 12866 24024
rect 13722 24012 13728 24024
rect 13780 24052 13786 24064
rect 18874 24052 18880 24064
rect 13780 24024 18880 24052
rect 13780 24012 13786 24024
rect 18874 24012 18880 24024
rect 18932 24012 18938 24064
rect 19518 24012 19524 24064
rect 19576 24052 19582 24064
rect 20990 24052 20996 24064
rect 19576 24024 20996 24052
rect 19576 24012 19582 24024
rect 20990 24012 20996 24024
rect 21048 24012 21054 24064
rect 21266 24012 21272 24064
rect 21324 24012 21330 24064
rect 21652 24052 21680 24083
rect 23566 24080 23572 24132
rect 23624 24080 23630 24132
rect 23750 24080 23756 24132
rect 23808 24080 23814 24132
rect 24670 24080 24676 24132
rect 24728 24120 24734 24132
rect 28077 24123 28135 24129
rect 28077 24120 28089 24123
rect 24728 24092 28089 24120
rect 24728 24080 24734 24092
rect 28077 24089 28089 24092
rect 28123 24089 28135 24123
rect 28077 24083 28135 24089
rect 28184 24120 28212 24151
rect 28810 24148 28816 24200
rect 28868 24148 28874 24200
rect 29012 24197 29040 24228
rect 29362 24216 29368 24228
rect 29420 24216 29426 24268
rect 31726 24256 31754 24296
rect 32122 24256 32128 24268
rect 31726 24228 32128 24256
rect 32122 24216 32128 24228
rect 32180 24216 32186 24268
rect 28997 24191 29055 24197
rect 28997 24157 29009 24191
rect 29043 24157 29055 24191
rect 28997 24151 29055 24157
rect 29178 24148 29184 24200
rect 29236 24148 29242 24200
rect 29638 24148 29644 24200
rect 29696 24188 29702 24200
rect 30009 24191 30067 24197
rect 30009 24188 30021 24191
rect 29696 24160 30021 24188
rect 29696 24148 29702 24160
rect 30009 24157 30021 24160
rect 30055 24157 30067 24191
rect 30009 24151 30067 24157
rect 30101 24191 30159 24197
rect 30101 24157 30113 24191
rect 30147 24188 30159 24191
rect 30650 24188 30656 24200
rect 30147 24160 30656 24188
rect 30147 24157 30159 24160
rect 30101 24151 30159 24157
rect 30650 24148 30656 24160
rect 30708 24188 30714 24200
rect 30926 24188 30932 24200
rect 30708 24160 30932 24188
rect 30708 24148 30714 24160
rect 30926 24148 30932 24160
rect 30984 24148 30990 24200
rect 29089 24123 29147 24129
rect 28184 24092 29040 24120
rect 21910 24052 21916 24064
rect 21652 24024 21916 24052
rect 21910 24012 21916 24024
rect 21968 24012 21974 24064
rect 23017 24055 23075 24061
rect 23017 24021 23029 24055
rect 23063 24052 23075 24055
rect 23106 24052 23112 24064
rect 23063 24024 23112 24052
rect 23063 24021 23075 24024
rect 23017 24015 23075 24021
rect 23106 24012 23112 24024
rect 23164 24012 23170 24064
rect 25130 24012 25136 24064
rect 25188 24052 25194 24064
rect 25682 24052 25688 24064
rect 25188 24024 25688 24052
rect 25188 24012 25194 24024
rect 25682 24012 25688 24024
rect 25740 24012 25746 24064
rect 27617 24055 27675 24061
rect 27617 24021 27629 24055
rect 27663 24052 27675 24055
rect 27706 24052 27712 24064
rect 27663 24024 27712 24052
rect 27663 24021 27675 24024
rect 27617 24015 27675 24021
rect 27706 24012 27712 24024
rect 27764 24012 27770 24064
rect 27798 24012 27804 24064
rect 27856 24052 27862 24064
rect 28184 24052 28212 24092
rect 27856 24024 28212 24052
rect 27856 24012 27862 24024
rect 28534 24012 28540 24064
rect 28592 24012 28598 24064
rect 29012 24052 29040 24092
rect 29089 24089 29101 24123
rect 29135 24120 29147 24123
rect 29656 24120 29684 24148
rect 29135 24092 29684 24120
rect 30368 24123 30426 24129
rect 29135 24089 29147 24092
rect 29089 24083 29147 24089
rect 30368 24089 30380 24123
rect 30414 24120 30426 24123
rect 30466 24120 30472 24132
rect 30414 24092 30472 24120
rect 30414 24089 30426 24092
rect 30368 24083 30426 24089
rect 30466 24080 30472 24092
rect 30524 24080 30530 24132
rect 29178 24052 29184 24064
rect 29012 24024 29184 24052
rect 29178 24012 29184 24024
rect 29236 24012 29242 24064
rect 29362 24012 29368 24064
rect 29420 24012 29426 24064
rect 30282 24012 30288 24064
rect 30340 24052 30346 24064
rect 31573 24055 31631 24061
rect 31573 24052 31585 24055
rect 30340 24024 31585 24052
rect 30340 24012 30346 24024
rect 31573 24021 31585 24024
rect 31619 24021 31631 24055
rect 31573 24015 31631 24021
rect 1104 23962 32844 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 32844 23962
rect 1104 23888 32844 23910
rect 2406 23808 2412 23860
rect 2464 23848 2470 23860
rect 2958 23848 2964 23860
rect 2464 23820 2964 23848
rect 2464 23808 2470 23820
rect 2958 23808 2964 23820
rect 3016 23808 3022 23860
rect 3050 23808 3056 23860
rect 3108 23808 3114 23860
rect 3881 23851 3939 23857
rect 3252 23820 3740 23848
rect 1854 23740 1860 23792
rect 1912 23780 1918 23792
rect 3252 23780 3280 23820
rect 1912 23752 3280 23780
rect 1912 23740 1918 23752
rect 3326 23740 3332 23792
rect 3384 23780 3390 23792
rect 3421 23783 3479 23789
rect 3421 23780 3433 23783
rect 3384 23752 3433 23780
rect 3384 23740 3390 23752
rect 3421 23749 3433 23752
rect 3467 23749 3479 23783
rect 3712 23780 3740 23820
rect 3881 23817 3893 23851
rect 3927 23848 3939 23851
rect 3970 23848 3976 23860
rect 3927 23820 3976 23848
rect 3927 23817 3939 23820
rect 3881 23811 3939 23817
rect 3970 23808 3976 23820
rect 4028 23808 4034 23860
rect 4157 23851 4215 23857
rect 4157 23817 4169 23851
rect 4203 23848 4215 23851
rect 5442 23848 5448 23860
rect 4203 23820 5448 23848
rect 4203 23817 4215 23820
rect 4157 23811 4215 23817
rect 5442 23808 5448 23820
rect 5500 23808 5506 23860
rect 5902 23808 5908 23860
rect 5960 23848 5966 23860
rect 5997 23851 6055 23857
rect 5997 23848 6009 23851
rect 5960 23820 6009 23848
rect 5960 23808 5966 23820
rect 5997 23817 6009 23820
rect 6043 23817 6055 23851
rect 5997 23811 6055 23817
rect 10686 23808 10692 23860
rect 10744 23848 10750 23860
rect 10965 23851 11023 23857
rect 10744 23820 10824 23848
rect 10744 23808 10750 23820
rect 4338 23780 4344 23792
rect 3712 23752 4344 23780
rect 3421 23743 3479 23749
rect 4338 23740 4344 23752
rect 4396 23740 4402 23792
rect 4614 23740 4620 23792
rect 4672 23740 4678 23792
rect 4706 23740 4712 23792
rect 4764 23780 4770 23792
rect 4764 23752 6224 23780
rect 4764 23740 4770 23752
rect 2222 23672 2228 23724
rect 2280 23712 2286 23724
rect 2685 23715 2743 23721
rect 2685 23712 2697 23715
rect 2280 23684 2697 23712
rect 2280 23672 2286 23684
rect 2685 23681 2697 23684
rect 2731 23681 2743 23715
rect 2685 23675 2743 23681
rect 2777 23715 2835 23721
rect 2777 23681 2789 23715
rect 2823 23681 2835 23715
rect 2777 23675 2835 23681
rect 934 23604 940 23656
rect 992 23644 998 23656
rect 1302 23644 1308 23656
rect 992 23616 1308 23644
rect 992 23604 998 23616
rect 1302 23604 1308 23616
rect 1360 23604 1366 23656
rect 2406 23604 2412 23656
rect 2464 23644 2470 23656
rect 2792 23644 2820 23675
rect 2866 23672 2872 23724
rect 2924 23712 2930 23724
rect 3237 23715 3295 23721
rect 3237 23712 3249 23715
rect 2924 23684 3249 23712
rect 2924 23672 2930 23684
rect 3237 23681 3249 23684
rect 3283 23681 3295 23715
rect 3237 23675 3295 23681
rect 4062 23672 4068 23724
rect 4120 23712 4126 23724
rect 4433 23715 4491 23721
rect 4433 23712 4445 23715
rect 4120 23684 4445 23712
rect 4120 23672 4126 23684
rect 4433 23681 4445 23684
rect 4479 23681 4491 23715
rect 4433 23675 4491 23681
rect 4525 23715 4583 23721
rect 4525 23681 4537 23715
rect 4571 23712 4583 23715
rect 4632 23712 4660 23740
rect 4571 23684 4660 23712
rect 5077 23715 5135 23721
rect 4571 23681 4583 23684
rect 4525 23675 4583 23681
rect 5077 23681 5089 23715
rect 5123 23681 5135 23715
rect 5077 23675 5135 23681
rect 2464 23616 2820 23644
rect 3973 23647 4031 23653
rect 2464 23604 2470 23616
rect 3973 23613 3985 23647
rect 4019 23613 4031 23647
rect 3973 23607 4031 23613
rect 2314 23536 2320 23588
rect 2372 23576 2378 23588
rect 2501 23579 2559 23585
rect 2501 23576 2513 23579
rect 2372 23548 2513 23576
rect 2372 23536 2378 23548
rect 2501 23545 2513 23548
rect 2547 23576 2559 23579
rect 2774 23576 2780 23588
rect 2547 23548 2780 23576
rect 2547 23545 2559 23548
rect 2501 23539 2559 23545
rect 2774 23536 2780 23548
rect 2832 23536 2838 23588
rect 3418 23536 3424 23588
rect 3476 23536 3482 23588
rect 3988 23576 4016 23607
rect 4338 23604 4344 23656
rect 4396 23604 4402 23656
rect 4617 23647 4675 23653
rect 4617 23613 4629 23647
rect 4663 23644 4675 23647
rect 4798 23644 4804 23656
rect 4663 23616 4804 23644
rect 4663 23613 4675 23616
rect 4617 23607 4675 23613
rect 4154 23576 4160 23588
rect 3988 23548 4160 23576
rect 4154 23536 4160 23548
rect 4212 23576 4218 23588
rect 4632 23576 4660 23607
rect 4798 23604 4804 23616
rect 4856 23604 4862 23656
rect 5092 23644 5120 23675
rect 5166 23672 5172 23724
rect 5224 23672 5230 23724
rect 5350 23672 5356 23724
rect 5408 23712 5414 23724
rect 5629 23715 5687 23721
rect 5629 23712 5641 23715
rect 5408 23684 5641 23712
rect 5408 23672 5414 23684
rect 5629 23681 5641 23684
rect 5675 23681 5687 23715
rect 5629 23675 5687 23681
rect 5902 23672 5908 23724
rect 5960 23672 5966 23724
rect 6196 23721 6224 23752
rect 10134 23740 10140 23792
rect 10192 23780 10198 23792
rect 10597 23783 10655 23789
rect 10597 23780 10609 23783
rect 10192 23752 10609 23780
rect 10192 23740 10198 23752
rect 10597 23749 10609 23752
rect 10643 23749 10655 23783
rect 10597 23743 10655 23749
rect 6181 23715 6239 23721
rect 6181 23681 6193 23715
rect 6227 23681 6239 23715
rect 6181 23675 6239 23681
rect 6362 23672 6368 23724
rect 6420 23712 6426 23724
rect 6549 23715 6607 23721
rect 6549 23712 6561 23715
rect 6420 23684 6561 23712
rect 6420 23672 6426 23684
rect 6549 23681 6561 23684
rect 6595 23681 6607 23715
rect 6549 23675 6607 23681
rect 6914 23672 6920 23724
rect 6972 23712 6978 23724
rect 7558 23712 7564 23724
rect 6972 23684 7564 23712
rect 6972 23672 6978 23684
rect 7558 23672 7564 23684
rect 7616 23672 7622 23724
rect 8478 23672 8484 23724
rect 8536 23712 8542 23724
rect 8757 23715 8815 23721
rect 8757 23712 8769 23715
rect 8536 23684 8769 23712
rect 8536 23672 8542 23684
rect 8757 23681 8769 23684
rect 8803 23681 8815 23715
rect 8757 23675 8815 23681
rect 8846 23672 8852 23724
rect 8904 23712 8910 23724
rect 8941 23715 8999 23721
rect 8941 23712 8953 23715
rect 8904 23684 8953 23712
rect 8904 23672 8910 23684
rect 8941 23681 8953 23684
rect 8987 23681 8999 23715
rect 8941 23675 8999 23681
rect 9030 23672 9036 23724
rect 9088 23672 9094 23724
rect 9125 23715 9183 23721
rect 9125 23681 9137 23715
rect 9171 23712 9183 23715
rect 9398 23712 9404 23724
rect 9171 23684 9404 23712
rect 9171 23681 9183 23684
rect 9125 23675 9183 23681
rect 9398 23672 9404 23684
rect 9456 23672 9462 23724
rect 10413 23715 10471 23721
rect 10413 23681 10425 23715
rect 10459 23712 10471 23715
rect 10502 23712 10508 23724
rect 10459 23684 10508 23712
rect 10459 23681 10471 23684
rect 10413 23675 10471 23681
rect 10502 23672 10508 23684
rect 10560 23672 10566 23724
rect 10796 23721 10824 23820
rect 10965 23817 10977 23851
rect 11011 23817 11023 23851
rect 10965 23811 11023 23817
rect 10980 23724 11008 23811
rect 11698 23808 11704 23860
rect 11756 23848 11762 23860
rect 11756 23820 12020 23848
rect 11756 23808 11762 23820
rect 11422 23740 11428 23792
rect 11480 23780 11486 23792
rect 11793 23783 11851 23789
rect 11793 23780 11805 23783
rect 11480 23752 11805 23780
rect 11480 23740 11486 23752
rect 11793 23749 11805 23752
rect 11839 23749 11851 23783
rect 11992 23780 12020 23820
rect 12066 23808 12072 23860
rect 12124 23808 12130 23860
rect 12345 23851 12403 23857
rect 12345 23817 12357 23851
rect 12391 23817 12403 23851
rect 12345 23811 12403 23817
rect 12360 23780 12388 23811
rect 12986 23808 12992 23860
rect 13044 23848 13050 23860
rect 14826 23848 14832 23860
rect 13044 23820 14832 23848
rect 13044 23808 13050 23820
rect 14826 23808 14832 23820
rect 14884 23848 14890 23860
rect 14884 23820 18092 23848
rect 14884 23808 14890 23820
rect 11992 23752 12388 23780
rect 11793 23743 11851 23749
rect 12434 23740 12440 23792
rect 12492 23780 12498 23792
rect 15197 23783 15255 23789
rect 15197 23780 15209 23783
rect 12492 23752 15209 23780
rect 12492 23740 12498 23752
rect 15197 23749 15209 23752
rect 15243 23749 15255 23783
rect 15197 23743 15255 23749
rect 16482 23740 16488 23792
rect 16540 23780 16546 23792
rect 16540 23752 16896 23780
rect 16540 23740 16546 23752
rect 10689 23715 10747 23721
rect 10689 23681 10701 23715
rect 10735 23681 10747 23715
rect 10689 23675 10747 23681
rect 10781 23715 10839 23721
rect 10781 23681 10793 23715
rect 10827 23681 10839 23715
rect 10781 23675 10839 23681
rect 5258 23644 5264 23656
rect 5092 23616 5264 23644
rect 5258 23604 5264 23616
rect 5316 23604 5322 23656
rect 9766 23644 9772 23656
rect 5484 23616 9772 23644
rect 5484 23576 5512 23616
rect 9766 23604 9772 23616
rect 9824 23604 9830 23656
rect 9950 23604 9956 23656
rect 10008 23644 10014 23656
rect 10318 23644 10324 23656
rect 10008 23616 10324 23644
rect 10008 23604 10014 23616
rect 10318 23604 10324 23616
rect 10376 23604 10382 23656
rect 10704 23644 10732 23675
rect 10962 23672 10968 23724
rect 11020 23672 11026 23724
rect 11440 23644 11468 23740
rect 16868 23724 16896 23752
rect 17678 23740 17684 23792
rect 17736 23780 17742 23792
rect 17957 23783 18015 23789
rect 17957 23780 17969 23783
rect 17736 23752 17969 23780
rect 17736 23740 17742 23752
rect 17957 23749 17969 23752
rect 18003 23749 18015 23783
rect 18064 23780 18092 23820
rect 18138 23808 18144 23860
rect 18196 23848 18202 23860
rect 20714 23848 20720 23860
rect 18196 23820 20720 23848
rect 18196 23808 18202 23820
rect 20714 23808 20720 23820
rect 20772 23808 20778 23860
rect 24581 23851 24639 23857
rect 24581 23848 24593 23851
rect 24320 23820 24593 23848
rect 21726 23780 21732 23792
rect 18064 23752 21732 23780
rect 17957 23743 18015 23749
rect 21726 23740 21732 23752
rect 21784 23740 21790 23792
rect 24320 23789 24348 23820
rect 24581 23817 24593 23820
rect 24627 23848 24639 23851
rect 25222 23848 25228 23860
rect 24627 23820 25228 23848
rect 24627 23817 24639 23820
rect 24581 23811 24639 23817
rect 25222 23808 25228 23820
rect 25280 23808 25286 23860
rect 27798 23848 27804 23860
rect 26160 23820 27804 23848
rect 24305 23783 24363 23789
rect 22112 23752 24072 23780
rect 11517 23715 11575 23721
rect 11517 23681 11529 23715
rect 11563 23712 11575 23715
rect 11606 23712 11612 23724
rect 11563 23684 11612 23712
rect 11563 23681 11575 23684
rect 11517 23675 11575 23681
rect 11606 23672 11612 23684
rect 11664 23672 11670 23724
rect 11698 23672 11704 23724
rect 11756 23672 11762 23724
rect 11882 23672 11888 23724
rect 11940 23672 11946 23724
rect 11974 23672 11980 23724
rect 12032 23712 12038 23724
rect 12161 23715 12219 23721
rect 12161 23712 12173 23715
rect 12032 23684 12173 23712
rect 12032 23672 12038 23684
rect 12161 23681 12173 23684
rect 12207 23681 12219 23715
rect 12161 23675 12219 23681
rect 12529 23715 12587 23721
rect 12529 23681 12541 23715
rect 12575 23712 12587 23715
rect 12618 23712 12624 23724
rect 12575 23684 12624 23712
rect 12575 23681 12587 23684
rect 12529 23675 12587 23681
rect 12618 23672 12624 23684
rect 12676 23672 12682 23724
rect 12713 23715 12771 23721
rect 12713 23681 12725 23715
rect 12759 23712 12771 23715
rect 12986 23712 12992 23724
rect 12759 23684 12992 23712
rect 12759 23681 12771 23684
rect 12713 23675 12771 23681
rect 12986 23672 12992 23684
rect 13044 23672 13050 23724
rect 13170 23672 13176 23724
rect 13228 23672 13234 23724
rect 13722 23672 13728 23724
rect 13780 23712 13786 23724
rect 13817 23715 13875 23721
rect 13817 23712 13829 23715
rect 13780 23684 13829 23712
rect 13780 23672 13786 23684
rect 13817 23681 13829 23684
rect 13863 23681 13875 23715
rect 13817 23675 13875 23681
rect 14001 23715 14059 23721
rect 14001 23681 14013 23715
rect 14047 23712 14059 23715
rect 14182 23712 14188 23724
rect 14047 23684 14188 23712
rect 14047 23681 14059 23684
rect 14001 23675 14059 23681
rect 14182 23672 14188 23684
rect 14240 23672 14246 23724
rect 14274 23672 14280 23724
rect 14332 23672 14338 23724
rect 15013 23715 15071 23721
rect 15013 23681 15025 23715
rect 15059 23712 15071 23715
rect 15102 23712 15108 23724
rect 15059 23684 15108 23712
rect 15059 23681 15071 23684
rect 15013 23675 15071 23681
rect 15102 23672 15108 23684
rect 15160 23672 15166 23724
rect 15654 23672 15660 23724
rect 15712 23672 15718 23724
rect 16114 23672 16120 23724
rect 16172 23712 16178 23724
rect 16669 23715 16727 23721
rect 16669 23712 16681 23715
rect 16172 23684 16681 23712
rect 16172 23672 16178 23684
rect 16669 23681 16681 23684
rect 16715 23681 16727 23715
rect 16669 23675 16727 23681
rect 16850 23672 16856 23724
rect 16908 23672 16914 23724
rect 18233 23715 18291 23721
rect 18233 23681 18245 23715
rect 18279 23712 18291 23715
rect 18966 23712 18972 23724
rect 18279 23684 18972 23712
rect 18279 23681 18291 23684
rect 18233 23675 18291 23681
rect 18966 23672 18972 23684
rect 19024 23672 19030 23724
rect 19058 23672 19064 23724
rect 19116 23712 19122 23724
rect 19705 23715 19763 23721
rect 19705 23712 19717 23715
rect 19116 23684 19717 23712
rect 19116 23672 19122 23684
rect 19705 23681 19717 23684
rect 19751 23681 19763 23715
rect 22005 23715 22063 23721
rect 22005 23712 22017 23715
rect 19705 23675 19763 23681
rect 20640 23684 22017 23712
rect 14292 23644 14320 23672
rect 10704 23616 11468 23644
rect 11624 23616 11836 23644
rect 4212 23548 4660 23576
rect 4816 23548 5512 23576
rect 4212 23536 4218 23548
rect 4816 23517 4844 23548
rect 6362 23536 6368 23588
rect 6420 23536 6426 23588
rect 7466 23536 7472 23588
rect 7524 23576 7530 23588
rect 11624 23576 11652 23616
rect 7524 23548 11652 23576
rect 7524 23536 7530 23548
rect 4801 23511 4859 23517
rect 4801 23477 4813 23511
rect 4847 23477 4859 23511
rect 4801 23471 4859 23477
rect 4890 23468 4896 23520
rect 4948 23508 4954 23520
rect 5074 23508 5080 23520
rect 4948 23480 5080 23508
rect 4948 23468 4954 23480
rect 5074 23468 5080 23480
rect 5132 23468 5138 23520
rect 5350 23468 5356 23520
rect 5408 23468 5414 23520
rect 5442 23468 5448 23520
rect 5500 23468 5506 23520
rect 5718 23468 5724 23520
rect 5776 23468 5782 23520
rect 6730 23468 6736 23520
rect 6788 23508 6794 23520
rect 7558 23508 7564 23520
rect 6788 23480 7564 23508
rect 6788 23468 6794 23480
rect 7558 23468 7564 23480
rect 7616 23468 7622 23520
rect 8294 23468 8300 23520
rect 8352 23508 8358 23520
rect 8754 23508 8760 23520
rect 8352 23480 8760 23508
rect 8352 23468 8358 23480
rect 8754 23468 8760 23480
rect 8812 23468 8818 23520
rect 9030 23468 9036 23520
rect 9088 23508 9094 23520
rect 9309 23511 9367 23517
rect 9309 23508 9321 23511
rect 9088 23480 9321 23508
rect 9088 23468 9094 23480
rect 9309 23477 9321 23480
rect 9355 23477 9367 23511
rect 9309 23471 9367 23477
rect 9766 23468 9772 23520
rect 9824 23508 9830 23520
rect 11698 23508 11704 23520
rect 9824 23480 11704 23508
rect 9824 23468 9830 23480
rect 11698 23468 11704 23480
rect 11756 23468 11762 23520
rect 11808 23508 11836 23616
rect 12820 23616 14320 23644
rect 17037 23647 17095 23653
rect 12820 23508 12848 23616
rect 17037 23613 17049 23647
rect 17083 23644 17095 23647
rect 18141 23647 18199 23653
rect 18141 23644 18153 23647
rect 17083 23616 18153 23644
rect 17083 23613 17095 23616
rect 17037 23607 17095 23613
rect 18141 23613 18153 23616
rect 18187 23644 18199 23647
rect 18598 23644 18604 23656
rect 18187 23616 18604 23644
rect 18187 23613 18199 23616
rect 18141 23607 18199 23613
rect 18598 23604 18604 23616
rect 18656 23604 18662 23656
rect 18690 23604 18696 23656
rect 18748 23644 18754 23656
rect 20640 23644 20668 23684
rect 22005 23681 22017 23684
rect 22051 23681 22063 23715
rect 22005 23675 22063 23681
rect 22112 23644 22140 23752
rect 22278 23672 22284 23724
rect 22336 23712 22342 23724
rect 22925 23715 22983 23721
rect 22925 23712 22937 23715
rect 22336 23684 22937 23712
rect 22336 23672 22342 23684
rect 22925 23681 22937 23684
rect 22971 23681 22983 23715
rect 23934 23712 23940 23724
rect 22925 23675 22983 23681
rect 23032 23684 23940 23712
rect 18748 23616 20668 23644
rect 21652 23616 22140 23644
rect 18748 23604 18754 23616
rect 13633 23579 13691 23585
rect 13633 23545 13645 23579
rect 13679 23576 13691 23579
rect 14458 23576 14464 23588
rect 13679 23548 14464 23576
rect 13679 23545 13691 23548
rect 13633 23539 13691 23545
rect 14458 23536 14464 23548
rect 14516 23536 14522 23588
rect 15102 23536 15108 23588
rect 15160 23576 15166 23588
rect 15473 23579 15531 23585
rect 15473 23576 15485 23579
rect 15160 23548 15485 23576
rect 15160 23536 15166 23548
rect 15473 23545 15485 23548
rect 15519 23545 15531 23579
rect 15473 23539 15531 23545
rect 15562 23536 15568 23588
rect 15620 23576 15626 23588
rect 18046 23576 18052 23588
rect 15620 23548 18052 23576
rect 15620 23536 15626 23548
rect 18046 23536 18052 23548
rect 18104 23536 18110 23588
rect 18782 23576 18788 23588
rect 18248 23548 18788 23576
rect 11808 23480 12848 23508
rect 12897 23511 12955 23517
rect 12897 23477 12909 23511
rect 12943 23508 12955 23511
rect 13722 23508 13728 23520
rect 12943 23480 13728 23508
rect 12943 23477 12955 23480
rect 12897 23471 12955 23477
rect 13722 23468 13728 23480
rect 13780 23468 13786 23520
rect 14093 23511 14151 23517
rect 14093 23477 14105 23511
rect 14139 23508 14151 23511
rect 14182 23508 14188 23520
rect 14139 23480 14188 23508
rect 14139 23477 14151 23480
rect 14093 23471 14151 23477
rect 14182 23468 14188 23480
rect 14240 23468 14246 23520
rect 15286 23468 15292 23520
rect 15344 23508 15350 23520
rect 15381 23511 15439 23517
rect 15381 23508 15393 23511
rect 15344 23480 15393 23508
rect 15344 23468 15350 23480
rect 15381 23477 15393 23480
rect 15427 23477 15439 23511
rect 15381 23471 15439 23477
rect 15746 23468 15752 23520
rect 15804 23508 15810 23520
rect 17494 23508 17500 23520
rect 15804 23480 17500 23508
rect 15804 23468 15810 23480
rect 17494 23468 17500 23480
rect 17552 23468 17558 23520
rect 18248 23517 18276 23548
rect 18782 23536 18788 23548
rect 18840 23536 18846 23588
rect 18874 23536 18880 23588
rect 18932 23576 18938 23588
rect 21652 23576 21680 23616
rect 23032 23576 23060 23684
rect 23934 23672 23940 23684
rect 23992 23672 23998 23724
rect 24044 23721 24072 23752
rect 24305 23749 24317 23783
rect 24351 23749 24363 23783
rect 24305 23743 24363 23749
rect 24854 23740 24860 23792
rect 24912 23780 24918 23792
rect 26160 23780 26188 23820
rect 27798 23808 27804 23820
rect 27856 23808 27862 23860
rect 28074 23808 28080 23860
rect 28132 23848 28138 23860
rect 28350 23848 28356 23860
rect 28132 23820 28356 23848
rect 28132 23808 28138 23820
rect 28350 23808 28356 23820
rect 28408 23808 28414 23860
rect 30466 23808 30472 23860
rect 30524 23808 30530 23860
rect 31846 23808 31852 23860
rect 31904 23848 31910 23860
rect 31941 23851 31999 23857
rect 31941 23848 31953 23851
rect 31904 23820 31953 23848
rect 31904 23808 31910 23820
rect 31941 23817 31953 23820
rect 31987 23817 31999 23851
rect 31941 23811 31999 23817
rect 24912 23752 26188 23780
rect 24912 23740 24918 23752
rect 26234 23740 26240 23792
rect 26292 23780 26298 23792
rect 28810 23780 28816 23792
rect 26292 23752 28816 23780
rect 26292 23740 26298 23752
rect 28810 23740 28816 23752
rect 28868 23740 28874 23792
rect 29362 23740 29368 23792
rect 29420 23780 29426 23792
rect 30806 23783 30864 23789
rect 30806 23780 30818 23783
rect 29420 23752 30818 23780
rect 29420 23740 29426 23752
rect 30806 23749 30818 23752
rect 30852 23749 30864 23783
rect 30806 23743 30864 23749
rect 24029 23715 24087 23721
rect 24029 23681 24041 23715
rect 24075 23681 24087 23715
rect 24029 23675 24087 23681
rect 24397 23715 24455 23721
rect 24397 23681 24409 23715
rect 24443 23681 24455 23715
rect 24397 23675 24455 23681
rect 23290 23644 23296 23656
rect 23124 23616 23296 23644
rect 23124 23585 23152 23616
rect 23290 23604 23296 23616
rect 23348 23644 23354 23656
rect 24121 23647 24179 23653
rect 24121 23644 24133 23647
rect 23348 23616 24133 23644
rect 23348 23604 23354 23616
rect 24121 23613 24133 23616
rect 24167 23613 24179 23647
rect 24121 23607 24179 23613
rect 18932 23548 21680 23576
rect 22066 23548 23060 23576
rect 23109 23579 23167 23585
rect 18932 23536 18938 23548
rect 18233 23511 18291 23517
rect 18233 23477 18245 23511
rect 18279 23477 18291 23511
rect 18233 23471 18291 23477
rect 18417 23511 18475 23517
rect 18417 23477 18429 23511
rect 18463 23508 18475 23511
rect 18506 23508 18512 23520
rect 18463 23480 18512 23508
rect 18463 23477 18475 23480
rect 18417 23471 18475 23477
rect 18506 23468 18512 23480
rect 18564 23468 18570 23520
rect 19334 23468 19340 23520
rect 19392 23508 19398 23520
rect 19889 23511 19947 23517
rect 19889 23508 19901 23511
rect 19392 23480 19901 23508
rect 19392 23468 19398 23480
rect 19889 23477 19901 23480
rect 19935 23508 19947 23511
rect 19978 23508 19984 23520
rect 19935 23480 19984 23508
rect 19935 23477 19947 23480
rect 19889 23471 19947 23477
rect 19978 23468 19984 23480
rect 20036 23468 20042 23520
rect 20714 23468 20720 23520
rect 20772 23508 20778 23520
rect 22066 23508 22094 23548
rect 23109 23545 23121 23579
rect 23155 23545 23167 23579
rect 23109 23539 23167 23545
rect 23382 23536 23388 23588
rect 23440 23576 23446 23588
rect 24412 23576 24440 23675
rect 26050 23672 26056 23724
rect 26108 23672 26114 23724
rect 29917 23715 29975 23721
rect 29917 23681 29929 23715
rect 29963 23712 29975 23715
rect 30101 23715 30159 23721
rect 29963 23684 30052 23712
rect 29963 23681 29975 23684
rect 29917 23675 29975 23681
rect 25958 23604 25964 23656
rect 26016 23644 26022 23656
rect 26145 23647 26203 23653
rect 26145 23644 26157 23647
rect 26016 23616 26157 23644
rect 26016 23604 26022 23616
rect 26145 23613 26157 23616
rect 26191 23613 26203 23647
rect 26145 23607 26203 23613
rect 23440 23548 24440 23576
rect 23440 23536 23446 23548
rect 20772 23480 22094 23508
rect 20772 23468 20778 23480
rect 22186 23468 22192 23520
rect 22244 23468 22250 23520
rect 23842 23468 23848 23520
rect 23900 23468 23906 23520
rect 24026 23468 24032 23520
rect 24084 23468 24090 23520
rect 25774 23468 25780 23520
rect 25832 23508 25838 23520
rect 26053 23511 26111 23517
rect 26053 23508 26065 23511
rect 25832 23480 26065 23508
rect 25832 23468 25838 23480
rect 26053 23477 26065 23480
rect 26099 23477 26111 23511
rect 26053 23471 26111 23477
rect 26421 23511 26479 23517
rect 26421 23477 26433 23511
rect 26467 23508 26479 23511
rect 27798 23508 27804 23520
rect 26467 23480 27804 23508
rect 26467 23477 26479 23480
rect 26421 23471 26479 23477
rect 27798 23468 27804 23480
rect 27856 23468 27862 23520
rect 27890 23468 27896 23520
rect 27948 23508 27954 23520
rect 28718 23508 28724 23520
rect 27948 23480 28724 23508
rect 27948 23468 27954 23480
rect 28718 23468 28724 23480
rect 28776 23468 28782 23520
rect 28994 23468 29000 23520
rect 29052 23508 29058 23520
rect 29454 23508 29460 23520
rect 29052 23480 29460 23508
rect 29052 23468 29058 23480
rect 29454 23468 29460 23480
rect 29512 23468 29518 23520
rect 30024 23508 30052 23684
rect 30101 23681 30113 23715
rect 30147 23681 30159 23715
rect 30101 23675 30159 23681
rect 30116 23576 30144 23675
rect 30190 23672 30196 23724
rect 30248 23672 30254 23724
rect 30282 23672 30288 23724
rect 30340 23672 30346 23724
rect 30561 23715 30619 23721
rect 30561 23681 30573 23715
rect 30607 23712 30619 23715
rect 30650 23712 30656 23724
rect 30607 23684 30656 23712
rect 30607 23681 30619 23684
rect 30561 23675 30619 23681
rect 30650 23672 30656 23684
rect 30708 23672 30714 23724
rect 32217 23715 32275 23721
rect 32217 23681 32229 23715
rect 32263 23712 32275 23715
rect 32582 23712 32588 23724
rect 32263 23684 32588 23712
rect 32263 23681 32275 23684
rect 32217 23675 32275 23681
rect 32582 23672 32588 23684
rect 32640 23672 32646 23724
rect 30374 23576 30380 23588
rect 30116 23548 30380 23576
rect 30374 23536 30380 23548
rect 30432 23536 30438 23588
rect 30558 23508 30564 23520
rect 30024 23480 30564 23508
rect 30558 23468 30564 23480
rect 30616 23468 30622 23520
rect 32398 23468 32404 23520
rect 32456 23468 32462 23520
rect 1104 23418 32844 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 32844 23418
rect 1104 23344 32844 23366
rect 2038 23264 2044 23316
rect 2096 23304 2102 23316
rect 2133 23307 2191 23313
rect 2133 23304 2145 23307
rect 2096 23276 2145 23304
rect 2096 23264 2102 23276
rect 2133 23273 2145 23276
rect 2179 23273 2191 23307
rect 3786 23304 3792 23316
rect 2133 23267 2191 23273
rect 2746 23276 3792 23304
rect 2148 23168 2176 23267
rect 2593 23239 2651 23245
rect 2593 23205 2605 23239
rect 2639 23236 2651 23239
rect 2746 23236 2774 23276
rect 3786 23264 3792 23276
rect 3844 23304 3850 23316
rect 4341 23307 4399 23313
rect 3844 23276 4016 23304
rect 3844 23264 3850 23276
rect 2639 23208 2774 23236
rect 2869 23239 2927 23245
rect 2639 23205 2651 23208
rect 2593 23199 2651 23205
rect 2869 23205 2881 23239
rect 2915 23236 2927 23239
rect 3878 23236 3884 23248
rect 2915 23208 3884 23236
rect 2915 23205 2927 23208
rect 2869 23199 2927 23205
rect 3878 23196 3884 23208
rect 3936 23196 3942 23248
rect 2148 23140 2452 23168
rect 2314 23060 2320 23112
rect 2372 23060 2378 23112
rect 2424 23109 2452 23140
rect 2774 23128 2780 23180
rect 2832 23168 2838 23180
rect 3988 23168 4016 23276
rect 4341 23273 4353 23307
rect 4387 23304 4399 23307
rect 5166 23304 5172 23316
rect 4387 23276 5172 23304
rect 4387 23273 4399 23276
rect 4341 23267 4399 23273
rect 5166 23264 5172 23276
rect 5224 23264 5230 23316
rect 5902 23304 5908 23316
rect 5644 23276 5908 23304
rect 4430 23196 4436 23248
rect 4488 23236 4494 23248
rect 4890 23236 4896 23248
rect 4488 23208 4896 23236
rect 4488 23196 4494 23208
rect 4890 23196 4896 23208
rect 4948 23196 4954 23248
rect 5350 23236 5356 23248
rect 5276 23208 5356 23236
rect 4065 23171 4123 23177
rect 4065 23168 4077 23171
rect 2832 23140 3924 23168
rect 3988 23140 4077 23168
rect 2832 23128 2838 23140
rect 2409 23103 2467 23109
rect 2409 23069 2421 23103
rect 2455 23100 2467 23103
rect 2685 23103 2743 23109
rect 2685 23100 2697 23103
rect 2455 23072 2697 23100
rect 2455 23069 2467 23072
rect 2409 23063 2467 23069
rect 2685 23069 2697 23072
rect 2731 23069 2743 23103
rect 2685 23063 2743 23069
rect 2961 23103 3019 23109
rect 2961 23069 2973 23103
rect 3007 23100 3019 23103
rect 3142 23100 3148 23112
rect 3007 23072 3148 23100
rect 3007 23069 3019 23072
rect 2961 23063 3019 23069
rect 3142 23060 3148 23072
rect 3200 23060 3206 23112
rect 3896 23109 3924 23140
rect 4065 23137 4077 23140
rect 4111 23137 4123 23171
rect 4065 23131 4123 23137
rect 4522 23128 4528 23180
rect 4580 23168 4586 23180
rect 5276 23168 5304 23208
rect 5350 23196 5356 23208
rect 5408 23196 5414 23248
rect 4580 23140 5304 23168
rect 4580 23128 4586 23140
rect 3237 23103 3295 23109
rect 3237 23069 3249 23103
rect 3283 23069 3295 23103
rect 3237 23063 3295 23069
rect 3881 23103 3939 23109
rect 3881 23069 3893 23103
rect 3927 23069 3939 23103
rect 3881 23063 3939 23069
rect 2222 22992 2228 23044
rect 2280 23032 2286 23044
rect 3252 23032 3280 23063
rect 3970 23060 3976 23112
rect 4028 23060 4034 23112
rect 4157 23103 4215 23109
rect 4157 23069 4169 23103
rect 4203 23069 4215 23103
rect 4157 23063 4215 23069
rect 2280 23004 3280 23032
rect 2280 22992 2286 23004
rect 3786 22992 3792 23044
rect 3844 23032 3850 23044
rect 4172 23032 4200 23063
rect 4614 23060 4620 23112
rect 4672 23060 4678 23112
rect 4893 23103 4951 23109
rect 4893 23069 4905 23103
rect 4939 23100 4951 23103
rect 4982 23100 4988 23112
rect 4939 23072 4988 23100
rect 4939 23069 4951 23072
rect 4893 23063 4951 23069
rect 4982 23060 4988 23072
rect 5040 23060 5046 23112
rect 5077 23103 5135 23109
rect 5077 23069 5089 23103
rect 5123 23100 5135 23103
rect 5258 23100 5264 23112
rect 5123 23072 5264 23100
rect 5123 23069 5135 23072
rect 5077 23063 5135 23069
rect 5258 23060 5264 23072
rect 5316 23060 5322 23112
rect 5350 23060 5356 23112
rect 5408 23060 5414 23112
rect 5445 23103 5503 23109
rect 5445 23069 5457 23103
rect 5491 23100 5503 23103
rect 5644 23100 5672 23276
rect 5902 23264 5908 23276
rect 5960 23264 5966 23316
rect 5997 23307 6055 23313
rect 5997 23273 6009 23307
rect 6043 23304 6055 23307
rect 6730 23304 6736 23316
rect 6043 23276 6736 23304
rect 6043 23273 6055 23276
rect 5997 23267 6055 23273
rect 6730 23264 6736 23276
rect 6788 23264 6794 23316
rect 7101 23307 7159 23313
rect 7101 23273 7113 23307
rect 7147 23304 7159 23307
rect 7147 23276 7328 23304
rect 7147 23273 7159 23276
rect 7101 23267 7159 23273
rect 6914 23236 6920 23248
rect 5491 23072 5672 23100
rect 5736 23208 6920 23236
rect 5491 23069 5503 23072
rect 5445 23063 5503 23069
rect 3844 23004 4200 23032
rect 3844 22992 3850 23004
rect 4798 22992 4804 23044
rect 4856 23032 4862 23044
rect 5736 23041 5764 23208
rect 6914 23196 6920 23208
rect 6972 23236 6978 23248
rect 7190 23236 7196 23248
rect 6972 23208 7196 23236
rect 6972 23196 6978 23208
rect 7190 23196 7196 23208
rect 7248 23196 7254 23248
rect 7300 23236 7328 23276
rect 7558 23264 7564 23316
rect 7616 23304 7622 23316
rect 9674 23304 9680 23316
rect 7616 23276 9680 23304
rect 7616 23264 7622 23276
rect 9674 23264 9680 23276
rect 9732 23264 9738 23316
rect 11606 23264 11612 23316
rect 11664 23304 11670 23316
rect 13814 23304 13820 23316
rect 11664 23276 13820 23304
rect 11664 23264 11670 23276
rect 13814 23264 13820 23276
rect 13872 23264 13878 23316
rect 14093 23307 14151 23313
rect 14093 23273 14105 23307
rect 14139 23273 14151 23307
rect 14093 23267 14151 23273
rect 16209 23307 16267 23313
rect 16209 23273 16221 23307
rect 16255 23304 16267 23307
rect 16298 23304 16304 23316
rect 16255 23276 16304 23304
rect 16255 23273 16267 23276
rect 16209 23267 16267 23273
rect 10965 23239 11023 23245
rect 7300 23208 9812 23236
rect 7282 23128 7288 23180
rect 7340 23128 7346 23180
rect 7392 23140 7696 23168
rect 5813 23103 5871 23109
rect 5813 23069 5825 23103
rect 5859 23100 5871 23103
rect 6086 23100 6092 23112
rect 5859 23072 6092 23100
rect 5859 23069 5871 23072
rect 5813 23063 5871 23069
rect 5629 23035 5687 23041
rect 5629 23032 5641 23035
rect 4856 23004 5641 23032
rect 4856 22992 4862 23004
rect 5629 23001 5641 23004
rect 5675 23001 5687 23035
rect 5629 22995 5687 23001
rect 5721 23035 5779 23041
rect 5721 23001 5733 23035
rect 5767 23001 5779 23035
rect 5721 22995 5779 23001
rect 3142 22924 3148 22976
rect 3200 22924 3206 22976
rect 3234 22924 3240 22976
rect 3292 22964 3298 22976
rect 3421 22967 3479 22973
rect 3421 22964 3433 22967
rect 3292 22936 3433 22964
rect 3292 22924 3298 22936
rect 3421 22933 3433 22936
rect 3467 22933 3479 22967
rect 3421 22927 3479 22933
rect 4433 22967 4491 22973
rect 4433 22933 4445 22967
rect 4479 22964 4491 22967
rect 4890 22964 4896 22976
rect 4479 22936 4896 22964
rect 4479 22933 4491 22936
rect 4433 22927 4491 22933
rect 4890 22924 4896 22936
rect 4948 22924 4954 22976
rect 5169 22967 5227 22973
rect 5169 22933 5181 22967
rect 5215 22964 5227 22967
rect 5534 22964 5540 22976
rect 5215 22936 5540 22964
rect 5215 22933 5227 22936
rect 5169 22927 5227 22933
rect 5534 22924 5540 22936
rect 5592 22964 5598 22976
rect 5828 22964 5856 23063
rect 6086 23060 6092 23072
rect 6144 23060 6150 23112
rect 6178 23060 6184 23112
rect 6236 23100 6242 23112
rect 6273 23103 6331 23109
rect 6273 23100 6285 23103
rect 6236 23072 6285 23100
rect 6236 23060 6242 23072
rect 6273 23069 6285 23072
rect 6319 23069 6331 23103
rect 6273 23063 6331 23069
rect 6546 23060 6552 23112
rect 6604 23060 6610 23112
rect 6730 23060 6736 23112
rect 6788 23060 6794 23112
rect 6822 23060 6828 23112
rect 6880 23060 6886 23112
rect 6914 23060 6920 23112
rect 6972 23060 6978 23112
rect 7193 23103 7251 23109
rect 7193 23069 7205 23103
rect 7239 23100 7251 23103
rect 7300 23100 7328 23128
rect 7239 23072 7328 23100
rect 7239 23069 7251 23072
rect 7193 23063 7251 23069
rect 7392 23041 7420 23140
rect 7469 23103 7527 23109
rect 7469 23069 7481 23103
rect 7515 23069 7527 23103
rect 7469 23063 7527 23069
rect 7377 23035 7435 23041
rect 7377 23001 7389 23035
rect 7423 23001 7435 23035
rect 7377 22995 7435 23001
rect 5592 22936 5856 22964
rect 5592 22924 5598 22936
rect 5902 22924 5908 22976
rect 5960 22964 5966 22976
rect 6089 22967 6147 22973
rect 6089 22964 6101 22967
rect 5960 22936 6101 22964
rect 5960 22924 5966 22936
rect 6089 22933 6101 22936
rect 6135 22933 6147 22967
rect 6089 22927 6147 22933
rect 6730 22924 6736 22976
rect 6788 22964 6794 22976
rect 7392 22964 7420 22995
rect 6788 22936 7420 22964
rect 7484 22964 7512 23063
rect 7558 23060 7564 23112
rect 7616 23060 7622 23112
rect 7668 23032 7696 23140
rect 7926 23128 7932 23180
rect 7984 23168 7990 23180
rect 9784 23168 9812 23208
rect 10965 23205 10977 23239
rect 11011 23236 11023 23239
rect 11790 23236 11796 23248
rect 11011 23208 11796 23236
rect 11011 23205 11023 23208
rect 10965 23199 11023 23205
rect 11790 23196 11796 23208
rect 11848 23236 11854 23248
rect 13998 23236 14004 23248
rect 11848 23208 14004 23236
rect 11848 23196 11854 23208
rect 13998 23196 14004 23208
rect 14056 23196 14062 23248
rect 7984 23140 8340 23168
rect 9784 23140 13400 23168
rect 7984 23128 7990 23140
rect 7834 23060 7840 23112
rect 7892 23060 7898 23112
rect 8110 23060 8116 23112
rect 8168 23060 8174 23112
rect 8202 23060 8208 23112
rect 8260 23060 8266 23112
rect 8021 23035 8079 23041
rect 8021 23032 8033 23035
rect 7668 23004 8033 23032
rect 8021 23001 8033 23004
rect 8067 23001 8079 23035
rect 8312 23032 8340 23140
rect 10778 23060 10784 23112
rect 10836 23060 10842 23112
rect 11054 23060 11060 23112
rect 11112 23060 11118 23112
rect 11333 23103 11391 23109
rect 11333 23069 11345 23103
rect 11379 23100 11391 23103
rect 11974 23100 11980 23112
rect 11379 23072 11980 23100
rect 11379 23069 11391 23072
rect 11333 23063 11391 23069
rect 11974 23060 11980 23072
rect 12032 23100 12038 23112
rect 12345 23103 12403 23109
rect 12345 23100 12357 23103
rect 12032 23072 12357 23100
rect 12032 23060 12038 23072
rect 12345 23069 12357 23072
rect 12391 23069 12403 23103
rect 12345 23063 12403 23069
rect 12621 23103 12679 23109
rect 12621 23069 12633 23103
rect 12667 23100 12679 23103
rect 12802 23100 12808 23112
rect 12667 23072 12808 23100
rect 12667 23069 12679 23072
rect 12621 23063 12679 23069
rect 12802 23060 12808 23072
rect 12860 23060 12866 23112
rect 8312 23004 11376 23032
rect 8021 22995 8079 23001
rect 7650 22964 7656 22976
rect 7484 22936 7656 22964
rect 6788 22924 6794 22936
rect 7650 22924 7656 22936
rect 7708 22924 7714 22976
rect 7745 22967 7803 22973
rect 7745 22933 7757 22967
rect 7791 22964 7803 22967
rect 8294 22964 8300 22976
rect 7791 22936 8300 22964
rect 7791 22933 7803 22936
rect 7745 22927 7803 22933
rect 8294 22924 8300 22936
rect 8352 22924 8358 22976
rect 8389 22967 8447 22973
rect 8389 22933 8401 22967
rect 8435 22964 8447 22967
rect 11054 22964 11060 22976
rect 8435 22936 11060 22964
rect 8435 22933 8447 22936
rect 8389 22927 8447 22933
rect 11054 22924 11060 22936
rect 11112 22924 11118 22976
rect 11238 22924 11244 22976
rect 11296 22924 11302 22976
rect 11348 22964 11376 23004
rect 11514 22992 11520 23044
rect 11572 22992 11578 23044
rect 12066 23032 12072 23044
rect 11624 23004 12072 23032
rect 11624 22964 11652 23004
rect 12066 22992 12072 23004
rect 12124 22992 12130 23044
rect 11348 22936 11652 22964
rect 11698 22924 11704 22976
rect 11756 22924 11762 22976
rect 11882 22924 11888 22976
rect 11940 22964 11946 22976
rect 12618 22964 12624 22976
rect 11940 22936 12624 22964
rect 11940 22924 11946 22936
rect 12618 22924 12624 22936
rect 12676 22924 12682 22976
rect 13372 22964 13400 23140
rect 13446 23060 13452 23112
rect 13504 23100 13510 23112
rect 14108 23100 14136 23267
rect 16298 23264 16304 23276
rect 16356 23264 16362 23316
rect 16393 23307 16451 23313
rect 16393 23273 16405 23307
rect 16439 23304 16451 23307
rect 16574 23304 16580 23316
rect 16439 23276 16580 23304
rect 16439 23273 16451 23276
rect 16393 23267 16451 23273
rect 16574 23264 16580 23276
rect 16632 23264 16638 23316
rect 17770 23264 17776 23316
rect 17828 23264 17834 23316
rect 18046 23264 18052 23316
rect 18104 23304 18110 23316
rect 18693 23307 18751 23313
rect 18104 23276 18644 23304
rect 18104 23264 18110 23276
rect 14553 23239 14611 23245
rect 14553 23205 14565 23239
rect 14599 23236 14611 23239
rect 14599 23208 18460 23236
rect 14599 23205 14611 23208
rect 14553 23199 14611 23205
rect 16574 23128 16580 23180
rect 16632 23168 16638 23180
rect 16850 23168 16856 23180
rect 16632 23140 16856 23168
rect 16632 23128 16638 23140
rect 16850 23128 16856 23140
rect 16908 23128 16914 23180
rect 17586 23128 17592 23180
rect 17644 23168 17650 23180
rect 17957 23171 18015 23177
rect 17957 23168 17969 23171
rect 17644 23140 17969 23168
rect 17644 23128 17650 23140
rect 17957 23137 17969 23140
rect 18003 23137 18015 23171
rect 17957 23131 18015 23137
rect 13504 23072 14136 23100
rect 14277 23103 14335 23109
rect 13504 23060 13510 23072
rect 14277 23069 14289 23103
rect 14323 23069 14335 23103
rect 14277 23063 14335 23069
rect 13998 22992 14004 23044
rect 14056 23032 14062 23044
rect 14093 23035 14151 23041
rect 14093 23032 14105 23035
rect 14056 23004 14105 23032
rect 14056 22992 14062 23004
rect 14093 23001 14105 23004
rect 14139 23001 14151 23035
rect 14292 23032 14320 23063
rect 14366 23060 14372 23112
rect 14424 23100 14430 23112
rect 15010 23100 15016 23112
rect 14424 23072 15016 23100
rect 14424 23060 14430 23072
rect 15010 23060 15016 23072
rect 15068 23060 15074 23112
rect 15378 23060 15384 23112
rect 15436 23100 15442 23112
rect 16025 23103 16083 23109
rect 16025 23100 16037 23103
rect 15436 23072 16037 23100
rect 15436 23060 15442 23072
rect 16025 23069 16037 23072
rect 16071 23069 16083 23103
rect 16025 23063 16083 23069
rect 16209 23103 16267 23109
rect 16209 23069 16221 23103
rect 16255 23100 16267 23103
rect 16390 23100 16396 23112
rect 16255 23072 16396 23100
rect 16255 23069 16267 23072
rect 16209 23063 16267 23069
rect 14550 23032 14556 23044
rect 14292 23004 14556 23032
rect 14093 22995 14151 23001
rect 14550 22992 14556 23004
rect 14608 22992 14614 23044
rect 15194 22992 15200 23044
rect 15252 23032 15258 23044
rect 16224 23032 16252 23063
rect 16390 23060 16396 23072
rect 16448 23060 16454 23112
rect 18432 23109 18460 23208
rect 18506 23128 18512 23180
rect 18564 23128 18570 23180
rect 18616 23168 18644 23276
rect 18693 23273 18705 23307
rect 18739 23273 18751 23307
rect 18693 23267 18751 23273
rect 18708 23236 18736 23267
rect 19702 23264 19708 23316
rect 19760 23304 19766 23316
rect 20073 23307 20131 23313
rect 20073 23304 20085 23307
rect 19760 23276 20085 23304
rect 19760 23264 19766 23276
rect 20073 23273 20085 23276
rect 20119 23273 20131 23307
rect 20073 23267 20131 23273
rect 20346 23264 20352 23316
rect 20404 23304 20410 23316
rect 20714 23304 20720 23316
rect 20404 23276 20720 23304
rect 20404 23264 20410 23276
rect 20714 23264 20720 23276
rect 20772 23264 20778 23316
rect 21726 23264 21732 23316
rect 21784 23264 21790 23316
rect 22554 23304 22560 23316
rect 21836 23276 22560 23304
rect 19889 23239 19947 23245
rect 19889 23236 19901 23239
rect 18708 23208 19901 23236
rect 19889 23205 19901 23208
rect 19935 23236 19947 23239
rect 20806 23236 20812 23248
rect 19935 23208 20812 23236
rect 19935 23205 19947 23208
rect 19889 23199 19947 23205
rect 20806 23196 20812 23208
rect 20864 23196 20870 23248
rect 20898 23196 20904 23248
rect 20956 23236 20962 23248
rect 21836 23236 21864 23276
rect 22554 23264 22560 23276
rect 22612 23264 22618 23316
rect 22830 23264 22836 23316
rect 22888 23304 22894 23316
rect 23566 23304 23572 23316
rect 22888 23276 23572 23304
rect 22888 23264 22894 23276
rect 23566 23264 23572 23276
rect 23624 23264 23630 23316
rect 24670 23264 24676 23316
rect 24728 23264 24734 23316
rect 25038 23304 25044 23316
rect 24780 23276 25044 23304
rect 24780 23236 24808 23276
rect 25038 23264 25044 23276
rect 25096 23264 25102 23316
rect 25774 23264 25780 23316
rect 25832 23264 25838 23316
rect 25961 23307 26019 23313
rect 25961 23273 25973 23307
rect 26007 23304 26019 23307
rect 26234 23304 26240 23316
rect 26007 23276 26240 23304
rect 26007 23273 26019 23276
rect 25961 23267 26019 23273
rect 26234 23264 26240 23276
rect 26292 23264 26298 23316
rect 26418 23264 26424 23316
rect 26476 23264 26482 23316
rect 26881 23307 26939 23313
rect 26881 23273 26893 23307
rect 26927 23304 26939 23307
rect 28629 23307 28687 23313
rect 28629 23304 28641 23307
rect 26927 23276 28641 23304
rect 26927 23273 26939 23276
rect 26881 23267 26939 23273
rect 28629 23273 28641 23276
rect 28675 23273 28687 23307
rect 32674 23304 32680 23316
rect 28629 23267 28687 23273
rect 28828 23276 32680 23304
rect 20956 23208 21864 23236
rect 21928 23208 24808 23236
rect 24857 23239 24915 23245
rect 20956 23196 20962 23208
rect 19518 23168 19524 23180
rect 18616 23140 19524 23168
rect 19518 23128 19524 23140
rect 19576 23128 19582 23180
rect 21928 23168 21956 23208
rect 24857 23205 24869 23239
rect 24903 23236 24915 23239
rect 24903 23208 28672 23236
rect 24903 23205 24915 23208
rect 24857 23199 24915 23205
rect 19628 23140 21956 23168
rect 18049 23103 18107 23109
rect 18049 23100 18061 23103
rect 17604 23072 18061 23100
rect 17604 23044 17632 23072
rect 18049 23069 18061 23072
rect 18095 23069 18107 23103
rect 18049 23063 18107 23069
rect 18417 23103 18475 23109
rect 18417 23069 18429 23103
rect 18463 23069 18475 23103
rect 18417 23063 18475 23069
rect 18693 23103 18751 23109
rect 18693 23069 18705 23103
rect 18739 23100 18751 23103
rect 19058 23100 19064 23112
rect 18739 23072 19064 23100
rect 18739 23069 18751 23072
rect 18693 23063 18751 23069
rect 19058 23060 19064 23072
rect 19116 23060 19122 23112
rect 19150 23060 19156 23112
rect 19208 23100 19214 23112
rect 19628 23100 19656 23140
rect 22370 23128 22376 23180
rect 22428 23168 22434 23180
rect 24581 23171 24639 23177
rect 22428 23140 24440 23168
rect 22428 23128 22434 23140
rect 20073 23103 20131 23109
rect 20073 23100 20085 23103
rect 19208 23072 19656 23100
rect 19720 23072 20085 23100
rect 19208 23060 19214 23072
rect 15252 23004 16252 23032
rect 15252 22992 15258 23004
rect 17586 22992 17592 23044
rect 17644 22992 17650 23044
rect 17678 22992 17684 23044
rect 17736 23032 17742 23044
rect 17773 23035 17831 23041
rect 17773 23032 17785 23035
rect 17736 23004 17785 23032
rect 17736 22992 17742 23004
rect 17773 23001 17785 23004
rect 17819 23001 17831 23035
rect 19720 23032 19748 23072
rect 20073 23069 20085 23072
rect 20119 23069 20131 23103
rect 20073 23063 20131 23069
rect 20165 23103 20223 23109
rect 20165 23069 20177 23103
rect 20211 23069 20223 23103
rect 20165 23063 20223 23069
rect 20180 23032 20208 23063
rect 20254 23060 20260 23112
rect 20312 23100 20318 23112
rect 21174 23100 21180 23112
rect 20312 23072 21180 23100
rect 20312 23060 20318 23072
rect 21174 23060 21180 23072
rect 21232 23060 21238 23112
rect 21729 23103 21787 23109
rect 21729 23069 21741 23103
rect 21775 23069 21787 23103
rect 21729 23063 21787 23069
rect 17773 22995 17831 23001
rect 17880 23004 19748 23032
rect 19904 23004 20208 23032
rect 20349 23035 20407 23041
rect 15654 22964 15660 22976
rect 13372 22936 15660 22964
rect 15654 22924 15660 22936
rect 15712 22924 15718 22976
rect 16022 22924 16028 22976
rect 16080 22964 16086 22976
rect 16390 22964 16396 22976
rect 16080 22936 16396 22964
rect 16080 22924 16086 22936
rect 16390 22924 16396 22936
rect 16448 22924 16454 22976
rect 16942 22924 16948 22976
rect 17000 22964 17006 22976
rect 17880 22964 17908 23004
rect 17000 22936 17908 22964
rect 17000 22924 17006 22936
rect 18230 22924 18236 22976
rect 18288 22924 18294 22976
rect 18874 22924 18880 22976
rect 18932 22924 18938 22976
rect 18966 22924 18972 22976
rect 19024 22964 19030 22976
rect 19904 22964 19932 23004
rect 20349 23001 20361 23035
rect 20395 23032 20407 23035
rect 20441 23035 20499 23041
rect 20441 23032 20453 23035
rect 20395 23004 20453 23032
rect 20395 23001 20407 23004
rect 20349 22995 20407 23001
rect 20441 23001 20453 23004
rect 20487 23001 20499 23035
rect 20441 22995 20499 23001
rect 20625 23035 20683 23041
rect 20625 23001 20637 23035
rect 20671 23032 20683 23035
rect 20714 23032 20720 23044
rect 20671 23004 20720 23032
rect 20671 23001 20683 23004
rect 20625 22995 20683 23001
rect 20714 22992 20720 23004
rect 20772 22992 20778 23044
rect 20809 23035 20867 23041
rect 20809 23001 20821 23035
rect 20855 23001 20867 23035
rect 20809 22995 20867 23001
rect 21545 23035 21603 23041
rect 21545 23001 21557 23035
rect 21591 23001 21603 23035
rect 21744 23032 21772 23063
rect 21818 23060 21824 23112
rect 21876 23060 21882 23112
rect 22186 23060 22192 23112
rect 22244 23100 22250 23112
rect 22465 23103 22523 23109
rect 22465 23100 22477 23103
rect 22244 23072 22477 23100
rect 22244 23060 22250 23072
rect 22465 23069 22477 23072
rect 22511 23100 22523 23103
rect 23109 23103 23167 23109
rect 23109 23100 23121 23103
rect 22511 23072 23121 23100
rect 22511 23069 22523 23072
rect 22465 23063 22523 23069
rect 23109 23069 23121 23072
rect 23155 23069 23167 23103
rect 23109 23063 23167 23069
rect 23290 23060 23296 23112
rect 23348 23060 23354 23112
rect 24412 23109 24440 23140
rect 24581 23137 24593 23171
rect 24627 23168 24639 23171
rect 25038 23168 25044 23180
rect 24627 23140 25044 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 25038 23128 25044 23140
rect 25096 23128 25102 23180
rect 26050 23128 26056 23180
rect 26108 23168 26114 23180
rect 26510 23168 26516 23180
rect 26108 23140 26516 23168
rect 26108 23128 26114 23140
rect 26510 23128 26516 23140
rect 26568 23128 26574 23180
rect 24397 23103 24455 23109
rect 24397 23069 24409 23103
rect 24443 23069 24455 23103
rect 24397 23063 24455 23069
rect 24486 23060 24492 23112
rect 24544 23100 24550 23112
rect 24673 23103 24731 23109
rect 24673 23100 24685 23103
rect 24544 23072 24685 23100
rect 24544 23060 24550 23072
rect 24673 23069 24685 23072
rect 24719 23069 24731 23103
rect 24673 23063 24731 23069
rect 22281 23035 22339 23041
rect 21744 23004 22232 23032
rect 21545 22995 21603 23001
rect 19024 22936 19932 22964
rect 19024 22924 19030 22936
rect 19978 22924 19984 22976
rect 20036 22964 20042 22976
rect 20824 22964 20852 22995
rect 20036 22936 20852 22964
rect 21560 22964 21588 22995
rect 21910 22964 21916 22976
rect 21560 22936 21916 22964
rect 20036 22924 20042 22936
rect 21910 22924 21916 22936
rect 21968 22924 21974 22976
rect 22002 22924 22008 22976
rect 22060 22924 22066 22976
rect 22094 22924 22100 22976
rect 22152 22924 22158 22976
rect 22204 22964 22232 23004
rect 22281 23001 22293 23035
rect 22327 23032 22339 23035
rect 22554 23032 22560 23044
rect 22327 23004 22560 23032
rect 22327 23001 22339 23004
rect 22281 22995 22339 23001
rect 22554 22992 22560 23004
rect 22612 22992 22618 23044
rect 22646 22992 22652 23044
rect 22704 22992 22710 23044
rect 24688 23032 24716 23063
rect 24854 23060 24860 23112
rect 24912 23100 24918 23112
rect 25685 23103 25743 23109
rect 25685 23100 25697 23103
rect 24912 23072 25697 23100
rect 24912 23060 24918 23072
rect 25685 23069 25697 23072
rect 25731 23069 25743 23103
rect 25685 23063 25743 23069
rect 25777 23103 25835 23109
rect 25777 23069 25789 23103
rect 25823 23100 25835 23103
rect 25958 23100 25964 23112
rect 25823 23072 25964 23100
rect 25823 23069 25835 23072
rect 25777 23063 25835 23069
rect 24949 23035 25007 23041
rect 24949 23032 24961 23035
rect 24688 23004 24961 23032
rect 24949 23001 24961 23004
rect 24995 23001 25007 23035
rect 24949 22995 25007 23001
rect 25498 22992 25504 23044
rect 25556 22992 25562 23044
rect 25590 22992 25596 23044
rect 25648 23032 25654 23044
rect 25792 23032 25820 23063
rect 25958 23060 25964 23072
rect 26016 23060 26022 23112
rect 26142 23060 26148 23112
rect 26200 23100 26206 23112
rect 26421 23103 26479 23109
rect 26421 23100 26433 23103
rect 26200 23072 26433 23100
rect 26200 23060 26206 23072
rect 26421 23069 26433 23072
rect 26467 23069 26479 23103
rect 26421 23063 26479 23069
rect 26697 23103 26755 23109
rect 26697 23069 26709 23103
rect 26743 23100 26755 23103
rect 27154 23100 27160 23112
rect 26743 23072 27160 23100
rect 26743 23069 26755 23072
rect 26697 23063 26755 23069
rect 27154 23060 27160 23072
rect 27212 23060 27218 23112
rect 28644 23109 28672 23208
rect 28828 23177 28856 23276
rect 32674 23264 32680 23276
rect 32732 23264 32738 23316
rect 28813 23171 28871 23177
rect 28813 23137 28825 23171
rect 28859 23137 28871 23171
rect 28813 23131 28871 23137
rect 30650 23128 30656 23180
rect 30708 23168 30714 23180
rect 31113 23171 31171 23177
rect 31113 23168 31125 23171
rect 30708 23140 31125 23168
rect 30708 23128 30714 23140
rect 31113 23137 31125 23140
rect 31159 23137 31171 23171
rect 31113 23131 31171 23137
rect 28629 23103 28687 23109
rect 28629 23069 28641 23103
rect 28675 23069 28687 23103
rect 28629 23063 28687 23069
rect 28902 23060 28908 23112
rect 28960 23060 28966 23112
rect 31021 23103 31079 23109
rect 31021 23069 31033 23103
rect 31067 23100 31079 23103
rect 31754 23100 31760 23112
rect 31067 23072 31760 23100
rect 31067 23069 31079 23072
rect 31021 23063 31079 23069
rect 31754 23060 31760 23072
rect 31812 23060 31818 23112
rect 25648 23004 25820 23032
rect 25648 22992 25654 23004
rect 26234 22992 26240 23044
rect 26292 23032 26298 23044
rect 29549 23035 29607 23041
rect 29549 23032 29561 23035
rect 26292 23004 29561 23032
rect 26292 22992 26298 23004
rect 29549 23001 29561 23004
rect 29595 23001 29607 23035
rect 29549 22995 29607 23001
rect 29733 23035 29791 23041
rect 29733 23001 29745 23035
rect 29779 23001 29791 23035
rect 29733 22995 29791 23001
rect 31380 23035 31438 23041
rect 31380 23001 31392 23035
rect 31426 23032 31438 23035
rect 31478 23032 31484 23044
rect 31426 23004 31484 23032
rect 31426 23001 31438 23004
rect 31380 22995 31438 23001
rect 22738 22964 22744 22976
rect 22204 22936 22744 22964
rect 22738 22924 22744 22936
rect 22796 22924 22802 22976
rect 22830 22924 22836 22976
rect 22888 22964 22894 22976
rect 22925 22967 22983 22973
rect 22925 22964 22937 22967
rect 22888 22936 22937 22964
rect 22888 22924 22894 22936
rect 22925 22933 22937 22936
rect 22971 22933 22983 22967
rect 22925 22927 22983 22933
rect 29089 22967 29147 22973
rect 29089 22933 29101 22967
rect 29135 22964 29147 22967
rect 29748 22964 29776 22995
rect 31478 22992 31484 23004
rect 31536 22992 31542 23044
rect 29135 22936 29776 22964
rect 29135 22933 29147 22936
rect 29089 22927 29147 22933
rect 29822 22924 29828 22976
rect 29880 22964 29886 22976
rect 29917 22967 29975 22973
rect 29917 22964 29929 22967
rect 29880 22936 29929 22964
rect 29880 22924 29886 22936
rect 29917 22933 29929 22936
rect 29963 22933 29975 22967
rect 29917 22927 29975 22933
rect 30098 22924 30104 22976
rect 30156 22964 30162 22976
rect 30377 22967 30435 22973
rect 30377 22964 30389 22967
rect 30156 22936 30389 22964
rect 30156 22924 30162 22936
rect 30377 22933 30389 22936
rect 30423 22933 30435 22967
rect 30377 22927 30435 22933
rect 32493 22967 32551 22973
rect 32493 22933 32505 22967
rect 32539 22964 32551 22967
rect 32582 22964 32588 22976
rect 32539 22936 32588 22964
rect 32539 22933 32551 22936
rect 32493 22927 32551 22933
rect 32582 22924 32588 22936
rect 32640 22924 32646 22976
rect 1104 22874 32844 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 32844 22874
rect 1104 22800 32844 22822
rect 2314 22720 2320 22772
rect 2372 22760 2378 22772
rect 2777 22763 2835 22769
rect 2777 22760 2789 22763
rect 2372 22732 2789 22760
rect 2372 22720 2378 22732
rect 2777 22729 2789 22732
rect 2823 22729 2835 22763
rect 2777 22723 2835 22729
rect 2958 22720 2964 22772
rect 3016 22760 3022 22772
rect 3237 22763 3295 22769
rect 3237 22760 3249 22763
rect 3016 22732 3249 22760
rect 3016 22720 3022 22732
rect 3237 22729 3249 22732
rect 3283 22729 3295 22763
rect 3237 22723 3295 22729
rect 3513 22763 3571 22769
rect 3513 22729 3525 22763
rect 3559 22760 3571 22763
rect 6181 22763 6239 22769
rect 3559 22732 5856 22760
rect 3559 22729 3571 22732
rect 3513 22723 3571 22729
rect 3050 22652 3056 22704
rect 3108 22692 3114 22704
rect 3354 22695 3412 22701
rect 3354 22692 3366 22695
rect 3108 22664 3366 22692
rect 3108 22652 3114 22664
rect 3354 22661 3366 22664
rect 3400 22692 3412 22695
rect 3970 22692 3976 22704
rect 3400 22664 3976 22692
rect 3400 22661 3412 22664
rect 3354 22655 3412 22661
rect 3970 22652 3976 22664
rect 4028 22652 4034 22704
rect 4430 22652 4436 22704
rect 4488 22692 4494 22704
rect 4709 22695 4767 22701
rect 4709 22692 4721 22695
rect 4488 22664 4721 22692
rect 4488 22652 4494 22664
rect 4709 22661 4721 22664
rect 4755 22661 4767 22695
rect 4709 22655 4767 22661
rect 5721 22651 5779 22657
rect 1670 22633 1676 22636
rect 1664 22587 1676 22633
rect 1670 22584 1676 22587
rect 1728 22584 1734 22636
rect 2774 22584 2780 22636
rect 2832 22624 2838 22636
rect 2869 22627 2927 22633
rect 2869 22624 2881 22627
rect 2832 22596 2881 22624
rect 2832 22584 2838 22596
rect 2869 22593 2881 22596
rect 2915 22624 2927 22627
rect 4090 22627 4148 22633
rect 4090 22624 4102 22627
rect 2915 22596 4102 22624
rect 2915 22593 2927 22596
rect 2869 22587 2927 22593
rect 4090 22593 4102 22596
rect 4136 22593 4148 22627
rect 4090 22587 4148 22593
rect 4617 22627 4675 22633
rect 4617 22593 4629 22627
rect 4663 22593 4675 22627
rect 4617 22587 4675 22593
rect 1394 22516 1400 22568
rect 1452 22516 1458 22568
rect 3145 22559 3203 22565
rect 3145 22525 3157 22559
rect 3191 22556 3203 22559
rect 3605 22559 3663 22565
rect 3605 22556 3617 22559
rect 3191 22528 3617 22556
rect 3191 22525 3203 22528
rect 3145 22519 3203 22525
rect 3605 22525 3617 22528
rect 3651 22556 3663 22559
rect 3694 22556 3700 22568
rect 3651 22528 3700 22556
rect 3651 22525 3663 22528
rect 3605 22519 3663 22525
rect 3694 22516 3700 22528
rect 3752 22516 3758 22568
rect 3881 22559 3939 22565
rect 3881 22525 3893 22559
rect 3927 22525 3939 22559
rect 4632 22556 4660 22587
rect 4798 22584 4804 22636
rect 4856 22584 4862 22636
rect 4982 22584 4988 22636
rect 5040 22584 5046 22636
rect 5074 22584 5080 22636
rect 5132 22624 5138 22636
rect 5169 22627 5227 22633
rect 5620 22631 5678 22637
rect 5620 22628 5632 22631
rect 5169 22624 5181 22627
rect 5132 22596 5181 22624
rect 5132 22584 5138 22596
rect 5169 22593 5181 22596
rect 5215 22593 5227 22627
rect 5169 22587 5227 22593
rect 5552 22600 5632 22628
rect 4890 22556 4896 22568
rect 4632 22528 4896 22556
rect 3881 22519 3939 22525
rect 2958 22448 2964 22500
rect 3016 22488 3022 22500
rect 3786 22488 3792 22500
rect 3016 22460 3792 22488
rect 3016 22448 3022 22460
rect 3786 22448 3792 22460
rect 3844 22488 3850 22500
rect 3896 22488 3924 22519
rect 4890 22516 4896 22528
rect 4948 22516 4954 22568
rect 3844 22460 3924 22488
rect 4249 22491 4307 22497
rect 3844 22448 3850 22460
rect 4249 22457 4261 22491
rect 4295 22488 4307 22491
rect 4706 22488 4712 22500
rect 4295 22460 4712 22488
rect 4295 22457 4307 22460
rect 4249 22451 4307 22457
rect 4706 22448 4712 22460
rect 4764 22448 4770 22500
rect 4798 22448 4804 22500
rect 4856 22488 4862 22500
rect 5445 22491 5503 22497
rect 5445 22488 5457 22491
rect 4856 22460 5457 22488
rect 4856 22448 4862 22460
rect 5445 22457 5457 22460
rect 5491 22457 5503 22491
rect 5552 22488 5580 22600
rect 5620 22597 5632 22600
rect 5666 22597 5678 22631
rect 5721 22617 5733 22651
rect 5767 22648 5779 22651
rect 5828 22648 5856 22732
rect 6181 22729 6193 22763
rect 6227 22729 6239 22763
rect 6181 22723 6239 22729
rect 6086 22652 6092 22704
rect 6144 22652 6150 22704
rect 6196 22692 6224 22723
rect 6638 22720 6644 22772
rect 6696 22720 6702 22772
rect 6730 22720 6736 22772
rect 6788 22760 6794 22772
rect 7193 22763 7251 22769
rect 7193 22760 7205 22763
rect 6788 22732 7205 22760
rect 6788 22720 6794 22732
rect 7193 22729 7205 22732
rect 7239 22729 7251 22763
rect 7193 22723 7251 22729
rect 7469 22763 7527 22769
rect 7469 22729 7481 22763
rect 7515 22760 7527 22763
rect 7558 22760 7564 22772
rect 7515 22732 7564 22760
rect 7515 22729 7527 22732
rect 7469 22723 7527 22729
rect 7558 22720 7564 22732
rect 7616 22720 7622 22772
rect 7834 22720 7840 22772
rect 7892 22760 7898 22772
rect 9398 22760 9404 22772
rect 7892 22732 9404 22760
rect 7892 22720 7898 22732
rect 9398 22720 9404 22732
rect 9456 22720 9462 22772
rect 10686 22720 10692 22772
rect 10744 22760 10750 22772
rect 11103 22763 11161 22769
rect 11103 22760 11115 22763
rect 10744 22732 11115 22760
rect 10744 22720 10750 22732
rect 11103 22729 11115 22732
rect 11149 22760 11161 22763
rect 11606 22760 11612 22772
rect 11149 22732 11612 22760
rect 11149 22729 11161 22732
rect 11103 22723 11161 22729
rect 11606 22720 11612 22732
rect 11664 22720 11670 22772
rect 12342 22720 12348 22772
rect 12400 22760 12406 22772
rect 12529 22763 12587 22769
rect 12529 22760 12541 22763
rect 12400 22732 12541 22760
rect 12400 22720 12406 22732
rect 12529 22729 12541 22732
rect 12575 22760 12587 22763
rect 12894 22760 12900 22772
rect 12575 22732 12900 22760
rect 12575 22729 12587 22732
rect 12529 22723 12587 22729
rect 12894 22720 12900 22732
rect 12952 22720 12958 22772
rect 13173 22763 13231 22769
rect 13173 22729 13185 22763
rect 13219 22760 13231 22763
rect 13354 22760 13360 22772
rect 13219 22732 13360 22760
rect 13219 22729 13231 22732
rect 13173 22723 13231 22729
rect 13354 22720 13360 22732
rect 13412 22720 13418 22772
rect 13446 22720 13452 22772
rect 13504 22760 13510 22772
rect 13814 22760 13820 22772
rect 13504 22732 13820 22760
rect 13504 22720 13510 22732
rect 13814 22720 13820 22732
rect 13872 22760 13878 22772
rect 18138 22760 18144 22772
rect 13872 22732 18144 22760
rect 13872 22720 13878 22732
rect 18138 22720 18144 22732
rect 18196 22720 18202 22772
rect 19061 22763 19119 22769
rect 19061 22729 19073 22763
rect 19107 22760 19119 22763
rect 19150 22760 19156 22772
rect 19107 22732 19156 22760
rect 19107 22729 19119 22732
rect 19061 22723 19119 22729
rect 19150 22720 19156 22732
rect 19208 22720 19214 22772
rect 19337 22763 19395 22769
rect 19337 22729 19349 22763
rect 19383 22760 19395 22763
rect 19426 22760 19432 22772
rect 19383 22732 19432 22760
rect 19383 22729 19395 22732
rect 19337 22723 19395 22729
rect 19426 22720 19432 22732
rect 19484 22720 19490 22772
rect 19610 22720 19616 22772
rect 19668 22760 19674 22772
rect 20254 22760 20260 22772
rect 19668 22732 20260 22760
rect 19668 22720 19674 22732
rect 20254 22720 20260 22732
rect 20312 22720 20318 22772
rect 20533 22763 20591 22769
rect 20533 22729 20545 22763
rect 20579 22729 20591 22763
rect 20533 22723 20591 22729
rect 6546 22692 6552 22704
rect 6196 22664 6552 22692
rect 6546 22652 6552 22664
rect 6604 22652 6610 22704
rect 5767 22620 5856 22648
rect 5767 22617 5779 22620
rect 5721 22611 5779 22617
rect 5620 22591 5678 22597
rect 5902 22584 5908 22636
rect 5960 22624 5966 22636
rect 5997 22627 6055 22633
rect 5997 22624 6009 22627
rect 5960 22596 6009 22624
rect 5960 22584 5966 22596
rect 5997 22593 6009 22596
rect 6043 22593 6055 22627
rect 5997 22587 6055 22593
rect 6104 22556 6132 22652
rect 6270 22584 6276 22636
rect 6328 22624 6334 22636
rect 6656 22633 6684 22720
rect 9766 22692 9772 22704
rect 6748 22664 7144 22692
rect 6748 22633 6776 22664
rect 6365 22627 6423 22633
rect 6365 22624 6377 22627
rect 6328 22596 6377 22624
rect 6328 22584 6334 22596
rect 6365 22593 6377 22596
rect 6411 22593 6423 22627
rect 6365 22587 6423 22593
rect 6641 22627 6699 22633
rect 6641 22593 6653 22627
rect 6687 22593 6699 22627
rect 6641 22587 6699 22593
rect 6733 22627 6791 22633
rect 6733 22593 6745 22627
rect 6779 22593 6791 22627
rect 7009 22627 7067 22633
rect 7009 22624 7021 22627
rect 6733 22587 6791 22593
rect 6840 22596 7021 22624
rect 6748 22556 6776 22587
rect 6104 22528 6776 22556
rect 5905 22491 5963 22497
rect 5905 22488 5917 22491
rect 5552 22460 5917 22488
rect 5445 22451 5503 22457
rect 5905 22457 5917 22460
rect 5951 22488 5963 22491
rect 6086 22488 6092 22500
rect 5951 22460 6092 22488
rect 5951 22457 5963 22460
rect 5905 22451 5963 22457
rect 4433 22423 4491 22429
rect 4433 22389 4445 22423
rect 4479 22420 4491 22423
rect 5258 22420 5264 22432
rect 4479 22392 5264 22420
rect 4479 22389 4491 22392
rect 4433 22383 4491 22389
rect 5258 22380 5264 22392
rect 5316 22380 5322 22432
rect 5350 22380 5356 22432
rect 5408 22380 5414 22432
rect 5460 22420 5488 22451
rect 6086 22448 6092 22460
rect 6144 22448 6150 22500
rect 6840 22420 6868 22596
rect 7009 22593 7021 22596
rect 7055 22593 7067 22627
rect 7009 22587 7067 22593
rect 7116 22556 7144 22664
rect 8588 22664 9772 22692
rect 7190 22584 7196 22636
rect 7248 22624 7254 22636
rect 7285 22627 7343 22633
rect 7285 22624 7297 22627
rect 7248 22596 7297 22624
rect 7248 22584 7254 22596
rect 7285 22593 7297 22596
rect 7331 22593 7343 22627
rect 7285 22587 7343 22593
rect 7374 22584 7380 22636
rect 7432 22624 7438 22636
rect 7561 22627 7619 22633
rect 7561 22624 7573 22627
rect 7432 22596 7573 22624
rect 7432 22584 7438 22596
rect 7561 22593 7573 22596
rect 7607 22593 7619 22627
rect 7561 22587 7619 22593
rect 7834 22584 7840 22636
rect 7892 22624 7898 22636
rect 8588 22633 8616 22664
rect 9766 22652 9772 22664
rect 9824 22652 9830 22704
rect 9861 22695 9919 22701
rect 9861 22661 9873 22695
rect 9907 22692 9919 22695
rect 10502 22692 10508 22704
rect 9907 22664 10508 22692
rect 9907 22661 9919 22664
rect 9861 22655 9919 22661
rect 10502 22652 10508 22664
rect 10560 22652 10566 22704
rect 12713 22695 12771 22701
rect 11808 22664 12480 22692
rect 8573 22627 8631 22633
rect 8573 22624 8585 22627
rect 7892 22596 8585 22624
rect 7892 22584 7898 22596
rect 8573 22593 8585 22596
rect 8619 22593 8631 22627
rect 8573 22587 8631 22593
rect 8662 22584 8668 22636
rect 8720 22624 8726 22636
rect 8757 22627 8815 22633
rect 8757 22624 8769 22627
rect 8720 22596 8769 22624
rect 8720 22584 8726 22596
rect 8757 22593 8769 22596
rect 8803 22593 8815 22627
rect 8757 22587 8815 22593
rect 8846 22584 8852 22636
rect 8904 22584 8910 22636
rect 8938 22584 8944 22636
rect 8996 22633 9002 22636
rect 8996 22627 9023 22633
rect 9011 22593 9023 22627
rect 8996 22587 9023 22593
rect 10045 22627 10103 22633
rect 10045 22593 10057 22627
rect 10091 22593 10103 22627
rect 10045 22587 10103 22593
rect 8996 22584 9002 22587
rect 9677 22559 9735 22565
rect 7116 22528 8294 22556
rect 8266 22488 8294 22528
rect 9677 22525 9689 22559
rect 9723 22556 9735 22559
rect 9950 22556 9956 22568
rect 9723 22528 9956 22556
rect 9723 22525 9735 22528
rect 9677 22519 9735 22525
rect 9950 22516 9956 22528
rect 10008 22516 10014 22568
rect 10060 22556 10088 22587
rect 10226 22584 10232 22636
rect 10284 22584 10290 22636
rect 11238 22584 11244 22636
rect 11296 22624 11302 22636
rect 11808 22633 11836 22664
rect 11793 22627 11851 22633
rect 11793 22624 11805 22627
rect 11296 22596 11805 22624
rect 11296 22584 11302 22596
rect 11793 22593 11805 22596
rect 11839 22593 11851 22627
rect 11793 22587 11851 22593
rect 11882 22584 11888 22636
rect 11940 22584 11946 22636
rect 12066 22584 12072 22636
rect 12124 22584 12130 22636
rect 12250 22584 12256 22636
rect 12308 22624 12314 22636
rect 12345 22627 12403 22633
rect 12345 22624 12357 22627
rect 12308 22596 12357 22624
rect 12308 22584 12314 22596
rect 12345 22593 12357 22596
rect 12391 22593 12403 22627
rect 12452 22624 12480 22664
rect 12713 22661 12725 22695
rect 12759 22692 12771 22695
rect 13078 22692 13084 22704
rect 12759 22664 13084 22692
rect 12759 22661 12771 22664
rect 12713 22655 12771 22661
rect 13078 22652 13084 22664
rect 13136 22652 13142 22704
rect 14274 22652 14280 22704
rect 14332 22692 14338 22704
rect 16025 22695 16083 22701
rect 16025 22692 16037 22695
rect 14332 22664 16037 22692
rect 14332 22652 14338 22664
rect 16025 22661 16037 22664
rect 16071 22661 16083 22695
rect 20548 22692 20576 22723
rect 20714 22720 20720 22772
rect 20772 22760 20778 22772
rect 22462 22760 22468 22772
rect 20772 22732 22468 22760
rect 20772 22720 20778 22732
rect 22462 22720 22468 22732
rect 22520 22720 22526 22772
rect 23382 22720 23388 22772
rect 23440 22760 23446 22772
rect 24762 22760 24768 22772
rect 23440 22732 24768 22760
rect 23440 22720 23446 22732
rect 24762 22720 24768 22732
rect 24820 22720 24826 22772
rect 25409 22763 25467 22769
rect 25409 22729 25421 22763
rect 25455 22760 25467 22763
rect 25774 22760 25780 22772
rect 25455 22732 25780 22760
rect 25455 22729 25467 22732
rect 25409 22723 25467 22729
rect 25774 22720 25780 22732
rect 25832 22720 25838 22772
rect 30285 22763 30343 22769
rect 30285 22729 30297 22763
rect 30331 22729 30343 22763
rect 30285 22723 30343 22729
rect 20622 22692 20628 22704
rect 16025 22655 16083 22661
rect 16224 22664 19334 22692
rect 20548 22664 20628 22692
rect 12989 22627 13047 22633
rect 12989 22624 13001 22627
rect 12452 22596 13001 22624
rect 12345 22587 12403 22593
rect 12989 22593 13001 22596
rect 13035 22624 13047 22627
rect 13035 22596 14504 22624
rect 13035 22593 13047 22596
rect 12989 22587 13047 22593
rect 10962 22556 10968 22568
rect 10060 22528 10968 22556
rect 10962 22516 10968 22528
rect 11020 22516 11026 22568
rect 11333 22559 11391 22565
rect 11333 22525 11345 22559
rect 11379 22556 11391 22559
rect 11422 22556 11428 22568
rect 11379 22528 11428 22556
rect 11379 22525 11391 22528
rect 11333 22519 11391 22525
rect 11422 22516 11428 22528
rect 11480 22516 11486 22568
rect 8938 22488 8944 22500
rect 8266 22460 8944 22488
rect 8938 22448 8944 22460
rect 8996 22448 9002 22500
rect 9122 22448 9128 22500
rect 9180 22448 9186 22500
rect 10413 22491 10471 22497
rect 10413 22457 10425 22491
rect 10459 22488 10471 22491
rect 11900 22488 11928 22584
rect 12268 22556 12296 22584
rect 12084 22528 12296 22556
rect 12084 22500 12112 22528
rect 12618 22516 12624 22568
rect 12676 22556 12682 22568
rect 12805 22559 12863 22565
rect 12805 22556 12817 22559
rect 12676 22528 12817 22556
rect 12676 22516 12682 22528
rect 12805 22525 12817 22528
rect 12851 22525 12863 22559
rect 12805 22519 12863 22525
rect 13262 22516 13268 22568
rect 13320 22556 13326 22568
rect 14366 22556 14372 22568
rect 13320 22528 14372 22556
rect 13320 22516 13326 22528
rect 14366 22516 14372 22528
rect 14424 22516 14430 22568
rect 10459 22460 11928 22488
rect 10459 22457 10471 22460
rect 10413 22451 10471 22457
rect 12066 22448 12072 22500
rect 12124 22448 12130 22500
rect 12250 22448 12256 22500
rect 12308 22488 12314 22500
rect 12526 22488 12532 22500
rect 12308 22460 12532 22488
rect 12308 22448 12314 22460
rect 12526 22448 12532 22460
rect 12584 22448 12590 22500
rect 12894 22448 12900 22500
rect 12952 22488 12958 22500
rect 14274 22488 14280 22500
rect 12952 22460 14280 22488
rect 12952 22448 12958 22460
rect 14274 22448 14280 22460
rect 14332 22448 14338 22500
rect 14476 22488 14504 22596
rect 15948 22596 16160 22624
rect 14550 22516 14556 22568
rect 14608 22556 14614 22568
rect 15948 22556 15976 22596
rect 16132 22565 16160 22596
rect 14608 22528 15976 22556
rect 16117 22559 16175 22565
rect 14608 22516 14614 22528
rect 16117 22525 16129 22559
rect 16163 22525 16175 22559
rect 16117 22519 16175 22525
rect 16224 22488 16252 22664
rect 19306 22636 19334 22664
rect 20622 22652 20628 22664
rect 20680 22652 20686 22704
rect 20990 22652 20996 22704
rect 21048 22692 21054 22704
rect 27890 22692 27896 22704
rect 21048 22664 27896 22692
rect 21048 22652 21054 22664
rect 27890 22652 27896 22664
rect 27948 22652 27954 22704
rect 30009 22695 30067 22701
rect 30009 22661 30021 22695
rect 30055 22692 30067 22695
rect 30300 22692 30328 22723
rect 30622 22695 30680 22701
rect 30622 22692 30634 22695
rect 30055 22664 30236 22692
rect 30300 22664 30634 22692
rect 30055 22661 30067 22664
rect 30009 22655 30067 22661
rect 16301 22627 16359 22633
rect 16301 22593 16313 22627
rect 16347 22624 16359 22627
rect 16482 22624 16488 22636
rect 16347 22596 16488 22624
rect 16347 22593 16359 22596
rect 16301 22587 16359 22593
rect 16482 22584 16488 22596
rect 16540 22624 16546 22636
rect 17218 22624 17224 22636
rect 16540 22596 17224 22624
rect 16540 22584 16546 22596
rect 17218 22584 17224 22596
rect 17276 22584 17282 22636
rect 17494 22584 17500 22636
rect 17552 22624 17558 22636
rect 17589 22627 17647 22633
rect 17589 22624 17601 22627
rect 17552 22596 17601 22624
rect 17552 22584 17558 22596
rect 17589 22593 17601 22596
rect 17635 22593 17647 22627
rect 17589 22587 17647 22593
rect 17678 22584 17684 22636
rect 17736 22624 17742 22636
rect 18690 22624 18696 22636
rect 17736 22596 18696 22624
rect 17736 22584 17742 22596
rect 18690 22584 18696 22596
rect 18748 22624 18754 22636
rect 18877 22627 18935 22633
rect 18877 22624 18889 22627
rect 18748 22596 18889 22624
rect 18748 22584 18754 22596
rect 18877 22593 18889 22596
rect 18923 22593 18935 22627
rect 19153 22627 19211 22633
rect 19153 22624 19165 22627
rect 18877 22587 18935 22593
rect 18984 22596 19165 22624
rect 16390 22516 16396 22568
rect 16448 22556 16454 22568
rect 18984 22556 19012 22596
rect 19153 22593 19165 22596
rect 19199 22593 19211 22627
rect 19306 22596 19340 22636
rect 19153 22587 19211 22593
rect 19334 22584 19340 22596
rect 19392 22584 19398 22636
rect 19426 22584 19432 22636
rect 19484 22584 19490 22636
rect 19518 22584 19524 22636
rect 19576 22624 19582 22636
rect 19576 22596 19748 22624
rect 19576 22584 19582 22596
rect 19610 22556 19616 22568
rect 16448 22528 19012 22556
rect 19306 22528 19616 22556
rect 16448 22516 16454 22528
rect 14476 22460 16252 22488
rect 18782 22448 18788 22500
rect 18840 22488 18846 22500
rect 19306 22488 19334 22528
rect 19610 22516 19616 22528
rect 19668 22516 19674 22568
rect 19720 22556 19748 22596
rect 19794 22584 19800 22636
rect 19852 22584 19858 22636
rect 20073 22627 20131 22633
rect 20073 22593 20085 22627
rect 20119 22624 20131 22627
rect 20162 22624 20168 22636
rect 20119 22596 20168 22624
rect 20119 22593 20131 22596
rect 20073 22587 20131 22593
rect 20162 22584 20168 22596
rect 20220 22624 20226 22636
rect 20717 22627 20775 22633
rect 20717 22624 20729 22627
rect 20220 22596 20729 22624
rect 20220 22584 20226 22596
rect 20717 22593 20729 22596
rect 20763 22593 20775 22627
rect 20717 22587 20775 22593
rect 20809 22627 20867 22633
rect 20809 22593 20821 22627
rect 20855 22624 20867 22627
rect 20855 22596 21128 22624
rect 20855 22593 20867 22596
rect 20809 22587 20867 22593
rect 19720 22528 19840 22556
rect 18840 22460 19334 22488
rect 18840 22448 18846 22460
rect 5460 22392 6868 22420
rect 6917 22423 6975 22429
rect 6917 22389 6929 22423
rect 6963 22420 6975 22423
rect 7098 22420 7104 22432
rect 6963 22392 7104 22420
rect 6963 22389 6975 22392
rect 6917 22383 6975 22389
rect 7098 22380 7104 22392
rect 7156 22380 7162 22432
rect 7190 22380 7196 22432
rect 7248 22420 7254 22432
rect 7745 22423 7803 22429
rect 7745 22420 7757 22423
rect 7248 22392 7757 22420
rect 7248 22380 7254 22392
rect 7745 22389 7757 22392
rect 7791 22420 7803 22423
rect 8202 22420 8208 22432
rect 7791 22392 8208 22420
rect 7791 22389 7803 22392
rect 7745 22383 7803 22389
rect 8202 22380 8208 22392
rect 8260 22380 8266 22432
rect 9674 22380 9680 22432
rect 9732 22420 9738 22432
rect 9858 22420 9864 22432
rect 9732 22392 9864 22420
rect 9732 22380 9738 22392
rect 9858 22380 9864 22392
rect 9916 22380 9922 22432
rect 10778 22380 10784 22432
rect 10836 22420 10842 22432
rect 11517 22423 11575 22429
rect 11517 22420 11529 22423
rect 10836 22392 11529 22420
rect 10836 22380 10842 22392
rect 11517 22389 11529 22392
rect 11563 22389 11575 22423
rect 11517 22383 11575 22389
rect 11790 22380 11796 22432
rect 11848 22380 11854 22432
rect 11974 22380 11980 22432
rect 12032 22420 12038 22432
rect 12158 22420 12164 22432
rect 12032 22392 12164 22420
rect 12032 22380 12038 22392
rect 12158 22380 12164 22392
rect 12216 22380 12222 22432
rect 12710 22380 12716 22432
rect 12768 22380 12774 22432
rect 12986 22380 12992 22432
rect 13044 22420 13050 22432
rect 13354 22420 13360 22432
rect 13044 22392 13360 22420
rect 13044 22380 13050 22392
rect 13354 22380 13360 22392
rect 13412 22380 13418 22432
rect 14366 22380 14372 22432
rect 14424 22420 14430 22432
rect 15470 22420 15476 22432
rect 14424 22392 15476 22420
rect 14424 22380 14430 22392
rect 15470 22380 15476 22392
rect 15528 22380 15534 22432
rect 16206 22380 16212 22432
rect 16264 22380 16270 22432
rect 16390 22380 16396 22432
rect 16448 22420 16454 22432
rect 16485 22423 16543 22429
rect 16485 22420 16497 22423
rect 16448 22392 16497 22420
rect 16448 22380 16454 22392
rect 16485 22389 16497 22392
rect 16531 22389 16543 22423
rect 16485 22383 16543 22389
rect 17770 22380 17776 22432
rect 17828 22380 17834 22432
rect 19518 22380 19524 22432
rect 19576 22420 19582 22432
rect 19812 22429 19840 22528
rect 19886 22516 19892 22568
rect 19944 22516 19950 22568
rect 19978 22516 19984 22568
rect 20036 22556 20042 22568
rect 20824 22556 20852 22587
rect 20036 22528 20852 22556
rect 20036 22516 20042 22528
rect 20898 22516 20904 22568
rect 20956 22556 20962 22568
rect 21100 22556 21128 22596
rect 21174 22584 21180 22636
rect 21232 22624 21238 22636
rect 21821 22627 21879 22633
rect 21821 22624 21833 22627
rect 21232 22596 21833 22624
rect 21232 22584 21238 22596
rect 21821 22593 21833 22596
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 22097 22627 22155 22633
rect 22097 22593 22109 22627
rect 22143 22624 22155 22627
rect 22370 22624 22376 22636
rect 22143 22596 22376 22624
rect 22143 22593 22155 22596
rect 22097 22587 22155 22593
rect 22370 22584 22376 22596
rect 22428 22584 22434 22636
rect 22738 22584 22744 22636
rect 22796 22624 22802 22636
rect 22833 22627 22891 22633
rect 22833 22624 22845 22627
rect 22796 22596 22845 22624
rect 22796 22584 22802 22596
rect 22833 22593 22845 22596
rect 22879 22593 22891 22627
rect 22833 22587 22891 22593
rect 25038 22584 25044 22636
rect 25096 22584 25102 22636
rect 25222 22584 25228 22636
rect 25280 22584 25286 22636
rect 27614 22584 27620 22636
rect 27672 22584 27678 22636
rect 27801 22627 27859 22633
rect 27801 22593 27813 22627
rect 27847 22624 27859 22627
rect 27982 22624 27988 22636
rect 27847 22596 27988 22624
rect 27847 22593 27859 22596
rect 27801 22587 27859 22593
rect 27982 22584 27988 22596
rect 28040 22584 28046 22636
rect 29733 22627 29791 22633
rect 29733 22593 29745 22627
rect 29779 22624 29791 22627
rect 29822 22624 29828 22636
rect 29779 22596 29828 22624
rect 29779 22593 29791 22596
rect 29733 22587 29791 22593
rect 29822 22584 29828 22596
rect 29880 22584 29886 22636
rect 29917 22627 29975 22633
rect 29917 22593 29929 22627
rect 29963 22593 29975 22627
rect 29917 22587 29975 22593
rect 20956 22528 21036 22556
rect 21100 22528 21220 22556
rect 20956 22516 20962 22528
rect 21008 22488 21036 22528
rect 20548 22460 21036 22488
rect 21192 22488 21220 22528
rect 21634 22516 21640 22568
rect 21692 22556 21698 22568
rect 21913 22559 21971 22565
rect 21913 22556 21925 22559
rect 21692 22528 21925 22556
rect 21692 22516 21698 22528
rect 21913 22525 21925 22528
rect 21959 22525 21971 22559
rect 21913 22519 21971 22525
rect 22554 22488 22560 22500
rect 21192 22460 22560 22488
rect 19613 22423 19671 22429
rect 19613 22420 19625 22423
rect 19576 22392 19625 22420
rect 19576 22380 19582 22392
rect 19613 22389 19625 22392
rect 19659 22389 19671 22423
rect 19613 22383 19671 22389
rect 19797 22423 19855 22429
rect 19797 22389 19809 22423
rect 19843 22389 19855 22423
rect 19797 22383 19855 22389
rect 20254 22380 20260 22432
rect 20312 22380 20318 22432
rect 20441 22423 20499 22429
rect 20441 22389 20453 22423
rect 20487 22420 20499 22423
rect 20548 22420 20576 22460
rect 22554 22448 22560 22460
rect 22612 22448 22618 22500
rect 20487 22392 20576 22420
rect 20487 22389 20499 22392
rect 20441 22383 20499 22389
rect 20898 22380 20904 22432
rect 20956 22380 20962 22432
rect 21266 22380 21272 22432
rect 21324 22420 21330 22432
rect 21821 22423 21879 22429
rect 21821 22420 21833 22423
rect 21324 22392 21833 22420
rect 21324 22380 21330 22392
rect 21821 22389 21833 22392
rect 21867 22389 21879 22423
rect 21821 22383 21879 22389
rect 22278 22380 22284 22432
rect 22336 22380 22342 22432
rect 23014 22380 23020 22432
rect 23072 22380 23078 22432
rect 27798 22380 27804 22432
rect 27856 22380 27862 22432
rect 27985 22423 28043 22429
rect 27985 22389 27997 22423
rect 28031 22420 28043 22423
rect 29822 22420 29828 22432
rect 28031 22392 29828 22420
rect 28031 22389 28043 22392
rect 27985 22383 28043 22389
rect 29822 22380 29828 22392
rect 29880 22380 29886 22432
rect 29932 22420 29960 22587
rect 30098 22584 30104 22636
rect 30156 22584 30162 22636
rect 30208 22624 30236 22664
rect 30622 22661 30634 22664
rect 30668 22661 30680 22695
rect 30622 22655 30680 22661
rect 30926 22624 30932 22636
rect 30208 22596 30932 22624
rect 30926 22584 30932 22596
rect 30984 22584 30990 22636
rect 32214 22584 32220 22636
rect 32272 22584 32278 22636
rect 30374 22516 30380 22568
rect 30432 22516 30438 22568
rect 31018 22420 31024 22432
rect 29932 22392 31024 22420
rect 31018 22380 31024 22392
rect 31076 22380 31082 22432
rect 31754 22380 31760 22432
rect 31812 22380 31818 22432
rect 32401 22423 32459 22429
rect 32401 22389 32413 22423
rect 32447 22420 32459 22423
rect 32490 22420 32496 22432
rect 32447 22392 32496 22420
rect 32447 22389 32459 22392
rect 32401 22383 32459 22389
rect 32490 22380 32496 22392
rect 32548 22380 32554 22432
rect 1104 22330 32844 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 32844 22330
rect 1104 22256 32844 22278
rect 2222 22176 2228 22228
rect 2280 22176 2286 22228
rect 4430 22176 4436 22228
rect 4488 22216 4494 22228
rect 4488 22188 4936 22216
rect 4488 22176 4494 22188
rect 3142 22108 3148 22160
rect 3200 22148 3206 22160
rect 4341 22151 4399 22157
rect 3200 22120 4200 22148
rect 3200 22108 3206 22120
rect 3234 22080 3240 22092
rect 2516 22052 3240 22080
rect 2038 21972 2044 22024
rect 2096 21972 2102 22024
rect 2516 22021 2544 22052
rect 2501 22015 2559 22021
rect 2501 21981 2513 22015
rect 2547 21981 2559 22015
rect 2501 21975 2559 21981
rect 2593 22015 2651 22021
rect 2593 21981 2605 22015
rect 2639 22012 2651 22015
rect 2682 22012 2688 22024
rect 2639 21984 2688 22012
rect 2639 21981 2651 21984
rect 2593 21975 2651 21981
rect 2682 21972 2688 21984
rect 2740 21972 2746 22024
rect 2884 22021 2912 22052
rect 3234 22040 3240 22052
rect 3292 22080 3298 22092
rect 4172 22089 4200 22120
rect 4341 22117 4353 22151
rect 4387 22148 4399 22151
rect 4706 22148 4712 22160
rect 4387 22120 4712 22148
rect 4387 22117 4399 22120
rect 4341 22111 4399 22117
rect 4706 22108 4712 22120
rect 4764 22108 4770 22160
rect 4065 22083 4123 22089
rect 4065 22080 4077 22083
rect 3292 22052 4077 22080
rect 3292 22040 3298 22052
rect 4065 22049 4077 22052
rect 4111 22049 4123 22083
rect 4065 22043 4123 22049
rect 4157 22083 4215 22089
rect 4157 22049 4169 22083
rect 4203 22049 4215 22083
rect 4157 22043 4215 22049
rect 2869 22015 2927 22021
rect 2869 21981 2881 22015
rect 2915 21981 2927 22015
rect 2869 21975 2927 21981
rect 3326 21972 3332 22024
rect 3384 21972 3390 22024
rect 3421 22015 3479 22021
rect 3421 21981 3433 22015
rect 3467 21981 3479 22015
rect 3421 21975 3479 21981
rect 3436 21944 3464 21975
rect 3878 21972 3884 22024
rect 3936 21972 3942 22024
rect 3970 21972 3976 22024
rect 4028 21972 4034 22024
rect 4522 21972 4528 22024
rect 4580 22008 4586 22024
rect 4617 22015 4675 22021
rect 4617 22008 4629 22015
rect 4580 21981 4629 22008
rect 4663 21981 4675 22015
rect 4580 21980 4675 21981
rect 4580 21972 4586 21980
rect 4617 21975 4675 21980
rect 4709 22015 4767 22021
rect 4709 21981 4721 22015
rect 4755 21981 4767 22015
rect 4908 22012 4936 22188
rect 4982 22176 4988 22228
rect 5040 22216 5046 22228
rect 5534 22216 5540 22228
rect 5040 22188 5540 22216
rect 5040 22176 5046 22188
rect 5534 22176 5540 22188
rect 5592 22176 5598 22228
rect 5629 22219 5687 22225
rect 5629 22185 5641 22219
rect 5675 22216 5687 22219
rect 5718 22216 5724 22228
rect 5675 22188 5724 22216
rect 5675 22185 5687 22188
rect 5629 22179 5687 22185
rect 5718 22176 5724 22188
rect 5776 22216 5782 22228
rect 7834 22216 7840 22228
rect 5776 22188 7840 22216
rect 5776 22176 5782 22188
rect 7834 22176 7840 22188
rect 7892 22176 7898 22228
rect 8481 22219 8539 22225
rect 8481 22185 8493 22219
rect 8527 22216 8539 22219
rect 8662 22216 8668 22228
rect 8527 22188 8668 22216
rect 8527 22185 8539 22188
rect 8481 22179 8539 22185
rect 8662 22176 8668 22188
rect 8720 22176 8726 22228
rect 9398 22176 9404 22228
rect 9456 22216 9462 22228
rect 12710 22216 12716 22228
rect 9456 22188 12716 22216
rect 9456 22176 9462 22188
rect 12710 22176 12716 22188
rect 12768 22176 12774 22228
rect 12802 22176 12808 22228
rect 12860 22216 12866 22228
rect 13357 22219 13415 22225
rect 13357 22216 13369 22219
rect 12860 22188 13369 22216
rect 12860 22176 12866 22188
rect 13357 22185 13369 22188
rect 13403 22185 13415 22219
rect 13357 22179 13415 22185
rect 13722 22176 13728 22228
rect 13780 22216 13786 22228
rect 18966 22216 18972 22228
rect 13780 22188 18972 22216
rect 13780 22176 13786 22188
rect 18966 22176 18972 22188
rect 19024 22176 19030 22228
rect 20162 22176 20168 22228
rect 20220 22216 20226 22228
rect 21085 22219 21143 22225
rect 21085 22216 21097 22219
rect 20220 22188 21097 22216
rect 20220 22176 20226 22188
rect 21085 22185 21097 22188
rect 21131 22216 21143 22219
rect 21174 22216 21180 22228
rect 21131 22188 21180 22216
rect 21131 22185 21143 22188
rect 21085 22179 21143 22185
rect 21174 22176 21180 22188
rect 21232 22176 21238 22228
rect 22002 22176 22008 22228
rect 22060 22216 22066 22228
rect 22097 22219 22155 22225
rect 22097 22216 22109 22219
rect 22060 22188 22109 22216
rect 22060 22176 22066 22188
rect 22097 22185 22109 22188
rect 22143 22185 22155 22219
rect 22097 22179 22155 22185
rect 22646 22176 22652 22228
rect 22704 22216 22710 22228
rect 22925 22219 22983 22225
rect 22925 22216 22937 22219
rect 22704 22188 22937 22216
rect 22704 22176 22710 22188
rect 22925 22185 22937 22188
rect 22971 22216 22983 22219
rect 23014 22216 23020 22228
rect 22971 22188 23020 22216
rect 22971 22185 22983 22188
rect 22925 22179 22983 22185
rect 23014 22176 23020 22188
rect 23072 22176 23078 22228
rect 24029 22219 24087 22225
rect 24029 22185 24041 22219
rect 24075 22216 24087 22219
rect 24946 22216 24952 22228
rect 24075 22188 24952 22216
rect 24075 22185 24087 22188
rect 24029 22179 24087 22185
rect 24946 22176 24952 22188
rect 25004 22176 25010 22228
rect 25777 22219 25835 22225
rect 25777 22185 25789 22219
rect 25823 22185 25835 22219
rect 25777 22179 25835 22185
rect 5902 22108 5908 22160
rect 5960 22108 5966 22160
rect 6914 22108 6920 22160
rect 6972 22148 6978 22160
rect 8680 22148 8708 22176
rect 8846 22148 8852 22160
rect 6972 22120 8340 22148
rect 8680 22120 8852 22148
rect 6972 22108 6978 22120
rect 5368 22052 7144 22080
rect 4985 22015 5043 22021
rect 4985 22012 4997 22015
rect 4908 21984 4997 22012
rect 4709 21975 4767 21981
rect 4985 21981 4997 21984
rect 5031 21981 5043 22015
rect 4985 21975 5043 21981
rect 3344 21916 3464 21944
rect 3344 21888 3372 21916
rect 3786 21904 3792 21956
rect 3844 21944 3850 21956
rect 4724 21944 4752 21975
rect 3844 21916 4752 21944
rect 3844 21904 3850 21916
rect 2314 21836 2320 21888
rect 2372 21836 2378 21888
rect 2777 21879 2835 21885
rect 2777 21845 2789 21879
rect 2823 21876 2835 21879
rect 2958 21876 2964 21888
rect 2823 21848 2964 21876
rect 2823 21845 2835 21848
rect 2777 21839 2835 21845
rect 2958 21836 2964 21848
rect 3016 21836 3022 21888
rect 3050 21836 3056 21888
rect 3108 21836 3114 21888
rect 3142 21836 3148 21888
rect 3200 21836 3206 21888
rect 3326 21836 3332 21888
rect 3384 21836 3390 21888
rect 3418 21836 3424 21888
rect 3476 21876 3482 21888
rect 3605 21879 3663 21885
rect 3605 21876 3617 21879
rect 3476 21848 3617 21876
rect 3476 21836 3482 21848
rect 3605 21845 3617 21848
rect 3651 21845 3663 21879
rect 3605 21839 3663 21845
rect 3694 21836 3700 21888
rect 3752 21876 3758 21888
rect 4433 21879 4491 21885
rect 4433 21876 4445 21879
rect 3752 21848 4445 21876
rect 3752 21836 3758 21848
rect 4433 21845 4445 21848
rect 4479 21845 4491 21879
rect 4433 21839 4491 21845
rect 4522 21836 4528 21888
rect 4580 21876 4586 21888
rect 4893 21879 4951 21885
rect 4893 21876 4905 21879
rect 4580 21848 4905 21876
rect 4580 21836 4586 21848
rect 4893 21845 4905 21848
rect 4939 21845 4951 21879
rect 4893 21839 4951 21845
rect 5169 21879 5227 21885
rect 5169 21845 5181 21879
rect 5215 21876 5227 21879
rect 5258 21876 5264 21888
rect 5215 21848 5264 21876
rect 5215 21845 5227 21848
rect 5169 21839 5227 21845
rect 5258 21836 5264 21848
rect 5316 21876 5322 21888
rect 5368 21876 5396 22052
rect 5445 22015 5503 22021
rect 5445 21981 5457 22015
rect 5491 21981 5503 22015
rect 5445 21975 5503 21981
rect 5460 21944 5488 21975
rect 5626 21972 5632 22024
rect 5684 22012 5690 22024
rect 5721 22015 5779 22021
rect 5721 22012 5733 22015
rect 5684 21984 5733 22012
rect 5684 21972 5690 21984
rect 5721 21981 5733 21984
rect 5767 21981 5779 22015
rect 5721 21975 5779 21981
rect 5994 21972 6000 22024
rect 6052 21972 6058 22024
rect 6822 21972 6828 22024
rect 6880 21972 6886 22024
rect 7116 22021 7144 22052
rect 7101 22015 7159 22021
rect 7101 21981 7113 22015
rect 7147 21981 7159 22015
rect 7101 21975 7159 21981
rect 7190 21972 7196 22024
rect 7248 21972 7254 22024
rect 8312 22021 8340 22120
rect 8846 22108 8852 22120
rect 8904 22108 8910 22160
rect 9585 22151 9643 22157
rect 9585 22117 9597 22151
rect 9631 22148 9643 22151
rect 10134 22148 10140 22160
rect 9631 22120 10140 22148
rect 9631 22117 9643 22120
rect 9585 22111 9643 22117
rect 10134 22108 10140 22120
rect 10192 22148 10198 22160
rect 10192 22120 12112 22148
rect 10192 22108 10198 22120
rect 8864 22080 8892 22108
rect 8864 22052 9168 22080
rect 8297 22015 8355 22021
rect 8297 21981 8309 22015
rect 8343 21981 8355 22015
rect 8297 21975 8355 21981
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 22012 8631 22015
rect 8662 22012 8668 22024
rect 8619 21984 8668 22012
rect 8619 21981 8631 21984
rect 8573 21975 8631 21981
rect 8662 21972 8668 21984
rect 8720 21972 8726 22024
rect 8938 21972 8944 22024
rect 8996 21972 9002 22024
rect 9140 22021 9168 22052
rect 11146 22040 11152 22092
rect 11204 22040 11210 22092
rect 11974 22040 11980 22092
rect 12032 22040 12038 22092
rect 12084 22080 12112 22120
rect 12986 22108 12992 22160
rect 13044 22148 13050 22160
rect 13740 22148 13768 22176
rect 13044 22120 13768 22148
rect 13044 22108 13050 22120
rect 17126 22108 17132 22160
rect 17184 22108 17190 22160
rect 19705 22151 19763 22157
rect 19705 22148 19717 22151
rect 18984 22120 19717 22148
rect 15381 22083 15439 22089
rect 12084 22052 15240 22080
rect 11885 22031 11943 22037
rect 11885 22024 11897 22031
rect 11931 22024 11943 22031
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 21981 9183 22015
rect 9125 21975 9183 21981
rect 9401 22015 9459 22021
rect 9401 21981 9413 22015
rect 9447 22012 9459 22015
rect 9582 22012 9588 22024
rect 9447 21984 9588 22012
rect 9447 21981 9459 21984
rect 9401 21975 9459 21981
rect 9582 21972 9588 21984
rect 9640 21972 9646 22024
rect 9674 21972 9680 22024
rect 9732 22012 9738 22024
rect 9858 22012 9864 22024
rect 9732 21984 9864 22012
rect 9732 21972 9738 21984
rect 9858 21972 9864 21984
rect 9916 21972 9922 22024
rect 9950 21972 9956 22024
rect 10008 22012 10014 22024
rect 10229 22015 10287 22021
rect 10008 21984 10088 22012
rect 10008 21972 10014 21984
rect 5902 21944 5908 21956
rect 5460 21916 5908 21944
rect 5902 21904 5908 21916
rect 5960 21904 5966 21956
rect 6086 21904 6092 21956
rect 6144 21944 6150 21956
rect 7009 21947 7067 21953
rect 7009 21944 7021 21947
rect 6144 21916 7021 21944
rect 6144 21904 6150 21916
rect 7009 21913 7021 21916
rect 7055 21913 7067 21947
rect 7009 21907 7067 21913
rect 9214 21904 9220 21956
rect 9272 21944 9278 21956
rect 10060 21953 10088 21984
rect 10229 21981 10241 22015
rect 10275 22012 10287 22015
rect 10870 22012 10876 22024
rect 10275 21984 10876 22012
rect 10275 21981 10287 21984
rect 10229 21975 10287 21981
rect 10870 21972 10876 21984
rect 10928 21972 10934 22024
rect 11606 21972 11612 22024
rect 11664 21972 11670 22024
rect 11882 21972 11888 22024
rect 11940 21972 11946 22024
rect 12158 21972 12164 22024
rect 12216 22012 12222 22024
rect 12253 22015 12311 22021
rect 12253 22012 12265 22015
rect 12216 21984 12265 22012
rect 12216 21972 12222 21984
rect 12253 21981 12265 21984
rect 12299 21981 12311 22015
rect 12253 21975 12311 21981
rect 12618 21972 12624 22024
rect 12676 22012 12682 22024
rect 13541 22015 13599 22021
rect 13541 22012 13553 22015
rect 12676 21984 13553 22012
rect 12676 21972 12682 21984
rect 13541 21981 13553 21984
rect 13587 21981 13599 22015
rect 13541 21975 13599 21981
rect 13630 21972 13636 22024
rect 13688 22012 13694 22024
rect 14274 22012 14280 22024
rect 13688 21984 14280 22012
rect 13688 21972 13694 21984
rect 14274 21972 14280 21984
rect 14332 21972 14338 22024
rect 15212 22021 15240 22052
rect 15381 22049 15393 22083
rect 15427 22080 15439 22083
rect 15746 22080 15752 22092
rect 15427 22052 15752 22080
rect 15427 22049 15439 22052
rect 15381 22043 15439 22049
rect 15746 22040 15752 22052
rect 15804 22080 15810 22092
rect 18782 22080 18788 22092
rect 15804 22052 18788 22080
rect 15804 22040 15810 22052
rect 18782 22040 18788 22052
rect 18840 22040 18846 22092
rect 15197 22015 15255 22021
rect 15197 21981 15209 22015
rect 15243 21981 15255 22015
rect 15197 21975 15255 21981
rect 15654 21972 15660 22024
rect 15712 22012 15718 22024
rect 16945 22015 17003 22021
rect 16945 22012 16957 22015
rect 15712 21984 16957 22012
rect 15712 21972 15718 21984
rect 16945 21981 16957 21984
rect 16991 21981 17003 22015
rect 16945 21975 17003 21981
rect 17497 22015 17555 22021
rect 17497 21981 17509 22015
rect 17543 22012 17555 22015
rect 17678 22012 17684 22024
rect 17543 21984 17684 22012
rect 17543 21981 17555 21984
rect 17497 21975 17555 21981
rect 17678 21972 17684 21984
rect 17736 21972 17742 22024
rect 18984 22021 19012 22120
rect 19705 22117 19717 22120
rect 19751 22117 19763 22151
rect 19705 22111 19763 22117
rect 19610 22080 19616 22092
rect 19306 22052 19616 22080
rect 17773 22015 17831 22021
rect 17773 21981 17785 22015
rect 17819 21981 17831 22015
rect 17773 21975 17831 21981
rect 18969 22015 19027 22021
rect 18969 21981 18981 22015
rect 19015 21981 19027 22015
rect 18969 21975 19027 21981
rect 10045 21947 10103 21953
rect 9272 21916 9996 21944
rect 9272 21904 9278 21916
rect 5316 21848 5396 21876
rect 5316 21836 5322 21848
rect 6178 21836 6184 21888
rect 6236 21836 6242 21888
rect 7377 21879 7435 21885
rect 7377 21845 7389 21879
rect 7423 21876 7435 21879
rect 8662 21876 8668 21888
rect 7423 21848 8668 21876
rect 7423 21845 7435 21848
rect 7377 21839 7435 21845
rect 8662 21836 8668 21848
rect 8720 21836 8726 21888
rect 8757 21879 8815 21885
rect 8757 21845 8769 21879
rect 8803 21876 8815 21879
rect 9306 21876 9312 21888
rect 8803 21848 9312 21876
rect 8803 21845 8815 21848
rect 8757 21839 8815 21845
rect 9306 21836 9312 21848
rect 9364 21836 9370 21888
rect 9858 21836 9864 21888
rect 9916 21836 9922 21888
rect 9968 21876 9996 21916
rect 10045 21913 10057 21947
rect 10091 21944 10103 21947
rect 10686 21944 10692 21956
rect 10091 21916 10692 21944
rect 10091 21913 10103 21916
rect 10045 21907 10103 21913
rect 10686 21904 10692 21916
rect 10744 21904 10750 21956
rect 10962 21904 10968 21956
rect 11020 21944 11026 21956
rect 11425 21947 11483 21953
rect 11020 21916 11376 21944
rect 11020 21904 11026 21916
rect 10502 21876 10508 21888
rect 9968 21848 10508 21876
rect 10502 21836 10508 21848
rect 10560 21836 10566 21888
rect 11238 21836 11244 21888
rect 11296 21836 11302 21888
rect 11348 21876 11376 21916
rect 11425 21913 11437 21947
rect 11471 21944 11483 21947
rect 12342 21944 12348 21956
rect 11471 21916 12348 21944
rect 11471 21913 11483 21916
rect 11425 21907 11483 21913
rect 12342 21904 12348 21916
rect 12400 21904 12406 21956
rect 13170 21904 13176 21956
rect 13228 21944 13234 21956
rect 13357 21947 13415 21953
rect 13357 21944 13369 21947
rect 13228 21916 13369 21944
rect 13228 21904 13234 21916
rect 13357 21913 13369 21916
rect 13403 21913 13415 21947
rect 13357 21907 13415 21913
rect 13464 21916 13952 21944
rect 11514 21876 11520 21888
rect 11348 21848 11520 21876
rect 11514 21836 11520 21848
rect 11572 21876 11578 21888
rect 11701 21879 11759 21885
rect 11701 21876 11713 21879
rect 11572 21848 11713 21876
rect 11572 21836 11578 21848
rect 11701 21845 11713 21848
rect 11747 21845 11759 21879
rect 11701 21839 11759 21845
rect 12158 21836 12164 21888
rect 12216 21876 12222 21888
rect 13464 21876 13492 21916
rect 12216 21848 13492 21876
rect 12216 21836 12222 21848
rect 13814 21836 13820 21888
rect 13872 21836 13878 21888
rect 13924 21876 13952 21916
rect 15010 21904 15016 21956
rect 15068 21904 15074 21956
rect 17313 21947 17371 21953
rect 17313 21913 17325 21947
rect 17359 21913 17371 21947
rect 17313 21907 17371 21913
rect 17328 21876 17356 21907
rect 17586 21904 17592 21956
rect 17644 21944 17650 21956
rect 17788 21944 17816 21975
rect 19150 21972 19156 22024
rect 19208 22012 19214 22024
rect 19306 22012 19334 22052
rect 19610 22040 19616 22052
rect 19668 22040 19674 22092
rect 19720 22080 19748 22111
rect 19978 22108 19984 22160
rect 20036 22148 20042 22160
rect 25792 22148 25820 22179
rect 29822 22176 29828 22228
rect 29880 22216 29886 22228
rect 30742 22216 30748 22228
rect 29880 22188 30748 22216
rect 29880 22176 29886 22188
rect 30742 22176 30748 22188
rect 30800 22176 30806 22228
rect 31478 22176 31484 22228
rect 31536 22176 31542 22228
rect 20036 22120 25820 22148
rect 20036 22108 20042 22120
rect 20162 22080 20168 22092
rect 19720 22052 20168 22080
rect 20162 22040 20168 22052
rect 20220 22040 20226 22092
rect 20254 22040 20260 22092
rect 20312 22080 20318 22092
rect 20714 22080 20720 22092
rect 20312 22052 20720 22080
rect 20312 22040 20318 22052
rect 20714 22040 20720 22052
rect 20772 22040 20778 22092
rect 21174 22040 21180 22092
rect 21232 22080 21238 22092
rect 21818 22080 21824 22092
rect 21232 22052 21824 22080
rect 21232 22040 21238 22052
rect 21818 22040 21824 22052
rect 21876 22080 21882 22092
rect 22741 22083 22799 22089
rect 22741 22080 22753 22083
rect 21876 22052 22753 22080
rect 21876 22040 21882 22052
rect 22741 22049 22753 22052
rect 22787 22049 22799 22083
rect 22741 22043 22799 22049
rect 25406 22040 25412 22092
rect 25464 22080 25470 22092
rect 25682 22080 25688 22092
rect 25464 22052 25688 22080
rect 25464 22040 25470 22052
rect 25682 22040 25688 22052
rect 25740 22040 25746 22092
rect 25866 22040 25872 22092
rect 25924 22040 25930 22092
rect 32493 22083 32551 22089
rect 32493 22049 32505 22083
rect 32539 22080 32551 22083
rect 32582 22080 32588 22092
rect 32539 22052 32588 22080
rect 32539 22049 32551 22052
rect 32493 22043 32551 22049
rect 32582 22040 32588 22052
rect 32640 22040 32646 22092
rect 19208 21984 19334 22012
rect 19208 21972 19214 21984
rect 19886 21972 19892 22024
rect 19944 22012 19950 22024
rect 20622 22012 20628 22024
rect 19944 21984 20628 22012
rect 19944 21972 19950 21984
rect 20622 21972 20628 21984
rect 20680 21972 20686 22024
rect 21269 22015 21327 22021
rect 21269 21981 21281 22015
rect 21315 22012 21327 22015
rect 21358 22012 21364 22024
rect 21315 21984 21364 22012
rect 21315 21981 21327 21984
rect 21269 21975 21327 21981
rect 21358 21972 21364 21984
rect 21416 21972 21422 22024
rect 22097 22015 22155 22021
rect 22097 21981 22109 22015
rect 22143 21981 22155 22015
rect 22097 21975 22155 21981
rect 17644 21916 17816 21944
rect 17644 21904 17650 21916
rect 17862 21904 17868 21956
rect 17920 21944 17926 21956
rect 20993 21947 21051 21953
rect 20993 21944 21005 21947
rect 17920 21916 21005 21944
rect 17920 21904 17926 21916
rect 20993 21913 21005 21916
rect 21039 21913 21051 21947
rect 22112 21944 22140 21975
rect 22186 21972 22192 22024
rect 22244 21972 22250 22024
rect 22278 21972 22284 22024
rect 22336 22012 22342 22024
rect 22373 22015 22431 22021
rect 22373 22012 22385 22015
rect 22336 21984 22385 22012
rect 22336 21972 22342 21984
rect 22373 21981 22385 21984
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 22554 21972 22560 22024
rect 22612 22012 22618 22024
rect 22649 22015 22707 22021
rect 22649 22012 22661 22015
rect 22612 21984 22661 22012
rect 22612 21972 22618 21984
rect 22649 21981 22661 21984
rect 22695 21981 22707 22015
rect 22649 21975 22707 21981
rect 22925 22015 22983 22021
rect 22925 21981 22937 22015
rect 22971 22012 22983 22015
rect 23198 22012 23204 22024
rect 22971 21984 23204 22012
rect 22971 21981 22983 21984
rect 22925 21975 22983 21981
rect 23198 21972 23204 21984
rect 23256 21972 23262 22024
rect 23934 21972 23940 22024
rect 23992 21972 23998 22024
rect 24029 22015 24087 22021
rect 24029 21981 24041 22015
rect 24075 22012 24087 22015
rect 25130 22012 25136 22024
rect 24075 21984 25136 22012
rect 24075 21981 24087 21984
rect 24029 21975 24087 21981
rect 25130 21972 25136 21984
rect 25188 21972 25194 22024
rect 26053 22015 26111 22021
rect 26053 21981 26065 22015
rect 26099 22012 26111 22015
rect 27062 22012 27068 22024
rect 26099 21984 27068 22012
rect 26099 21981 26111 21984
rect 26053 21975 26111 21981
rect 27062 21972 27068 21984
rect 27120 21972 27126 22024
rect 30742 21972 30748 22024
rect 30800 22012 30806 22024
rect 30929 22015 30987 22021
rect 30929 22012 30941 22015
rect 30800 21984 30941 22012
rect 30800 21972 30806 21984
rect 30929 21981 30941 21984
rect 30975 21981 30987 22015
rect 30929 21975 30987 21981
rect 31297 22015 31355 22021
rect 31297 21981 31309 22015
rect 31343 22012 31355 22015
rect 31849 22015 31907 22021
rect 31849 22012 31861 22015
rect 31343 21984 31861 22012
rect 31343 21981 31355 21984
rect 31297 21975 31355 21981
rect 31849 21981 31861 21984
rect 31895 21981 31907 22015
rect 31849 21975 31907 21981
rect 20993 21907 21051 21913
rect 21284 21916 22048 21944
rect 22112 21916 23704 21944
rect 13924 21848 17356 21876
rect 17678 21836 17684 21888
rect 17736 21836 17742 21888
rect 17770 21836 17776 21888
rect 17828 21876 17834 21888
rect 17957 21879 18015 21885
rect 17957 21876 17969 21879
rect 17828 21848 17969 21876
rect 17828 21836 17834 21848
rect 17957 21845 17969 21848
rect 18003 21876 18015 21879
rect 21284 21876 21312 21916
rect 18003 21848 21312 21876
rect 18003 21845 18015 21848
rect 17957 21839 18015 21845
rect 21358 21836 21364 21888
rect 21416 21876 21422 21888
rect 21913 21879 21971 21885
rect 21913 21876 21925 21879
rect 21416 21848 21925 21876
rect 21416 21836 21422 21848
rect 21913 21845 21925 21848
rect 21959 21845 21971 21879
rect 22020 21876 22048 21916
rect 22554 21876 22560 21888
rect 22020 21848 22560 21876
rect 21913 21839 21971 21845
rect 22554 21836 22560 21848
rect 22612 21836 22618 21888
rect 23106 21836 23112 21888
rect 23164 21836 23170 21888
rect 23676 21876 23704 21916
rect 23750 21904 23756 21956
rect 23808 21904 23814 21956
rect 24136 21916 24532 21944
rect 24136 21876 24164 21916
rect 23676 21848 24164 21876
rect 24213 21879 24271 21885
rect 24213 21845 24225 21879
rect 24259 21876 24271 21879
rect 24394 21876 24400 21888
rect 24259 21848 24400 21876
rect 24259 21845 24271 21848
rect 24213 21839 24271 21845
rect 24394 21836 24400 21848
rect 24452 21836 24458 21888
rect 24504 21876 24532 21916
rect 25682 21904 25688 21956
rect 25740 21944 25746 21956
rect 25777 21947 25835 21953
rect 25777 21944 25789 21947
rect 25740 21916 25789 21944
rect 25740 21904 25746 21916
rect 25777 21913 25789 21916
rect 25823 21913 25835 21947
rect 25777 21907 25835 21913
rect 31113 21947 31171 21953
rect 31113 21913 31125 21947
rect 31159 21913 31171 21947
rect 31113 21907 31171 21913
rect 26237 21879 26295 21885
rect 26237 21876 26249 21879
rect 24504 21848 26249 21876
rect 26237 21845 26249 21848
rect 26283 21845 26295 21879
rect 26237 21839 26295 21845
rect 30742 21836 30748 21888
rect 30800 21876 30806 21888
rect 31128 21876 31156 21907
rect 31202 21904 31208 21956
rect 31260 21904 31266 21956
rect 30800 21848 31156 21876
rect 30800 21836 30806 21848
rect 1104 21786 32844 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 32844 21786
rect 1104 21712 32844 21734
rect 2038 21632 2044 21684
rect 2096 21672 2102 21684
rect 2777 21675 2835 21681
rect 2777 21672 2789 21675
rect 2096 21644 2789 21672
rect 2096 21632 2102 21644
rect 2777 21641 2789 21644
rect 2823 21641 2835 21675
rect 2777 21635 2835 21641
rect 2958 21632 2964 21684
rect 3016 21672 3022 21684
rect 3329 21675 3387 21681
rect 3329 21672 3341 21675
rect 3016 21644 3341 21672
rect 3016 21632 3022 21644
rect 3329 21641 3341 21644
rect 3375 21672 3387 21675
rect 3697 21675 3755 21681
rect 3375 21644 3648 21672
rect 3375 21641 3387 21644
rect 3329 21635 3387 21641
rect 2314 21564 2320 21616
rect 2372 21604 2378 21616
rect 3145 21607 3203 21613
rect 3145 21604 3157 21607
rect 2372 21576 3157 21604
rect 2372 21564 2378 21576
rect 3145 21573 3157 21576
rect 3191 21573 3203 21607
rect 3145 21567 3203 21573
rect 3237 21607 3295 21613
rect 3237 21573 3249 21607
rect 3283 21604 3295 21607
rect 3510 21604 3516 21616
rect 3283 21576 3516 21604
rect 3283 21573 3295 21576
rect 3237 21567 3295 21573
rect 3510 21564 3516 21576
rect 3568 21564 3574 21616
rect 3620 21613 3648 21644
rect 3697 21641 3709 21675
rect 3743 21672 3755 21675
rect 3786 21672 3792 21684
rect 3743 21644 3792 21672
rect 3743 21641 3755 21644
rect 3697 21635 3755 21641
rect 3786 21632 3792 21644
rect 3844 21632 3850 21684
rect 4430 21632 4436 21684
rect 4488 21672 4494 21684
rect 4525 21675 4583 21681
rect 4525 21672 4537 21675
rect 4488 21644 4537 21672
rect 4488 21632 4494 21644
rect 4525 21641 4537 21644
rect 4571 21672 4583 21675
rect 5626 21672 5632 21684
rect 4571 21644 5632 21672
rect 4571 21641 4583 21644
rect 4525 21635 4583 21641
rect 5626 21632 5632 21644
rect 5684 21632 5690 21684
rect 5905 21675 5963 21681
rect 5905 21672 5917 21675
rect 5736 21644 5917 21672
rect 3605 21607 3663 21613
rect 3605 21573 3617 21607
rect 3651 21573 3663 21607
rect 3605 21567 3663 21573
rect 3970 21564 3976 21616
rect 4028 21564 4034 21616
rect 5736 21604 5764 21644
rect 5905 21641 5917 21644
rect 5951 21672 5963 21675
rect 6822 21672 6828 21684
rect 5951 21644 6828 21672
rect 5951 21641 5963 21644
rect 5905 21635 5963 21641
rect 6822 21632 6828 21644
rect 6880 21632 6886 21684
rect 7837 21675 7895 21681
rect 7837 21641 7849 21675
rect 7883 21672 7895 21675
rect 7926 21672 7932 21684
rect 7883 21644 7932 21672
rect 7883 21641 7895 21644
rect 7837 21635 7895 21641
rect 7926 21632 7932 21644
rect 7984 21632 7990 21684
rect 9217 21675 9275 21681
rect 9217 21641 9229 21675
rect 9263 21672 9275 21675
rect 11054 21672 11060 21684
rect 9263 21644 11060 21672
rect 9263 21641 9275 21644
rect 9217 21635 9275 21641
rect 4172 21576 4752 21604
rect 1394 21496 1400 21548
rect 1452 21496 1458 21548
rect 1486 21496 1492 21548
rect 1544 21536 1550 21548
rect 1653 21539 1711 21545
rect 1653 21536 1665 21539
rect 1544 21508 1665 21536
rect 1544 21496 1550 21508
rect 1653 21505 1665 21508
rect 1699 21505 1711 21539
rect 1653 21499 1711 21505
rect 2961 21539 3019 21545
rect 2961 21505 2973 21539
rect 3007 21536 3019 21539
rect 3988 21536 4016 21564
rect 3007 21508 4016 21536
rect 3007 21505 3019 21508
rect 2961 21499 3019 21505
rect 2406 21360 2412 21412
rect 2464 21400 2470 21412
rect 2976 21400 3004 21499
rect 4062 21496 4068 21548
rect 4120 21496 4126 21548
rect 3050 21428 3056 21480
rect 3108 21468 3114 21480
rect 3881 21471 3939 21477
rect 3881 21468 3893 21471
rect 3108 21440 3893 21468
rect 3108 21428 3114 21440
rect 3881 21437 3893 21440
rect 3927 21437 3939 21471
rect 3881 21431 3939 21437
rect 3970 21428 3976 21480
rect 4028 21468 4034 21480
rect 4172 21468 4200 21576
rect 4338 21496 4344 21548
rect 4396 21496 4402 21548
rect 4617 21539 4675 21545
rect 4617 21505 4629 21539
rect 4663 21505 4675 21539
rect 4617 21499 4675 21505
rect 4028 21440 4200 21468
rect 4028 21428 4034 21440
rect 4632 21400 4660 21499
rect 4724 21468 4752 21576
rect 5368 21576 5764 21604
rect 5077 21539 5135 21545
rect 5077 21505 5089 21539
rect 5123 21536 5135 21539
rect 5258 21536 5264 21548
rect 5123 21508 5264 21536
rect 5123 21505 5135 21508
rect 5077 21499 5135 21505
rect 5258 21496 5264 21508
rect 5316 21496 5322 21548
rect 5368 21545 5396 21576
rect 6730 21564 6736 21616
rect 6788 21564 6794 21616
rect 8018 21604 8024 21616
rect 6840 21576 8024 21604
rect 5353 21539 5411 21545
rect 5353 21505 5365 21539
rect 5399 21505 5411 21539
rect 5353 21499 5411 21505
rect 5445 21539 5503 21545
rect 5445 21505 5457 21539
rect 5491 21505 5503 21539
rect 5445 21499 5503 21505
rect 5460 21468 5488 21499
rect 5718 21496 5724 21548
rect 5776 21496 5782 21548
rect 5997 21539 6055 21545
rect 5997 21505 6009 21539
rect 6043 21505 6055 21539
rect 5997 21499 6055 21505
rect 4724 21440 5488 21468
rect 5534 21428 5540 21480
rect 5592 21428 5598 21480
rect 6012 21468 6040 21499
rect 6454 21496 6460 21548
rect 6512 21536 6518 21548
rect 6840 21545 6868 21576
rect 8018 21564 8024 21576
rect 8076 21564 8082 21616
rect 9674 21604 9680 21616
rect 9048 21576 9680 21604
rect 6549 21539 6607 21545
rect 6549 21536 6561 21539
rect 6512 21508 6561 21536
rect 6512 21496 6518 21508
rect 6549 21505 6561 21508
rect 6595 21505 6607 21539
rect 6549 21499 6607 21505
rect 6825 21539 6883 21545
rect 6825 21505 6837 21539
rect 6871 21505 6883 21539
rect 6825 21499 6883 21505
rect 6917 21539 6975 21545
rect 6917 21505 6929 21539
rect 6963 21536 6975 21539
rect 7006 21536 7012 21548
rect 6963 21508 7012 21536
rect 6963 21505 6975 21508
rect 6917 21499 6975 21505
rect 7006 21496 7012 21508
rect 7064 21536 7070 21548
rect 7193 21539 7251 21545
rect 7193 21536 7205 21539
rect 7064 21508 7205 21536
rect 7064 21496 7070 21508
rect 7193 21505 7205 21508
rect 7239 21505 7251 21539
rect 7193 21499 7251 21505
rect 7377 21539 7435 21545
rect 7377 21505 7389 21539
rect 7423 21536 7435 21539
rect 7558 21536 7564 21548
rect 7423 21508 7564 21536
rect 7423 21505 7435 21508
rect 7377 21499 7435 21505
rect 7558 21496 7564 21508
rect 7616 21496 7622 21548
rect 7653 21539 7711 21545
rect 7653 21505 7665 21539
rect 7699 21505 7711 21539
rect 7653 21499 7711 21505
rect 5644 21440 6040 21468
rect 2464 21372 3004 21400
rect 3436 21372 4660 21400
rect 4893 21403 4951 21409
rect 2464 21360 2470 21372
rect 658 21292 664 21344
rect 716 21332 722 21344
rect 1762 21332 1768 21344
rect 716 21304 1768 21332
rect 716 21292 722 21304
rect 1762 21292 1768 21304
rect 1820 21292 1826 21344
rect 2682 21292 2688 21344
rect 2740 21332 2746 21344
rect 3436 21332 3464 21372
rect 4893 21369 4905 21403
rect 4939 21400 4951 21403
rect 5074 21400 5080 21412
rect 4939 21372 5080 21400
rect 4939 21369 4951 21372
rect 4893 21363 4951 21369
rect 5074 21360 5080 21372
rect 5132 21400 5138 21412
rect 5552 21400 5580 21428
rect 5132 21372 5580 21400
rect 5132 21360 5138 21372
rect 2740 21304 3464 21332
rect 2740 21292 2746 21304
rect 3510 21292 3516 21344
rect 3568 21292 3574 21344
rect 3602 21292 3608 21344
rect 3660 21332 3666 21344
rect 3789 21335 3847 21341
rect 3789 21332 3801 21335
rect 3660 21304 3801 21332
rect 3660 21292 3666 21304
rect 3789 21301 3801 21304
rect 3835 21332 3847 21335
rect 4062 21332 4068 21344
rect 3835 21304 4068 21332
rect 3835 21301 3847 21304
rect 3789 21295 3847 21301
rect 4062 21292 4068 21304
rect 4120 21292 4126 21344
rect 4246 21292 4252 21344
rect 4304 21292 4310 21344
rect 4706 21292 4712 21344
rect 4764 21332 4770 21344
rect 4801 21335 4859 21341
rect 4801 21332 4813 21335
rect 4764 21304 4813 21332
rect 4764 21292 4770 21304
rect 4801 21301 4813 21304
rect 4847 21301 4859 21335
rect 4801 21295 4859 21301
rect 5169 21335 5227 21341
rect 5169 21301 5181 21335
rect 5215 21332 5227 21335
rect 5350 21332 5356 21344
rect 5215 21304 5356 21332
rect 5215 21301 5227 21304
rect 5169 21295 5227 21301
rect 5350 21292 5356 21304
rect 5408 21292 5414 21344
rect 5442 21292 5448 21344
rect 5500 21332 5506 21344
rect 5644 21341 5672 21440
rect 6730 21428 6736 21480
rect 6788 21468 6794 21480
rect 7668 21468 7696 21499
rect 7834 21496 7840 21548
rect 7892 21536 7898 21548
rect 9048 21545 9076 21576
rect 9674 21564 9680 21576
rect 9732 21564 9738 21616
rect 10244 21613 10272 21644
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 11698 21632 11704 21684
rect 11756 21672 11762 21684
rect 13262 21672 13268 21684
rect 11756 21644 13268 21672
rect 11756 21632 11762 21644
rect 13262 21632 13268 21644
rect 13320 21632 13326 21684
rect 13541 21675 13599 21681
rect 13541 21641 13553 21675
rect 13587 21672 13599 21675
rect 13814 21672 13820 21684
rect 13587 21644 13820 21672
rect 13587 21641 13599 21644
rect 13541 21635 13599 21641
rect 13814 21632 13820 21644
rect 13872 21632 13878 21684
rect 17221 21675 17279 21681
rect 17221 21641 17233 21675
rect 17267 21672 17279 21675
rect 19153 21675 19211 21681
rect 17267 21644 19104 21672
rect 17267 21641 17279 21644
rect 17221 21635 17279 21641
rect 10229 21607 10287 21613
rect 10229 21573 10241 21607
rect 10275 21573 10287 21607
rect 10229 21567 10287 21573
rect 10502 21564 10508 21616
rect 10560 21604 10566 21616
rect 16761 21607 16819 21613
rect 16761 21604 16773 21607
rect 10560 21576 14872 21604
rect 10560 21564 10566 21576
rect 7929 21539 7987 21545
rect 7929 21536 7941 21539
rect 7892 21508 7941 21536
rect 7892 21496 7898 21508
rect 7929 21505 7941 21508
rect 7975 21505 7987 21539
rect 7929 21499 7987 21505
rect 9033 21539 9091 21545
rect 9033 21505 9045 21539
rect 9079 21505 9091 21539
rect 9033 21499 9091 21505
rect 9306 21496 9312 21548
rect 9364 21496 9370 21548
rect 9493 21539 9551 21545
rect 9493 21505 9505 21539
rect 9539 21536 9551 21539
rect 9582 21536 9588 21548
rect 9539 21508 9588 21536
rect 9539 21505 9551 21508
rect 9493 21499 9551 21505
rect 9582 21496 9588 21508
rect 9640 21496 9646 21548
rect 9953 21539 10011 21545
rect 9953 21505 9965 21539
rect 9999 21536 10011 21539
rect 10686 21536 10692 21548
rect 9999 21508 10692 21536
rect 9999 21505 10011 21508
rect 9953 21499 10011 21505
rect 10686 21496 10692 21508
rect 10744 21496 10750 21548
rect 10781 21539 10839 21545
rect 10781 21505 10793 21539
rect 10827 21505 10839 21539
rect 10781 21499 10839 21505
rect 8570 21468 8576 21480
rect 6788 21440 8576 21468
rect 6788 21428 6794 21440
rect 8570 21428 8576 21440
rect 8628 21428 8634 21480
rect 9677 21471 9735 21477
rect 9677 21437 9689 21471
rect 9723 21468 9735 21471
rect 10137 21471 10195 21477
rect 10137 21468 10149 21471
rect 9723 21440 10149 21468
rect 9723 21437 9735 21440
rect 9677 21431 9735 21437
rect 10137 21437 10149 21440
rect 10183 21437 10195 21471
rect 10137 21431 10195 21437
rect 5718 21360 5724 21412
rect 5776 21400 5782 21412
rect 8754 21400 8760 21412
rect 5776 21372 8760 21400
rect 5776 21360 5782 21372
rect 8754 21360 8760 21372
rect 8812 21360 8818 21412
rect 9490 21360 9496 21412
rect 9548 21400 9554 21412
rect 9769 21403 9827 21409
rect 9769 21400 9781 21403
rect 9548 21372 9781 21400
rect 9548 21360 9554 21372
rect 9769 21369 9781 21372
rect 9815 21369 9827 21403
rect 10152 21400 10180 21431
rect 10410 21428 10416 21480
rect 10468 21468 10474 21480
rect 10796 21468 10824 21499
rect 10962 21496 10968 21548
rect 11020 21496 11026 21548
rect 11149 21539 11207 21545
rect 11149 21505 11161 21539
rect 11195 21536 11207 21539
rect 11606 21536 11612 21548
rect 11195 21508 11612 21536
rect 11195 21505 11207 21508
rect 11149 21499 11207 21505
rect 11606 21496 11612 21508
rect 11664 21496 11670 21548
rect 11701 21539 11759 21545
rect 11701 21505 11713 21539
rect 11747 21536 11759 21539
rect 11790 21536 11796 21548
rect 11747 21508 11796 21536
rect 11747 21505 11759 21508
rect 11701 21499 11759 21505
rect 11790 21496 11796 21508
rect 11848 21496 11854 21548
rect 11885 21539 11943 21545
rect 11885 21505 11897 21539
rect 11931 21536 11943 21539
rect 12066 21536 12072 21548
rect 11931 21508 12072 21536
rect 11931 21505 11943 21508
rect 11885 21499 11943 21505
rect 12066 21496 12072 21508
rect 12124 21496 12130 21548
rect 12894 21536 12900 21548
rect 12176 21508 12900 21536
rect 12176 21468 12204 21508
rect 12894 21496 12900 21508
rect 12952 21496 12958 21548
rect 12986 21496 12992 21548
rect 13044 21496 13050 21548
rect 13081 21539 13139 21545
rect 13081 21505 13093 21539
rect 13127 21536 13139 21539
rect 13262 21536 13268 21548
rect 13127 21508 13268 21536
rect 13127 21505 13139 21508
rect 13081 21499 13139 21505
rect 13262 21496 13268 21508
rect 13320 21496 13326 21548
rect 13354 21496 13360 21548
rect 13412 21496 13418 21548
rect 14844 21545 14872 21576
rect 16132 21576 16773 21604
rect 14829 21539 14887 21545
rect 14829 21505 14841 21539
rect 14875 21536 14887 21539
rect 15470 21536 15476 21548
rect 14875 21508 15476 21536
rect 14875 21505 14887 21508
rect 14829 21499 14887 21505
rect 15470 21496 15476 21508
rect 15528 21496 15534 21548
rect 15838 21496 15844 21548
rect 15896 21536 15902 21548
rect 16132 21545 16160 21576
rect 16761 21573 16773 21576
rect 16807 21573 16819 21607
rect 17770 21604 17776 21616
rect 16761 21567 16819 21573
rect 17052 21576 17776 21604
rect 17052 21545 17080 21576
rect 17770 21564 17776 21576
rect 17828 21564 17834 21616
rect 18782 21564 18788 21616
rect 18840 21604 18846 21616
rect 18840 21576 19012 21604
rect 18840 21564 18846 21576
rect 16117 21539 16175 21545
rect 16117 21536 16129 21539
rect 15896 21508 16129 21536
rect 15896 21496 15902 21508
rect 16117 21505 16129 21508
rect 16163 21505 16175 21539
rect 16301 21539 16359 21545
rect 16301 21536 16313 21539
rect 16117 21499 16175 21505
rect 16224 21508 16313 21536
rect 10468 21440 10824 21468
rect 10888 21440 12204 21468
rect 10468 21428 10474 21440
rect 10888 21400 10916 21440
rect 12618 21428 12624 21480
rect 12676 21468 12682 21480
rect 12713 21471 12771 21477
rect 12713 21468 12725 21471
rect 12676 21440 12725 21468
rect 12676 21428 12682 21440
rect 12713 21437 12725 21440
rect 12759 21437 12771 21471
rect 12713 21431 12771 21437
rect 13173 21471 13231 21477
rect 13173 21437 13185 21471
rect 13219 21437 13231 21471
rect 13173 21431 13231 21437
rect 10152 21372 10916 21400
rect 9769 21363 9827 21369
rect 11422 21360 11428 21412
rect 11480 21400 11486 21412
rect 11480 21372 11919 21400
rect 11480 21360 11486 21372
rect 5629 21335 5687 21341
rect 5629 21332 5641 21335
rect 5500 21304 5641 21332
rect 5500 21292 5506 21304
rect 5629 21301 5641 21304
rect 5675 21301 5687 21335
rect 5629 21295 5687 21301
rect 6181 21335 6239 21341
rect 6181 21301 6193 21335
rect 6227 21332 6239 21335
rect 6362 21332 6368 21344
rect 6227 21304 6368 21332
rect 6227 21301 6239 21304
rect 6181 21295 6239 21301
rect 6362 21292 6368 21304
rect 6420 21292 6426 21344
rect 7101 21335 7159 21341
rect 7101 21301 7113 21335
rect 7147 21332 7159 21335
rect 7282 21332 7288 21344
rect 7147 21304 7288 21332
rect 7147 21301 7159 21304
rect 7101 21295 7159 21301
rect 7282 21292 7288 21304
rect 7340 21292 7346 21344
rect 7558 21292 7564 21344
rect 7616 21332 7622 21344
rect 8018 21332 8024 21344
rect 7616 21304 8024 21332
rect 7616 21292 7622 21304
rect 8018 21292 8024 21304
rect 8076 21332 8082 21344
rect 8113 21335 8171 21341
rect 8113 21332 8125 21335
rect 8076 21304 8125 21332
rect 8076 21292 8082 21304
rect 8113 21301 8125 21304
rect 8159 21301 8171 21335
rect 8113 21295 8171 21301
rect 8202 21292 8208 21344
rect 8260 21332 8266 21344
rect 9674 21332 9680 21344
rect 8260 21304 9680 21332
rect 8260 21292 8266 21304
rect 9674 21292 9680 21304
rect 9732 21292 9738 21344
rect 9858 21292 9864 21344
rect 9916 21332 9922 21344
rect 10226 21332 10232 21344
rect 9916 21304 10232 21332
rect 9916 21292 9922 21304
rect 10226 21292 10232 21304
rect 10284 21292 10290 21344
rect 11333 21335 11391 21341
rect 11333 21301 11345 21335
rect 11379 21332 11391 21335
rect 11790 21332 11796 21344
rect 11379 21304 11796 21332
rect 11379 21301 11391 21304
rect 11333 21295 11391 21301
rect 11790 21292 11796 21304
rect 11848 21292 11854 21344
rect 11891 21332 11919 21372
rect 11974 21360 11980 21412
rect 12032 21400 12038 21412
rect 12069 21403 12127 21409
rect 12069 21400 12081 21403
rect 12032 21372 12081 21400
rect 12032 21360 12038 21372
rect 12069 21369 12081 21372
rect 12115 21400 12127 21403
rect 13188 21400 13216 21431
rect 13722 21428 13728 21480
rect 13780 21468 13786 21480
rect 15194 21468 15200 21480
rect 13780 21440 15200 21468
rect 13780 21428 13786 21440
rect 15194 21428 15200 21440
rect 15252 21428 15258 21480
rect 14918 21400 14924 21412
rect 12115 21372 13216 21400
rect 13287 21372 14924 21400
rect 12115 21369 12127 21372
rect 12069 21363 12127 21369
rect 12710 21332 12716 21344
rect 11891 21304 12716 21332
rect 12710 21292 12716 21304
rect 12768 21292 12774 21344
rect 13170 21292 13176 21344
rect 13228 21332 13234 21344
rect 13287 21332 13315 21372
rect 14918 21360 14924 21372
rect 14976 21400 14982 21412
rect 16224 21400 16252 21508
rect 16301 21505 16313 21508
rect 16347 21505 16359 21539
rect 16301 21499 16359 21505
rect 17037 21539 17095 21545
rect 17037 21505 17049 21539
rect 17083 21505 17095 21539
rect 17037 21499 17095 21505
rect 17402 21496 17408 21548
rect 17460 21536 17466 21548
rect 17589 21539 17647 21545
rect 17589 21536 17601 21539
rect 17460 21508 17601 21536
rect 17460 21496 17466 21508
rect 17589 21505 17601 21508
rect 17635 21505 17647 21539
rect 17589 21499 17647 21505
rect 17865 21539 17923 21545
rect 17865 21505 17877 21539
rect 17911 21505 17923 21539
rect 17865 21499 17923 21505
rect 17957 21539 18015 21545
rect 17957 21505 17969 21539
rect 18003 21536 18015 21539
rect 18046 21536 18052 21548
rect 18003 21508 18052 21536
rect 18003 21505 18015 21508
rect 17957 21499 18015 21505
rect 16945 21471 17003 21477
rect 16945 21437 16957 21471
rect 16991 21468 17003 21471
rect 17126 21468 17132 21480
rect 16991 21440 17132 21468
rect 16991 21437 17003 21440
rect 16945 21431 17003 21437
rect 17126 21428 17132 21440
rect 17184 21428 17190 21480
rect 17770 21428 17776 21480
rect 17828 21428 17834 21480
rect 17880 21468 17908 21499
rect 18046 21496 18052 21508
rect 18104 21496 18110 21548
rect 18230 21496 18236 21548
rect 18288 21496 18294 21548
rect 18506 21496 18512 21548
rect 18564 21536 18570 21548
rect 18984 21545 19012 21576
rect 18693 21539 18751 21545
rect 18693 21536 18705 21539
rect 18564 21508 18705 21536
rect 18564 21496 18570 21508
rect 18693 21505 18705 21508
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 18969 21539 19027 21545
rect 18969 21505 18981 21539
rect 19015 21505 19027 21539
rect 19076 21536 19104 21644
rect 19153 21641 19165 21675
rect 19199 21672 19211 21675
rect 19334 21672 19340 21684
rect 19199 21644 19340 21672
rect 19199 21641 19211 21644
rect 19153 21635 19211 21641
rect 19334 21632 19340 21644
rect 19392 21632 19398 21684
rect 19705 21675 19763 21681
rect 19705 21641 19717 21675
rect 19751 21672 19763 21675
rect 19794 21672 19800 21684
rect 19751 21644 19800 21672
rect 19751 21641 19763 21644
rect 19705 21635 19763 21641
rect 19794 21632 19800 21644
rect 19852 21632 19858 21684
rect 20346 21672 20352 21684
rect 20180 21644 20352 21672
rect 19150 21536 19156 21548
rect 19076 21508 19156 21536
rect 18969 21499 19027 21505
rect 19150 21496 19156 21508
rect 19208 21496 19214 21548
rect 19242 21496 19248 21548
rect 19300 21496 19306 21548
rect 19334 21496 19340 21548
rect 19392 21536 19398 21548
rect 19518 21536 19524 21548
rect 19392 21508 19524 21536
rect 19392 21496 19398 21508
rect 19518 21496 19524 21508
rect 19576 21496 19582 21548
rect 19886 21496 19892 21548
rect 19944 21536 19950 21548
rect 19981 21539 20039 21545
rect 19981 21536 19993 21539
rect 19944 21508 19993 21536
rect 19944 21496 19950 21508
rect 19981 21505 19993 21508
rect 20027 21505 20039 21539
rect 19981 21499 20039 21505
rect 20073 21539 20131 21545
rect 20073 21505 20085 21539
rect 20119 21536 20131 21539
rect 20180 21536 20208 21644
rect 20346 21632 20352 21644
rect 20404 21632 20410 21684
rect 23842 21632 23848 21684
rect 23900 21672 23906 21684
rect 23900 21644 24532 21672
rect 23900 21632 23906 21644
rect 20254 21564 20260 21616
rect 20312 21604 20318 21616
rect 20625 21607 20683 21613
rect 20625 21604 20637 21607
rect 20312 21576 20637 21604
rect 20312 21564 20318 21576
rect 20625 21573 20637 21576
rect 20671 21573 20683 21607
rect 20806 21604 20812 21616
rect 20625 21567 20683 21573
rect 20732 21576 20812 21604
rect 20119 21508 20208 21536
rect 20349 21540 20407 21545
rect 20349 21539 20484 21540
rect 20119 21505 20131 21508
rect 20073 21499 20131 21505
rect 20349 21505 20361 21539
rect 20395 21536 20484 21539
rect 20732 21536 20760 21576
rect 20806 21564 20812 21576
rect 20864 21564 20870 21616
rect 23106 21564 23112 21616
rect 23164 21604 23170 21616
rect 24504 21613 24532 21644
rect 27614 21632 27620 21684
rect 27672 21632 27678 21684
rect 27798 21632 27804 21684
rect 27856 21672 27862 21684
rect 27982 21672 27988 21684
rect 27856 21644 27988 21672
rect 27856 21632 27862 21644
rect 27982 21632 27988 21644
rect 28040 21632 28046 21684
rect 28629 21675 28687 21681
rect 28629 21672 28641 21675
rect 28092 21644 28641 21672
rect 28092 21613 28120 21644
rect 28629 21641 28641 21644
rect 28675 21641 28687 21675
rect 28629 21635 28687 21641
rect 29181 21675 29239 21681
rect 29181 21641 29193 21675
rect 29227 21672 29239 21675
rect 29546 21672 29552 21684
rect 29227 21644 29552 21672
rect 29227 21641 29239 21644
rect 29181 21635 29239 21641
rect 29546 21632 29552 21644
rect 29604 21632 29610 21684
rect 31941 21675 31999 21681
rect 31941 21641 31953 21675
rect 31987 21672 31999 21675
rect 32214 21672 32220 21684
rect 31987 21644 32220 21672
rect 31987 21641 31999 21644
rect 31941 21635 31999 21641
rect 32214 21632 32220 21644
rect 32272 21632 32278 21684
rect 23937 21607 23995 21613
rect 23937 21604 23949 21607
rect 23164 21576 23949 21604
rect 23164 21564 23170 21576
rect 23937 21573 23949 21576
rect 23983 21573 23995 21607
rect 23937 21567 23995 21573
rect 24489 21607 24547 21613
rect 24489 21573 24501 21607
rect 24535 21573 24547 21607
rect 28077 21607 28135 21613
rect 24489 21567 24547 21573
rect 26988 21576 27936 21604
rect 26988 21548 27016 21576
rect 20901 21539 20959 21545
rect 20901 21536 20913 21539
rect 20395 21512 20760 21536
rect 20395 21505 20407 21512
rect 20456 21508 20760 21512
rect 20824 21508 20913 21536
rect 20349 21499 20407 21505
rect 18414 21468 18420 21480
rect 17880 21440 18420 21468
rect 18414 21428 18420 21440
rect 18472 21428 18478 21480
rect 18785 21471 18843 21477
rect 18785 21437 18797 21471
rect 18831 21437 18843 21471
rect 18785 21431 18843 21437
rect 14976 21372 16252 21400
rect 16485 21403 16543 21409
rect 14976 21360 14982 21372
rect 16485 21369 16497 21403
rect 16531 21400 16543 21403
rect 18800 21400 18828 21431
rect 19426 21428 19432 21480
rect 19484 21428 19490 21480
rect 20165 21471 20223 21477
rect 20165 21468 20177 21471
rect 19904 21440 20177 21468
rect 19904 21412 19932 21440
rect 20165 21437 20177 21440
rect 20211 21437 20223 21471
rect 20165 21431 20223 21437
rect 20714 21428 20720 21480
rect 20772 21428 20778 21480
rect 16531 21372 18828 21400
rect 18984 21372 19840 21400
rect 16531 21369 16543 21372
rect 16485 21363 16543 21369
rect 13228 21304 13315 21332
rect 13357 21335 13415 21341
rect 13228 21292 13234 21304
rect 13357 21301 13369 21335
rect 13403 21332 13415 21335
rect 13630 21332 13636 21344
rect 13403 21304 13636 21332
rect 13403 21301 13415 21304
rect 13357 21295 13415 21301
rect 13630 21292 13636 21304
rect 13688 21332 13694 21344
rect 14274 21332 14280 21344
rect 13688 21304 14280 21332
rect 13688 21292 13694 21304
rect 14274 21292 14280 21304
rect 14332 21292 14338 21344
rect 14645 21335 14703 21341
rect 14645 21301 14657 21335
rect 14691 21332 14703 21335
rect 14734 21332 14740 21344
rect 14691 21304 14740 21332
rect 14691 21301 14703 21304
rect 14645 21295 14703 21301
rect 14734 21292 14740 21304
rect 14792 21292 14798 21344
rect 16850 21292 16856 21344
rect 16908 21292 16914 21344
rect 17402 21292 17408 21344
rect 17460 21292 17466 21344
rect 17678 21292 17684 21344
rect 17736 21292 17742 21344
rect 17770 21292 17776 21344
rect 17828 21332 17834 21344
rect 18138 21332 18144 21344
rect 17828 21304 18144 21332
rect 17828 21292 17834 21304
rect 18138 21292 18144 21304
rect 18196 21292 18202 21344
rect 18414 21292 18420 21344
rect 18472 21292 18478 21344
rect 18984 21341 19012 21372
rect 19812 21344 19840 21372
rect 19886 21360 19892 21412
rect 19944 21360 19950 21412
rect 20533 21403 20591 21409
rect 20533 21369 20545 21403
rect 20579 21400 20591 21403
rect 20824 21400 20852 21508
rect 20901 21505 20913 21508
rect 20947 21505 20959 21539
rect 20901 21499 20959 21505
rect 21174 21496 21180 21548
rect 21232 21536 21238 21548
rect 24213 21539 24271 21545
rect 24213 21536 24225 21539
rect 21232 21508 24225 21536
rect 21232 21496 21238 21508
rect 24213 21505 24225 21508
rect 24259 21505 24271 21539
rect 24213 21499 24271 21505
rect 24762 21496 24768 21548
rect 24820 21496 24826 21548
rect 26970 21496 26976 21548
rect 27028 21496 27034 21548
rect 27246 21496 27252 21548
rect 27304 21496 27310 21548
rect 27522 21496 27528 21548
rect 27580 21536 27586 21548
rect 27801 21539 27859 21545
rect 27801 21536 27813 21539
rect 27580 21508 27813 21536
rect 27580 21496 27586 21508
rect 27801 21505 27813 21508
rect 27847 21505 27859 21539
rect 27908 21536 27936 21576
rect 28077 21573 28089 21607
rect 28123 21573 28135 21607
rect 28077 21567 28135 21573
rect 30374 21564 30380 21616
rect 30432 21604 30438 21616
rect 31110 21604 31116 21616
rect 30432 21576 31116 21604
rect 30432 21564 30438 21576
rect 28169 21539 28227 21545
rect 28169 21536 28181 21539
rect 27908 21508 28181 21536
rect 27801 21499 27859 21505
rect 28169 21505 28181 21508
rect 28215 21505 28227 21539
rect 28169 21499 28227 21505
rect 28350 21496 28356 21548
rect 28408 21536 28414 21548
rect 28445 21539 28503 21545
rect 28445 21536 28457 21539
rect 28408 21508 28457 21536
rect 28408 21496 28414 21508
rect 28445 21505 28457 21508
rect 28491 21536 28503 21539
rect 28626 21536 28632 21548
rect 28491 21508 28632 21536
rect 28491 21505 28503 21508
rect 28445 21499 28503 21505
rect 28626 21496 28632 21508
rect 28684 21496 28690 21548
rect 28721 21539 28779 21545
rect 28721 21505 28733 21539
rect 28767 21505 28779 21539
rect 28721 21499 28779 21505
rect 28997 21539 29055 21545
rect 28997 21505 29009 21539
rect 29043 21536 29055 21539
rect 30282 21536 30288 21548
rect 29043 21508 30288 21536
rect 29043 21505 29055 21508
rect 28997 21499 29055 21505
rect 23474 21428 23480 21480
rect 23532 21428 23538 21480
rect 24026 21428 24032 21480
rect 24084 21428 24090 21480
rect 24673 21471 24731 21477
rect 24673 21468 24685 21471
rect 24136 21440 24685 21468
rect 20579 21372 20852 21400
rect 23492 21400 23520 21428
rect 24136 21400 24164 21440
rect 24673 21437 24685 21440
rect 24719 21437 24731 21471
rect 24673 21431 24731 21437
rect 26510 21428 26516 21480
rect 26568 21468 26574 21480
rect 27065 21471 27123 21477
rect 27065 21468 27077 21471
rect 26568 21440 27077 21468
rect 26568 21428 26574 21440
rect 27065 21437 27077 21440
rect 27111 21437 27123 21471
rect 27065 21431 27123 21437
rect 27614 21428 27620 21480
rect 27672 21468 27678 21480
rect 27893 21471 27951 21477
rect 27893 21468 27905 21471
rect 27672 21440 27905 21468
rect 27672 21428 27678 21440
rect 27893 21437 27905 21440
rect 27939 21437 27951 21471
rect 27893 21431 27951 21437
rect 27982 21428 27988 21480
rect 28040 21468 28046 21480
rect 28261 21471 28319 21477
rect 28261 21468 28273 21471
rect 28040 21440 28273 21468
rect 28040 21428 28046 21440
rect 28261 21437 28273 21440
rect 28307 21437 28319 21471
rect 28261 21431 28319 21437
rect 23492 21372 24164 21400
rect 20579 21369 20591 21372
rect 20533 21363 20591 21369
rect 24578 21360 24584 21412
rect 24636 21400 24642 21412
rect 24949 21403 25007 21409
rect 24949 21400 24961 21403
rect 24636 21372 24961 21400
rect 24636 21360 24642 21372
rect 24949 21369 24961 21372
rect 24995 21400 25007 21403
rect 28736 21400 28764 21499
rect 30282 21496 30288 21508
rect 30340 21496 30346 21548
rect 30576 21545 30604 21576
rect 31110 21564 31116 21576
rect 31168 21564 31174 21616
rect 30561 21539 30619 21545
rect 30561 21505 30573 21539
rect 30607 21505 30619 21539
rect 30561 21499 30619 21505
rect 30828 21539 30886 21545
rect 30828 21505 30840 21539
rect 30874 21536 30886 21539
rect 31294 21536 31300 21548
rect 30874 21508 31300 21536
rect 30874 21505 30886 21508
rect 30828 21499 30886 21505
rect 31294 21496 31300 21508
rect 31352 21496 31358 21548
rect 32122 21496 32128 21548
rect 32180 21536 32186 21548
rect 32217 21539 32275 21545
rect 32217 21536 32229 21539
rect 32180 21508 32229 21536
rect 32180 21496 32186 21508
rect 32217 21505 32229 21508
rect 32263 21505 32275 21539
rect 32217 21499 32275 21505
rect 28810 21428 28816 21480
rect 28868 21428 28874 21480
rect 24995 21372 28764 21400
rect 24995 21369 25007 21372
rect 24949 21363 25007 21369
rect 18969 21335 19027 21341
rect 18969 21301 18981 21335
rect 19015 21301 19027 21335
rect 18969 21295 19027 21301
rect 19518 21292 19524 21344
rect 19576 21292 19582 21344
rect 19794 21292 19800 21344
rect 19852 21292 19858 21344
rect 20254 21292 20260 21344
rect 20312 21292 20318 21344
rect 20806 21292 20812 21344
rect 20864 21292 20870 21344
rect 21085 21335 21143 21341
rect 21085 21301 21097 21335
rect 21131 21332 21143 21335
rect 23474 21332 23480 21344
rect 21131 21304 23480 21332
rect 21131 21301 21143 21304
rect 21085 21295 21143 21301
rect 23474 21292 23480 21304
rect 23532 21292 23538 21344
rect 23842 21292 23848 21344
rect 23900 21292 23906 21344
rect 24213 21335 24271 21341
rect 24213 21301 24225 21335
rect 24259 21332 24271 21335
rect 24302 21332 24308 21344
rect 24259 21304 24308 21332
rect 24259 21301 24271 21304
rect 24213 21295 24271 21301
rect 24302 21292 24308 21304
rect 24360 21292 24366 21344
rect 24394 21292 24400 21344
rect 24452 21292 24458 21344
rect 24486 21292 24492 21344
rect 24544 21292 24550 21344
rect 25498 21292 25504 21344
rect 25556 21332 25562 21344
rect 25866 21332 25872 21344
rect 25556 21304 25872 21332
rect 25556 21292 25562 21304
rect 25866 21292 25872 21304
rect 25924 21292 25930 21344
rect 26602 21292 26608 21344
rect 26660 21332 26666 21344
rect 26973 21335 27031 21341
rect 26973 21332 26985 21335
rect 26660 21304 26985 21332
rect 26660 21292 26666 21304
rect 26973 21301 26985 21304
rect 27019 21301 27031 21335
rect 26973 21295 27031 21301
rect 27154 21292 27160 21344
rect 27212 21332 27218 21344
rect 27433 21335 27491 21341
rect 27433 21332 27445 21335
rect 27212 21304 27445 21332
rect 27212 21292 27218 21304
rect 27433 21301 27445 21304
rect 27479 21301 27491 21335
rect 27433 21295 27491 21301
rect 28077 21335 28135 21341
rect 28077 21301 28089 21335
rect 28123 21332 28135 21335
rect 28166 21332 28172 21344
rect 28123 21304 28172 21332
rect 28123 21301 28135 21304
rect 28077 21295 28135 21301
rect 28166 21292 28172 21304
rect 28224 21292 28230 21344
rect 28258 21292 28264 21344
rect 28316 21292 28322 21344
rect 28718 21292 28724 21344
rect 28776 21292 28782 21344
rect 32398 21292 32404 21344
rect 32456 21292 32462 21344
rect 1104 21242 32844 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 32844 21242
rect 1104 21168 32844 21190
rect 2222 21088 2228 21140
rect 2280 21088 2286 21140
rect 2501 21131 2559 21137
rect 2501 21097 2513 21131
rect 2547 21128 2559 21131
rect 3234 21128 3240 21140
rect 2547 21100 3240 21128
rect 2547 21097 2559 21100
rect 2501 21091 2559 21097
rect 3234 21088 3240 21100
rect 3292 21128 3298 21140
rect 4430 21128 4436 21140
rect 3292 21100 4436 21128
rect 3292 21088 3298 21100
rect 4430 21088 4436 21100
rect 4488 21088 4494 21140
rect 4525 21131 4583 21137
rect 4525 21097 4537 21131
rect 4571 21128 4583 21131
rect 4890 21128 4896 21140
rect 4571 21100 4896 21128
rect 4571 21097 4583 21100
rect 4525 21091 4583 21097
rect 4890 21088 4896 21100
rect 4948 21088 4954 21140
rect 4982 21088 4988 21140
rect 5040 21128 5046 21140
rect 5994 21128 6000 21140
rect 5040 21100 6000 21128
rect 5040 21088 5046 21100
rect 5994 21088 6000 21100
rect 6052 21088 6058 21140
rect 6086 21088 6092 21140
rect 6144 21128 6150 21140
rect 6144 21100 8616 21128
rect 6144 21088 6150 21100
rect 1762 21020 1768 21072
rect 1820 21060 1826 21072
rect 1949 21063 2007 21069
rect 1949 21060 1961 21063
rect 1820 21032 1961 21060
rect 1820 21020 1826 21032
rect 1949 21029 1961 21032
rect 1995 21060 2007 21063
rect 2406 21060 2412 21072
rect 1995 21032 2412 21060
rect 1995 21029 2007 21032
rect 1949 21023 2007 21029
rect 2406 21020 2412 21032
rect 2464 21020 2470 21072
rect 2590 21020 2596 21072
rect 2648 21060 2654 21072
rect 2685 21063 2743 21069
rect 2685 21060 2697 21063
rect 2648 21032 2697 21060
rect 2648 21020 2654 21032
rect 2685 21029 2697 21032
rect 2731 21029 2743 21063
rect 2685 21023 2743 21029
rect 3142 21020 3148 21072
rect 3200 21060 3206 21072
rect 4338 21060 4344 21072
rect 3200 21032 4344 21060
rect 3200 21020 3206 21032
rect 4338 21020 4344 21032
rect 4396 21060 4402 21072
rect 5534 21060 5540 21072
rect 4396 21032 5540 21060
rect 4396 21020 4402 21032
rect 5534 21020 5540 21032
rect 5592 21020 5598 21072
rect 5629 21063 5687 21069
rect 5629 21029 5641 21063
rect 5675 21060 5687 21063
rect 6454 21060 6460 21072
rect 5675 21032 6460 21060
rect 5675 21029 5687 21032
rect 5629 21023 5687 21029
rect 3602 20992 3608 21004
rect 1504 20964 3608 20992
rect 1504 20933 1532 20964
rect 3602 20952 3608 20964
rect 3660 20952 3666 21004
rect 4982 20992 4988 21004
rect 4080 20964 4988 20992
rect 1489 20927 1547 20933
rect 1489 20893 1501 20927
rect 1535 20893 1547 20927
rect 1489 20887 1547 20893
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20893 1823 20927
rect 1765 20887 1823 20893
rect 1780 20856 1808 20887
rect 2038 20884 2044 20936
rect 2096 20884 2102 20936
rect 2222 20884 2228 20936
rect 2280 20924 2286 20936
rect 2317 20927 2375 20933
rect 2317 20924 2329 20927
rect 2280 20896 2329 20924
rect 2280 20884 2286 20896
rect 2317 20893 2329 20896
rect 2363 20893 2375 20927
rect 2317 20887 2375 20893
rect 2406 20884 2412 20936
rect 2464 20924 2470 20936
rect 2464 20896 2728 20924
rect 2464 20884 2470 20896
rect 2700 20865 2728 20896
rect 3786 20884 3792 20936
rect 3844 20924 3850 20936
rect 3973 20927 4031 20933
rect 3973 20924 3985 20927
rect 3844 20896 3985 20924
rect 3844 20884 3850 20896
rect 3973 20893 3985 20896
rect 4019 20893 4031 20927
rect 3973 20887 4031 20893
rect 2685 20859 2743 20865
rect 1780 20828 2268 20856
rect 1670 20748 1676 20800
rect 1728 20748 1734 20800
rect 2240 20788 2268 20828
rect 2685 20825 2697 20859
rect 2731 20825 2743 20859
rect 2685 20819 2743 20825
rect 3694 20816 3700 20868
rect 3752 20856 3758 20868
rect 4080 20865 4108 20964
rect 4982 20952 4988 20964
rect 5040 20952 5046 21004
rect 5074 20952 5080 21004
rect 5132 20952 5138 21004
rect 5644 20992 5672 21023
rect 6454 21020 6460 21032
rect 6512 21020 6518 21072
rect 7282 21020 7288 21072
rect 7340 21060 7346 21072
rect 8202 21060 8208 21072
rect 7340 21032 8208 21060
rect 7340 21020 7346 21032
rect 8202 21020 8208 21032
rect 8260 21020 8266 21072
rect 8588 20992 8616 21100
rect 8662 21088 8668 21140
rect 8720 21128 8726 21140
rect 8720 21100 9168 21128
rect 8720 21088 8726 21100
rect 8757 21063 8815 21069
rect 8757 21029 8769 21063
rect 8803 21060 8815 21063
rect 8938 21060 8944 21072
rect 8803 21032 8944 21060
rect 8803 21029 8815 21032
rect 8757 21023 8815 21029
rect 8938 21020 8944 21032
rect 8996 21020 9002 21072
rect 9140 21060 9168 21100
rect 9214 21088 9220 21140
rect 9272 21128 9278 21140
rect 9953 21131 10011 21137
rect 9272 21100 9904 21128
rect 9272 21088 9278 21100
rect 9876 21060 9904 21100
rect 9953 21097 9965 21131
rect 9999 21128 10011 21131
rect 10502 21128 10508 21140
rect 9999 21100 10508 21128
rect 9999 21097 10011 21100
rect 9953 21091 10011 21097
rect 10502 21088 10508 21100
rect 10560 21088 10566 21140
rect 11238 21088 11244 21140
rect 11296 21128 11302 21140
rect 12161 21131 12219 21137
rect 12161 21128 12173 21131
rect 11296 21100 12173 21128
rect 11296 21088 11302 21100
rect 12161 21097 12173 21100
rect 12207 21097 12219 21131
rect 12161 21091 12219 21097
rect 12621 21131 12679 21137
rect 12621 21097 12633 21131
rect 12667 21128 12679 21131
rect 12710 21128 12716 21140
rect 12667 21100 12716 21128
rect 12667 21097 12679 21100
rect 12621 21091 12679 21097
rect 12710 21088 12716 21100
rect 12768 21088 12774 21140
rect 12802 21088 12808 21140
rect 12860 21088 12866 21140
rect 12986 21088 12992 21140
rect 13044 21128 13050 21140
rect 13906 21128 13912 21140
rect 13044 21100 13912 21128
rect 13044 21088 13050 21100
rect 13906 21088 13912 21100
rect 13964 21088 13970 21140
rect 14734 21088 14740 21140
rect 14792 21088 14798 21140
rect 14921 21131 14979 21137
rect 14921 21097 14933 21131
rect 14967 21128 14979 21131
rect 15930 21128 15936 21140
rect 14967 21100 15936 21128
rect 14967 21097 14979 21100
rect 14921 21091 14979 21097
rect 15930 21088 15936 21100
rect 15988 21088 15994 21140
rect 19794 21088 19800 21140
rect 19852 21128 19858 21140
rect 20254 21128 20260 21140
rect 19852 21100 20260 21128
rect 19852 21088 19858 21100
rect 20254 21088 20260 21100
rect 20312 21128 20318 21140
rect 21174 21128 21180 21140
rect 20312 21100 21180 21128
rect 20312 21088 20318 21100
rect 21174 21088 21180 21100
rect 21232 21088 21238 21140
rect 21266 21088 21272 21140
rect 21324 21128 21330 21140
rect 21542 21128 21548 21140
rect 21324 21100 21548 21128
rect 21324 21088 21330 21100
rect 21542 21088 21548 21100
rect 21600 21088 21606 21140
rect 22005 21131 22063 21137
rect 22005 21097 22017 21131
rect 22051 21128 22063 21131
rect 22186 21128 22192 21140
rect 22051 21100 22192 21128
rect 22051 21097 22063 21100
rect 22005 21091 22063 21097
rect 22186 21088 22192 21100
rect 22244 21088 22250 21140
rect 23474 21088 23480 21140
rect 23532 21128 23538 21140
rect 24854 21128 24860 21140
rect 23532 21100 24860 21128
rect 23532 21088 23538 21100
rect 24854 21088 24860 21100
rect 24912 21088 24918 21140
rect 25314 21088 25320 21140
rect 25372 21128 25378 21140
rect 25774 21128 25780 21140
rect 25372 21100 25780 21128
rect 25372 21088 25378 21100
rect 25774 21088 25780 21100
rect 25832 21088 25838 21140
rect 25869 21131 25927 21137
rect 25869 21097 25881 21131
rect 25915 21128 25927 21131
rect 26970 21128 26976 21140
rect 25915 21100 26976 21128
rect 25915 21097 25927 21100
rect 25869 21091 25927 21097
rect 10045 21063 10103 21069
rect 10045 21060 10057 21063
rect 9140 21032 9536 21060
rect 9876 21032 10057 21060
rect 9214 20992 9220 21004
rect 5184 20964 5672 20992
rect 6012 20964 8248 20992
rect 4157 20927 4215 20933
rect 4157 20893 4169 20927
rect 4203 20924 4215 20927
rect 4246 20924 4252 20936
rect 4203 20896 4252 20924
rect 4203 20893 4215 20896
rect 4157 20887 4215 20893
rect 4246 20884 4252 20896
rect 4304 20884 4310 20936
rect 4338 20884 4344 20936
rect 4396 20884 4402 20936
rect 4706 20884 4712 20936
rect 4764 20884 4770 20936
rect 4801 20927 4859 20933
rect 4801 20893 4813 20927
rect 4847 20924 4859 20927
rect 5092 20924 5120 20952
rect 5184 20933 5212 20964
rect 4847 20896 5120 20924
rect 5169 20927 5227 20933
rect 4847 20893 4859 20896
rect 4801 20887 4859 20893
rect 5169 20893 5181 20927
rect 5215 20893 5227 20927
rect 5169 20887 5227 20893
rect 5350 20884 5356 20936
rect 5408 20884 5414 20936
rect 5442 20884 5448 20936
rect 5500 20884 5506 20936
rect 5534 20884 5540 20936
rect 5592 20924 5598 20936
rect 5721 20927 5779 20933
rect 5721 20924 5733 20927
rect 5592 20896 5733 20924
rect 5592 20884 5598 20896
rect 5721 20893 5733 20896
rect 5767 20893 5779 20927
rect 6012 20924 6040 20964
rect 8220 20936 8248 20964
rect 8588 20964 9220 20992
rect 5721 20887 5779 20893
rect 5828 20896 6040 20924
rect 4065 20859 4123 20865
rect 4065 20856 4077 20859
rect 3752 20828 4077 20856
rect 3752 20816 3758 20828
rect 4065 20825 4077 20828
rect 4111 20825 4123 20859
rect 4065 20819 4123 20825
rect 4890 20816 4896 20868
rect 4948 20856 4954 20868
rect 4985 20859 5043 20865
rect 4985 20856 4997 20859
rect 4948 20828 4997 20856
rect 4948 20816 4954 20828
rect 4985 20825 4997 20828
rect 5031 20825 5043 20859
rect 4985 20819 5043 20825
rect 5077 20859 5135 20865
rect 5077 20825 5089 20859
rect 5123 20856 5135 20859
rect 5368 20856 5396 20884
rect 5828 20856 5856 20896
rect 6086 20884 6092 20936
rect 6144 20924 6150 20936
rect 6362 20924 6368 20936
rect 6144 20896 6368 20924
rect 6144 20884 6150 20896
rect 6362 20884 6368 20896
rect 6420 20884 6426 20936
rect 8202 20884 8208 20936
rect 8260 20884 8266 20936
rect 8588 20933 8616 20964
rect 9214 20952 9220 20964
rect 9272 20952 9278 21004
rect 9508 20992 9536 21032
rect 10045 21029 10057 21032
rect 10091 21029 10103 21063
rect 10045 21023 10103 21029
rect 10686 21020 10692 21072
rect 10744 21060 10750 21072
rect 10744 21032 12296 21060
rect 10744 21020 10750 21032
rect 9508 20964 10272 20992
rect 9324 20933 9444 20940
rect 10244 20933 10272 20964
rect 10410 20952 10416 21004
rect 10468 20952 10474 21004
rect 10502 20952 10508 21004
rect 10560 20992 10566 21004
rect 11698 20992 11704 21004
rect 10560 20964 11704 20992
rect 10560 20952 10566 20964
rect 11698 20952 11704 20964
rect 11756 20952 11762 21004
rect 12158 20992 12164 21004
rect 11808 20964 12164 20992
rect 8573 20927 8631 20933
rect 8573 20893 8585 20927
rect 8619 20893 8631 20927
rect 9324 20927 9459 20933
rect 9324 20924 9413 20927
rect 8573 20887 8631 20893
rect 8772 20912 9413 20924
rect 8772 20896 9352 20912
rect 8772 20868 8800 20896
rect 9401 20893 9413 20912
rect 9447 20893 9459 20927
rect 9769 20927 9827 20933
rect 9769 20924 9781 20927
rect 9401 20887 9459 20893
rect 9508 20896 9781 20924
rect 5123 20828 5856 20856
rect 5123 20825 5135 20828
rect 5077 20819 5135 20825
rect 5902 20816 5908 20868
rect 5960 20816 5966 20868
rect 5994 20816 6000 20868
rect 6052 20816 6058 20868
rect 7834 20856 7840 20868
rect 6196 20828 7840 20856
rect 2958 20788 2964 20800
rect 2240 20760 2964 20788
rect 2958 20748 2964 20760
rect 3016 20748 3022 20800
rect 3142 20748 3148 20800
rect 3200 20748 3206 20800
rect 3234 20748 3240 20800
rect 3292 20748 3298 20800
rect 3418 20748 3424 20800
rect 3476 20748 3482 20800
rect 3786 20748 3792 20800
rect 3844 20748 3850 20800
rect 5258 20748 5264 20800
rect 5316 20788 5322 20800
rect 5353 20791 5411 20797
rect 5353 20788 5365 20791
rect 5316 20760 5365 20788
rect 5316 20748 5322 20760
rect 5353 20757 5365 20760
rect 5399 20757 5411 20791
rect 5353 20751 5411 20757
rect 5718 20748 5724 20800
rect 5776 20788 5782 20800
rect 6196 20788 6224 20828
rect 7834 20816 7840 20828
rect 7892 20816 7898 20868
rect 7926 20816 7932 20868
rect 7984 20856 7990 20868
rect 8389 20859 8447 20865
rect 8389 20856 8401 20859
rect 7984 20828 8401 20856
rect 7984 20816 7990 20828
rect 8389 20825 8401 20828
rect 8435 20825 8447 20859
rect 8389 20819 8447 20825
rect 8481 20859 8539 20865
rect 8481 20825 8493 20859
rect 8527 20856 8539 20859
rect 8754 20856 8760 20868
rect 8527 20828 8760 20856
rect 8527 20825 8539 20828
rect 8481 20819 8539 20825
rect 5776 20760 6224 20788
rect 5776 20748 5782 20760
rect 6270 20748 6276 20800
rect 6328 20748 6334 20800
rect 6362 20748 6368 20800
rect 6420 20788 6426 20800
rect 7374 20788 7380 20800
rect 6420 20760 7380 20788
rect 6420 20748 6426 20760
rect 7374 20748 7380 20760
rect 7432 20748 7438 20800
rect 8404 20788 8432 20819
rect 8754 20816 8760 20828
rect 8812 20816 8818 20868
rect 9214 20816 9220 20868
rect 9272 20856 9278 20868
rect 9508 20856 9536 20896
rect 9769 20893 9781 20896
rect 9815 20893 9827 20927
rect 9769 20887 9827 20893
rect 10229 20927 10287 20933
rect 10229 20893 10241 20927
rect 10275 20924 10287 20927
rect 11808 20924 11836 20964
rect 12158 20952 12164 20964
rect 12216 20952 12222 21004
rect 12268 21001 12296 21032
rect 13354 21020 13360 21072
rect 13412 21060 13418 21072
rect 13412 21032 14686 21060
rect 13412 21020 13418 21032
rect 12253 20995 12311 21001
rect 12253 20961 12265 20995
rect 12299 20961 12311 20995
rect 12253 20955 12311 20961
rect 12618 20952 12624 21004
rect 12676 20952 12682 21004
rect 12802 20952 12808 21004
rect 12860 20992 12866 21004
rect 14550 20992 14556 21004
rect 12860 20964 14556 20992
rect 12860 20952 12866 20964
rect 14550 20952 14556 20964
rect 14608 20952 14614 21004
rect 14658 20992 14686 21032
rect 15470 21020 15476 21072
rect 15528 21060 15534 21072
rect 15528 21032 21680 21060
rect 15528 21020 15534 21032
rect 14658 20964 15792 20992
rect 10275 20896 11836 20924
rect 11974 20920 11980 20936
rect 10275 20893 10287 20896
rect 10229 20887 10287 20893
rect 11900 20892 11980 20920
rect 9272 20828 9536 20856
rect 9585 20859 9643 20865
rect 9272 20816 9278 20828
rect 9585 20825 9597 20859
rect 9631 20825 9643 20859
rect 9585 20819 9643 20825
rect 9677 20859 9735 20865
rect 9677 20825 9689 20859
rect 9723 20856 9735 20859
rect 9858 20856 9864 20868
rect 9723 20828 9864 20856
rect 9723 20825 9735 20828
rect 9677 20819 9735 20825
rect 9600 20788 9628 20819
rect 9858 20816 9864 20828
rect 9916 20816 9922 20868
rect 11900 20856 11928 20892
rect 11974 20884 11980 20892
rect 12032 20884 12038 20936
rect 12069 20927 12127 20933
rect 12069 20893 12081 20927
rect 12115 20924 12127 20927
rect 12437 20927 12495 20933
rect 12115 20896 12388 20924
rect 12115 20893 12127 20896
rect 12069 20887 12127 20893
rect 12161 20859 12219 20865
rect 12161 20856 12173 20859
rect 11900 20828 12173 20856
rect 12161 20825 12173 20828
rect 12207 20825 12219 20859
rect 12360 20856 12388 20896
rect 12437 20893 12449 20927
rect 12483 20924 12495 20927
rect 12636 20924 12664 20952
rect 12483 20896 12664 20924
rect 12483 20893 12495 20896
rect 12437 20887 12495 20893
rect 12894 20884 12900 20936
rect 12952 20884 12958 20936
rect 13081 20927 13139 20933
rect 13081 20893 13093 20927
rect 13127 20924 13139 20927
rect 13354 20924 13360 20936
rect 13127 20896 13360 20924
rect 13127 20893 13139 20896
rect 13081 20887 13139 20893
rect 13354 20884 13360 20896
rect 13412 20884 13418 20936
rect 13906 20884 13912 20936
rect 13964 20924 13970 20936
rect 14458 20924 14464 20936
rect 13964 20896 14464 20924
rect 13964 20884 13970 20896
rect 14458 20884 14464 20896
rect 14516 20884 14522 20936
rect 14642 20884 14648 20936
rect 14700 20884 14706 20936
rect 14737 20927 14795 20933
rect 14737 20893 14749 20927
rect 14783 20924 14795 20927
rect 15764 20924 15792 20964
rect 15930 20952 15936 21004
rect 15988 20992 15994 21004
rect 16482 20992 16488 21004
rect 15988 20964 16488 20992
rect 15988 20952 15994 20964
rect 16482 20952 16488 20964
rect 16540 20952 16546 21004
rect 18414 20952 18420 21004
rect 18472 20992 18478 21004
rect 18472 20964 20300 20992
rect 18472 20952 18478 20964
rect 18506 20924 18512 20936
rect 14783 20896 15700 20924
rect 15764 20896 18512 20924
rect 14783 20893 14795 20896
rect 14737 20887 14795 20893
rect 13630 20856 13636 20868
rect 12360 20828 13636 20856
rect 12161 20819 12219 20825
rect 13630 20816 13636 20828
rect 13688 20816 13694 20868
rect 13814 20816 13820 20868
rect 13872 20856 13878 20868
rect 14752 20856 14780 20887
rect 13872 20828 14780 20856
rect 15672 20856 15700 20896
rect 18506 20884 18512 20896
rect 18564 20884 18570 20936
rect 19702 20884 19708 20936
rect 19760 20924 19766 20936
rect 19760 20918 20116 20924
rect 20165 20923 20223 20929
rect 20165 20918 20177 20923
rect 19760 20896 20177 20918
rect 19760 20884 19766 20896
rect 20088 20890 20177 20896
rect 20165 20889 20177 20890
rect 20211 20889 20223 20923
rect 20272 20924 20300 20964
rect 20806 20952 20812 21004
rect 20864 20992 20870 21004
rect 21174 20992 21180 21004
rect 20864 20964 21180 20992
rect 20864 20952 20870 20964
rect 21174 20952 21180 20964
rect 21232 20952 21238 21004
rect 21652 21001 21680 21032
rect 22370 21020 22376 21072
rect 22428 21060 22434 21072
rect 24302 21060 24308 21072
rect 22428 21032 24308 21060
rect 22428 21020 22434 21032
rect 24302 21020 24308 21032
rect 24360 21020 24366 21072
rect 25884 21060 25912 21091
rect 26970 21088 26976 21100
rect 27028 21088 27034 21140
rect 27062 21088 27068 21140
rect 27120 21128 27126 21140
rect 27157 21131 27215 21137
rect 27157 21128 27169 21131
rect 27120 21100 27169 21128
rect 27120 21088 27126 21100
rect 27157 21097 27169 21100
rect 27203 21128 27215 21131
rect 27522 21128 27528 21140
rect 27203 21100 27528 21128
rect 27203 21097 27215 21100
rect 27157 21091 27215 21097
rect 27522 21088 27528 21100
rect 27580 21088 27586 21140
rect 31294 21088 31300 21140
rect 31352 21088 31358 21140
rect 25792 21032 25912 21060
rect 26237 21063 26295 21069
rect 21637 20995 21695 21001
rect 21637 20961 21649 20995
rect 21683 20961 21695 20995
rect 21637 20955 21695 20961
rect 22554 20952 22560 21004
rect 22612 20992 22618 21004
rect 25792 20992 25820 21032
rect 26237 21029 26249 21063
rect 26283 21060 26295 21063
rect 26418 21060 26424 21072
rect 26283 21032 26424 21060
rect 26283 21029 26295 21032
rect 26237 21023 26295 21029
rect 26418 21020 26424 21032
rect 26476 21020 26482 21072
rect 27430 21060 27436 21072
rect 27356 21032 27436 21060
rect 27356 21001 27384 21032
rect 27430 21020 27436 21032
rect 27488 21020 27494 21072
rect 30742 21020 30748 21072
rect 30800 21020 30806 21072
rect 30834 21020 30840 21072
rect 30892 21060 30898 21072
rect 31018 21060 31024 21072
rect 30892 21032 31024 21060
rect 30892 21020 30898 21032
rect 31018 21020 31024 21032
rect 31076 21060 31082 21072
rect 32309 21063 32367 21069
rect 32309 21060 32321 21063
rect 31076 21032 32321 21060
rect 31076 21020 31082 21032
rect 32309 21029 32321 21032
rect 32355 21029 32367 21063
rect 32309 21023 32367 21029
rect 22612 20964 25820 20992
rect 27341 20995 27399 21001
rect 22612 20952 22618 20964
rect 27341 20961 27353 20995
rect 27387 20961 27399 20995
rect 27341 20955 27399 20961
rect 30466 20952 30472 21004
rect 30524 20992 30530 21004
rect 30760 20992 30788 21020
rect 30524 20964 30972 20992
rect 30524 20952 30530 20964
rect 21821 20927 21879 20933
rect 21821 20924 21833 20927
rect 20272 20896 21833 20924
rect 20165 20883 20223 20889
rect 21821 20893 21833 20896
rect 21867 20893 21879 20927
rect 21821 20887 21879 20893
rect 23106 20884 23112 20936
rect 23164 20924 23170 20936
rect 24762 20924 24768 20936
rect 23164 20896 24768 20924
rect 23164 20884 23170 20896
rect 24762 20884 24768 20896
rect 24820 20884 24826 20936
rect 24854 20884 24860 20936
rect 24912 20924 24918 20936
rect 25593 20927 25651 20933
rect 25593 20924 25605 20927
rect 24912 20896 25605 20924
rect 24912 20884 24918 20896
rect 25593 20893 25605 20896
rect 25639 20893 25651 20927
rect 25593 20887 25651 20893
rect 25866 20884 25872 20936
rect 25924 20884 25930 20936
rect 25958 20884 25964 20936
rect 26016 20924 26022 20936
rect 26053 20927 26111 20933
rect 26053 20924 26065 20927
rect 26016 20896 26065 20924
rect 26016 20884 26022 20896
rect 26053 20893 26065 20896
rect 26099 20893 26111 20927
rect 26053 20887 26111 20893
rect 26418 20884 26424 20936
rect 26476 20924 26482 20936
rect 27157 20927 27215 20933
rect 27157 20924 27169 20927
rect 26476 20896 27169 20924
rect 26476 20884 26482 20896
rect 27157 20893 27169 20896
rect 27203 20893 27215 20927
rect 27157 20887 27215 20893
rect 27430 20884 27436 20936
rect 27488 20884 27494 20936
rect 28350 20884 28356 20936
rect 28408 20924 28414 20936
rect 28810 20924 28816 20936
rect 28408 20896 28816 20924
rect 28408 20884 28414 20896
rect 28810 20884 28816 20896
rect 28868 20884 28874 20936
rect 30742 20884 30748 20936
rect 30800 20884 30806 20936
rect 30944 20933 30972 20964
rect 32214 20952 32220 21004
rect 32272 20952 32278 21004
rect 30929 20927 30987 20933
rect 30929 20893 30941 20927
rect 30975 20893 30987 20927
rect 30929 20887 30987 20893
rect 31113 20927 31171 20933
rect 31113 20893 31125 20927
rect 31159 20924 31171 20927
rect 31573 20927 31631 20933
rect 31573 20924 31585 20927
rect 31159 20896 31585 20924
rect 31159 20893 31171 20896
rect 31113 20887 31171 20893
rect 31573 20893 31585 20896
rect 31619 20893 31631 20927
rect 31573 20887 31631 20893
rect 31846 20884 31852 20936
rect 31904 20924 31910 20936
rect 32493 20927 32551 20933
rect 32493 20924 32505 20927
rect 31904 20896 32505 20924
rect 31904 20884 31910 20896
rect 32493 20893 32505 20896
rect 32539 20893 32551 20927
rect 32493 20887 32551 20893
rect 15672 20828 20116 20856
rect 13872 20816 13878 20828
rect 8404 20760 9628 20788
rect 10226 20748 10232 20800
rect 10284 20788 10290 20800
rect 11698 20788 11704 20800
rect 10284 20760 11704 20788
rect 10284 20748 10290 20760
rect 11698 20748 11704 20760
rect 11756 20748 11762 20800
rect 12066 20748 12072 20800
rect 12124 20788 12130 20800
rect 13265 20791 13323 20797
rect 13265 20788 13277 20791
rect 12124 20760 13277 20788
rect 12124 20748 12130 20760
rect 13265 20757 13277 20760
rect 13311 20757 13323 20791
rect 13265 20751 13323 20757
rect 14182 20748 14188 20800
rect 14240 20788 14246 20800
rect 14458 20788 14464 20800
rect 14240 20760 14464 20788
rect 14240 20748 14246 20760
rect 14458 20748 14464 20760
rect 14516 20748 14522 20800
rect 15378 20748 15384 20800
rect 15436 20788 15442 20800
rect 16114 20788 16120 20800
rect 15436 20760 16120 20788
rect 15436 20748 15442 20760
rect 16114 20748 16120 20760
rect 16172 20748 16178 20800
rect 18138 20748 18144 20800
rect 18196 20788 18202 20800
rect 19426 20788 19432 20800
rect 18196 20760 19432 20788
rect 18196 20748 18202 20760
rect 19426 20748 19432 20760
rect 19484 20748 19490 20800
rect 20088 20788 20116 20828
rect 20272 20828 21496 20856
rect 20272 20788 20300 20828
rect 20088 20760 20300 20788
rect 20349 20791 20407 20797
rect 20349 20757 20361 20791
rect 20395 20788 20407 20791
rect 20438 20788 20444 20800
rect 20395 20760 20444 20788
rect 20395 20757 20407 20760
rect 20349 20751 20407 20757
rect 20438 20748 20444 20760
rect 20496 20748 20502 20800
rect 21468 20788 21496 20828
rect 21542 20816 21548 20868
rect 21600 20816 21606 20868
rect 21634 20816 21640 20868
rect 21692 20856 21698 20868
rect 28718 20856 28724 20868
rect 21692 20828 28724 20856
rect 21692 20816 21698 20828
rect 28718 20816 28724 20828
rect 28776 20816 28782 20868
rect 31018 20816 31024 20868
rect 31076 20856 31082 20868
rect 31202 20856 31208 20868
rect 31076 20828 31208 20856
rect 31076 20816 31082 20828
rect 31202 20816 31208 20828
rect 31260 20816 31266 20868
rect 24210 20788 24216 20800
rect 21468 20760 24216 20788
rect 24210 20748 24216 20760
rect 24268 20748 24274 20800
rect 26602 20748 26608 20800
rect 26660 20788 26666 20800
rect 26973 20791 27031 20797
rect 26973 20788 26985 20791
rect 26660 20760 26985 20788
rect 26660 20748 26666 20760
rect 26973 20757 26985 20760
rect 27019 20757 27031 20791
rect 26973 20751 27031 20757
rect 27617 20791 27675 20797
rect 27617 20757 27629 20791
rect 27663 20788 27675 20791
rect 30006 20788 30012 20800
rect 27663 20760 30012 20788
rect 27663 20757 27675 20760
rect 27617 20751 27675 20757
rect 30006 20748 30012 20760
rect 30064 20748 30070 20800
rect 1104 20698 32844 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 32844 20698
rect 1104 20624 32844 20646
rect 1670 20544 1676 20596
rect 1728 20584 1734 20596
rect 2409 20587 2467 20593
rect 2409 20584 2421 20587
rect 1728 20556 2421 20584
rect 1728 20544 1734 20556
rect 2409 20553 2421 20556
rect 2455 20584 2467 20587
rect 3142 20584 3148 20596
rect 2455 20556 3148 20584
rect 2455 20553 2467 20556
rect 2409 20547 2467 20553
rect 3142 20544 3148 20556
rect 3200 20544 3206 20596
rect 3234 20544 3240 20596
rect 3292 20584 3298 20596
rect 3697 20587 3755 20593
rect 3697 20584 3709 20587
rect 3292 20556 3709 20584
rect 3292 20544 3298 20556
rect 3697 20553 3709 20556
rect 3743 20553 3755 20587
rect 3697 20547 3755 20553
rect 3878 20544 3884 20596
rect 3936 20584 3942 20596
rect 5721 20587 5779 20593
rect 3936 20556 4752 20584
rect 3936 20544 3942 20556
rect 2526 20519 2584 20525
rect 2526 20485 2538 20519
rect 2572 20516 2584 20519
rect 2869 20519 2927 20525
rect 2869 20516 2881 20519
rect 2572 20488 2881 20516
rect 2572 20485 2584 20488
rect 2526 20479 2584 20485
rect 2869 20485 2881 20488
rect 2915 20485 2927 20519
rect 2869 20479 2927 20485
rect 1762 20408 1768 20460
rect 1820 20408 1826 20460
rect 2041 20451 2099 20457
rect 2041 20417 2053 20451
rect 2087 20448 2099 20451
rect 2884 20448 2912 20479
rect 3050 20476 3056 20528
rect 3108 20516 3114 20528
rect 3421 20519 3479 20525
rect 3421 20516 3433 20519
rect 3108 20488 3433 20516
rect 3108 20476 3114 20488
rect 3421 20485 3433 20488
rect 3467 20485 3479 20519
rect 3421 20479 3479 20485
rect 3510 20476 3516 20528
rect 3568 20516 3574 20528
rect 3568 20488 4016 20516
rect 3568 20476 3574 20488
rect 3234 20448 3240 20460
rect 2087 20420 2636 20448
rect 2884 20420 3240 20448
rect 2087 20417 2099 20420
rect 2041 20411 2099 20417
rect 1949 20315 2007 20321
rect 1949 20281 1961 20315
rect 1995 20312 2007 20315
rect 2056 20312 2084 20411
rect 2608 20392 2636 20420
rect 3234 20408 3240 20420
rect 3292 20408 3298 20460
rect 3988 20457 4016 20488
rect 3881 20451 3939 20457
rect 3881 20417 3893 20451
rect 3927 20417 3939 20451
rect 3881 20411 3939 20417
rect 3973 20451 4031 20457
rect 3973 20417 3985 20451
rect 4019 20417 4031 20451
rect 3973 20411 4031 20417
rect 2314 20340 2320 20392
rect 2372 20340 2378 20392
rect 2590 20340 2596 20392
rect 2648 20380 2654 20392
rect 3329 20383 3387 20389
rect 3329 20380 3341 20383
rect 2648 20352 3341 20380
rect 2648 20340 2654 20352
rect 3329 20349 3341 20352
rect 3375 20349 3387 20383
rect 3329 20343 3387 20349
rect 1995 20284 2084 20312
rect 1995 20281 2007 20284
rect 1949 20275 2007 20281
rect 2682 20272 2688 20324
rect 2740 20272 2746 20324
rect 2869 20315 2927 20321
rect 2869 20281 2881 20315
rect 2915 20312 2927 20315
rect 3142 20312 3148 20324
rect 2915 20284 3148 20312
rect 2915 20281 2927 20284
rect 2869 20275 2927 20281
rect 3142 20272 3148 20284
rect 3200 20272 3206 20324
rect 3896 20312 3924 20411
rect 4430 20408 4436 20460
rect 4488 20408 4494 20460
rect 4724 20457 4752 20556
rect 5721 20553 5733 20587
rect 5767 20584 5779 20587
rect 5767 20556 8800 20584
rect 5767 20553 5779 20556
rect 5721 20547 5779 20553
rect 4798 20476 4804 20528
rect 4856 20516 4862 20528
rect 5353 20519 5411 20525
rect 5353 20516 5365 20519
rect 4856 20488 5365 20516
rect 4856 20476 4862 20488
rect 5353 20485 5365 20488
rect 5399 20485 5411 20519
rect 6362 20516 6368 20528
rect 5353 20479 5411 20485
rect 5552 20488 6368 20516
rect 4709 20451 4767 20457
rect 4709 20417 4721 20451
rect 4755 20417 4767 20451
rect 4709 20411 4767 20417
rect 5077 20451 5135 20457
rect 5077 20417 5089 20451
rect 5123 20417 5135 20451
rect 5077 20411 5135 20417
rect 5169 20451 5227 20457
rect 5169 20417 5181 20451
rect 5215 20417 5227 20451
rect 5169 20411 5227 20417
rect 4062 20340 4068 20392
rect 4120 20380 4126 20392
rect 4120 20352 4568 20380
rect 4120 20340 4126 20352
rect 4540 20321 4568 20352
rect 4249 20315 4307 20321
rect 4249 20312 4261 20315
rect 3252 20284 4261 20312
rect 2774 20204 2780 20256
rect 2832 20244 2838 20256
rect 3252 20244 3280 20284
rect 4249 20281 4261 20284
rect 4295 20281 4307 20315
rect 4249 20275 4307 20281
rect 4525 20315 4583 20321
rect 4525 20281 4537 20315
rect 4571 20281 4583 20315
rect 5092 20312 5120 20411
rect 5184 20380 5212 20411
rect 5442 20408 5448 20460
rect 5500 20408 5506 20460
rect 5552 20457 5580 20488
rect 6362 20476 6368 20488
rect 6420 20476 6426 20528
rect 6914 20476 6920 20528
rect 6972 20516 6978 20528
rect 8113 20519 8171 20525
rect 8113 20516 8125 20519
rect 6972 20488 8125 20516
rect 6972 20476 6978 20488
rect 8113 20485 8125 20488
rect 8159 20485 8171 20519
rect 8113 20479 8171 20485
rect 5537 20451 5595 20457
rect 5537 20417 5549 20451
rect 5583 20417 5595 20451
rect 5537 20411 5595 20417
rect 5626 20408 5632 20460
rect 5684 20448 5690 20460
rect 5813 20451 5871 20457
rect 5813 20448 5825 20451
rect 5684 20420 5825 20448
rect 5684 20408 5690 20420
rect 5813 20417 5825 20420
rect 5859 20448 5871 20451
rect 7929 20451 7987 20457
rect 7929 20448 7941 20451
rect 5859 20420 7941 20448
rect 5859 20417 5871 20420
rect 5813 20411 5871 20417
rect 7929 20417 7941 20420
rect 7975 20417 7987 20451
rect 7929 20411 7987 20417
rect 8128 20380 8156 20479
rect 8202 20476 8208 20528
rect 8260 20476 8266 20528
rect 8294 20408 8300 20460
rect 8352 20408 8358 20460
rect 8772 20448 8800 20556
rect 9766 20544 9772 20596
rect 9824 20584 9830 20596
rect 10502 20584 10508 20596
rect 9824 20556 10508 20584
rect 9824 20544 9830 20556
rect 10502 20544 10508 20556
rect 10560 20544 10566 20596
rect 12434 20584 12440 20596
rect 10980 20556 12440 20584
rect 10980 20525 11008 20556
rect 12434 20544 12440 20556
rect 12492 20544 12498 20596
rect 13354 20584 13360 20596
rect 12544 20556 13360 20584
rect 10965 20519 11023 20525
rect 10965 20485 10977 20519
rect 11011 20485 11023 20519
rect 11422 20516 11428 20528
rect 10965 20479 11023 20485
rect 11072 20488 11428 20516
rect 10410 20448 10416 20460
rect 8772 20420 10416 20448
rect 10410 20408 10416 20420
rect 10468 20448 10474 20460
rect 10505 20451 10563 20457
rect 10505 20448 10517 20451
rect 10468 20420 10517 20448
rect 10468 20408 10474 20420
rect 10505 20417 10517 20420
rect 10551 20417 10563 20451
rect 10781 20451 10839 20457
rect 10781 20448 10793 20451
rect 10505 20411 10563 20417
rect 10704 20420 10793 20448
rect 8846 20380 8852 20392
rect 5184 20352 6040 20380
rect 8128 20352 8852 20380
rect 5350 20312 5356 20324
rect 5092 20284 5356 20312
rect 4525 20275 4583 20281
rect 5350 20272 5356 20284
rect 5408 20272 5414 20324
rect 2832 20216 3280 20244
rect 2832 20204 2838 20216
rect 3326 20204 3332 20256
rect 3384 20244 3390 20256
rect 3605 20247 3663 20253
rect 3605 20244 3617 20247
rect 3384 20216 3617 20244
rect 3384 20204 3390 20216
rect 3605 20213 3617 20216
rect 3651 20213 3663 20247
rect 3605 20207 3663 20213
rect 3786 20204 3792 20256
rect 3844 20244 3850 20256
rect 4157 20247 4215 20253
rect 4157 20244 4169 20247
rect 3844 20216 4169 20244
rect 3844 20204 3850 20216
rect 4157 20213 4169 20216
rect 4203 20213 4215 20247
rect 4157 20207 4215 20213
rect 4893 20247 4951 20253
rect 4893 20213 4905 20247
rect 4939 20244 4951 20247
rect 5442 20244 5448 20256
rect 4939 20216 5448 20244
rect 4939 20213 4951 20216
rect 4893 20207 4951 20213
rect 5442 20204 5448 20216
rect 5500 20204 5506 20256
rect 6012 20253 6040 20352
rect 8846 20340 8852 20352
rect 8904 20340 8910 20392
rect 6270 20272 6276 20324
rect 6328 20312 6334 20324
rect 10502 20312 10508 20324
rect 6328 20284 10508 20312
rect 6328 20272 6334 20284
rect 10502 20272 10508 20284
rect 10560 20272 10566 20324
rect 5997 20247 6055 20253
rect 5997 20213 6009 20247
rect 6043 20244 6055 20247
rect 6362 20244 6368 20256
rect 6043 20216 6368 20244
rect 6043 20213 6055 20216
rect 5997 20207 6055 20213
rect 6362 20204 6368 20216
rect 6420 20204 6426 20256
rect 8481 20247 8539 20253
rect 8481 20213 8493 20247
rect 8527 20244 8539 20247
rect 8846 20244 8852 20256
rect 8527 20216 8852 20244
rect 8527 20213 8539 20216
rect 8481 20207 8539 20213
rect 8846 20204 8852 20216
rect 8904 20244 8910 20256
rect 9214 20244 9220 20256
rect 8904 20216 9220 20244
rect 8904 20204 8910 20216
rect 9214 20204 9220 20216
rect 9272 20204 9278 20256
rect 9858 20204 9864 20256
rect 9916 20244 9922 20256
rect 10704 20253 10732 20420
rect 10781 20417 10793 20420
rect 10827 20417 10839 20451
rect 10781 20411 10839 20417
rect 10870 20340 10876 20392
rect 10928 20380 10934 20392
rect 11072 20380 11100 20488
rect 11422 20476 11428 20488
rect 11480 20476 11486 20528
rect 12544 20516 12572 20556
rect 13354 20544 13360 20556
rect 13412 20584 13418 20596
rect 15102 20584 15108 20596
rect 13412 20556 13860 20584
rect 13412 20544 13418 20556
rect 13832 20525 13860 20556
rect 14108 20556 15108 20584
rect 11532 20488 12572 20516
rect 13817 20519 13875 20525
rect 11532 20457 11560 20488
rect 13817 20485 13829 20519
rect 13863 20485 13875 20519
rect 13817 20479 13875 20485
rect 11149 20451 11207 20457
rect 11149 20417 11161 20451
rect 11195 20448 11207 20451
rect 11517 20451 11575 20457
rect 11517 20448 11529 20451
rect 11195 20420 11529 20448
rect 11195 20417 11207 20420
rect 11149 20411 11207 20417
rect 11517 20417 11529 20420
rect 11563 20417 11575 20451
rect 11517 20411 11575 20417
rect 11698 20408 11704 20460
rect 11756 20408 11762 20460
rect 11790 20408 11796 20460
rect 11848 20408 11854 20460
rect 12250 20408 12256 20460
rect 12308 20408 12314 20460
rect 14108 20457 14136 20556
rect 15102 20544 15108 20556
rect 15160 20544 15166 20596
rect 15746 20544 15752 20596
rect 15804 20544 15810 20596
rect 16482 20584 16488 20596
rect 15948 20556 16488 20584
rect 14458 20476 14464 20528
rect 14516 20516 14522 20528
rect 14553 20519 14611 20525
rect 14553 20516 14565 20519
rect 14516 20488 14565 20516
rect 14516 20476 14522 20488
rect 14553 20485 14565 20488
rect 14599 20485 14611 20519
rect 14553 20479 14611 20485
rect 15194 20476 15200 20528
rect 15252 20516 15258 20528
rect 15473 20519 15531 20525
rect 15473 20516 15485 20519
rect 15252 20488 15485 20516
rect 15252 20476 15258 20488
rect 15473 20485 15485 20488
rect 15519 20516 15531 20519
rect 15764 20516 15792 20544
rect 15948 20525 15976 20556
rect 16482 20544 16488 20556
rect 16540 20544 16546 20596
rect 17034 20544 17040 20596
rect 17092 20584 17098 20596
rect 18417 20587 18475 20593
rect 17092 20556 18092 20584
rect 17092 20544 17098 20556
rect 15519 20488 15792 20516
rect 15933 20519 15991 20525
rect 15519 20485 15531 20488
rect 15473 20479 15531 20485
rect 15933 20485 15945 20519
rect 15979 20485 15991 20519
rect 15933 20479 15991 20485
rect 16022 20476 16028 20528
rect 16080 20516 16086 20528
rect 17957 20519 18015 20525
rect 17957 20516 17969 20519
rect 16080 20488 17969 20516
rect 16080 20476 16086 20488
rect 17957 20485 17969 20488
rect 18003 20485 18015 20519
rect 18064 20516 18092 20556
rect 18417 20553 18429 20587
rect 18463 20584 18475 20587
rect 21269 20587 21327 20593
rect 18463 20556 20852 20584
rect 18463 20553 18475 20556
rect 18417 20547 18475 20553
rect 20824 20525 20852 20556
rect 21269 20553 21281 20587
rect 21315 20584 21327 20587
rect 30377 20587 30435 20593
rect 21315 20556 26372 20584
rect 21315 20553 21327 20556
rect 21269 20547 21327 20553
rect 20809 20519 20867 20525
rect 18064 20488 20668 20516
rect 17957 20479 18015 20485
rect 12345 20451 12403 20457
rect 14093 20452 14151 20457
rect 12345 20417 12357 20451
rect 12391 20417 12403 20451
rect 12345 20411 12403 20417
rect 13924 20451 14151 20452
rect 13924 20424 14105 20451
rect 11422 20380 11428 20392
rect 10928 20352 11100 20380
rect 11164 20352 11428 20380
rect 10928 20340 10934 20352
rect 11164 20324 11192 20352
rect 11422 20340 11428 20352
rect 11480 20380 11486 20392
rect 12360 20380 12388 20411
rect 11480 20352 12388 20380
rect 11480 20340 11486 20352
rect 12710 20340 12716 20392
rect 12768 20380 12774 20392
rect 13924 20380 13952 20424
rect 14093 20417 14105 20424
rect 14139 20417 14151 20451
rect 14093 20411 14151 20417
rect 14642 20408 14648 20460
rect 14700 20448 14706 20460
rect 15289 20451 15347 20457
rect 15289 20448 15301 20451
rect 14700 20420 15301 20448
rect 14700 20408 14706 20420
rect 15289 20417 15301 20420
rect 15335 20417 15347 20451
rect 15289 20411 15347 20417
rect 15562 20408 15568 20460
rect 15620 20448 15626 20460
rect 15749 20451 15807 20457
rect 15749 20448 15761 20451
rect 15620 20420 15761 20448
rect 15620 20408 15626 20420
rect 15749 20417 15761 20420
rect 15795 20417 15807 20451
rect 15749 20411 15807 20417
rect 16482 20408 16488 20460
rect 16540 20448 16546 20460
rect 16669 20451 16727 20457
rect 16669 20448 16681 20451
rect 16540 20420 16681 20448
rect 16540 20408 16546 20420
rect 16669 20417 16681 20420
rect 16715 20417 16727 20451
rect 16669 20411 16727 20417
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 16853 20451 16911 20457
rect 16853 20448 16865 20451
rect 16816 20420 16865 20448
rect 16816 20408 16822 20420
rect 16853 20417 16865 20420
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 16942 20408 16948 20460
rect 17000 20408 17006 20460
rect 17218 20408 17224 20460
rect 17276 20448 17282 20460
rect 18233 20451 18291 20457
rect 18233 20448 18245 20451
rect 17276 20420 18245 20448
rect 17276 20408 17282 20420
rect 18233 20417 18245 20420
rect 18279 20417 18291 20451
rect 18233 20411 18291 20417
rect 18877 20451 18935 20457
rect 18877 20417 18889 20451
rect 18923 20448 18935 20451
rect 19334 20448 19340 20460
rect 18923 20420 19340 20448
rect 18923 20417 18935 20420
rect 18877 20411 18935 20417
rect 19334 20408 19340 20420
rect 19392 20408 19398 20460
rect 19978 20408 19984 20460
rect 20036 20408 20042 20460
rect 20254 20408 20260 20460
rect 20312 20408 20318 20460
rect 20640 20448 20668 20488
rect 20809 20485 20821 20519
rect 20855 20485 20867 20519
rect 20809 20479 20867 20485
rect 20898 20476 20904 20528
rect 20956 20516 20962 20528
rect 22741 20519 22799 20525
rect 22741 20516 22753 20519
rect 20956 20488 22753 20516
rect 20956 20476 20962 20488
rect 22741 20485 22753 20488
rect 22787 20485 22799 20519
rect 22741 20479 22799 20485
rect 23934 20476 23940 20528
rect 23992 20516 23998 20528
rect 26344 20516 26372 20556
rect 30377 20553 30389 20587
rect 30423 20584 30435 20587
rect 30742 20584 30748 20596
rect 30423 20556 30748 20584
rect 30423 20553 30435 20556
rect 30377 20547 30435 20553
rect 30742 20544 30748 20556
rect 30800 20544 30806 20596
rect 23992 20488 26280 20516
rect 26344 20488 30788 20516
rect 23992 20476 23998 20488
rect 20714 20448 20720 20460
rect 20640 20420 20720 20448
rect 20714 20408 20720 20420
rect 20772 20408 20778 20460
rect 21082 20408 21088 20460
rect 21140 20448 21146 20460
rect 21634 20448 21640 20460
rect 21140 20420 21640 20448
rect 21140 20408 21146 20420
rect 21634 20408 21640 20420
rect 21692 20408 21698 20460
rect 22554 20408 22560 20460
rect 22612 20408 22618 20460
rect 23290 20408 23296 20460
rect 23348 20448 23354 20460
rect 24213 20451 24271 20457
rect 24213 20448 24225 20451
rect 23348 20420 24225 20448
rect 23348 20408 23354 20420
rect 24213 20417 24225 20420
rect 24259 20417 24271 20451
rect 24213 20411 24271 20417
rect 24489 20451 24547 20457
rect 24489 20417 24501 20451
rect 24535 20417 24547 20451
rect 26252 20448 26280 20488
rect 30760 20460 30788 20488
rect 30834 20476 30840 20528
rect 30892 20476 30898 20528
rect 30926 20476 30932 20528
rect 30984 20476 30990 20528
rect 28718 20448 28724 20460
rect 26252 20420 28724 20448
rect 24489 20411 24547 20417
rect 12768 20352 13952 20380
rect 12768 20340 12774 20352
rect 13998 20340 14004 20392
rect 14056 20340 14062 20392
rect 14369 20383 14427 20389
rect 14108 20352 14320 20380
rect 11146 20272 11152 20324
rect 11204 20272 11210 20324
rect 11606 20272 11612 20324
rect 11664 20272 11670 20324
rect 11698 20272 11704 20324
rect 11756 20312 11762 20324
rect 11977 20315 12035 20321
rect 11977 20312 11989 20315
rect 11756 20284 11989 20312
rect 11756 20272 11762 20284
rect 11977 20281 11989 20284
rect 12023 20281 12035 20315
rect 11977 20275 12035 20281
rect 12069 20315 12127 20321
rect 12069 20281 12081 20315
rect 12115 20312 12127 20315
rect 12434 20312 12440 20324
rect 12115 20284 12440 20312
rect 12115 20281 12127 20284
rect 12069 20275 12127 20281
rect 10689 20247 10747 20253
rect 10689 20244 10701 20247
rect 9916 20216 10701 20244
rect 9916 20204 9922 20216
rect 10689 20213 10701 20216
rect 10735 20213 10747 20247
rect 10689 20207 10747 20213
rect 11238 20204 11244 20256
rect 11296 20244 11302 20256
rect 11517 20247 11575 20253
rect 11517 20244 11529 20247
rect 11296 20216 11529 20244
rect 11296 20204 11302 20216
rect 11517 20213 11529 20216
rect 11563 20213 11575 20247
rect 11624 20244 11652 20272
rect 12084 20244 12112 20275
rect 12434 20272 12440 20284
rect 12492 20272 12498 20324
rect 12526 20272 12532 20324
rect 12584 20312 12590 20324
rect 13630 20312 13636 20324
rect 12584 20284 13636 20312
rect 12584 20272 12590 20284
rect 13630 20272 13636 20284
rect 13688 20272 13694 20324
rect 14108 20312 14136 20352
rect 13740 20284 14136 20312
rect 14292 20312 14320 20352
rect 14369 20349 14381 20383
rect 14415 20380 14427 20383
rect 14458 20380 14464 20392
rect 14415 20352 14464 20380
rect 14415 20349 14427 20352
rect 14369 20343 14427 20349
rect 14458 20340 14464 20352
rect 14516 20340 14522 20392
rect 14734 20340 14740 20392
rect 14792 20380 14798 20392
rect 14918 20380 14924 20392
rect 14792 20352 14924 20380
rect 14792 20340 14798 20352
rect 14918 20340 14924 20352
rect 14976 20340 14982 20392
rect 16298 20340 16304 20392
rect 16356 20380 16362 20392
rect 18141 20383 18199 20389
rect 16356 20352 18092 20380
rect 16356 20340 16362 20352
rect 16758 20312 16764 20324
rect 14292 20284 16764 20312
rect 11624 20216 12112 20244
rect 11517 20207 11575 20213
rect 13078 20204 13084 20256
rect 13136 20244 13142 20256
rect 13740 20244 13768 20284
rect 16758 20272 16764 20284
rect 16816 20272 16822 20324
rect 17126 20272 17132 20324
rect 17184 20272 17190 20324
rect 18064 20312 18092 20352
rect 18141 20349 18153 20383
rect 18187 20380 18199 20383
rect 18322 20380 18328 20392
rect 18187 20352 18328 20380
rect 18187 20349 18199 20352
rect 18141 20343 18199 20349
rect 18322 20340 18328 20352
rect 18380 20340 18386 20392
rect 18969 20383 19027 20389
rect 18969 20349 18981 20383
rect 19015 20349 19027 20383
rect 18969 20343 19027 20349
rect 18984 20312 19012 20343
rect 19794 20340 19800 20392
rect 19852 20380 19858 20392
rect 20073 20383 20131 20389
rect 20073 20380 20085 20383
rect 19852 20352 20085 20380
rect 19852 20340 19858 20352
rect 20073 20349 20085 20352
rect 20119 20349 20131 20383
rect 20073 20343 20131 20349
rect 20901 20383 20959 20389
rect 20901 20349 20913 20383
rect 20947 20349 20959 20383
rect 20901 20343 20959 20349
rect 18064 20284 19012 20312
rect 19245 20315 19303 20321
rect 19245 20281 19257 20315
rect 19291 20312 19303 20315
rect 19886 20312 19892 20324
rect 19291 20284 19892 20312
rect 19291 20281 19303 20284
rect 19245 20275 19303 20281
rect 19886 20272 19892 20284
rect 19944 20272 19950 20324
rect 20441 20315 20499 20321
rect 20441 20281 20453 20315
rect 20487 20312 20499 20315
rect 20916 20312 20944 20343
rect 22278 20340 22284 20392
rect 22336 20380 22342 20392
rect 23014 20380 23020 20392
rect 22336 20352 23020 20380
rect 22336 20340 22342 20352
rect 23014 20340 23020 20352
rect 23072 20340 23078 20392
rect 24026 20340 24032 20392
rect 24084 20380 24090 20392
rect 24305 20383 24363 20389
rect 24305 20380 24317 20383
rect 24084 20352 24317 20380
rect 24084 20340 24090 20352
rect 24305 20349 24317 20352
rect 24351 20349 24363 20383
rect 24504 20380 24532 20411
rect 28718 20408 28724 20420
rect 28776 20408 28782 20460
rect 30009 20451 30067 20457
rect 30009 20417 30021 20451
rect 30055 20448 30067 20451
rect 30190 20448 30196 20460
rect 30055 20420 30196 20448
rect 30055 20417 30067 20420
rect 30009 20411 30067 20417
rect 30190 20408 30196 20420
rect 30248 20408 30254 20460
rect 30374 20408 30380 20460
rect 30432 20448 30438 20460
rect 30653 20451 30711 20457
rect 30653 20448 30665 20451
rect 30432 20420 30665 20448
rect 30432 20408 30438 20420
rect 30653 20417 30665 20420
rect 30699 20417 30711 20451
rect 30653 20411 30711 20417
rect 30742 20408 30748 20460
rect 30800 20408 30806 20460
rect 31021 20451 31079 20457
rect 31021 20417 31033 20451
rect 31067 20448 31079 20451
rect 31297 20451 31355 20457
rect 31297 20448 31309 20451
rect 31067 20420 31309 20448
rect 31067 20417 31079 20420
rect 31021 20411 31079 20417
rect 31297 20417 31309 20420
rect 31343 20417 31355 20451
rect 31297 20411 31355 20417
rect 31754 20408 31760 20460
rect 31812 20448 31818 20460
rect 32217 20451 32275 20457
rect 32217 20448 32229 20451
rect 31812 20420 32229 20448
rect 31812 20408 31818 20420
rect 32217 20417 32229 20420
rect 32263 20417 32275 20451
rect 32217 20411 32275 20417
rect 26418 20380 26424 20392
rect 24504 20352 26424 20380
rect 24305 20343 24363 20349
rect 26418 20340 26424 20352
rect 26476 20340 26482 20392
rect 29730 20340 29736 20392
rect 29788 20380 29794 20392
rect 29788 20352 30052 20380
rect 29788 20340 29794 20352
rect 20487 20284 20944 20312
rect 20487 20281 20499 20284
rect 20441 20275 20499 20281
rect 21450 20272 21456 20324
rect 21508 20312 21514 20324
rect 21634 20312 21640 20324
rect 21508 20284 21640 20312
rect 21508 20272 21514 20284
rect 21634 20272 21640 20284
rect 21692 20272 21698 20324
rect 24578 20312 24584 20324
rect 24412 20284 24584 20312
rect 13136 20216 13768 20244
rect 13136 20204 13142 20216
rect 13998 20204 14004 20256
rect 14056 20204 14062 20256
rect 14277 20247 14335 20253
rect 14277 20213 14289 20247
rect 14323 20244 14335 20247
rect 15378 20244 15384 20256
rect 14323 20216 15384 20244
rect 14323 20213 14335 20216
rect 14277 20207 14335 20213
rect 15378 20204 15384 20216
rect 15436 20204 15442 20256
rect 15654 20204 15660 20256
rect 15712 20204 15718 20256
rect 16117 20247 16175 20253
rect 16117 20213 16129 20247
rect 16163 20244 16175 20247
rect 16669 20247 16727 20253
rect 16669 20244 16681 20247
rect 16163 20216 16681 20244
rect 16163 20213 16175 20216
rect 16117 20207 16175 20213
rect 16669 20213 16681 20216
rect 16715 20213 16727 20247
rect 16669 20207 16727 20213
rect 17770 20204 17776 20256
rect 17828 20244 17834 20256
rect 17957 20247 18015 20253
rect 17957 20244 17969 20247
rect 17828 20216 17969 20244
rect 17828 20204 17834 20216
rect 17957 20213 17969 20216
rect 18003 20213 18015 20247
rect 17957 20207 18015 20213
rect 18785 20247 18843 20253
rect 18785 20213 18797 20247
rect 18831 20244 18843 20247
rect 18877 20247 18935 20253
rect 18877 20244 18889 20247
rect 18831 20216 18889 20244
rect 18831 20213 18843 20216
rect 18785 20207 18843 20213
rect 18877 20213 18889 20216
rect 18923 20244 18935 20247
rect 19150 20244 19156 20256
rect 18923 20216 19156 20244
rect 18923 20213 18935 20216
rect 18877 20207 18935 20213
rect 19150 20204 19156 20216
rect 19208 20204 19214 20256
rect 20257 20247 20315 20253
rect 20257 20213 20269 20247
rect 20303 20244 20315 20247
rect 20346 20244 20352 20256
rect 20303 20216 20352 20244
rect 20303 20213 20315 20216
rect 20257 20207 20315 20213
rect 20346 20204 20352 20216
rect 20404 20204 20410 20256
rect 20714 20204 20720 20256
rect 20772 20244 20778 20256
rect 20809 20247 20867 20253
rect 20809 20244 20821 20247
rect 20772 20216 20821 20244
rect 20772 20204 20778 20216
rect 20809 20213 20821 20216
rect 20855 20213 20867 20247
rect 20809 20207 20867 20213
rect 22925 20247 22983 20253
rect 22925 20213 22937 20247
rect 22971 20244 22983 20247
rect 23014 20244 23020 20256
rect 22971 20216 23020 20244
rect 22971 20213 22983 20216
rect 22925 20207 22983 20213
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 24412 20253 24440 20284
rect 24578 20272 24584 20284
rect 24636 20272 24642 20324
rect 29178 20272 29184 20324
rect 29236 20312 29242 20324
rect 29822 20312 29828 20324
rect 29236 20284 29828 20312
rect 29236 20272 29242 20284
rect 29822 20272 29828 20284
rect 29880 20272 29886 20324
rect 30024 20312 30052 20352
rect 30098 20340 30104 20392
rect 30156 20340 30162 20392
rect 31941 20383 31999 20389
rect 31941 20349 31953 20383
rect 31987 20380 31999 20383
rect 32122 20380 32128 20392
rect 31987 20352 32128 20380
rect 31987 20349 31999 20352
rect 31941 20343 31999 20349
rect 32122 20340 32128 20352
rect 32180 20380 32186 20392
rect 32490 20380 32496 20392
rect 32180 20352 32496 20380
rect 32180 20340 32186 20352
rect 32490 20340 32496 20352
rect 32548 20340 32554 20392
rect 30024 20284 30144 20312
rect 30116 20256 30144 20284
rect 24397 20247 24455 20253
rect 24397 20213 24409 20247
rect 24443 20213 24455 20247
rect 24397 20207 24455 20213
rect 24486 20204 24492 20256
rect 24544 20244 24550 20256
rect 24673 20247 24731 20253
rect 24673 20244 24685 20247
rect 24544 20216 24685 20244
rect 24544 20204 24550 20216
rect 24673 20213 24685 20216
rect 24719 20213 24731 20247
rect 24673 20207 24731 20213
rect 26878 20204 26884 20256
rect 26936 20244 26942 20256
rect 27430 20244 27436 20256
rect 26936 20216 27436 20244
rect 26936 20204 26942 20216
rect 27430 20204 27436 20216
rect 27488 20204 27494 20256
rect 29454 20204 29460 20256
rect 29512 20244 29518 20256
rect 29730 20244 29736 20256
rect 29512 20216 29736 20244
rect 29512 20204 29518 20216
rect 29730 20204 29736 20216
rect 29788 20204 29794 20256
rect 30006 20204 30012 20256
rect 30064 20204 30070 20256
rect 30098 20204 30104 20256
rect 30156 20204 30162 20256
rect 31202 20204 31208 20256
rect 31260 20204 31266 20256
rect 32398 20204 32404 20256
rect 32456 20204 32462 20256
rect 1104 20154 32844 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 32844 20154
rect 1104 20080 32844 20102
rect 3421 20043 3479 20049
rect 3421 20009 3433 20043
rect 3467 20040 3479 20043
rect 3970 20040 3976 20052
rect 3467 20012 3976 20040
rect 3467 20009 3479 20012
rect 3421 20003 3479 20009
rect 3970 20000 3976 20012
rect 4028 20000 4034 20052
rect 4890 20040 4896 20052
rect 4448 20012 4896 20040
rect 2777 19975 2835 19981
rect 2777 19941 2789 19975
rect 2823 19941 2835 19975
rect 2777 19935 2835 19941
rect 1394 19864 1400 19916
rect 1452 19864 1458 19916
rect 2792 19904 2820 19935
rect 2958 19932 2964 19984
rect 3016 19972 3022 19984
rect 3789 19975 3847 19981
rect 3789 19972 3801 19975
rect 3016 19944 3801 19972
rect 3016 19932 3022 19944
rect 3789 19941 3801 19944
rect 3835 19941 3847 19975
rect 3789 19935 3847 19941
rect 3878 19932 3884 19984
rect 3936 19972 3942 19984
rect 4448 19972 4476 20012
rect 4890 20000 4896 20012
rect 4948 20040 4954 20052
rect 5629 20043 5687 20049
rect 5629 20040 5641 20043
rect 4948 20012 5641 20040
rect 4948 20000 4954 20012
rect 5629 20009 5641 20012
rect 5675 20009 5687 20043
rect 5629 20003 5687 20009
rect 8202 20000 8208 20052
rect 8260 20000 8266 20052
rect 9398 20000 9404 20052
rect 9456 20000 9462 20052
rect 12802 20000 12808 20052
rect 12860 20040 12866 20052
rect 13630 20040 13636 20052
rect 12860 20012 13636 20040
rect 12860 20000 12866 20012
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 13725 20043 13783 20049
rect 13725 20009 13737 20043
rect 13771 20040 13783 20043
rect 13998 20040 14004 20052
rect 13771 20012 14004 20040
rect 13771 20009 13783 20012
rect 13725 20003 13783 20009
rect 5442 19972 5448 19984
rect 3936 19944 4476 19972
rect 4540 19944 5448 19972
rect 3936 19932 3942 19944
rect 2792 19876 4016 19904
rect 2590 19796 2596 19848
rect 2648 19836 2654 19848
rect 2961 19839 3019 19845
rect 2961 19836 2973 19839
rect 2648 19808 2973 19836
rect 2648 19796 2654 19808
rect 2961 19805 2973 19808
rect 3007 19805 3019 19839
rect 2961 19799 3019 19805
rect 3053 19839 3111 19845
rect 3053 19805 3065 19839
rect 3099 19805 3111 19839
rect 3053 19799 3111 19805
rect 1670 19777 1676 19780
rect 1664 19731 1676 19777
rect 1670 19728 1676 19731
rect 1728 19728 1734 19780
rect 2314 19728 2320 19780
rect 2372 19768 2378 19780
rect 3068 19768 3096 19799
rect 3142 19796 3148 19848
rect 3200 19796 3206 19848
rect 3234 19796 3240 19848
rect 3292 19796 3298 19848
rect 3988 19845 4016 19876
rect 3973 19839 4031 19845
rect 3973 19805 3985 19839
rect 4019 19805 4031 19839
rect 3973 19799 4031 19805
rect 4341 19839 4399 19845
rect 4341 19805 4353 19839
rect 4387 19836 4399 19839
rect 4540 19836 4568 19944
rect 5442 19932 5448 19944
rect 5500 19932 5506 19984
rect 5537 19975 5595 19981
rect 5537 19941 5549 19975
rect 5583 19972 5595 19975
rect 6270 19972 6276 19984
rect 5583 19944 6276 19972
rect 5583 19941 5595 19944
rect 5537 19935 5595 19941
rect 6270 19932 6276 19944
rect 6328 19932 6334 19984
rect 6546 19932 6552 19984
rect 6604 19972 6610 19984
rect 6604 19944 7328 19972
rect 6604 19932 6610 19944
rect 4632 19876 6408 19904
rect 4632 19845 4660 19876
rect 4387 19808 4568 19836
rect 4617 19839 4675 19845
rect 4387 19805 4399 19808
rect 4341 19799 4399 19805
rect 4617 19805 4629 19839
rect 4663 19805 4675 19839
rect 4617 19799 4675 19805
rect 4709 19839 4767 19845
rect 4709 19805 4721 19839
rect 4755 19836 4767 19839
rect 4890 19836 4896 19848
rect 4755 19808 4896 19836
rect 4755 19805 4767 19808
rect 4709 19799 4767 19805
rect 4890 19796 4896 19808
rect 4948 19796 4954 19848
rect 5000 19845 5028 19876
rect 6380 19848 6408 19876
rect 7190 19864 7196 19916
rect 7248 19864 7254 19916
rect 4985 19839 5043 19845
rect 4985 19805 4997 19839
rect 5031 19805 5043 19839
rect 4985 19799 5043 19805
rect 5350 19796 5356 19848
rect 5408 19796 5414 19848
rect 5718 19796 5724 19848
rect 5776 19836 5782 19848
rect 5813 19839 5871 19845
rect 5813 19836 5825 19839
rect 5776 19808 5825 19836
rect 5776 19796 5782 19808
rect 5813 19805 5825 19808
rect 5859 19805 5871 19839
rect 5813 19799 5871 19805
rect 6089 19839 6147 19845
rect 6089 19805 6101 19839
rect 6135 19805 6147 19839
rect 6089 19799 6147 19805
rect 2372 19740 3096 19768
rect 3712 19740 3924 19768
rect 2372 19728 2378 19740
rect 2406 19660 2412 19712
rect 2464 19700 2470 19712
rect 3712 19700 3740 19740
rect 2464 19672 3740 19700
rect 3896 19700 3924 19740
rect 4062 19728 4068 19780
rect 4120 19768 4126 19780
rect 4525 19771 4583 19777
rect 4525 19768 4537 19771
rect 4120 19740 4537 19768
rect 4120 19728 4126 19740
rect 4525 19737 4537 19740
rect 4571 19737 4583 19771
rect 4525 19731 4583 19737
rect 4798 19728 4804 19780
rect 4856 19768 4862 19780
rect 5169 19771 5227 19777
rect 5169 19768 5181 19771
rect 4856 19740 5181 19768
rect 4856 19728 4862 19740
rect 5169 19737 5181 19740
rect 5215 19737 5227 19771
rect 5169 19731 5227 19737
rect 5261 19771 5319 19777
rect 5261 19737 5273 19771
rect 5307 19768 5319 19771
rect 5442 19768 5448 19780
rect 5307 19740 5448 19768
rect 5307 19737 5319 19740
rect 5261 19731 5319 19737
rect 5442 19728 5448 19740
rect 5500 19768 5506 19780
rect 6104 19768 6132 19799
rect 6362 19796 6368 19848
rect 6420 19796 6426 19848
rect 6454 19796 6460 19848
rect 6512 19796 6518 19848
rect 7009 19839 7067 19845
rect 7009 19805 7021 19839
rect 7055 19836 7067 19839
rect 7208 19836 7236 19864
rect 7300 19845 7328 19944
rect 7558 19932 7564 19984
rect 7616 19972 7622 19984
rect 13740 19972 13768 20003
rect 13998 20000 14004 20012
rect 14056 20000 14062 20052
rect 14642 20000 14648 20052
rect 14700 20000 14706 20052
rect 14829 20043 14887 20049
rect 14829 20009 14841 20043
rect 14875 20040 14887 20043
rect 16022 20040 16028 20052
rect 14875 20012 16028 20040
rect 14875 20009 14887 20012
rect 14829 20003 14887 20009
rect 16022 20000 16028 20012
rect 16080 20000 16086 20052
rect 16482 20000 16488 20052
rect 16540 20000 16546 20052
rect 16945 20043 17003 20049
rect 16945 20009 16957 20043
rect 16991 20040 17003 20043
rect 17218 20040 17224 20052
rect 16991 20012 17224 20040
rect 16991 20009 17003 20012
rect 16945 20003 17003 20009
rect 17218 20000 17224 20012
rect 17276 20000 17282 20052
rect 19610 20000 19616 20052
rect 19668 20040 19674 20052
rect 20254 20040 20260 20052
rect 19668 20012 20260 20040
rect 19668 20000 19674 20012
rect 20254 20000 20260 20012
rect 20312 20000 20318 20052
rect 20714 20000 20720 20052
rect 20772 20000 20778 20052
rect 20898 20000 20904 20052
rect 20956 20000 20962 20052
rect 23658 20000 23664 20052
rect 23716 20040 23722 20052
rect 24397 20043 24455 20049
rect 24397 20040 24409 20043
rect 23716 20012 24409 20040
rect 23716 20000 23722 20012
rect 24397 20009 24409 20012
rect 24443 20009 24455 20043
rect 24397 20003 24455 20009
rect 24762 20000 24768 20052
rect 24820 20000 24826 20052
rect 26050 20000 26056 20052
rect 26108 20000 26114 20052
rect 26418 20000 26424 20052
rect 26476 20040 26482 20052
rect 26513 20043 26571 20049
rect 26513 20040 26525 20043
rect 26476 20012 26525 20040
rect 26476 20000 26482 20012
rect 26513 20009 26525 20012
rect 26559 20040 26571 20043
rect 26694 20040 26700 20052
rect 26559 20012 26700 20040
rect 26559 20009 26571 20012
rect 26513 20003 26571 20009
rect 26694 20000 26700 20012
rect 26752 20000 26758 20052
rect 26786 20000 26792 20052
rect 26844 20000 26850 20052
rect 27890 20000 27896 20052
rect 27948 20040 27954 20052
rect 27985 20043 28043 20049
rect 27985 20040 27997 20043
rect 27948 20012 27997 20040
rect 27948 20000 27954 20012
rect 27985 20009 27997 20012
rect 28031 20009 28043 20043
rect 27985 20003 28043 20009
rect 28994 20000 29000 20052
rect 29052 20040 29058 20052
rect 29549 20043 29607 20049
rect 29549 20040 29561 20043
rect 29052 20012 29561 20040
rect 29052 20000 29058 20012
rect 29549 20009 29561 20012
rect 29595 20009 29607 20043
rect 30193 20043 30251 20049
rect 30193 20040 30205 20043
rect 29549 20003 29607 20009
rect 29656 20012 30205 20040
rect 7616 19944 13768 19972
rect 14016 19944 15608 19972
rect 7616 19932 7622 19944
rect 8110 19864 8116 19916
rect 8168 19864 8174 19916
rect 9674 19904 9680 19916
rect 9232 19876 9680 19904
rect 7055 19808 7236 19836
rect 7285 19839 7343 19845
rect 7055 19805 7067 19808
rect 7009 19799 7067 19805
rect 7285 19805 7297 19839
rect 7331 19805 7343 19839
rect 7285 19799 7343 19805
rect 7374 19796 7380 19848
rect 7432 19796 7438 19848
rect 7653 19839 7711 19845
rect 7653 19805 7665 19839
rect 7699 19836 7711 19839
rect 8128 19836 8156 19864
rect 8389 19839 8447 19845
rect 8389 19836 8401 19839
rect 7699 19808 8156 19836
rect 8266 19808 8401 19836
rect 7699 19805 7711 19808
rect 7653 19799 7711 19805
rect 5500 19740 6132 19768
rect 6273 19771 6331 19777
rect 5500 19728 5506 19740
rect 6273 19737 6285 19771
rect 6319 19737 6331 19771
rect 6273 19731 6331 19737
rect 7193 19771 7251 19777
rect 7193 19737 7205 19771
rect 7239 19768 7251 19771
rect 7929 19771 7987 19777
rect 7239 19740 7420 19768
rect 7239 19737 7251 19740
rect 7193 19731 7251 19737
rect 4893 19703 4951 19709
rect 4893 19700 4905 19703
rect 3896 19672 4905 19700
rect 2464 19660 2470 19672
rect 4893 19669 4905 19672
rect 4939 19669 4951 19703
rect 4893 19663 4951 19669
rect 5994 19660 6000 19712
rect 6052 19700 6058 19712
rect 6288 19700 6316 19731
rect 7392 19712 7420 19740
rect 7929 19737 7941 19771
rect 7975 19737 7987 19771
rect 7929 19731 7987 19737
rect 8113 19771 8171 19777
rect 8113 19737 8125 19771
rect 8159 19768 8171 19771
rect 8266 19768 8294 19808
rect 8389 19805 8401 19808
rect 8435 19836 8447 19839
rect 8662 19836 8668 19848
rect 8435 19808 8668 19836
rect 8435 19805 8447 19808
rect 8389 19799 8447 19805
rect 8662 19796 8668 19808
rect 8720 19796 8726 19848
rect 8938 19796 8944 19848
rect 8996 19796 9002 19848
rect 9232 19845 9260 19876
rect 9674 19864 9680 19876
rect 9732 19864 9738 19916
rect 10226 19864 10232 19916
rect 10284 19864 10290 19916
rect 11146 19864 11152 19916
rect 11204 19904 11210 19916
rect 12066 19904 12072 19916
rect 11204 19876 12072 19904
rect 11204 19864 11210 19876
rect 12066 19864 12072 19876
rect 12124 19864 12130 19916
rect 12253 19907 12311 19913
rect 12253 19873 12265 19907
rect 12299 19904 12311 19907
rect 12342 19904 12348 19916
rect 12299 19876 12348 19904
rect 12299 19873 12311 19876
rect 12253 19867 12311 19873
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 13633 19907 13691 19913
rect 13633 19873 13645 19907
rect 13679 19904 13691 19907
rect 14016 19904 14044 19944
rect 13679 19876 14044 19904
rect 13679 19873 13691 19876
rect 13633 19867 13691 19873
rect 14458 19864 14464 19916
rect 14516 19864 14522 19916
rect 9217 19839 9275 19845
rect 9217 19805 9229 19839
rect 9263 19805 9275 19839
rect 9217 19799 9275 19805
rect 9401 19839 9459 19845
rect 9401 19805 9413 19839
rect 9447 19836 9459 19839
rect 10045 19839 10103 19845
rect 9447 19808 9674 19836
rect 9447 19805 9459 19808
rect 9401 19799 9459 19805
rect 8159 19740 8294 19768
rect 8573 19771 8631 19777
rect 8159 19737 8171 19740
rect 8113 19731 8171 19737
rect 8573 19737 8585 19771
rect 8619 19768 8631 19771
rect 8754 19768 8760 19780
rect 8619 19740 8760 19768
rect 8619 19737 8631 19740
rect 8573 19731 8631 19737
rect 6052 19672 6316 19700
rect 6052 19660 6058 19672
rect 6454 19660 6460 19712
rect 6512 19700 6518 19712
rect 6641 19703 6699 19709
rect 6641 19700 6653 19703
rect 6512 19672 6653 19700
rect 6512 19660 6518 19672
rect 6641 19669 6653 19672
rect 6687 19669 6699 19703
rect 6641 19663 6699 19669
rect 7374 19660 7380 19712
rect 7432 19660 7438 19712
rect 7558 19660 7564 19712
rect 7616 19660 7622 19712
rect 7837 19703 7895 19709
rect 7837 19669 7849 19703
rect 7883 19700 7895 19703
rect 7944 19700 7972 19731
rect 8754 19728 8760 19740
rect 8812 19728 8818 19780
rect 9232 19768 9260 19799
rect 8864 19740 9260 19768
rect 9646 19768 9674 19808
rect 10045 19805 10057 19839
rect 10091 19836 10103 19839
rect 10091 19808 10456 19836
rect 10091 19805 10103 19808
rect 10045 19799 10103 19805
rect 9646 19740 9720 19768
rect 8864 19700 8892 19740
rect 7883 19672 8892 19700
rect 9125 19703 9183 19709
rect 7883 19669 7895 19672
rect 7837 19663 7895 19669
rect 9125 19669 9137 19703
rect 9171 19700 9183 19703
rect 9398 19700 9404 19712
rect 9171 19672 9404 19700
rect 9171 19669 9183 19672
rect 9125 19663 9183 19669
rect 9398 19660 9404 19672
rect 9456 19660 9462 19712
rect 9582 19660 9588 19712
rect 9640 19660 9646 19712
rect 9692 19700 9720 19740
rect 9766 19728 9772 19780
rect 9824 19768 9830 19780
rect 9861 19771 9919 19777
rect 9861 19768 9873 19771
rect 9824 19740 9873 19768
rect 9824 19728 9830 19740
rect 9861 19737 9873 19740
rect 9907 19768 9919 19771
rect 9907 19740 10180 19768
rect 9907 19737 9919 19740
rect 9861 19731 9919 19737
rect 9950 19700 9956 19712
rect 9692 19672 9956 19700
rect 9950 19660 9956 19672
rect 10008 19660 10014 19712
rect 10152 19700 10180 19740
rect 10321 19703 10379 19709
rect 10321 19700 10333 19703
rect 10152 19672 10333 19700
rect 10321 19669 10333 19672
rect 10367 19669 10379 19703
rect 10428 19700 10456 19808
rect 10502 19796 10508 19848
rect 10560 19796 10566 19848
rect 11882 19796 11888 19848
rect 11940 19836 11946 19848
rect 11977 19839 12035 19845
rect 11977 19836 11989 19839
rect 11940 19808 11989 19836
rect 11940 19796 11946 19808
rect 11977 19805 11989 19808
rect 12023 19805 12035 19839
rect 11977 19799 12035 19805
rect 13354 19796 13360 19848
rect 13412 19836 13418 19848
rect 13449 19839 13507 19845
rect 13449 19836 13461 19839
rect 13412 19808 13461 19836
rect 13412 19796 13418 19808
rect 13449 19805 13461 19808
rect 13495 19805 13507 19839
rect 13449 19799 13507 19805
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19836 13783 19839
rect 13814 19836 13820 19848
rect 13771 19808 13820 19836
rect 13771 19805 13783 19808
rect 13725 19799 13783 19805
rect 13814 19796 13820 19808
rect 13872 19796 13878 19848
rect 14093 19839 14151 19845
rect 14093 19805 14105 19839
rect 14139 19836 14151 19839
rect 14182 19836 14188 19848
rect 14139 19808 14188 19836
rect 14139 19805 14151 19808
rect 14093 19799 14151 19805
rect 14182 19796 14188 19808
rect 14240 19796 14246 19848
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19836 14703 19839
rect 14918 19836 14924 19848
rect 14691 19808 14924 19836
rect 14691 19805 14703 19808
rect 14645 19799 14703 19805
rect 14918 19796 14924 19808
rect 14976 19796 14982 19848
rect 15580 19836 15608 19944
rect 17034 19932 17040 19984
rect 17092 19972 17098 19984
rect 17092 19944 26832 19972
rect 17092 19932 17098 19944
rect 15654 19864 15660 19916
rect 15712 19904 15718 19916
rect 15712 19876 16988 19904
rect 15712 19864 15718 19876
rect 16482 19836 16488 19848
rect 15580 19808 16488 19836
rect 16482 19796 16488 19808
rect 16540 19796 16546 19848
rect 16666 19796 16672 19848
rect 16724 19796 16730 19848
rect 16758 19796 16764 19848
rect 16816 19796 16822 19848
rect 16960 19845 16988 19876
rect 19426 19864 19432 19916
rect 19484 19904 19490 19916
rect 19886 19904 19892 19916
rect 19484 19876 19892 19904
rect 19484 19864 19490 19876
rect 19886 19864 19892 19876
rect 19944 19864 19950 19916
rect 22186 19904 22192 19916
rect 20088 19876 22192 19904
rect 16945 19839 17003 19845
rect 16945 19805 16957 19839
rect 16991 19836 17003 19839
rect 19978 19836 19984 19848
rect 16991 19808 19984 19836
rect 16991 19805 17003 19808
rect 16945 19799 17003 19805
rect 19978 19796 19984 19808
rect 20036 19796 20042 19848
rect 10505 19781 10517 19796
rect 10551 19781 10563 19796
rect 10505 19775 10563 19781
rect 11790 19728 11796 19780
rect 11848 19768 11854 19780
rect 12526 19768 12532 19780
rect 11848 19740 12532 19768
rect 11848 19728 11854 19740
rect 12526 19728 12532 19740
rect 12584 19728 12590 19780
rect 14369 19771 14427 19777
rect 14369 19768 14381 19771
rect 14108 19740 14381 19768
rect 14108 19712 14136 19740
rect 14369 19737 14381 19740
rect 14415 19737 14427 19771
rect 20088 19768 20116 19876
rect 22186 19864 22192 19876
rect 22244 19904 22250 19916
rect 23106 19904 23112 19916
rect 22244 19876 23112 19904
rect 22244 19864 22250 19876
rect 23106 19864 23112 19876
rect 23164 19864 23170 19916
rect 24486 19864 24492 19916
rect 24544 19864 24550 19916
rect 24578 19864 24584 19916
rect 24636 19904 24642 19916
rect 24946 19904 24952 19916
rect 24636 19876 24952 19904
rect 24636 19864 24642 19876
rect 24946 19864 24952 19876
rect 25004 19864 25010 19916
rect 25222 19864 25228 19916
rect 25280 19904 25286 19916
rect 25280 19876 26188 19904
rect 25280 19864 25286 19876
rect 20901 19839 20959 19845
rect 20901 19805 20913 19839
rect 20947 19836 20959 19839
rect 20990 19836 20996 19848
rect 20947 19808 20996 19836
rect 20947 19805 20959 19808
rect 20901 19799 20959 19805
rect 20990 19796 20996 19808
rect 21048 19796 21054 19848
rect 21082 19796 21088 19848
rect 21140 19796 21146 19848
rect 24118 19796 24124 19848
rect 24176 19836 24182 19848
rect 24397 19839 24455 19845
rect 24397 19836 24409 19839
rect 24176 19808 24409 19836
rect 24176 19796 24182 19808
rect 24397 19805 24409 19808
rect 24443 19805 24455 19839
rect 24397 19799 24455 19805
rect 25774 19796 25780 19848
rect 25832 19796 25838 19848
rect 26050 19796 26056 19848
rect 26108 19796 26114 19848
rect 26160 19836 26188 19876
rect 26234 19864 26240 19916
rect 26292 19864 26298 19916
rect 26694 19864 26700 19916
rect 26752 19864 26758 19916
rect 26804 19904 26832 19944
rect 26878 19932 26884 19984
rect 26936 19972 26942 19984
rect 29656 19972 29684 20012
rect 30193 20009 30205 20012
rect 30239 20009 30251 20043
rect 30193 20003 30251 20009
rect 30558 20000 30564 20052
rect 30616 20000 30622 20052
rect 30837 20043 30895 20049
rect 30837 20009 30849 20043
rect 30883 20040 30895 20043
rect 30926 20040 30932 20052
rect 30883 20012 30932 20040
rect 30883 20009 30895 20012
rect 30837 20003 30895 20009
rect 30926 20000 30932 20012
rect 30984 20000 30990 20052
rect 32490 20000 32496 20052
rect 32548 20000 32554 20052
rect 26936 19944 29684 19972
rect 29917 19975 29975 19981
rect 26936 19932 26942 19944
rect 29917 19941 29929 19975
rect 29963 19972 29975 19975
rect 29963 19944 30328 19972
rect 29963 19941 29975 19944
rect 29917 19935 29975 19941
rect 28077 19907 28135 19913
rect 28077 19904 28089 19907
rect 26804 19876 28089 19904
rect 28077 19873 28089 19876
rect 28123 19873 28135 19907
rect 28077 19867 28135 19873
rect 28166 19864 28172 19916
rect 28224 19904 28230 19916
rect 30300 19913 30328 19944
rect 30285 19907 30343 19913
rect 28224 19876 30236 19904
rect 28224 19864 28230 19876
rect 26329 19839 26387 19845
rect 26329 19836 26341 19839
rect 26160 19808 26341 19836
rect 26329 19805 26341 19808
rect 26375 19805 26387 19839
rect 26329 19799 26387 19805
rect 26418 19796 26424 19848
rect 26476 19836 26482 19848
rect 26605 19839 26663 19845
rect 26605 19836 26617 19839
rect 26476 19808 26617 19836
rect 26476 19796 26482 19808
rect 26605 19805 26617 19808
rect 26651 19805 26663 19839
rect 26605 19799 26663 19805
rect 26881 19839 26939 19845
rect 26881 19805 26893 19839
rect 26927 19836 26939 19839
rect 26927 19808 27936 19836
rect 26927 19805 26939 19808
rect 26881 19799 26939 19805
rect 14369 19731 14427 19737
rect 15764 19740 20116 19768
rect 10686 19700 10692 19712
rect 10428 19672 10692 19700
rect 10321 19663 10379 19669
rect 10686 19660 10692 19672
rect 10744 19660 10750 19712
rect 11974 19660 11980 19712
rect 12032 19700 12038 19712
rect 12710 19700 12716 19712
rect 12032 19672 12716 19700
rect 12032 19660 12038 19672
rect 12710 19660 12716 19672
rect 12768 19660 12774 19712
rect 13262 19660 13268 19712
rect 13320 19700 13326 19712
rect 13722 19700 13728 19712
rect 13320 19672 13728 19700
rect 13320 19660 13326 19672
rect 13722 19660 13728 19672
rect 13780 19660 13786 19712
rect 13909 19703 13967 19709
rect 13909 19669 13921 19703
rect 13955 19700 13967 19703
rect 13998 19700 14004 19712
rect 13955 19672 14004 19700
rect 13955 19669 13967 19672
rect 13909 19663 13967 19669
rect 13998 19660 14004 19672
rect 14056 19660 14062 19712
rect 14090 19660 14096 19712
rect 14148 19660 14154 19712
rect 14182 19660 14188 19712
rect 14240 19700 14246 19712
rect 14277 19703 14335 19709
rect 14277 19700 14289 19703
rect 14240 19672 14289 19700
rect 14240 19660 14246 19672
rect 14277 19669 14289 19672
rect 14323 19700 14335 19703
rect 14550 19700 14556 19712
rect 14323 19672 14556 19700
rect 14323 19669 14335 19672
rect 14277 19663 14335 19669
rect 14550 19660 14556 19672
rect 14608 19660 14614 19712
rect 14642 19660 14648 19712
rect 14700 19700 14706 19712
rect 15764 19700 15792 19740
rect 21174 19728 21180 19780
rect 21232 19768 21238 19780
rect 21232 19740 27108 19768
rect 21232 19728 21238 19740
rect 14700 19672 15792 19700
rect 14700 19660 14706 19672
rect 16666 19660 16672 19712
rect 16724 19700 16730 19712
rect 17770 19700 17776 19712
rect 16724 19672 17776 19700
rect 16724 19660 16730 19672
rect 17770 19660 17776 19672
rect 17828 19660 17834 19712
rect 19886 19660 19892 19712
rect 19944 19700 19950 19712
rect 25222 19700 25228 19712
rect 19944 19672 25228 19700
rect 19944 19660 19950 19672
rect 25222 19660 25228 19672
rect 25280 19660 25286 19712
rect 25314 19660 25320 19712
rect 25372 19700 25378 19712
rect 25961 19703 26019 19709
rect 25961 19700 25973 19703
rect 25372 19672 25973 19700
rect 25372 19660 25378 19672
rect 25961 19669 25973 19672
rect 26007 19700 26019 19703
rect 26050 19700 26056 19712
rect 26007 19672 26056 19700
rect 26007 19669 26019 19672
rect 25961 19663 26019 19669
rect 26050 19660 26056 19672
rect 26108 19660 26114 19712
rect 27080 19709 27108 19740
rect 27065 19703 27123 19709
rect 27065 19669 27077 19703
rect 27111 19669 27123 19703
rect 27908 19700 27936 19808
rect 27982 19796 27988 19848
rect 28040 19796 28046 19848
rect 28810 19796 28816 19848
rect 28868 19836 28874 19848
rect 28868 19808 29316 19836
rect 28868 19796 28874 19808
rect 28074 19728 28080 19780
rect 28132 19768 28138 19780
rect 28445 19771 28503 19777
rect 28445 19768 28457 19771
rect 28132 19740 28457 19768
rect 28132 19728 28138 19740
rect 28445 19737 28457 19740
rect 28491 19737 28503 19771
rect 28445 19731 28503 19737
rect 28626 19728 28632 19780
rect 28684 19728 28690 19780
rect 29178 19768 29184 19780
rect 28736 19740 29184 19768
rect 28353 19703 28411 19709
rect 28353 19700 28365 19703
rect 27908 19672 28365 19700
rect 27065 19663 27123 19669
rect 28353 19669 28365 19672
rect 28399 19700 28411 19703
rect 28736 19700 28764 19740
rect 29178 19728 29184 19740
rect 29236 19728 29242 19780
rect 29288 19768 29316 19808
rect 29362 19796 29368 19848
rect 29420 19836 29426 19848
rect 30208 19845 30236 19876
rect 30285 19873 30297 19907
rect 30331 19873 30343 19907
rect 30285 19867 30343 19873
rect 29549 19839 29607 19845
rect 29549 19836 29561 19839
rect 29420 19808 29561 19836
rect 29420 19796 29426 19808
rect 29549 19805 29561 19808
rect 29595 19805 29607 19839
rect 29549 19799 29607 19805
rect 29641 19839 29699 19845
rect 29641 19805 29653 19839
rect 29687 19805 29699 19839
rect 29641 19799 29699 19805
rect 30193 19839 30251 19845
rect 30193 19805 30205 19839
rect 30239 19805 30251 19839
rect 30193 19799 30251 19805
rect 29656 19768 29684 19799
rect 30374 19796 30380 19848
rect 30432 19836 30438 19848
rect 30653 19839 30711 19845
rect 30653 19836 30665 19839
rect 30432 19808 30665 19836
rect 30432 19796 30438 19808
rect 30653 19805 30665 19808
rect 30699 19805 30711 19839
rect 30653 19799 30711 19805
rect 31110 19796 31116 19848
rect 31168 19796 31174 19848
rect 31202 19796 31208 19848
rect 31260 19836 31266 19848
rect 31369 19839 31427 19845
rect 31369 19836 31381 19839
rect 31260 19808 31381 19836
rect 31260 19796 31266 19808
rect 31369 19805 31381 19808
rect 31415 19805 31427 19839
rect 31369 19799 31427 19805
rect 30009 19771 30067 19777
rect 30009 19768 30021 19771
rect 29288 19740 30021 19768
rect 30009 19737 30021 19740
rect 30055 19737 30067 19771
rect 30009 19731 30067 19737
rect 28399 19672 28764 19700
rect 28813 19703 28871 19709
rect 28399 19669 28411 19672
rect 28353 19663 28411 19669
rect 28813 19669 28825 19703
rect 28859 19700 28871 19703
rect 28994 19700 29000 19712
rect 28859 19672 29000 19700
rect 28859 19669 28871 19672
rect 28813 19663 28871 19669
rect 28994 19660 29000 19672
rect 29052 19660 29058 19712
rect 30098 19660 30104 19712
rect 30156 19700 30162 19712
rect 30558 19700 30564 19712
rect 30156 19672 30564 19700
rect 30156 19660 30162 19672
rect 30558 19660 30564 19672
rect 30616 19660 30622 19712
rect 1104 19610 32844 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 32844 19610
rect 1104 19536 32844 19558
rect 1581 19499 1639 19505
rect 1581 19465 1593 19499
rect 1627 19496 1639 19499
rect 1670 19496 1676 19508
rect 1627 19468 1676 19496
rect 1627 19465 1639 19468
rect 1581 19459 1639 19465
rect 1670 19456 1676 19468
rect 1728 19456 1734 19508
rect 2774 19456 2780 19508
rect 2832 19496 2838 19508
rect 3786 19496 3792 19508
rect 2832 19468 3792 19496
rect 2832 19456 2838 19468
rect 3786 19456 3792 19468
rect 3844 19456 3850 19508
rect 4338 19456 4344 19508
rect 4396 19496 4402 19508
rect 4525 19499 4583 19505
rect 4525 19496 4537 19499
rect 4396 19468 4537 19496
rect 4396 19456 4402 19468
rect 4525 19465 4537 19468
rect 4571 19496 4583 19499
rect 7374 19496 7380 19508
rect 4571 19468 7380 19496
rect 4571 19465 4583 19468
rect 4525 19459 4583 19465
rect 7374 19456 7380 19468
rect 7432 19456 7438 19508
rect 7650 19456 7656 19508
rect 7708 19496 7714 19508
rect 10502 19496 10508 19508
rect 7708 19468 10508 19496
rect 7708 19456 7714 19468
rect 10502 19456 10508 19468
rect 10560 19456 10566 19508
rect 11517 19499 11575 19505
rect 11517 19465 11529 19499
rect 11563 19496 11575 19499
rect 11563 19468 12020 19496
rect 11563 19465 11575 19468
rect 11517 19459 11575 19465
rect 4614 19428 4620 19440
rect 4448 19400 4620 19428
rect 1302 19320 1308 19372
rect 1360 19360 1366 19372
rect 1397 19363 1455 19369
rect 1397 19360 1409 19363
rect 1360 19332 1409 19360
rect 1360 19320 1366 19332
rect 1397 19329 1409 19332
rect 1443 19329 1455 19363
rect 1397 19323 1455 19329
rect 4062 19320 4068 19372
rect 4120 19320 4126 19372
rect 4448 19369 4476 19400
rect 4614 19388 4620 19400
rect 4672 19388 4678 19440
rect 7466 19388 7472 19440
rect 7524 19428 7530 19440
rect 7561 19431 7619 19437
rect 7561 19428 7573 19431
rect 7524 19400 7573 19428
rect 7524 19388 7530 19400
rect 7561 19397 7573 19400
rect 7607 19397 7619 19431
rect 7561 19391 7619 19397
rect 8110 19388 8116 19440
rect 8168 19428 8174 19440
rect 8570 19428 8576 19440
rect 8168 19400 8576 19428
rect 8168 19388 8174 19400
rect 8570 19388 8576 19400
rect 8628 19388 8634 19440
rect 8754 19388 8760 19440
rect 8812 19428 8818 19440
rect 9674 19428 9680 19440
rect 8812 19400 9680 19428
rect 8812 19388 8818 19400
rect 9674 19388 9680 19400
rect 9732 19388 9738 19440
rect 9950 19388 9956 19440
rect 10008 19428 10014 19440
rect 10870 19428 10876 19440
rect 10008 19400 10876 19428
rect 10008 19388 10014 19400
rect 10870 19388 10876 19400
rect 10928 19388 10934 19440
rect 11146 19388 11152 19440
rect 11204 19388 11210 19440
rect 11992 19437 12020 19468
rect 12802 19456 12808 19508
rect 12860 19496 12866 19508
rect 13262 19496 13268 19508
rect 12860 19468 13268 19496
rect 12860 19456 12866 19468
rect 13262 19456 13268 19468
rect 13320 19456 13326 19508
rect 13354 19456 13360 19508
rect 13412 19456 13418 19508
rect 13633 19499 13691 19505
rect 13633 19465 13645 19499
rect 13679 19496 13691 19499
rect 13814 19496 13820 19508
rect 13679 19468 13820 19496
rect 13679 19465 13691 19468
rect 13633 19459 13691 19465
rect 13814 19456 13820 19468
rect 13872 19496 13878 19508
rect 14918 19496 14924 19508
rect 13872 19468 14924 19496
rect 13872 19456 13878 19468
rect 14918 19456 14924 19468
rect 14976 19456 14982 19508
rect 16206 19456 16212 19508
rect 16264 19456 16270 19508
rect 16482 19456 16488 19508
rect 16540 19496 16546 19508
rect 17586 19496 17592 19508
rect 16540 19468 17592 19496
rect 16540 19456 16546 19468
rect 17586 19456 17592 19468
rect 17644 19456 17650 19508
rect 18966 19456 18972 19508
rect 19024 19496 19030 19508
rect 20625 19499 20683 19505
rect 20625 19496 20637 19499
rect 19024 19468 20637 19496
rect 19024 19456 19030 19468
rect 20625 19465 20637 19468
rect 20671 19496 20683 19499
rect 23934 19496 23940 19508
rect 20671 19468 23940 19496
rect 20671 19465 20683 19468
rect 20625 19459 20683 19465
rect 23934 19456 23940 19468
rect 23992 19456 23998 19508
rect 24121 19499 24179 19505
rect 24121 19465 24133 19499
rect 24167 19496 24179 19499
rect 24857 19499 24915 19505
rect 24167 19468 24624 19496
rect 24167 19465 24179 19468
rect 24121 19459 24179 19465
rect 11977 19431 12035 19437
rect 11977 19397 11989 19431
rect 12023 19397 12035 19431
rect 13372 19428 13400 19456
rect 14093 19431 14151 19437
rect 14093 19428 14105 19431
rect 13372 19400 14105 19428
rect 11977 19391 12035 19397
rect 14093 19397 14105 19400
rect 14139 19397 14151 19431
rect 14093 19391 14151 19397
rect 14642 19388 14648 19440
rect 14700 19428 14706 19440
rect 14700 19400 14872 19428
rect 14700 19388 14706 19400
rect 4433 19363 4491 19369
rect 4433 19329 4445 19363
rect 4479 19329 4491 19363
rect 4433 19323 4491 19329
rect 4709 19363 4767 19369
rect 4709 19329 4721 19363
rect 4755 19360 4767 19363
rect 5074 19360 5080 19372
rect 4755 19332 5080 19360
rect 4755 19329 4767 19332
rect 4709 19323 4767 19329
rect 5074 19320 5080 19332
rect 5132 19320 5138 19372
rect 5261 19347 5319 19353
rect 5261 19344 5273 19347
rect 5184 19316 5273 19344
rect 3970 19252 3976 19304
rect 4028 19292 4034 19304
rect 4028 19264 5120 19292
rect 4028 19252 4034 19264
rect 3602 19184 3608 19236
rect 3660 19224 3666 19236
rect 5092 19233 5120 19264
rect 5077 19227 5135 19233
rect 3660 19196 5028 19224
rect 3660 19184 3666 19196
rect 1210 19116 1216 19168
rect 1268 19156 1274 19168
rect 3142 19156 3148 19168
rect 1268 19128 3148 19156
rect 1268 19116 1274 19128
rect 3142 19116 3148 19128
rect 3200 19116 3206 19168
rect 3881 19159 3939 19165
rect 3881 19125 3893 19159
rect 3927 19156 3939 19159
rect 4062 19156 4068 19168
rect 3927 19128 4068 19156
rect 3927 19125 3939 19128
rect 3881 19119 3939 19125
rect 4062 19116 4068 19128
rect 4120 19116 4126 19168
rect 4249 19159 4307 19165
rect 4249 19125 4261 19159
rect 4295 19156 4307 19159
rect 4798 19156 4804 19168
rect 4295 19128 4804 19156
rect 4295 19125 4307 19128
rect 4249 19119 4307 19125
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 5000 19156 5028 19196
rect 5077 19193 5089 19227
rect 5123 19193 5135 19227
rect 5077 19187 5135 19193
rect 5184 19156 5212 19316
rect 5261 19313 5273 19316
rect 5307 19313 5319 19347
rect 5261 19307 5319 19313
rect 7484 19332 8064 19360
rect 5994 19252 6000 19304
rect 6052 19292 6058 19304
rect 7484 19292 7512 19332
rect 6052 19264 7512 19292
rect 6052 19252 6058 19264
rect 7558 19252 7564 19304
rect 7616 19292 7622 19304
rect 7926 19292 7932 19304
rect 7616 19264 7932 19292
rect 7616 19252 7622 19264
rect 7926 19252 7932 19264
rect 7984 19252 7990 19304
rect 8036 19292 8064 19332
rect 10226 19320 10232 19372
rect 10284 19360 10290 19372
rect 11164 19360 11192 19388
rect 11701 19363 11759 19369
rect 11701 19360 11713 19363
rect 10284 19332 11192 19360
rect 11532 19332 11713 19360
rect 10284 19320 10290 19332
rect 11532 19304 11560 19332
rect 11701 19329 11713 19332
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 11882 19320 11888 19372
rect 11940 19320 11946 19372
rect 12066 19320 12072 19372
rect 12124 19360 12130 19372
rect 12253 19363 12311 19369
rect 12253 19360 12265 19363
rect 12124 19332 12265 19360
rect 12124 19320 12130 19332
rect 12253 19329 12265 19332
rect 12299 19329 12311 19363
rect 12253 19323 12311 19329
rect 12526 19320 12532 19372
rect 12584 19360 12590 19372
rect 13357 19363 13415 19369
rect 13357 19360 13369 19363
rect 12584 19332 13369 19360
rect 12584 19320 12590 19332
rect 13357 19329 13369 19332
rect 13403 19329 13415 19363
rect 13817 19363 13875 19369
rect 13817 19360 13829 19363
rect 13357 19323 13415 19329
rect 13740 19332 13829 19360
rect 11146 19292 11152 19304
rect 8036 19264 11152 19292
rect 11146 19252 11152 19264
rect 11204 19252 11210 19304
rect 11514 19252 11520 19304
rect 11572 19252 11578 19304
rect 11974 19292 11980 19304
rect 11716 19264 11980 19292
rect 7466 19184 7472 19236
rect 7524 19224 7530 19236
rect 9950 19224 9956 19236
rect 7524 19196 9956 19224
rect 7524 19184 7530 19196
rect 9950 19184 9956 19196
rect 10008 19184 10014 19236
rect 11716 19224 11744 19264
rect 11974 19252 11980 19264
rect 12032 19252 12038 19304
rect 12161 19295 12219 19301
rect 12161 19292 12173 19295
rect 12084 19264 12173 19292
rect 12084 19236 12112 19264
rect 12161 19261 12173 19264
rect 12207 19261 12219 19295
rect 12161 19255 12219 19261
rect 13262 19252 13268 19304
rect 13320 19292 13326 19304
rect 13740 19292 13768 19332
rect 13817 19329 13829 19332
rect 13863 19329 13875 19363
rect 13817 19323 13875 19329
rect 14001 19363 14059 19369
rect 14001 19329 14013 19363
rect 14047 19360 14059 19363
rect 14182 19360 14188 19372
rect 14047 19332 14188 19360
rect 14047 19329 14059 19332
rect 14001 19323 14059 19329
rect 14182 19320 14188 19332
rect 14240 19320 14246 19372
rect 14277 19363 14335 19369
rect 14277 19329 14289 19363
rect 14323 19360 14335 19363
rect 14660 19360 14688 19388
rect 14323 19332 14688 19360
rect 14737 19363 14795 19369
rect 14323 19329 14335 19332
rect 14277 19323 14335 19329
rect 14737 19329 14749 19363
rect 14783 19329 14795 19363
rect 14737 19323 14795 19329
rect 13320 19264 13768 19292
rect 13320 19252 13326 19264
rect 13906 19252 13912 19304
rect 13964 19292 13970 19304
rect 14553 19295 14611 19301
rect 14553 19292 14565 19295
rect 13964 19264 14565 19292
rect 13964 19252 13970 19264
rect 14553 19261 14565 19264
rect 14599 19292 14611 19295
rect 14752 19292 14780 19323
rect 14599 19264 14780 19292
rect 14844 19292 14872 19400
rect 15010 19388 15016 19440
rect 15068 19388 15074 19440
rect 15194 19344 15200 19396
rect 15252 19344 15258 19396
rect 15746 19388 15752 19440
rect 15804 19437 15810 19440
rect 15804 19391 15814 19437
rect 19797 19431 19855 19437
rect 19797 19397 19809 19431
rect 19843 19428 19855 19431
rect 20162 19428 20168 19440
rect 19843 19400 20168 19428
rect 19843 19397 19855 19400
rect 19797 19391 19855 19397
rect 15804 19388 15810 19391
rect 20162 19388 20168 19400
rect 20220 19388 20226 19440
rect 20346 19388 20352 19440
rect 20404 19428 20410 19440
rect 20404 19400 23888 19428
rect 20404 19388 20410 19400
rect 15197 19329 15209 19344
rect 15243 19329 15255 19344
rect 15197 19323 15255 19329
rect 15286 19320 15292 19372
rect 15344 19369 15350 19372
rect 15344 19363 15363 19369
rect 15351 19329 15363 19363
rect 15933 19363 15991 19369
rect 15933 19360 15945 19363
rect 15344 19323 15363 19329
rect 15580 19332 15945 19360
rect 15344 19320 15350 19323
rect 14844 19264 14964 19292
rect 14599 19261 14611 19264
rect 14553 19255 14611 19261
rect 10888 19196 11744 19224
rect 5000 19128 5212 19156
rect 6546 19116 6552 19168
rect 6604 19156 6610 19168
rect 7653 19159 7711 19165
rect 7653 19156 7665 19159
rect 6604 19128 7665 19156
rect 6604 19116 6610 19128
rect 7653 19125 7665 19128
rect 7699 19125 7711 19159
rect 7653 19119 7711 19125
rect 8478 19116 8484 19168
rect 8536 19156 8542 19168
rect 10888 19156 10916 19196
rect 12066 19184 12072 19236
rect 12124 19184 12130 19236
rect 12437 19227 12495 19233
rect 12437 19193 12449 19227
rect 12483 19224 12495 19227
rect 13078 19224 13084 19236
rect 12483 19196 13084 19224
rect 12483 19193 12495 19196
rect 12437 19187 12495 19193
rect 13078 19184 13084 19196
rect 13136 19184 13142 19236
rect 13541 19227 13599 19233
rect 13541 19193 13553 19227
rect 13587 19224 13599 19227
rect 14182 19224 14188 19236
rect 13587 19196 14188 19224
rect 13587 19193 13599 19196
rect 13541 19187 13599 19193
rect 14182 19184 14188 19196
rect 14240 19184 14246 19236
rect 14826 19224 14832 19236
rect 14384 19196 14832 19224
rect 8536 19128 10916 19156
rect 8536 19116 8542 19128
rect 10962 19116 10968 19168
rect 11020 19156 11026 19168
rect 11885 19159 11943 19165
rect 11885 19156 11897 19159
rect 11020 19128 11897 19156
rect 11020 19116 11026 19128
rect 11885 19125 11897 19128
rect 11931 19156 11943 19159
rect 11974 19156 11980 19168
rect 11931 19128 11980 19156
rect 11931 19125 11943 19128
rect 11885 19119 11943 19125
rect 11974 19116 11980 19128
rect 12032 19116 12038 19168
rect 12253 19159 12311 19165
rect 12253 19125 12265 19159
rect 12299 19156 12311 19159
rect 12618 19156 12624 19168
rect 12299 19128 12624 19156
rect 12299 19125 12311 19128
rect 12253 19119 12311 19125
rect 12618 19116 12624 19128
rect 12676 19116 12682 19168
rect 13814 19116 13820 19168
rect 13872 19156 13878 19168
rect 14384 19156 14412 19196
rect 14826 19184 14832 19196
rect 14884 19184 14890 19236
rect 14936 19233 14964 19264
rect 14921 19227 14979 19233
rect 14921 19193 14933 19227
rect 14967 19193 14979 19227
rect 14921 19187 14979 19193
rect 15473 19227 15531 19233
rect 15473 19193 15485 19227
rect 15519 19224 15531 19227
rect 15580 19224 15608 19332
rect 15933 19329 15945 19332
rect 15979 19329 15991 19363
rect 15933 19323 15991 19329
rect 16022 19320 16028 19372
rect 16080 19320 16086 19372
rect 17678 19320 17684 19372
rect 17736 19360 17742 19372
rect 18046 19360 18052 19372
rect 17736 19332 18052 19360
rect 17736 19320 17742 19332
rect 18046 19320 18052 19332
rect 18104 19320 18110 19372
rect 19978 19320 19984 19372
rect 20036 19320 20042 19372
rect 20257 19363 20315 19369
rect 20257 19329 20269 19363
rect 20303 19360 20315 19363
rect 20438 19360 20444 19372
rect 20303 19332 20444 19360
rect 20303 19329 20315 19332
rect 20257 19323 20315 19329
rect 20438 19320 20444 19332
rect 20496 19320 20502 19372
rect 22554 19320 22560 19372
rect 22612 19360 22618 19372
rect 22741 19363 22799 19369
rect 22741 19360 22753 19363
rect 22612 19332 22753 19360
rect 22612 19320 22618 19332
rect 22741 19329 22753 19332
rect 22787 19329 22799 19363
rect 22741 19323 22799 19329
rect 23014 19320 23020 19372
rect 23072 19360 23078 19372
rect 23860 19369 23888 19400
rect 23661 19363 23719 19369
rect 23661 19360 23673 19363
rect 23072 19332 23673 19360
rect 23072 19320 23078 19332
rect 23661 19329 23673 19332
rect 23707 19329 23719 19363
rect 23661 19323 23719 19329
rect 23845 19363 23903 19369
rect 23845 19329 23857 19363
rect 23891 19329 23903 19363
rect 23845 19323 23903 19329
rect 23937 19363 23995 19369
rect 23937 19329 23949 19363
rect 23983 19360 23995 19363
rect 24397 19363 24455 19369
rect 23983 19332 24348 19360
rect 23983 19329 23995 19332
rect 23937 19323 23995 19329
rect 15657 19295 15715 19301
rect 15657 19261 15669 19295
rect 15703 19292 15715 19295
rect 16040 19292 16068 19320
rect 15703 19264 16068 19292
rect 15703 19261 15715 19264
rect 15657 19255 15715 19261
rect 16574 19252 16580 19304
rect 16632 19292 16638 19304
rect 20162 19292 20168 19304
rect 16632 19264 20168 19292
rect 16632 19252 16638 19264
rect 20162 19252 20168 19264
rect 20220 19252 20226 19304
rect 20349 19295 20407 19301
rect 20349 19261 20361 19295
rect 20395 19292 20407 19295
rect 20806 19292 20812 19304
rect 20395 19264 20812 19292
rect 20395 19261 20407 19264
rect 20349 19255 20407 19261
rect 20456 19236 20484 19264
rect 20806 19252 20812 19264
rect 20864 19252 20870 19304
rect 24320 19292 24348 19332
rect 24397 19329 24409 19363
rect 24443 19360 24455 19363
rect 24486 19360 24492 19372
rect 24443 19332 24492 19360
rect 24443 19329 24455 19332
rect 24397 19323 24455 19329
rect 24486 19320 24492 19332
rect 24544 19320 24550 19372
rect 24596 19369 24624 19468
rect 24857 19465 24869 19499
rect 24903 19496 24915 19499
rect 26605 19499 26663 19505
rect 24903 19468 26556 19496
rect 24903 19465 24915 19468
rect 24857 19459 24915 19465
rect 25038 19388 25044 19440
rect 25096 19428 25102 19440
rect 25222 19428 25228 19440
rect 25096 19400 25228 19428
rect 25096 19388 25102 19400
rect 25222 19388 25228 19400
rect 25280 19388 25286 19440
rect 26528 19428 26556 19468
rect 26605 19465 26617 19499
rect 26651 19496 26663 19499
rect 28166 19496 28172 19508
rect 26651 19468 28172 19496
rect 26651 19465 26663 19468
rect 26605 19459 26663 19465
rect 28166 19456 28172 19468
rect 28224 19456 28230 19508
rect 29362 19456 29368 19508
rect 29420 19456 29426 19508
rect 30285 19499 30343 19505
rect 30285 19465 30297 19499
rect 30331 19496 30343 19499
rect 30374 19496 30380 19508
rect 30331 19468 30380 19496
rect 30331 19465 30343 19468
rect 30285 19459 30343 19465
rect 30374 19456 30380 19468
rect 30432 19456 30438 19508
rect 31018 19496 31024 19508
rect 30944 19468 31024 19496
rect 26878 19428 26884 19440
rect 26528 19400 26884 19428
rect 26878 19388 26884 19400
rect 26936 19388 26942 19440
rect 28718 19388 28724 19440
rect 28776 19428 28782 19440
rect 28905 19431 28963 19437
rect 28905 19428 28917 19431
rect 28776 19400 28917 19428
rect 28776 19388 28782 19400
rect 28905 19397 28917 19400
rect 28951 19397 28963 19431
rect 29454 19428 29460 19440
rect 28905 19391 28963 19397
rect 29104 19400 29460 19428
rect 24581 19363 24639 19369
rect 24581 19329 24593 19363
rect 24627 19329 24639 19363
rect 24581 19323 24639 19329
rect 24673 19363 24731 19369
rect 24673 19329 24685 19363
rect 24719 19360 24731 19363
rect 24762 19360 24768 19372
rect 24719 19332 24768 19360
rect 24719 19329 24731 19332
rect 24673 19323 24731 19329
rect 24762 19320 24768 19332
rect 24820 19320 24826 19372
rect 25593 19363 25651 19369
rect 25593 19329 25605 19363
rect 25639 19360 25651 19363
rect 25639 19332 25728 19360
rect 25639 19329 25651 19332
rect 25593 19323 25651 19329
rect 25038 19292 25044 19304
rect 24320 19264 25044 19292
rect 25038 19252 25044 19264
rect 25096 19252 25102 19304
rect 25700 19292 25728 19332
rect 25774 19320 25780 19372
rect 25832 19320 25838 19372
rect 25869 19363 25927 19369
rect 25869 19329 25881 19363
rect 25915 19360 25927 19363
rect 25958 19360 25964 19372
rect 25915 19332 25964 19360
rect 25915 19329 25927 19332
rect 25869 19323 25927 19329
rect 25958 19320 25964 19332
rect 26016 19320 26022 19372
rect 26050 19320 26056 19372
rect 26108 19360 26114 19372
rect 26145 19363 26203 19369
rect 26145 19360 26157 19363
rect 26108 19332 26157 19360
rect 26108 19320 26114 19332
rect 26145 19329 26157 19332
rect 26191 19329 26203 19363
rect 26145 19323 26203 19329
rect 26234 19320 26240 19372
rect 26292 19360 26298 19372
rect 26329 19363 26387 19369
rect 26329 19360 26341 19363
rect 26292 19332 26341 19360
rect 26292 19320 26298 19332
rect 26329 19329 26341 19332
rect 26375 19329 26387 19363
rect 26329 19323 26387 19329
rect 26418 19320 26424 19372
rect 26476 19320 26482 19372
rect 26786 19360 26792 19372
rect 26528 19332 26792 19360
rect 26528 19292 26556 19332
rect 26786 19320 26792 19332
rect 26844 19320 26850 19372
rect 27709 19363 27767 19369
rect 27709 19329 27721 19363
rect 27755 19360 27767 19363
rect 28074 19360 28080 19372
rect 27755 19332 28080 19360
rect 27755 19329 27767 19332
rect 27709 19323 27767 19329
rect 28074 19320 28080 19332
rect 28132 19320 28138 19372
rect 25700 19264 26556 19292
rect 27522 19252 27528 19304
rect 27580 19292 27586 19304
rect 27801 19295 27859 19301
rect 27801 19292 27813 19295
rect 27580 19264 27813 19292
rect 27580 19252 27586 19264
rect 27801 19261 27813 19264
rect 27847 19261 27859 19295
rect 28920 19292 28948 19391
rect 28994 19320 29000 19372
rect 29052 19360 29058 19372
rect 29104 19369 29132 19400
rect 29454 19388 29460 19400
rect 29512 19388 29518 19440
rect 30466 19388 30472 19440
rect 30524 19428 30530 19440
rect 30944 19437 30972 19468
rect 31018 19456 31024 19468
rect 31076 19456 31082 19508
rect 32398 19456 32404 19508
rect 32456 19456 32462 19508
rect 30837 19431 30895 19437
rect 30837 19428 30849 19431
rect 30524 19400 30849 19428
rect 30524 19388 30530 19400
rect 30837 19397 30849 19400
rect 30883 19397 30895 19431
rect 30837 19391 30895 19397
rect 30929 19431 30987 19437
rect 30929 19397 30941 19431
rect 30975 19397 30987 19431
rect 30929 19391 30987 19397
rect 29089 19363 29147 19369
rect 29089 19360 29101 19363
rect 29052 19332 29101 19360
rect 29052 19320 29058 19332
rect 29089 19329 29101 19332
rect 29135 19329 29147 19363
rect 29089 19323 29147 19329
rect 29178 19320 29184 19372
rect 29236 19320 29242 19372
rect 29638 19320 29644 19372
rect 29696 19360 29702 19372
rect 30101 19363 30159 19369
rect 30101 19360 30113 19363
rect 29696 19332 30113 19360
rect 29696 19320 29702 19332
rect 30101 19329 30113 19332
rect 30147 19360 30159 19363
rect 30147 19332 30420 19360
rect 30147 19329 30159 19332
rect 30101 19323 30159 19329
rect 28920 19264 29040 19292
rect 27801 19255 27859 19261
rect 29012 19236 29040 19264
rect 16301 19227 16359 19233
rect 16301 19224 16313 19227
rect 15519 19196 15608 19224
rect 15764 19196 16313 19224
rect 15519 19193 15531 19196
rect 15473 19187 15531 19193
rect 13872 19128 14412 19156
rect 13872 19116 13878 19128
rect 14458 19116 14464 19168
rect 14516 19156 14522 19168
rect 15102 19156 15108 19168
rect 14516 19128 15108 19156
rect 14516 19116 14522 19128
rect 15102 19116 15108 19128
rect 15160 19116 15166 19168
rect 15194 19116 15200 19168
rect 15252 19156 15258 19168
rect 15764 19165 15792 19196
rect 16301 19193 16313 19196
rect 16347 19193 16359 19227
rect 16301 19187 16359 19193
rect 17770 19184 17776 19236
rect 17828 19224 17834 19236
rect 17828 19196 17954 19224
rect 17828 19184 17834 19196
rect 15749 19159 15807 19165
rect 15749 19156 15761 19159
rect 15252 19128 15761 19156
rect 15252 19116 15258 19128
rect 15749 19125 15761 19128
rect 15795 19125 15807 19159
rect 15749 19119 15807 19125
rect 16114 19116 16120 19168
rect 16172 19156 16178 19168
rect 17034 19156 17040 19168
rect 16172 19128 17040 19156
rect 16172 19116 16178 19128
rect 17034 19116 17040 19128
rect 17092 19116 17098 19168
rect 17926 19156 17954 19196
rect 18874 19184 18880 19236
rect 18932 19224 18938 19236
rect 19610 19224 19616 19236
rect 18932 19196 19616 19224
rect 18932 19184 18938 19196
rect 19610 19184 19616 19196
rect 19668 19184 19674 19236
rect 20070 19184 20076 19236
rect 20128 19224 20134 19236
rect 20128 19196 20300 19224
rect 20128 19184 20134 19196
rect 19886 19156 19892 19168
rect 17926 19128 19892 19156
rect 19886 19116 19892 19128
rect 19944 19116 19950 19168
rect 20162 19116 20168 19168
rect 20220 19116 20226 19168
rect 20272 19165 20300 19196
rect 20438 19184 20444 19236
rect 20496 19184 20502 19236
rect 20990 19184 20996 19236
rect 21048 19224 21054 19236
rect 28626 19224 28632 19236
rect 21048 19196 26372 19224
rect 21048 19184 21054 19196
rect 20257 19159 20315 19165
rect 20257 19125 20269 19159
rect 20303 19125 20315 19159
rect 20257 19119 20315 19125
rect 22370 19116 22376 19168
rect 22428 19156 22434 19168
rect 22738 19156 22744 19168
rect 22428 19128 22744 19156
rect 22428 19116 22434 19128
rect 22738 19116 22744 19128
rect 22796 19116 22802 19168
rect 22925 19159 22983 19165
rect 22925 19125 22937 19159
rect 22971 19156 22983 19159
rect 23566 19156 23572 19168
rect 22971 19128 23572 19156
rect 22971 19125 22983 19128
rect 22925 19119 22983 19125
rect 23566 19116 23572 19128
rect 23624 19116 23630 19168
rect 23934 19116 23940 19168
rect 23992 19116 23998 19168
rect 24394 19116 24400 19168
rect 24452 19116 24458 19168
rect 25866 19116 25872 19168
rect 25924 19116 25930 19168
rect 26053 19159 26111 19165
rect 26053 19125 26065 19159
rect 26099 19156 26111 19159
rect 26234 19156 26240 19168
rect 26099 19128 26240 19156
rect 26099 19125 26111 19128
rect 26053 19119 26111 19125
rect 26234 19116 26240 19128
rect 26292 19116 26298 19168
rect 26344 19165 26372 19196
rect 27816 19196 28632 19224
rect 27816 19165 27844 19196
rect 28626 19184 28632 19196
rect 28684 19184 28690 19236
rect 28994 19184 29000 19236
rect 29052 19184 29058 19236
rect 30392 19233 30420 19332
rect 30558 19320 30564 19372
rect 30616 19320 30622 19372
rect 30653 19363 30711 19369
rect 30653 19329 30665 19363
rect 30699 19360 30711 19363
rect 30742 19360 30748 19372
rect 30699 19332 30748 19360
rect 30699 19329 30711 19332
rect 30653 19323 30711 19329
rect 30742 19320 30748 19332
rect 30800 19320 30806 19372
rect 31021 19363 31079 19369
rect 31021 19329 31033 19363
rect 31067 19360 31079 19363
rect 31297 19363 31355 19369
rect 31297 19360 31309 19363
rect 31067 19332 31309 19360
rect 31067 19329 31079 19332
rect 31021 19323 31079 19329
rect 31297 19329 31309 19332
rect 31343 19329 31355 19363
rect 31297 19323 31355 19329
rect 32214 19320 32220 19372
rect 32272 19320 32278 19372
rect 31941 19295 31999 19301
rect 31941 19261 31953 19295
rect 31987 19292 31999 19295
rect 31987 19264 32904 19292
rect 31987 19261 31999 19264
rect 31941 19255 31999 19261
rect 30377 19227 30435 19233
rect 30377 19193 30389 19227
rect 30423 19193 30435 19227
rect 30377 19187 30435 19193
rect 26329 19159 26387 19165
rect 26329 19125 26341 19159
rect 26375 19125 26387 19159
rect 26329 19119 26387 19125
rect 27801 19159 27859 19165
rect 27801 19125 27813 19159
rect 27847 19125 27859 19159
rect 27801 19119 27859 19125
rect 27890 19116 27896 19168
rect 27948 19156 27954 19168
rect 28077 19159 28135 19165
rect 28077 19156 28089 19159
rect 27948 19128 28089 19156
rect 27948 19116 27954 19128
rect 28077 19125 28089 19128
rect 28123 19125 28135 19159
rect 28077 19119 28135 19125
rect 29181 19159 29239 19165
rect 29181 19125 29193 19159
rect 29227 19156 29239 19159
rect 29362 19156 29368 19168
rect 29227 19128 29368 19156
rect 29227 19125 29239 19128
rect 29181 19119 29239 19125
rect 29362 19116 29368 19128
rect 29420 19156 29426 19168
rect 29822 19156 29828 19168
rect 29420 19128 29828 19156
rect 29420 19116 29426 19128
rect 29822 19116 29828 19128
rect 29880 19116 29886 19168
rect 31202 19116 31208 19168
rect 31260 19116 31266 19168
rect 1104 19066 32844 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 32844 19066
rect 1104 18992 32844 19014
rect 2038 18912 2044 18964
rect 2096 18952 2102 18964
rect 2777 18955 2835 18961
rect 2777 18952 2789 18955
rect 2096 18924 2789 18952
rect 2096 18912 2102 18924
rect 2777 18921 2789 18924
rect 2823 18921 2835 18955
rect 2777 18915 2835 18921
rect 6825 18955 6883 18961
rect 6825 18921 6837 18955
rect 6871 18952 6883 18955
rect 7466 18952 7472 18964
rect 6871 18924 7472 18952
rect 6871 18921 6883 18924
rect 6825 18915 6883 18921
rect 7466 18912 7472 18924
rect 7524 18912 7530 18964
rect 7650 18912 7656 18964
rect 7708 18952 7714 18964
rect 7929 18955 7987 18961
rect 7929 18952 7941 18955
rect 7708 18924 7941 18952
rect 7708 18912 7714 18924
rect 7929 18921 7941 18924
rect 7975 18921 7987 18955
rect 9217 18955 9275 18961
rect 9217 18952 9229 18955
rect 7929 18915 7987 18921
rect 8036 18924 9229 18952
rect 8036 18884 8064 18924
rect 9217 18921 9229 18924
rect 9263 18921 9275 18955
rect 9217 18915 9275 18921
rect 9953 18955 10011 18961
rect 9953 18921 9965 18955
rect 9999 18952 10011 18955
rect 9999 18924 10180 18952
rect 9999 18921 10011 18924
rect 9953 18915 10011 18921
rect 2746 18856 8064 18884
rect 8297 18887 8355 18893
rect 1394 18776 1400 18828
rect 1452 18776 1458 18828
rect 1302 18708 1308 18760
rect 1360 18748 1366 18760
rect 2746 18748 2774 18856
rect 8297 18853 8309 18887
rect 8343 18884 8355 18887
rect 9677 18887 9735 18893
rect 8343 18856 9352 18884
rect 8343 18853 8355 18856
rect 8297 18847 8355 18853
rect 4338 18816 4344 18828
rect 4264 18788 4344 18816
rect 1360 18720 2774 18748
rect 1360 18708 1366 18720
rect 3326 18708 3332 18760
rect 3384 18708 3390 18760
rect 3418 18708 3424 18760
rect 3476 18708 3482 18760
rect 3973 18751 4031 18757
rect 3973 18717 3985 18751
rect 4019 18748 4031 18751
rect 4062 18748 4068 18760
rect 4019 18720 4068 18748
rect 4019 18717 4031 18720
rect 3973 18711 4031 18717
rect 4062 18708 4068 18720
rect 4120 18708 4126 18760
rect 4264 18757 4292 18788
rect 4338 18776 4344 18788
rect 4396 18816 4402 18828
rect 4706 18816 4712 18828
rect 4396 18788 4712 18816
rect 4396 18776 4402 18788
rect 4706 18776 4712 18788
rect 4764 18776 4770 18828
rect 5074 18776 5080 18828
rect 5132 18816 5138 18828
rect 6178 18816 6184 18828
rect 5132 18788 6184 18816
rect 5132 18776 5138 18788
rect 4249 18751 4307 18757
rect 4249 18717 4261 18751
rect 4295 18717 4307 18751
rect 4249 18711 4307 18717
rect 4433 18751 4491 18757
rect 4433 18717 4445 18751
rect 4479 18748 4491 18751
rect 4798 18748 4804 18760
rect 4479 18720 4804 18748
rect 4479 18717 4491 18720
rect 4433 18711 4491 18717
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 5353 18751 5411 18757
rect 5353 18717 5365 18751
rect 5399 18748 5411 18751
rect 5442 18748 5448 18760
rect 5399 18720 5448 18748
rect 5399 18717 5411 18720
rect 5353 18711 5411 18717
rect 5442 18708 5448 18720
rect 5500 18708 5506 18760
rect 5920 18757 5948 18788
rect 6178 18776 6184 18788
rect 6236 18776 6242 18828
rect 6730 18816 6736 18828
rect 6380 18788 6736 18816
rect 5905 18751 5963 18757
rect 5905 18717 5917 18751
rect 5951 18717 5963 18751
rect 5905 18711 5963 18717
rect 6086 18708 6092 18760
rect 6144 18708 6150 18760
rect 6380 18757 6408 18788
rect 6730 18776 6736 18788
rect 6788 18776 6794 18828
rect 8021 18819 8079 18825
rect 8021 18785 8033 18819
rect 8067 18816 8079 18819
rect 8202 18816 8208 18828
rect 8067 18788 8208 18816
rect 8067 18785 8079 18788
rect 8021 18779 8079 18785
rect 8202 18776 8208 18788
rect 8260 18776 8266 18828
rect 9324 18825 9352 18856
rect 9677 18853 9689 18887
rect 9723 18884 9735 18887
rect 10042 18884 10048 18896
rect 9723 18856 10048 18884
rect 9723 18853 9735 18856
rect 9677 18847 9735 18853
rect 10042 18844 10048 18856
rect 10100 18844 10106 18896
rect 10152 18884 10180 18924
rect 10226 18912 10232 18964
rect 10284 18912 10290 18964
rect 10502 18912 10508 18964
rect 10560 18912 10566 18964
rect 11146 18912 11152 18964
rect 11204 18952 11210 18964
rect 11609 18955 11667 18961
rect 11609 18952 11621 18955
rect 11204 18924 11621 18952
rect 11204 18912 11210 18924
rect 11609 18921 11621 18924
rect 11655 18921 11667 18955
rect 11609 18915 11667 18921
rect 11882 18912 11888 18964
rect 11940 18952 11946 18964
rect 11940 18924 12020 18952
rect 11940 18912 11946 18924
rect 10520 18884 10548 18912
rect 10152 18856 10548 18884
rect 10594 18844 10600 18896
rect 10652 18884 10658 18896
rect 11992 18884 12020 18924
rect 12066 18912 12072 18964
rect 12124 18912 12130 18964
rect 12618 18912 12624 18964
rect 12676 18952 12682 18964
rect 13262 18952 13268 18964
rect 12676 18924 13268 18952
rect 12676 18912 12682 18924
rect 13262 18912 13268 18924
rect 13320 18912 13326 18964
rect 14090 18912 14096 18964
rect 14148 18952 14154 18964
rect 14458 18952 14464 18964
rect 14148 18924 14464 18952
rect 14148 18912 14154 18924
rect 14458 18912 14464 18924
rect 14516 18912 14522 18964
rect 14553 18955 14611 18961
rect 14553 18921 14565 18955
rect 14599 18952 14611 18955
rect 15010 18952 15016 18964
rect 14599 18924 15016 18952
rect 14599 18921 14611 18924
rect 14553 18915 14611 18921
rect 15010 18912 15016 18924
rect 15068 18912 15074 18964
rect 16482 18912 16488 18964
rect 16540 18952 16546 18964
rect 16758 18952 16764 18964
rect 16540 18924 16764 18952
rect 16540 18912 16546 18924
rect 16758 18912 16764 18924
rect 16816 18952 16822 18964
rect 17221 18955 17279 18961
rect 17221 18952 17233 18955
rect 16816 18924 17233 18952
rect 16816 18912 16822 18924
rect 17221 18921 17233 18924
rect 17267 18921 17279 18955
rect 17770 18952 17776 18964
rect 17221 18915 17279 18921
rect 17604 18924 17776 18952
rect 12526 18884 12532 18896
rect 10652 18856 10916 18884
rect 11992 18856 12532 18884
rect 10652 18844 10658 18856
rect 9309 18819 9367 18825
rect 9309 18785 9321 18819
rect 9355 18785 9367 18819
rect 9861 18819 9919 18825
rect 9861 18816 9873 18819
rect 9309 18779 9367 18785
rect 9416 18788 9873 18816
rect 6365 18751 6423 18757
rect 6365 18717 6377 18751
rect 6411 18717 6423 18751
rect 6365 18711 6423 18717
rect 6641 18751 6699 18757
rect 6641 18717 6653 18751
rect 6687 18717 6699 18751
rect 6641 18711 6699 18717
rect 1670 18689 1676 18692
rect 1664 18643 1676 18689
rect 1670 18640 1676 18643
rect 1728 18640 1734 18692
rect 5718 18680 5724 18692
rect 3344 18652 5724 18680
rect 3344 18624 3372 18652
rect 5718 18640 5724 18652
rect 5776 18640 5782 18692
rect 6656 18680 6684 18711
rect 7006 18708 7012 18760
rect 7064 18708 7070 18760
rect 7116 18720 7420 18748
rect 6730 18680 6736 18692
rect 6656 18652 6736 18680
rect 6730 18640 6736 18652
rect 6788 18640 6794 18692
rect 3145 18615 3203 18621
rect 3145 18581 3157 18615
rect 3191 18612 3203 18615
rect 3326 18612 3332 18624
rect 3191 18584 3332 18612
rect 3191 18581 3203 18584
rect 3145 18575 3203 18581
rect 3326 18572 3332 18584
rect 3384 18572 3390 18624
rect 3602 18572 3608 18624
rect 3660 18572 3666 18624
rect 3786 18572 3792 18624
rect 3844 18572 3850 18624
rect 5169 18615 5227 18621
rect 5169 18581 5181 18615
rect 5215 18612 5227 18615
rect 5350 18612 5356 18624
rect 5215 18584 5356 18612
rect 5215 18581 5227 18584
rect 5169 18575 5227 18581
rect 5350 18572 5356 18584
rect 5408 18572 5414 18624
rect 6549 18615 6607 18621
rect 6549 18581 6561 18615
rect 6595 18612 6607 18615
rect 7116 18612 7144 18720
rect 7193 18683 7251 18689
rect 7193 18649 7205 18683
rect 7239 18680 7251 18683
rect 7285 18683 7343 18689
rect 7285 18680 7297 18683
rect 7239 18652 7297 18680
rect 7239 18649 7251 18652
rect 7193 18643 7251 18649
rect 7285 18649 7297 18652
rect 7331 18649 7343 18683
rect 7392 18680 7420 18720
rect 7466 18708 7472 18760
rect 7524 18708 7530 18760
rect 7926 18708 7932 18760
rect 7984 18708 7990 18760
rect 8938 18708 8944 18760
rect 8996 18748 9002 18760
rect 9416 18748 9444 18788
rect 9861 18785 9873 18788
rect 9907 18785 9919 18819
rect 10888 18816 10916 18856
rect 12526 18844 12532 18856
rect 12584 18844 12590 18896
rect 16574 18884 16580 18896
rect 13924 18856 16580 18884
rect 11701 18819 11759 18825
rect 11701 18816 11713 18819
rect 9861 18779 9919 18785
rect 10060 18788 10824 18816
rect 10888 18788 11713 18816
rect 8996 18720 9444 18748
rect 8996 18708 9002 18720
rect 9490 18708 9496 18760
rect 9548 18708 9554 18760
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 10060 18757 10088 18788
rect 10045 18751 10103 18757
rect 10045 18748 10057 18751
rect 9732 18720 10057 18748
rect 9732 18708 9738 18720
rect 10045 18717 10057 18720
rect 10091 18717 10103 18751
rect 10045 18711 10103 18717
rect 10318 18708 10324 18760
rect 10376 18708 10382 18760
rect 10597 18751 10655 18757
rect 10597 18717 10609 18751
rect 10643 18717 10655 18751
rect 10597 18711 10655 18717
rect 8754 18680 8760 18692
rect 7392 18652 8760 18680
rect 7285 18643 7343 18649
rect 6595 18584 7144 18612
rect 7208 18612 7236 18643
rect 8754 18640 8760 18652
rect 8812 18640 8818 18692
rect 9214 18640 9220 18692
rect 9272 18640 9278 18692
rect 9769 18683 9827 18689
rect 9769 18649 9781 18683
rect 9815 18680 9827 18683
rect 9950 18680 9956 18692
rect 9815 18652 9956 18680
rect 9815 18649 9827 18652
rect 9769 18643 9827 18649
rect 9950 18640 9956 18652
rect 10008 18640 10014 18692
rect 7466 18612 7472 18624
rect 7208 18584 7472 18612
rect 6595 18581 6607 18584
rect 6549 18575 6607 18581
rect 7466 18572 7472 18584
rect 7524 18572 7530 18624
rect 7650 18572 7656 18624
rect 7708 18572 7714 18624
rect 7742 18572 7748 18624
rect 7800 18612 7806 18624
rect 10612 18612 10640 18711
rect 10796 18621 10824 18788
rect 11701 18785 11713 18788
rect 11747 18785 11759 18819
rect 11701 18779 11759 18785
rect 12066 18776 12072 18828
rect 12124 18816 12130 18828
rect 13262 18816 13268 18828
rect 12124 18788 13268 18816
rect 12124 18776 12130 18788
rect 13262 18776 13268 18788
rect 13320 18776 13326 18828
rect 11238 18708 11244 18760
rect 11296 18748 11302 18760
rect 11333 18751 11391 18757
rect 11333 18748 11345 18751
rect 11296 18720 11345 18748
rect 11296 18708 11302 18720
rect 11333 18717 11345 18720
rect 11379 18717 11391 18751
rect 11333 18711 11391 18717
rect 11517 18751 11575 18757
rect 11517 18717 11529 18751
rect 11563 18748 11575 18751
rect 11925 18751 11983 18757
rect 11563 18720 11836 18748
rect 11563 18717 11575 18720
rect 11517 18711 11575 18717
rect 11054 18640 11060 18692
rect 11112 18680 11118 18692
rect 11598 18683 11656 18689
rect 11598 18680 11610 18683
rect 11112 18652 11610 18680
rect 11112 18640 11118 18652
rect 11598 18649 11610 18652
rect 11644 18649 11656 18683
rect 11808 18680 11836 18720
rect 11925 18717 11937 18751
rect 11971 18748 11983 18751
rect 12250 18748 12256 18760
rect 11971 18720 12256 18748
rect 11971 18717 11983 18720
rect 11925 18711 11983 18717
rect 12250 18708 12256 18720
rect 12308 18708 12314 18760
rect 12345 18751 12403 18757
rect 12345 18717 12357 18751
rect 12391 18748 12403 18751
rect 12618 18748 12624 18760
rect 12391 18720 12624 18748
rect 12391 18717 12403 18720
rect 12345 18711 12403 18717
rect 12618 18708 12624 18720
rect 12676 18708 12682 18760
rect 12802 18708 12808 18760
rect 12860 18708 12866 18760
rect 13924 18748 13952 18856
rect 16574 18844 16580 18856
rect 16632 18844 16638 18896
rect 17494 18884 17500 18896
rect 16960 18856 17500 18884
rect 14274 18776 14280 18828
rect 14332 18816 14338 18828
rect 16298 18816 16304 18828
rect 14332 18788 16304 18816
rect 14332 18776 14338 18788
rect 16298 18776 16304 18788
rect 16356 18776 16362 18828
rect 13556 18720 13952 18748
rect 12529 18683 12587 18689
rect 12529 18680 12541 18683
rect 11808 18652 12541 18680
rect 11598 18643 11656 18649
rect 12529 18649 12541 18652
rect 12575 18680 12587 18683
rect 13556 18680 13584 18720
rect 14182 18708 14188 18760
rect 14240 18708 14246 18760
rect 16960 18757 16988 18856
rect 17494 18844 17500 18856
rect 17552 18844 17558 18896
rect 17129 18819 17187 18825
rect 17129 18785 17141 18819
rect 17175 18816 17187 18819
rect 17313 18819 17371 18825
rect 17313 18816 17325 18819
rect 17175 18788 17325 18816
rect 17175 18785 17187 18788
rect 17129 18779 17187 18785
rect 17313 18785 17325 18788
rect 17359 18816 17371 18819
rect 17604 18816 17632 18924
rect 17770 18912 17776 18924
rect 17828 18912 17834 18964
rect 18690 18912 18696 18964
rect 18748 18952 18754 18964
rect 19245 18955 19303 18961
rect 19245 18952 19257 18955
rect 18748 18924 19257 18952
rect 18748 18912 18754 18924
rect 19245 18921 19257 18924
rect 19291 18921 19303 18955
rect 19245 18915 19303 18921
rect 21266 18912 21272 18964
rect 21324 18912 21330 18964
rect 21453 18955 21511 18961
rect 21453 18921 21465 18955
rect 21499 18952 21511 18955
rect 21821 18955 21879 18961
rect 21821 18952 21833 18955
rect 21499 18924 21833 18952
rect 21499 18921 21511 18924
rect 21453 18915 21511 18921
rect 21821 18921 21833 18924
rect 21867 18952 21879 18955
rect 21910 18952 21916 18964
rect 21867 18924 21916 18952
rect 21867 18921 21879 18924
rect 21821 18915 21879 18921
rect 21910 18912 21916 18924
rect 21968 18912 21974 18964
rect 22097 18955 22155 18961
rect 22097 18921 22109 18955
rect 22143 18921 22155 18955
rect 22097 18915 22155 18921
rect 17681 18887 17739 18893
rect 17681 18853 17693 18887
rect 17727 18884 17739 18887
rect 19705 18887 19763 18893
rect 17727 18856 19656 18884
rect 17727 18853 17739 18856
rect 17681 18847 17739 18853
rect 19337 18819 19395 18825
rect 19337 18816 19349 18819
rect 17359 18788 17448 18816
rect 17604 18788 19349 18816
rect 17359 18785 17371 18788
rect 17313 18779 17371 18785
rect 16945 18751 17003 18757
rect 16945 18717 16957 18751
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 14369 18683 14427 18689
rect 14369 18680 14381 18683
rect 12575 18652 13584 18680
rect 13648 18652 14381 18680
rect 12575 18649 12587 18652
rect 12529 18643 12587 18649
rect 7800 18584 10640 18612
rect 10781 18615 10839 18621
rect 7800 18572 7806 18584
rect 10781 18581 10793 18615
rect 10827 18581 10839 18615
rect 10781 18575 10839 18581
rect 11882 18572 11888 18624
rect 11940 18612 11946 18624
rect 12161 18615 12219 18621
rect 12161 18612 12173 18615
rect 11940 18584 12173 18612
rect 11940 18572 11946 18584
rect 12161 18581 12173 18584
rect 12207 18581 12219 18615
rect 12161 18575 12219 18581
rect 12618 18572 12624 18624
rect 12676 18612 12682 18624
rect 13648 18612 13676 18652
rect 14369 18649 14381 18652
rect 14415 18680 14427 18683
rect 14642 18680 14648 18692
rect 14415 18652 14648 18680
rect 14415 18649 14427 18652
rect 14369 18643 14427 18649
rect 14642 18640 14648 18652
rect 14700 18640 14706 18692
rect 17221 18683 17279 18689
rect 17221 18680 17233 18683
rect 14752 18652 17233 18680
rect 12676 18584 13676 18612
rect 12676 18572 12682 18584
rect 13722 18572 13728 18624
rect 13780 18612 13786 18624
rect 14752 18612 14780 18652
rect 17221 18649 17233 18652
rect 17267 18649 17279 18683
rect 17420 18680 17448 18788
rect 19337 18785 19349 18788
rect 19383 18785 19395 18819
rect 19628 18816 19656 18856
rect 19705 18853 19717 18887
rect 19751 18884 19763 18887
rect 22112 18884 22140 18915
rect 22462 18912 22468 18964
rect 22520 18912 22526 18964
rect 22646 18912 22652 18964
rect 22704 18952 22710 18964
rect 22922 18952 22928 18964
rect 22704 18924 22928 18952
rect 22704 18912 22710 18924
rect 22922 18912 22928 18924
rect 22980 18912 22986 18964
rect 23017 18955 23075 18961
rect 23017 18921 23029 18955
rect 23063 18952 23075 18955
rect 23382 18952 23388 18964
rect 23063 18924 23388 18952
rect 23063 18921 23075 18924
rect 23017 18915 23075 18921
rect 23382 18912 23388 18924
rect 23440 18912 23446 18964
rect 23753 18955 23811 18961
rect 23753 18921 23765 18955
rect 23799 18921 23811 18955
rect 23753 18915 23811 18921
rect 19751 18856 22140 18884
rect 19751 18853 19763 18856
rect 19705 18847 19763 18853
rect 22738 18844 22744 18896
rect 22796 18884 22802 18896
rect 23768 18884 23796 18915
rect 24118 18912 24124 18964
rect 24176 18912 24182 18964
rect 24302 18912 24308 18964
rect 24360 18952 24366 18964
rect 24949 18955 25007 18961
rect 24949 18952 24961 18955
rect 24360 18924 24961 18952
rect 24360 18912 24366 18924
rect 24949 18921 24961 18924
rect 24995 18921 25007 18955
rect 24949 18915 25007 18921
rect 25866 18912 25872 18964
rect 25924 18952 25930 18964
rect 26142 18952 26148 18964
rect 25924 18924 26148 18952
rect 25924 18912 25930 18924
rect 26142 18912 26148 18924
rect 26200 18912 26206 18964
rect 29822 18912 29828 18964
rect 29880 18952 29886 18964
rect 30190 18952 30196 18964
rect 29880 18924 30196 18952
rect 29880 18912 29886 18924
rect 30190 18912 30196 18924
rect 30248 18912 30254 18964
rect 30282 18912 30288 18964
rect 30340 18952 30346 18964
rect 30745 18955 30803 18961
rect 30745 18952 30757 18955
rect 30340 18924 30757 18952
rect 30340 18912 30346 18924
rect 30745 18921 30757 18924
rect 30791 18952 30803 18955
rect 31846 18952 31852 18964
rect 30791 18924 31852 18952
rect 30791 18921 30803 18924
rect 30745 18915 30803 18921
rect 31846 18912 31852 18924
rect 31904 18912 31910 18964
rect 32493 18955 32551 18961
rect 32493 18921 32505 18955
rect 32539 18952 32551 18955
rect 32876 18952 32904 19264
rect 32539 18924 32904 18952
rect 32539 18921 32551 18924
rect 32493 18915 32551 18921
rect 22796 18856 23796 18884
rect 22796 18844 22802 18856
rect 19628 18788 21680 18816
rect 19337 18779 19395 18785
rect 17494 18708 17500 18760
rect 17552 18708 17558 18760
rect 17770 18708 17776 18760
rect 17828 18708 17834 18760
rect 19521 18751 19579 18757
rect 19521 18717 19533 18751
rect 19567 18717 19579 18751
rect 19521 18711 19579 18717
rect 17420 18652 18184 18680
rect 17221 18643 17279 18649
rect 13780 18584 14780 18612
rect 13780 18572 13786 18584
rect 16758 18572 16764 18624
rect 16816 18572 16822 18624
rect 17126 18572 17132 18624
rect 17184 18612 17190 18624
rect 17494 18612 17500 18624
rect 17184 18584 17500 18612
rect 17184 18572 17190 18584
rect 17494 18572 17500 18584
rect 17552 18572 17558 18624
rect 17957 18615 18015 18621
rect 17957 18581 17969 18615
rect 18003 18612 18015 18615
rect 18046 18612 18052 18624
rect 18003 18584 18052 18612
rect 18003 18581 18015 18584
rect 17957 18575 18015 18581
rect 18046 18572 18052 18584
rect 18104 18572 18110 18624
rect 18156 18612 18184 18652
rect 19242 18640 19248 18692
rect 19300 18640 19306 18692
rect 19334 18640 19340 18692
rect 19392 18680 19398 18692
rect 19536 18680 19564 18711
rect 19886 18708 19892 18760
rect 19944 18748 19950 18760
rect 20990 18748 20996 18760
rect 19944 18720 20996 18748
rect 19944 18708 19950 18720
rect 20990 18708 20996 18720
rect 21048 18748 21054 18760
rect 21085 18751 21143 18757
rect 21085 18748 21097 18751
rect 21048 18720 21097 18748
rect 21048 18708 21054 18720
rect 21085 18717 21097 18720
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 21269 18751 21327 18757
rect 21269 18717 21281 18751
rect 21315 18748 21327 18751
rect 21450 18748 21456 18760
rect 21315 18720 21456 18748
rect 21315 18717 21327 18720
rect 21269 18711 21327 18717
rect 21450 18708 21456 18720
rect 21508 18708 21514 18760
rect 20346 18680 20352 18692
rect 19392 18652 20352 18680
rect 19392 18640 19398 18652
rect 20346 18640 20352 18652
rect 20404 18640 20410 18692
rect 20530 18640 20536 18692
rect 20588 18680 20594 18692
rect 21545 18683 21603 18689
rect 21545 18680 21557 18683
rect 20588 18652 21557 18680
rect 20588 18640 20594 18652
rect 21545 18649 21557 18652
rect 21591 18649 21603 18683
rect 21652 18680 21680 18788
rect 21726 18776 21732 18828
rect 21784 18776 21790 18828
rect 22189 18819 22247 18825
rect 22189 18816 22201 18819
rect 21928 18788 22201 18816
rect 21818 18708 21824 18760
rect 21876 18708 21882 18760
rect 21928 18680 21956 18788
rect 22189 18785 22201 18788
rect 22235 18785 22247 18819
rect 22189 18779 22247 18785
rect 22833 18819 22891 18825
rect 22833 18785 22845 18819
rect 22879 18785 22891 18819
rect 23293 18819 23351 18825
rect 23293 18816 23305 18819
rect 22833 18779 22891 18785
rect 22940 18788 23305 18816
rect 22097 18751 22155 18757
rect 22097 18748 22109 18751
rect 21652 18652 21956 18680
rect 22020 18720 22109 18748
rect 21545 18643 21603 18649
rect 20714 18612 20720 18624
rect 18156 18584 20720 18612
rect 20714 18572 20720 18584
rect 20772 18572 20778 18624
rect 22020 18621 22048 18720
rect 22097 18717 22109 18720
rect 22143 18717 22155 18751
rect 22097 18711 22155 18717
rect 22462 18708 22468 18760
rect 22520 18748 22526 18760
rect 22649 18751 22707 18757
rect 22649 18748 22661 18751
rect 22520 18720 22661 18748
rect 22520 18708 22526 18720
rect 22649 18717 22661 18720
rect 22695 18748 22707 18751
rect 22848 18748 22876 18779
rect 22695 18720 22876 18748
rect 22695 18717 22707 18720
rect 22649 18711 22707 18717
rect 22940 18692 22968 18788
rect 23293 18785 23305 18788
rect 23339 18785 23351 18819
rect 23293 18779 23351 18785
rect 23474 18776 23480 18828
rect 23532 18816 23538 18828
rect 27522 18816 27528 18828
rect 23532 18788 27528 18816
rect 23532 18776 23538 18788
rect 27522 18776 27528 18788
rect 27580 18776 27586 18828
rect 30650 18776 30656 18828
rect 30708 18816 30714 18828
rect 31113 18819 31171 18825
rect 31113 18816 31125 18819
rect 30708 18788 31125 18816
rect 30708 18776 30714 18788
rect 31113 18785 31125 18788
rect 31159 18785 31171 18819
rect 31113 18779 31171 18785
rect 23017 18751 23075 18757
rect 23017 18717 23029 18751
rect 23063 18748 23075 18751
rect 23106 18748 23112 18760
rect 23063 18720 23112 18748
rect 23063 18717 23075 18720
rect 23017 18711 23075 18717
rect 23106 18708 23112 18720
rect 23164 18708 23170 18760
rect 23753 18751 23811 18757
rect 23753 18748 23765 18751
rect 23216 18720 23765 18748
rect 22741 18683 22799 18689
rect 22741 18649 22753 18683
rect 22787 18680 22799 18683
rect 22922 18680 22928 18692
rect 22787 18652 22928 18680
rect 22787 18649 22799 18652
rect 22741 18643 22799 18649
rect 22922 18640 22928 18652
rect 22980 18640 22986 18692
rect 23216 18621 23244 18720
rect 23753 18717 23765 18720
rect 23799 18717 23811 18751
rect 23753 18711 23811 18717
rect 23842 18708 23848 18760
rect 23900 18708 23906 18760
rect 24949 18751 25007 18757
rect 24949 18717 24961 18751
rect 24995 18748 25007 18751
rect 24995 18720 25029 18748
rect 24995 18717 25007 18720
rect 24949 18711 25007 18717
rect 23474 18640 23480 18692
rect 23532 18640 23538 18692
rect 23566 18640 23572 18692
rect 23624 18680 23630 18692
rect 23661 18683 23719 18689
rect 23661 18680 23673 18683
rect 23624 18652 23673 18680
rect 23624 18640 23630 18652
rect 23661 18649 23673 18652
rect 23707 18649 23719 18683
rect 23661 18643 23719 18649
rect 24857 18683 24915 18689
rect 24857 18649 24869 18683
rect 24903 18680 24915 18683
rect 24964 18680 24992 18711
rect 25130 18708 25136 18760
rect 25188 18708 25194 18760
rect 28994 18708 29000 18760
rect 29052 18748 29058 18760
rect 29089 18751 29147 18757
rect 29089 18748 29101 18751
rect 29052 18720 29101 18748
rect 29052 18708 29058 18720
rect 29089 18717 29101 18720
rect 29135 18717 29147 18751
rect 29089 18711 29147 18717
rect 29178 18708 29184 18760
rect 29236 18748 29242 18760
rect 29273 18751 29331 18757
rect 29273 18748 29285 18751
rect 29236 18720 29285 18748
rect 29236 18708 29242 18720
rect 29273 18717 29285 18720
rect 29319 18717 29331 18751
rect 29273 18711 29331 18717
rect 30561 18751 30619 18757
rect 30561 18717 30573 18751
rect 30607 18748 30619 18751
rect 30607 18720 30880 18748
rect 30607 18717 30619 18720
rect 30561 18711 30619 18717
rect 30098 18680 30104 18692
rect 24903 18652 30104 18680
rect 24903 18649 24915 18652
rect 24857 18643 24915 18649
rect 30098 18640 30104 18652
rect 30156 18640 30162 18692
rect 22005 18615 22063 18621
rect 22005 18581 22017 18615
rect 22051 18581 22063 18615
rect 22005 18575 22063 18581
rect 23201 18615 23259 18621
rect 23201 18581 23213 18615
rect 23247 18581 23259 18615
rect 23201 18575 23259 18581
rect 25317 18615 25375 18621
rect 25317 18581 25329 18615
rect 25363 18612 25375 18615
rect 28166 18612 28172 18624
rect 25363 18584 28172 18612
rect 25363 18581 25375 18584
rect 25317 18575 25375 18581
rect 28166 18572 28172 18584
rect 28224 18572 28230 18624
rect 29178 18572 29184 18624
rect 29236 18572 29242 18624
rect 30852 18621 30880 18720
rect 30926 18708 30932 18760
rect 30984 18748 30990 18760
rect 31021 18751 31079 18757
rect 31021 18748 31033 18751
rect 30984 18720 31033 18748
rect 30984 18708 30990 18720
rect 31021 18717 31033 18720
rect 31067 18717 31079 18751
rect 31021 18711 31079 18717
rect 31202 18708 31208 18760
rect 31260 18748 31266 18760
rect 31369 18751 31427 18757
rect 31369 18748 31381 18751
rect 31260 18720 31381 18748
rect 31260 18708 31266 18720
rect 31369 18717 31381 18720
rect 31415 18717 31427 18751
rect 31369 18711 31427 18717
rect 30837 18615 30895 18621
rect 30837 18581 30849 18615
rect 30883 18612 30895 18615
rect 31386 18612 31392 18624
rect 30883 18584 31392 18612
rect 30883 18581 30895 18584
rect 30837 18575 30895 18581
rect 31386 18572 31392 18584
rect 31444 18572 31450 18624
rect 1104 18522 32844 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 32844 18522
rect 1104 18448 32844 18470
rect 2409 18411 2467 18417
rect 2409 18377 2421 18411
rect 2455 18408 2467 18411
rect 2590 18408 2596 18420
rect 2455 18380 2596 18408
rect 2455 18377 2467 18380
rect 2409 18371 2467 18377
rect 2424 18340 2452 18371
rect 2590 18368 2596 18380
rect 2648 18368 2654 18420
rect 3510 18368 3516 18420
rect 3568 18368 3574 18420
rect 3605 18411 3663 18417
rect 3605 18377 3617 18411
rect 3651 18377 3663 18411
rect 3605 18371 3663 18377
rect 2866 18340 2872 18352
rect 2424 18312 2872 18340
rect 2866 18300 2872 18312
rect 2924 18300 2930 18352
rect 2961 18343 3019 18349
rect 2961 18309 2973 18343
rect 3007 18340 3019 18343
rect 3620 18340 3648 18371
rect 4614 18368 4620 18420
rect 4672 18368 4678 18420
rect 7285 18411 7343 18417
rect 7285 18377 7297 18411
rect 7331 18408 7343 18411
rect 7926 18408 7932 18420
rect 7331 18380 7932 18408
rect 7331 18377 7343 18380
rect 7285 18371 7343 18377
rect 7926 18368 7932 18380
rect 7984 18368 7990 18420
rect 8110 18368 8116 18420
rect 8168 18408 8174 18420
rect 8168 18380 8892 18408
rect 8168 18368 8174 18380
rect 4632 18340 4660 18368
rect 5077 18343 5135 18349
rect 3007 18312 4476 18340
rect 4632 18312 5028 18340
rect 3007 18309 3019 18312
rect 2961 18303 3019 18309
rect 2593 18275 2651 18281
rect 2593 18241 2605 18275
rect 2639 18241 2651 18275
rect 2593 18235 2651 18241
rect 2608 18204 2636 18235
rect 2682 18232 2688 18284
rect 2740 18232 2746 18284
rect 3050 18232 3056 18284
rect 3108 18281 3114 18284
rect 3108 18275 3157 18281
rect 3108 18241 3111 18275
rect 3145 18272 3157 18275
rect 3145 18244 3280 18272
rect 3145 18241 3157 18244
rect 3108 18235 3157 18241
rect 3108 18232 3114 18235
rect 3252 18204 3280 18244
rect 3326 18232 3332 18284
rect 3384 18232 3390 18284
rect 3694 18232 3700 18284
rect 3752 18272 3758 18284
rect 3789 18275 3847 18281
rect 3789 18272 3801 18275
rect 3752 18244 3801 18272
rect 3752 18232 3758 18244
rect 3789 18241 3801 18244
rect 3835 18241 3847 18275
rect 3789 18235 3847 18241
rect 4338 18232 4344 18284
rect 4396 18232 4402 18284
rect 4448 18272 4476 18312
rect 4614 18272 4620 18284
rect 4448 18244 4620 18272
rect 4614 18232 4620 18244
rect 4672 18272 4678 18284
rect 4801 18275 4859 18281
rect 4801 18272 4813 18275
rect 4672 18244 4813 18272
rect 4672 18232 4678 18244
rect 4801 18241 4813 18244
rect 4847 18272 4859 18275
rect 4890 18272 4896 18284
rect 4847 18244 4896 18272
rect 4847 18241 4859 18244
rect 4801 18235 4859 18241
rect 4890 18232 4896 18244
rect 4948 18232 4954 18284
rect 5000 18281 5028 18312
rect 5077 18309 5089 18343
rect 5123 18340 5135 18343
rect 5350 18340 5356 18352
rect 5123 18312 5356 18340
rect 5123 18309 5135 18312
rect 5077 18303 5135 18309
rect 4985 18275 5043 18281
rect 4985 18241 4997 18275
rect 5031 18241 5043 18275
rect 4985 18235 5043 18241
rect 3510 18204 3516 18216
rect 2608 18176 2774 18204
rect 3252 18176 3516 18204
rect 2746 18068 2774 18176
rect 3510 18164 3516 18176
rect 3568 18164 3574 18216
rect 4706 18164 4712 18216
rect 4764 18204 4770 18216
rect 5092 18204 5120 18303
rect 5350 18300 5356 18312
rect 5408 18300 5414 18352
rect 6454 18300 6460 18352
rect 6512 18340 6518 18352
rect 8864 18340 8892 18380
rect 8938 18368 8944 18420
rect 8996 18408 9002 18420
rect 9401 18411 9459 18417
rect 9401 18408 9413 18411
rect 8996 18380 9413 18408
rect 8996 18368 9002 18380
rect 9401 18377 9413 18380
rect 9447 18408 9459 18411
rect 9858 18408 9864 18420
rect 9447 18380 9864 18408
rect 9447 18377 9459 18380
rect 9401 18371 9459 18377
rect 9858 18368 9864 18380
rect 9916 18368 9922 18420
rect 11698 18368 11704 18420
rect 11756 18408 11762 18420
rect 11882 18408 11888 18420
rect 11756 18380 11888 18408
rect 11756 18368 11762 18380
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 12158 18368 12164 18420
rect 12216 18368 12222 18420
rect 12434 18368 12440 18420
rect 12492 18408 12498 18420
rect 12529 18411 12587 18417
rect 12529 18408 12541 18411
rect 12492 18380 12541 18408
rect 12492 18368 12498 18380
rect 12529 18377 12541 18380
rect 12575 18408 12587 18411
rect 12710 18408 12716 18420
rect 12575 18380 12716 18408
rect 12575 18377 12587 18380
rect 12529 18371 12587 18377
rect 12710 18368 12716 18380
rect 12768 18368 12774 18420
rect 12894 18368 12900 18420
rect 12952 18408 12958 18420
rect 14274 18408 14280 18420
rect 12952 18380 14280 18408
rect 12952 18368 12958 18380
rect 14274 18368 14280 18380
rect 14332 18368 14338 18420
rect 15286 18368 15292 18420
rect 15344 18408 15350 18420
rect 17218 18408 17224 18420
rect 15344 18380 17224 18408
rect 15344 18368 15350 18380
rect 17218 18368 17224 18380
rect 17276 18368 17282 18420
rect 17310 18368 17316 18420
rect 17368 18408 17374 18420
rect 20254 18408 20260 18420
rect 17368 18380 20260 18408
rect 17368 18368 17374 18380
rect 20254 18368 20260 18380
rect 20312 18368 20318 18420
rect 21450 18408 21456 18420
rect 21100 18380 21456 18408
rect 9769 18343 9827 18349
rect 6512 18312 8248 18340
rect 8864 18312 9720 18340
rect 6512 18300 6518 18312
rect 5169 18275 5227 18281
rect 5169 18241 5181 18275
rect 5215 18272 5227 18275
rect 5626 18272 5632 18284
rect 5215 18244 5632 18272
rect 5215 18241 5227 18244
rect 5169 18235 5227 18241
rect 5626 18232 5632 18244
rect 5684 18232 5690 18284
rect 7469 18275 7527 18281
rect 7469 18241 7481 18275
rect 7515 18272 7527 18275
rect 7515 18244 7696 18272
rect 7515 18241 7527 18244
rect 7469 18235 7527 18241
rect 4764 18176 5120 18204
rect 4764 18164 4770 18176
rect 6270 18164 6276 18216
rect 6328 18204 6334 18216
rect 6546 18204 6552 18216
rect 6328 18176 6552 18204
rect 6328 18164 6334 18176
rect 6546 18164 6552 18176
rect 6604 18204 6610 18216
rect 7561 18207 7619 18213
rect 7561 18204 7573 18207
rect 6604 18176 7573 18204
rect 6604 18164 6610 18176
rect 7561 18173 7573 18176
rect 7607 18173 7619 18207
rect 7668 18204 7696 18244
rect 7742 18232 7748 18284
rect 7800 18232 7806 18284
rect 7834 18232 7840 18284
rect 7892 18232 7898 18284
rect 7926 18204 7932 18216
rect 7668 18176 7932 18204
rect 7561 18167 7619 18173
rect 7926 18164 7932 18176
rect 7984 18204 7990 18216
rect 8110 18204 8116 18216
rect 7984 18176 8116 18204
rect 7984 18164 7990 18176
rect 8110 18164 8116 18176
rect 8168 18164 8174 18216
rect 3237 18139 3295 18145
rect 3237 18105 3249 18139
rect 3283 18136 3295 18139
rect 7006 18136 7012 18148
rect 3283 18108 7012 18136
rect 3283 18105 3295 18108
rect 3237 18099 3295 18105
rect 7006 18096 7012 18108
rect 7064 18096 7070 18148
rect 7466 18096 7472 18148
rect 7524 18136 7530 18148
rect 7524 18108 7696 18136
rect 7524 18096 7530 18108
rect 3602 18068 3608 18080
rect 2746 18040 3608 18068
rect 3602 18028 3608 18040
rect 3660 18028 3666 18080
rect 3694 18028 3700 18080
rect 3752 18068 3758 18080
rect 4157 18071 4215 18077
rect 4157 18068 4169 18071
rect 3752 18040 4169 18068
rect 3752 18028 3758 18040
rect 4157 18037 4169 18040
rect 4203 18037 4215 18071
rect 4157 18031 4215 18037
rect 5353 18071 5411 18077
rect 5353 18037 5365 18071
rect 5399 18068 5411 18071
rect 6086 18068 6092 18080
rect 5399 18040 6092 18068
rect 5399 18037 5411 18040
rect 5353 18031 5411 18037
rect 6086 18028 6092 18040
rect 6144 18028 6150 18080
rect 7668 18077 7696 18108
rect 7834 18096 7840 18148
rect 7892 18136 7898 18148
rect 8021 18139 8079 18145
rect 8021 18136 8033 18139
rect 7892 18108 8033 18136
rect 7892 18096 7898 18108
rect 8021 18105 8033 18108
rect 8067 18105 8079 18139
rect 8220 18136 8248 18312
rect 9398 18232 9404 18284
rect 9456 18272 9462 18284
rect 9585 18275 9643 18281
rect 9585 18272 9597 18275
rect 9456 18244 9597 18272
rect 9456 18232 9462 18244
rect 9585 18241 9597 18244
rect 9631 18241 9643 18275
rect 9692 18272 9720 18312
rect 9769 18309 9781 18343
rect 9815 18340 9827 18343
rect 10870 18340 10876 18352
rect 9815 18312 10876 18340
rect 9815 18309 9827 18312
rect 9769 18303 9827 18309
rect 10870 18300 10876 18312
rect 10928 18300 10934 18352
rect 16114 18340 16120 18352
rect 10980 18312 13400 18340
rect 10980 18272 11008 18312
rect 13372 18296 13400 18312
rect 13556 18312 16120 18340
rect 13449 18299 13507 18305
rect 13449 18296 13461 18299
rect 9692 18244 11008 18272
rect 9585 18235 9643 18241
rect 11514 18232 11520 18284
rect 11572 18272 11578 18284
rect 11790 18272 11796 18284
rect 11572 18244 11796 18272
rect 11572 18232 11578 18244
rect 11790 18232 11796 18244
rect 11848 18232 11854 18284
rect 11882 18232 11888 18284
rect 11940 18272 11946 18284
rect 12158 18272 12164 18284
rect 11940 18244 12164 18272
rect 11940 18232 11946 18244
rect 12158 18232 12164 18244
rect 12216 18272 12222 18284
rect 12345 18275 12403 18281
rect 12345 18272 12357 18275
rect 12216 18244 12357 18272
rect 12216 18232 12222 18244
rect 12345 18241 12357 18244
rect 12391 18241 12403 18275
rect 13372 18268 13461 18296
rect 13449 18265 13461 18268
rect 13495 18265 13507 18299
rect 13449 18259 13507 18265
rect 12345 18235 12403 18241
rect 8662 18164 8668 18216
rect 8720 18204 8726 18216
rect 11238 18204 11244 18216
rect 8720 18176 11244 18204
rect 8720 18164 8726 18176
rect 11238 18164 11244 18176
rect 11296 18204 11302 18216
rect 12250 18204 12256 18216
rect 11296 18176 12256 18204
rect 11296 18164 11302 18176
rect 12250 18164 12256 18176
rect 12308 18164 12314 18216
rect 12526 18164 12532 18216
rect 12584 18204 12590 18216
rect 13556 18204 13584 18312
rect 16114 18300 16120 18312
rect 16172 18300 16178 18352
rect 16850 18300 16856 18352
rect 16908 18340 16914 18352
rect 16945 18343 17003 18349
rect 16945 18340 16957 18343
rect 16908 18312 16957 18340
rect 16908 18300 16914 18312
rect 16945 18309 16957 18312
rect 16991 18309 17003 18343
rect 16945 18303 17003 18309
rect 17052 18312 17356 18340
rect 14553 18275 14611 18281
rect 14553 18241 14565 18275
rect 14599 18272 14611 18275
rect 14734 18272 14740 18284
rect 14599 18244 14740 18272
rect 14599 18241 14611 18244
rect 14553 18235 14611 18241
rect 14734 18232 14740 18244
rect 14792 18232 14798 18284
rect 14826 18232 14832 18284
rect 14884 18232 14890 18284
rect 15381 18275 15439 18281
rect 15381 18241 15393 18275
rect 15427 18272 15439 18275
rect 15470 18272 15476 18284
rect 15427 18244 15476 18272
rect 15427 18241 15439 18244
rect 15381 18235 15439 18241
rect 15470 18232 15476 18244
rect 15528 18232 15534 18284
rect 15654 18232 15660 18284
rect 15712 18272 15718 18284
rect 17052 18272 17080 18312
rect 15712 18244 17080 18272
rect 15712 18232 15718 18244
rect 17218 18232 17224 18284
rect 17276 18232 17282 18284
rect 17328 18272 17356 18312
rect 18598 18300 18604 18352
rect 18656 18340 18662 18352
rect 19153 18343 19211 18349
rect 19153 18340 19165 18343
rect 18656 18312 19165 18340
rect 18656 18300 18662 18312
rect 19153 18309 19165 18312
rect 19199 18309 19211 18343
rect 19153 18303 19211 18309
rect 18782 18272 18788 18284
rect 17328 18244 18788 18272
rect 18782 18232 18788 18244
rect 18840 18232 18846 18284
rect 18877 18275 18935 18281
rect 18877 18241 18889 18275
rect 18923 18241 18935 18275
rect 18877 18235 18935 18241
rect 12584 18176 13584 18204
rect 14277 18207 14335 18213
rect 12584 18164 12590 18176
rect 14277 18173 14289 18207
rect 14323 18204 14335 18207
rect 14642 18204 14648 18216
rect 14323 18176 14648 18204
rect 14323 18173 14335 18176
rect 14277 18167 14335 18173
rect 14642 18164 14648 18176
rect 14700 18164 14706 18216
rect 16758 18164 16764 18216
rect 16816 18204 16822 18216
rect 17037 18207 17095 18213
rect 17037 18204 17049 18207
rect 16816 18176 17049 18204
rect 16816 18164 16822 18176
rect 17037 18173 17049 18176
rect 17083 18173 17095 18207
rect 17770 18204 17776 18216
rect 17037 18167 17095 18173
rect 17144 18176 17776 18204
rect 10502 18136 10508 18148
rect 8220 18108 10508 18136
rect 8021 18099 8079 18105
rect 10502 18096 10508 18108
rect 10560 18096 10566 18148
rect 11514 18096 11520 18148
rect 11572 18136 11578 18148
rect 12342 18136 12348 18148
rect 11572 18108 12348 18136
rect 11572 18096 11578 18108
rect 12342 18096 12348 18108
rect 12400 18096 12406 18148
rect 17144 18136 17172 18176
rect 17770 18164 17776 18176
rect 17828 18164 17834 18216
rect 12544 18108 17172 18136
rect 17405 18139 17463 18145
rect 7653 18071 7711 18077
rect 7653 18037 7665 18071
rect 7699 18037 7711 18071
rect 7653 18031 7711 18037
rect 8754 18028 8760 18080
rect 8812 18068 8818 18080
rect 10594 18068 10600 18080
rect 8812 18040 10600 18068
rect 8812 18028 8818 18040
rect 10594 18028 10600 18040
rect 10652 18068 10658 18080
rect 12544 18068 12572 18108
rect 17405 18105 17417 18139
rect 17451 18136 17463 18139
rect 17494 18136 17500 18148
rect 17451 18108 17500 18136
rect 17451 18105 17463 18108
rect 17405 18099 17463 18105
rect 17494 18096 17500 18108
rect 17552 18136 17558 18148
rect 18892 18136 18920 18235
rect 18966 18232 18972 18284
rect 19024 18232 19030 18284
rect 19168 18204 19196 18303
rect 19886 18300 19892 18352
rect 19944 18340 19950 18352
rect 21100 18340 21128 18380
rect 21450 18368 21456 18380
rect 21508 18368 21514 18420
rect 21818 18368 21824 18420
rect 21876 18408 21882 18420
rect 23842 18408 23848 18420
rect 21876 18380 23848 18408
rect 21876 18368 21882 18380
rect 23842 18368 23848 18380
rect 23900 18368 23906 18420
rect 28353 18411 28411 18417
rect 28353 18377 28365 18411
rect 28399 18408 28411 18411
rect 28902 18408 28908 18420
rect 28399 18380 28908 18408
rect 28399 18377 28411 18380
rect 28353 18371 28411 18377
rect 28902 18368 28908 18380
rect 28960 18368 28966 18420
rect 30466 18368 30472 18420
rect 30524 18368 30530 18420
rect 31941 18411 31999 18417
rect 31941 18377 31953 18411
rect 31987 18408 31999 18411
rect 32214 18408 32220 18420
rect 31987 18380 32220 18408
rect 31987 18377 31999 18380
rect 31941 18371 31999 18377
rect 32214 18368 32220 18380
rect 32272 18368 32278 18420
rect 19944 18312 21128 18340
rect 19944 18300 19950 18312
rect 21174 18300 21180 18352
rect 21232 18340 21238 18352
rect 22738 18340 22744 18352
rect 21232 18312 22744 18340
rect 21232 18300 21238 18312
rect 22738 18300 22744 18312
rect 22796 18300 22802 18352
rect 23661 18343 23719 18349
rect 23661 18340 23673 18343
rect 22848 18312 23673 18340
rect 19518 18232 19524 18284
rect 19576 18272 19582 18284
rect 20070 18272 20076 18284
rect 19576 18244 20076 18272
rect 19576 18232 19582 18244
rect 20070 18232 20076 18244
rect 20128 18232 20134 18284
rect 20254 18232 20260 18284
rect 20312 18272 20318 18284
rect 22848 18272 22876 18312
rect 23661 18309 23673 18312
rect 23707 18309 23719 18343
rect 23661 18303 23719 18309
rect 26436 18312 30604 18340
rect 20312 18244 22876 18272
rect 20312 18232 20318 18244
rect 23474 18232 23480 18284
rect 23532 18232 23538 18284
rect 26142 18232 26148 18284
rect 26200 18272 26206 18284
rect 26436 18281 26464 18312
rect 26421 18275 26479 18281
rect 26421 18272 26433 18275
rect 26200 18244 26433 18272
rect 26200 18232 26206 18244
rect 26421 18241 26433 18244
rect 26467 18241 26479 18275
rect 26421 18235 26479 18241
rect 27522 18232 27528 18284
rect 27580 18272 27586 18284
rect 27706 18272 27712 18284
rect 27580 18244 27712 18272
rect 27580 18232 27586 18244
rect 27706 18232 27712 18244
rect 27764 18232 27770 18284
rect 27890 18232 27896 18284
rect 27948 18232 27954 18284
rect 28169 18275 28227 18281
rect 28169 18241 28181 18275
rect 28215 18241 28227 18275
rect 28169 18235 28227 18241
rect 27985 18207 28043 18213
rect 27985 18204 27997 18207
rect 19168 18176 27997 18204
rect 27985 18173 27997 18176
rect 28031 18173 28043 18207
rect 27985 18167 28043 18173
rect 17552 18108 18920 18136
rect 17552 18096 17558 18108
rect 21450 18096 21456 18148
rect 21508 18136 21514 18148
rect 22186 18136 22192 18148
rect 21508 18108 22192 18136
rect 21508 18096 21514 18108
rect 22186 18096 22192 18108
rect 22244 18096 22250 18148
rect 28184 18136 28212 18235
rect 28258 18232 28264 18284
rect 28316 18272 28322 18284
rect 29733 18275 29791 18281
rect 29733 18272 29745 18275
rect 28316 18244 29745 18272
rect 28316 18232 28322 18244
rect 29733 18241 29745 18244
rect 29779 18241 29791 18275
rect 29733 18235 29791 18241
rect 29917 18275 29975 18281
rect 29917 18241 29929 18275
rect 29963 18241 29975 18275
rect 29917 18235 29975 18241
rect 29270 18164 29276 18216
rect 29328 18204 29334 18216
rect 29932 18204 29960 18235
rect 30282 18232 30288 18284
rect 30340 18232 30346 18284
rect 30576 18281 30604 18312
rect 30561 18275 30619 18281
rect 30561 18241 30573 18275
rect 30607 18272 30619 18275
rect 30650 18272 30656 18284
rect 30607 18244 30656 18272
rect 30607 18241 30619 18244
rect 30561 18235 30619 18241
rect 30650 18232 30656 18244
rect 30708 18232 30714 18284
rect 30828 18275 30886 18281
rect 30828 18241 30840 18275
rect 30874 18272 30886 18275
rect 31386 18272 31392 18284
rect 30874 18244 31392 18272
rect 30874 18241 30886 18244
rect 30828 18235 30886 18241
rect 31386 18232 31392 18244
rect 31444 18232 31450 18284
rect 32217 18275 32275 18281
rect 32217 18241 32229 18275
rect 32263 18272 32275 18275
rect 32876 18272 32904 18924
rect 32263 18244 32904 18272
rect 32263 18241 32275 18244
rect 32217 18235 32275 18241
rect 29328 18176 29960 18204
rect 29328 18164 29334 18176
rect 22388 18108 28212 18136
rect 22388 18080 22416 18108
rect 10652 18040 12572 18068
rect 10652 18028 10658 18040
rect 13354 18028 13360 18080
rect 13412 18068 13418 18080
rect 13633 18071 13691 18077
rect 13633 18068 13645 18071
rect 13412 18040 13645 18068
rect 13412 18028 13418 18040
rect 13633 18037 13645 18040
rect 13679 18037 13691 18071
rect 13633 18031 13691 18037
rect 14369 18071 14427 18077
rect 14369 18037 14381 18071
rect 14415 18068 14427 18071
rect 14458 18068 14464 18080
rect 14415 18040 14464 18068
rect 14415 18037 14427 18040
rect 14369 18031 14427 18037
rect 14458 18028 14464 18040
rect 14516 18028 14522 18080
rect 14829 18071 14887 18077
rect 14829 18037 14841 18071
rect 14875 18068 14887 18071
rect 15010 18068 15016 18080
rect 14875 18040 15016 18068
rect 14875 18037 14887 18040
rect 14829 18031 14887 18037
rect 15010 18028 15016 18040
rect 15068 18028 15074 18080
rect 15194 18028 15200 18080
rect 15252 18028 15258 18080
rect 17221 18071 17279 18077
rect 17221 18037 17233 18071
rect 17267 18068 17279 18071
rect 18046 18068 18052 18080
rect 17267 18040 18052 18068
rect 17267 18037 17279 18040
rect 17221 18031 17279 18037
rect 18046 18028 18052 18040
rect 18104 18028 18110 18080
rect 18690 18028 18696 18080
rect 18748 18028 18754 18080
rect 19153 18071 19211 18077
rect 19153 18037 19165 18071
rect 19199 18068 19211 18071
rect 19518 18068 19524 18080
rect 19199 18040 19524 18068
rect 19199 18037 19211 18040
rect 19153 18031 19211 18037
rect 19518 18028 19524 18040
rect 19576 18028 19582 18080
rect 19978 18028 19984 18080
rect 20036 18068 20042 18080
rect 20622 18068 20628 18080
rect 20036 18040 20628 18068
rect 20036 18028 20042 18040
rect 20622 18028 20628 18040
rect 20680 18028 20686 18080
rect 20990 18028 20996 18080
rect 21048 18068 21054 18080
rect 22370 18068 22376 18080
rect 21048 18040 22376 18068
rect 21048 18028 21054 18040
rect 22370 18028 22376 18040
rect 22428 18028 22434 18080
rect 25406 18028 25412 18080
rect 25464 18068 25470 18080
rect 26694 18068 26700 18080
rect 25464 18040 26700 18068
rect 25464 18028 25470 18040
rect 26694 18028 26700 18040
rect 26752 18028 26758 18080
rect 27890 18028 27896 18080
rect 27948 18028 27954 18080
rect 29638 18028 29644 18080
rect 29696 18068 29702 18080
rect 30101 18071 30159 18077
rect 30101 18068 30113 18071
rect 29696 18040 30113 18068
rect 29696 18028 29702 18040
rect 30101 18037 30113 18040
rect 30147 18037 30159 18071
rect 30101 18031 30159 18037
rect 32398 18028 32404 18080
rect 32456 18028 32462 18080
rect 1104 17978 32844 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 32844 17978
rect 1104 17904 32844 17926
rect 2682 17824 2688 17876
rect 2740 17824 2746 17876
rect 5350 17864 5356 17876
rect 2884 17836 5356 17864
rect 2884 17669 2912 17836
rect 5350 17824 5356 17836
rect 5408 17824 5414 17876
rect 7834 17824 7840 17876
rect 7892 17864 7898 17876
rect 11146 17864 11152 17876
rect 7892 17836 11152 17864
rect 7892 17824 7898 17836
rect 11146 17824 11152 17836
rect 11204 17824 11210 17876
rect 11422 17824 11428 17876
rect 11480 17864 11486 17876
rect 11606 17864 11612 17876
rect 11480 17836 11612 17864
rect 11480 17824 11486 17836
rect 11606 17824 11612 17836
rect 11664 17824 11670 17876
rect 12066 17824 12072 17876
rect 12124 17864 12130 17876
rect 12434 17864 12440 17876
rect 12124 17836 12440 17864
rect 12124 17824 12130 17836
rect 12434 17824 12440 17836
rect 12492 17824 12498 17876
rect 12710 17824 12716 17876
rect 12768 17864 12774 17876
rect 13078 17864 13084 17876
rect 12768 17836 13084 17864
rect 12768 17824 12774 17836
rect 13078 17824 13084 17836
rect 13136 17824 13142 17876
rect 14093 17867 14151 17873
rect 14093 17864 14105 17867
rect 13372 17836 14105 17864
rect 4525 17799 4583 17805
rect 4525 17765 4537 17799
rect 4571 17796 4583 17799
rect 5442 17796 5448 17808
rect 4571 17768 5448 17796
rect 4571 17765 4583 17768
rect 4525 17759 4583 17765
rect 5442 17756 5448 17768
rect 5500 17756 5506 17808
rect 6362 17756 6368 17808
rect 6420 17796 6426 17808
rect 7561 17799 7619 17805
rect 6420 17768 7420 17796
rect 6420 17756 6426 17768
rect 3694 17688 3700 17740
rect 3752 17728 3758 17740
rect 4982 17728 4988 17740
rect 3752 17700 4200 17728
rect 3752 17688 3758 17700
rect 4172 17672 4200 17700
rect 4816 17700 4988 17728
rect 2869 17663 2927 17669
rect 2869 17629 2881 17663
rect 2915 17629 2927 17663
rect 2869 17623 2927 17629
rect 3142 17620 3148 17672
rect 3200 17620 3206 17672
rect 3418 17620 3424 17672
rect 3476 17620 3482 17672
rect 3973 17663 4031 17669
rect 3973 17629 3985 17663
rect 4019 17629 4031 17663
rect 3973 17623 4031 17629
rect 3694 17592 3700 17604
rect 2746 17564 3700 17592
rect 2746 17536 2774 17564
rect 3694 17552 3700 17564
rect 3752 17592 3758 17604
rect 3988 17592 4016 17623
rect 4154 17620 4160 17672
rect 4212 17620 4218 17672
rect 4341 17663 4399 17669
rect 4341 17629 4353 17663
rect 4387 17660 4399 17663
rect 4614 17660 4620 17672
rect 4387 17632 4620 17660
rect 4387 17629 4399 17632
rect 4341 17623 4399 17629
rect 4614 17620 4620 17632
rect 4672 17620 4678 17672
rect 4816 17669 4844 17700
rect 4982 17688 4988 17700
rect 5040 17728 5046 17740
rect 7282 17728 7288 17740
rect 5040 17700 7288 17728
rect 5040 17688 5046 17700
rect 7282 17688 7288 17700
rect 7340 17688 7346 17740
rect 7392 17728 7420 17768
rect 7561 17765 7573 17799
rect 7607 17796 7619 17799
rect 7650 17796 7656 17808
rect 7607 17768 7656 17796
rect 7607 17765 7619 17768
rect 7561 17759 7619 17765
rect 7650 17756 7656 17768
rect 7708 17756 7714 17808
rect 8018 17756 8024 17808
rect 8076 17796 8082 17808
rect 8754 17796 8760 17808
rect 8076 17768 8760 17796
rect 8076 17756 8082 17768
rect 8754 17756 8760 17768
rect 8812 17756 8818 17808
rect 9953 17799 10011 17805
rect 9953 17765 9965 17799
rect 9999 17796 10011 17799
rect 10502 17796 10508 17808
rect 9999 17768 10508 17796
rect 9999 17765 10011 17768
rect 9953 17759 10011 17765
rect 10502 17756 10508 17768
rect 10560 17756 10566 17808
rect 10870 17756 10876 17808
rect 10928 17796 10934 17808
rect 11974 17796 11980 17808
rect 10928 17768 11980 17796
rect 10928 17756 10934 17768
rect 11974 17756 11980 17768
rect 12032 17756 12038 17808
rect 12526 17796 12532 17808
rect 12268 17768 12532 17796
rect 9674 17728 9680 17740
rect 7392 17700 9680 17728
rect 9674 17688 9680 17700
rect 9732 17688 9738 17740
rect 11606 17688 11612 17740
rect 11664 17728 11670 17740
rect 12268 17737 12296 17768
rect 12526 17756 12532 17768
rect 12584 17756 12590 17808
rect 12621 17799 12679 17805
rect 12621 17765 12633 17799
rect 12667 17796 12679 17799
rect 12986 17796 12992 17808
rect 12667 17768 12992 17796
rect 12667 17765 12679 17768
rect 12621 17759 12679 17765
rect 12986 17756 12992 17768
rect 13044 17756 13050 17808
rect 12253 17731 12311 17737
rect 12253 17728 12265 17731
rect 11664 17700 12265 17728
rect 11664 17688 11670 17700
rect 12253 17697 12265 17700
rect 12299 17697 12311 17731
rect 12253 17691 12311 17697
rect 12342 17688 12348 17740
rect 12400 17728 12406 17740
rect 13372 17728 13400 17836
rect 14093 17833 14105 17836
rect 14139 17833 14151 17867
rect 14093 17827 14151 17833
rect 14642 17824 14648 17876
rect 14700 17864 14706 17876
rect 15105 17867 15163 17873
rect 14700 17836 15056 17864
rect 14700 17824 14706 17836
rect 13541 17799 13599 17805
rect 13541 17765 13553 17799
rect 13587 17796 13599 17799
rect 14734 17796 14740 17808
rect 13587 17768 14740 17796
rect 13587 17765 13599 17768
rect 13541 17759 13599 17765
rect 14734 17756 14740 17768
rect 14792 17756 14798 17808
rect 14826 17756 14832 17808
rect 14884 17756 14890 17808
rect 12400 17700 13400 17728
rect 12400 17688 12406 17700
rect 4801 17663 4859 17669
rect 4801 17629 4813 17663
rect 4847 17629 4859 17663
rect 4801 17623 4859 17629
rect 4890 17620 4896 17672
rect 4948 17660 4954 17672
rect 5077 17663 5135 17669
rect 5077 17660 5089 17663
rect 4948 17632 5089 17660
rect 4948 17620 4954 17632
rect 5077 17629 5089 17632
rect 5123 17629 5135 17663
rect 5077 17623 5135 17629
rect 5534 17620 5540 17672
rect 5592 17620 5598 17672
rect 5813 17663 5871 17669
rect 5813 17629 5825 17663
rect 5859 17660 5871 17663
rect 6454 17660 6460 17672
rect 5859 17632 6460 17660
rect 5859 17629 5871 17632
rect 5813 17623 5871 17629
rect 6454 17620 6460 17632
rect 6512 17620 6518 17672
rect 6546 17620 6552 17672
rect 6604 17660 6610 17672
rect 7745 17663 7803 17669
rect 7745 17660 7757 17663
rect 6604 17632 7757 17660
rect 6604 17620 6610 17632
rect 7745 17629 7757 17632
rect 7791 17660 7803 17663
rect 7834 17660 7840 17672
rect 7791 17632 7840 17660
rect 7791 17629 7803 17632
rect 7745 17623 7803 17629
rect 7834 17620 7840 17632
rect 7892 17620 7898 17672
rect 8570 17620 8576 17672
rect 8628 17660 8634 17672
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 8628 17632 9781 17660
rect 8628 17620 8634 17632
rect 9769 17629 9781 17632
rect 9815 17629 9827 17663
rect 9769 17623 9827 17629
rect 10045 17663 10103 17669
rect 10045 17629 10057 17663
rect 10091 17660 10103 17663
rect 10410 17660 10416 17672
rect 10091 17632 10416 17660
rect 10091 17629 10103 17632
rect 10045 17623 10103 17629
rect 10410 17620 10416 17632
rect 10468 17620 10474 17672
rect 10502 17620 10508 17672
rect 10560 17620 10566 17672
rect 11790 17620 11796 17672
rect 11848 17660 11854 17672
rect 12437 17663 12495 17669
rect 11848 17632 12204 17660
rect 11848 17620 11854 17632
rect 3752 17564 4016 17592
rect 3752 17552 3758 17564
rect 4246 17552 4252 17604
rect 4304 17592 4310 17604
rect 4304 17564 4936 17592
rect 4304 17552 4310 17564
rect 2682 17484 2688 17536
rect 2740 17496 2774 17536
rect 2961 17527 3019 17533
rect 2740 17484 2746 17496
rect 2961 17493 2973 17527
rect 3007 17524 3019 17527
rect 3142 17524 3148 17536
rect 3007 17496 3148 17524
rect 3007 17493 3019 17496
rect 2961 17487 3019 17493
rect 3142 17484 3148 17496
rect 3200 17484 3206 17536
rect 3234 17484 3240 17536
rect 3292 17484 3298 17536
rect 4614 17484 4620 17536
rect 4672 17484 4678 17536
rect 4908 17533 4936 17564
rect 7190 17552 7196 17604
rect 7248 17592 7254 17604
rect 12176 17601 12204 17632
rect 12437 17629 12449 17663
rect 12483 17660 12495 17663
rect 12483 17632 12664 17660
rect 12483 17629 12495 17632
rect 12437 17623 12495 17629
rect 12161 17595 12219 17601
rect 7248 17564 10824 17592
rect 7248 17552 7254 17564
rect 4893 17527 4951 17533
rect 4893 17493 4905 17527
rect 4939 17493 4951 17527
rect 4893 17487 4951 17493
rect 5350 17484 5356 17536
rect 5408 17484 5414 17536
rect 5626 17484 5632 17536
rect 5684 17484 5690 17536
rect 6454 17484 6460 17536
rect 6512 17524 6518 17536
rect 9122 17524 9128 17536
rect 6512 17496 9128 17524
rect 6512 17484 6518 17496
rect 9122 17484 9128 17496
rect 9180 17484 9186 17536
rect 10226 17484 10232 17536
rect 10284 17484 10290 17536
rect 10318 17484 10324 17536
rect 10376 17484 10382 17536
rect 10796 17524 10824 17564
rect 12161 17561 12173 17595
rect 12207 17592 12219 17595
rect 12636 17592 12664 17632
rect 12710 17620 12716 17672
rect 12768 17620 12774 17672
rect 13004 17632 13216 17660
rect 12802 17592 12808 17604
rect 12207 17564 12572 17592
rect 12636 17564 12808 17592
rect 12207 17561 12219 17564
rect 12161 17555 12219 17561
rect 12342 17524 12348 17536
rect 10796 17496 12348 17524
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 12544 17524 12572 17564
rect 12802 17552 12808 17564
rect 12860 17552 12866 17604
rect 12897 17527 12955 17533
rect 12897 17524 12909 17527
rect 12544 17496 12909 17524
rect 12897 17493 12909 17496
rect 12943 17524 12955 17527
rect 13004 17524 13032 17632
rect 13081 17595 13139 17601
rect 13081 17561 13093 17595
rect 13127 17561 13139 17595
rect 13188 17592 13216 17632
rect 13262 17620 13268 17672
rect 13320 17620 13326 17672
rect 13372 17660 13400 17700
rect 13449 17731 13507 17737
rect 13449 17697 13461 17731
rect 13495 17728 13507 17731
rect 13495 17700 14412 17728
rect 13495 17697 13507 17700
rect 13449 17691 13507 17697
rect 13725 17663 13783 17669
rect 13725 17660 13737 17663
rect 13372 17632 13737 17660
rect 13725 17629 13737 17632
rect 13771 17629 13783 17663
rect 13725 17623 13783 17629
rect 14274 17620 14280 17672
rect 14332 17620 14338 17672
rect 14384 17660 14412 17700
rect 14458 17688 14464 17740
rect 14516 17688 14522 17740
rect 14645 17663 14703 17669
rect 14645 17660 14657 17663
rect 14384 17632 14657 17660
rect 14645 17629 14657 17632
rect 14691 17629 14703 17663
rect 14752 17660 14780 17756
rect 15028 17728 15056 17836
rect 15105 17833 15117 17867
rect 15151 17833 15163 17867
rect 15105 17827 15163 17833
rect 15120 17796 15148 17827
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 17310 17864 17316 17876
rect 15252 17836 17316 17864
rect 15252 17824 15258 17836
rect 17310 17824 17316 17836
rect 17368 17824 17374 17876
rect 18046 17824 18052 17876
rect 18104 17864 18110 17876
rect 18104 17836 20116 17864
rect 18104 17824 18110 17836
rect 15286 17796 15292 17808
rect 15120 17768 15292 17796
rect 15286 17756 15292 17768
rect 15344 17796 15350 17808
rect 20088 17796 20116 17836
rect 20254 17824 20260 17876
rect 20312 17864 20318 17876
rect 21821 17867 21879 17873
rect 21821 17864 21833 17867
rect 20312 17836 21833 17864
rect 20312 17824 20318 17836
rect 21821 17833 21833 17836
rect 21867 17833 21879 17867
rect 21821 17827 21879 17833
rect 22186 17824 22192 17876
rect 22244 17864 22250 17876
rect 22646 17864 22652 17876
rect 22244 17836 22652 17864
rect 22244 17824 22250 17836
rect 22646 17824 22652 17836
rect 22704 17864 22710 17876
rect 22925 17867 22983 17873
rect 22925 17864 22937 17867
rect 22704 17836 22937 17864
rect 22704 17824 22710 17836
rect 22925 17833 22937 17836
rect 22971 17833 22983 17867
rect 22925 17827 22983 17833
rect 23385 17867 23443 17873
rect 23385 17833 23397 17867
rect 23431 17864 23443 17867
rect 23474 17864 23480 17876
rect 23431 17836 23480 17864
rect 23431 17833 23443 17836
rect 23385 17827 23443 17833
rect 23474 17824 23480 17836
rect 23532 17824 23538 17876
rect 26237 17867 26295 17873
rect 26237 17833 26249 17867
rect 26283 17833 26295 17867
rect 26237 17827 26295 17833
rect 24302 17796 24308 17808
rect 15344 17768 20024 17796
rect 20088 17768 24308 17796
rect 15344 17756 15350 17768
rect 16298 17728 16304 17740
rect 15028 17700 16304 17728
rect 16298 17688 16304 17700
rect 16356 17688 16362 17740
rect 17218 17688 17224 17740
rect 17276 17728 17282 17740
rect 17405 17731 17463 17737
rect 17405 17728 17417 17731
rect 17276 17700 17417 17728
rect 17276 17688 17282 17700
rect 17405 17697 17417 17700
rect 17451 17697 17463 17731
rect 17405 17691 17463 17697
rect 15013 17663 15071 17669
rect 15013 17660 15025 17663
rect 14752 17632 15025 17660
rect 14645 17623 14703 17629
rect 15013 17629 15025 17632
rect 15059 17629 15071 17663
rect 15013 17623 15071 17629
rect 15105 17663 15163 17669
rect 15105 17629 15117 17663
rect 15151 17660 15163 17663
rect 15194 17660 15200 17672
rect 15151 17632 15200 17660
rect 15151 17629 15163 17632
rect 15105 17623 15163 17629
rect 13188 17564 13860 17592
rect 13081 17555 13139 17561
rect 12943 17496 13032 17524
rect 13096 17524 13124 17555
rect 13354 17524 13360 17536
rect 13096 17496 13360 17524
rect 12943 17493 12955 17496
rect 12897 17487 12955 17493
rect 13354 17484 13360 17496
rect 13412 17484 13418 17536
rect 13832 17524 13860 17564
rect 13906 17552 13912 17604
rect 13964 17552 13970 17604
rect 14182 17552 14188 17604
rect 14240 17592 14246 17604
rect 14369 17595 14427 17601
rect 14369 17592 14381 17595
rect 14240 17564 14381 17592
rect 14240 17552 14246 17564
rect 14369 17561 14381 17564
rect 14415 17561 14427 17595
rect 14369 17555 14427 17561
rect 14734 17552 14740 17604
rect 14792 17592 14798 17604
rect 15120 17592 15148 17623
rect 15194 17620 15200 17632
rect 15252 17620 15258 17672
rect 16850 17620 16856 17672
rect 16908 17660 16914 17672
rect 17313 17663 17371 17669
rect 17313 17660 17325 17663
rect 16908 17632 17325 17660
rect 16908 17620 16914 17632
rect 17313 17629 17325 17632
rect 17359 17629 17371 17663
rect 19426 17660 19432 17672
rect 17313 17623 17371 17629
rect 19306 17632 19432 17660
rect 19306 17592 19334 17632
rect 19426 17620 19432 17632
rect 19484 17660 19490 17672
rect 19886 17660 19892 17672
rect 19484 17632 19892 17660
rect 19484 17620 19490 17632
rect 19886 17620 19892 17632
rect 19944 17620 19950 17672
rect 19996 17669 20024 17768
rect 24302 17756 24308 17768
rect 24360 17756 24366 17808
rect 26252 17740 26280 17827
rect 26694 17824 26700 17876
rect 26752 17864 26758 17876
rect 26789 17867 26847 17873
rect 26789 17864 26801 17867
rect 26752 17836 26801 17864
rect 26752 17824 26758 17836
rect 26789 17833 26801 17836
rect 26835 17864 26847 17867
rect 27249 17867 27307 17873
rect 26835 17836 27200 17864
rect 26835 17833 26847 17836
rect 26789 17827 26847 17833
rect 26510 17756 26516 17808
rect 26568 17796 26574 17808
rect 26568 17768 27016 17796
rect 26568 17756 26574 17768
rect 20622 17688 20628 17740
rect 20680 17688 20686 17740
rect 21910 17688 21916 17740
rect 21968 17688 21974 17740
rect 22278 17688 22284 17740
rect 22336 17728 22342 17740
rect 22646 17728 22652 17740
rect 22336 17700 22652 17728
rect 22336 17688 22342 17700
rect 22646 17688 22652 17700
rect 22704 17728 22710 17740
rect 23017 17731 23075 17737
rect 23017 17728 23029 17731
rect 22704 17700 23029 17728
rect 22704 17688 22710 17700
rect 23017 17697 23029 17700
rect 23063 17697 23075 17731
rect 23017 17691 23075 17697
rect 26142 17688 26148 17740
rect 26200 17688 26206 17740
rect 26234 17688 26240 17740
rect 26292 17688 26298 17740
rect 26988 17737 27016 17768
rect 26421 17731 26479 17737
rect 26421 17697 26433 17731
rect 26467 17728 26479 17731
rect 26973 17731 27031 17737
rect 26467 17700 26924 17728
rect 26467 17697 26479 17700
rect 26421 17691 26479 17697
rect 19981 17663 20039 17669
rect 19981 17629 19993 17663
rect 20027 17629 20039 17663
rect 20640 17660 20668 17688
rect 20809 17663 20867 17669
rect 20809 17660 20821 17663
rect 20640 17632 20821 17660
rect 19981 17623 20039 17629
rect 20809 17629 20821 17632
rect 20855 17629 20867 17663
rect 20809 17623 20867 17629
rect 14792 17564 15148 17592
rect 15212 17564 19334 17592
rect 20165 17595 20223 17601
rect 14792 17552 14798 17564
rect 15212 17524 15240 17564
rect 20165 17561 20177 17595
rect 20211 17592 20223 17595
rect 20530 17592 20536 17604
rect 20211 17564 20536 17592
rect 20211 17561 20223 17564
rect 20165 17555 20223 17561
rect 20530 17552 20536 17564
rect 20588 17552 20594 17604
rect 20622 17552 20628 17604
rect 20680 17552 20686 17604
rect 13832 17496 15240 17524
rect 15381 17527 15439 17533
rect 15381 17493 15393 17527
rect 15427 17524 15439 17527
rect 15470 17524 15476 17536
rect 15427 17496 15476 17524
rect 15427 17493 15439 17496
rect 15381 17487 15439 17493
rect 15470 17484 15476 17496
rect 15528 17484 15534 17536
rect 16114 17484 16120 17536
rect 16172 17524 16178 17536
rect 16666 17524 16672 17536
rect 16172 17496 16672 17524
rect 16172 17484 16178 17496
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 17681 17527 17739 17533
rect 17681 17493 17693 17527
rect 17727 17524 17739 17527
rect 18046 17524 18052 17536
rect 17727 17496 18052 17524
rect 17727 17493 17739 17496
rect 17681 17487 17739 17493
rect 18046 17484 18052 17496
rect 18104 17484 18110 17536
rect 19797 17527 19855 17533
rect 19797 17493 19809 17527
rect 19843 17524 19855 17527
rect 19886 17524 19892 17536
rect 19843 17496 19892 17524
rect 19843 17493 19855 17496
rect 19797 17487 19855 17493
rect 19886 17484 19892 17496
rect 19944 17484 19950 17536
rect 19978 17484 19984 17536
rect 20036 17524 20042 17536
rect 20441 17527 20499 17533
rect 20441 17524 20453 17527
rect 20036 17496 20453 17524
rect 20036 17484 20042 17496
rect 20441 17493 20453 17496
rect 20487 17493 20499 17527
rect 20824 17524 20852 17623
rect 21542 17620 21548 17672
rect 21600 17660 21606 17672
rect 22097 17663 22155 17669
rect 21600 17632 21956 17660
rect 21600 17620 21606 17632
rect 21818 17552 21824 17604
rect 21876 17552 21882 17604
rect 21928 17592 21956 17632
rect 22097 17629 22109 17663
rect 22143 17660 22155 17663
rect 22143 17632 22416 17660
rect 22143 17629 22155 17632
rect 22097 17623 22155 17629
rect 22388 17592 22416 17632
rect 22462 17620 22468 17672
rect 22520 17660 22526 17672
rect 22925 17663 22983 17669
rect 22925 17660 22937 17663
rect 22520 17632 22937 17660
rect 22520 17620 22526 17632
rect 22925 17629 22937 17632
rect 22971 17629 22983 17663
rect 22925 17623 22983 17629
rect 23198 17620 23204 17672
rect 23256 17620 23262 17672
rect 24320 17632 25084 17660
rect 24320 17592 24348 17632
rect 21928 17564 22324 17592
rect 22388 17564 24348 17592
rect 22186 17524 22192 17536
rect 20824 17496 22192 17524
rect 20441 17487 20499 17493
rect 22186 17484 22192 17496
rect 22244 17484 22250 17536
rect 22296 17533 22324 17564
rect 24394 17552 24400 17604
rect 24452 17552 24458 17604
rect 25056 17592 25084 17632
rect 25130 17620 25136 17672
rect 25188 17660 25194 17672
rect 26513 17663 26571 17669
rect 26513 17660 26525 17663
rect 25188 17632 26525 17660
rect 25188 17620 25194 17632
rect 26513 17629 26525 17632
rect 26559 17629 26571 17663
rect 26513 17623 26571 17629
rect 26142 17592 26148 17604
rect 25056 17564 26148 17592
rect 26142 17552 26148 17564
rect 26200 17552 26206 17604
rect 26237 17595 26295 17601
rect 26237 17561 26249 17595
rect 26283 17561 26295 17595
rect 26237 17555 26295 17561
rect 26789 17595 26847 17601
rect 26789 17561 26801 17595
rect 26835 17561 26847 17595
rect 26896 17592 26924 17700
rect 26973 17697 26985 17731
rect 27019 17697 27031 17731
rect 27172 17728 27200 17836
rect 27249 17833 27261 17867
rect 27295 17864 27307 17867
rect 27798 17864 27804 17876
rect 27295 17836 27804 17864
rect 27295 17833 27307 17836
rect 27249 17827 27307 17833
rect 27798 17824 27804 17836
rect 27856 17824 27862 17876
rect 30837 17867 30895 17873
rect 30837 17833 30849 17867
rect 30883 17864 30895 17867
rect 31018 17864 31024 17876
rect 30883 17836 31024 17864
rect 30883 17833 30895 17836
rect 30837 17827 30895 17833
rect 31018 17824 31024 17836
rect 31076 17824 31082 17876
rect 31386 17824 31392 17876
rect 31444 17864 31450 17876
rect 31481 17867 31539 17873
rect 31481 17864 31493 17867
rect 31444 17836 31493 17864
rect 31444 17824 31450 17836
rect 31481 17833 31493 17836
rect 31527 17833 31539 17867
rect 31481 17827 31539 17833
rect 27172 17700 28948 17728
rect 26973 17691 27031 17697
rect 28920 17672 28948 17700
rect 32214 17688 32220 17740
rect 32272 17688 32278 17740
rect 27065 17663 27123 17669
rect 27065 17629 27077 17663
rect 27111 17660 27123 17663
rect 27154 17660 27160 17672
rect 27111 17632 27160 17660
rect 27111 17629 27123 17632
rect 27065 17623 27123 17629
rect 27154 17620 27160 17632
rect 27212 17620 27218 17672
rect 28442 17620 28448 17672
rect 28500 17660 28506 17672
rect 28721 17663 28779 17669
rect 28721 17660 28733 17663
rect 28500 17632 28733 17660
rect 28500 17620 28506 17632
rect 28721 17629 28733 17632
rect 28767 17629 28779 17663
rect 28721 17623 28779 17629
rect 28902 17620 28908 17672
rect 28960 17620 28966 17672
rect 30374 17620 30380 17672
rect 30432 17660 30438 17672
rect 30653 17663 30711 17669
rect 30653 17660 30665 17663
rect 30432 17632 30665 17660
rect 30432 17620 30438 17632
rect 30653 17629 30665 17632
rect 30699 17629 30711 17663
rect 30653 17623 30711 17629
rect 30926 17620 30932 17672
rect 30984 17620 30990 17672
rect 31018 17620 31024 17672
rect 31076 17660 31082 17672
rect 31205 17663 31263 17669
rect 31205 17660 31217 17663
rect 31076 17632 31217 17660
rect 31076 17620 31082 17632
rect 31205 17629 31217 17632
rect 31251 17629 31263 17663
rect 31205 17623 31263 17629
rect 31297 17663 31355 17669
rect 31297 17629 31309 17663
rect 31343 17660 31355 17663
rect 31665 17663 31723 17669
rect 31665 17660 31677 17663
rect 31343 17632 31677 17660
rect 31343 17629 31355 17632
rect 31297 17623 31355 17629
rect 31665 17629 31677 17632
rect 31711 17629 31723 17663
rect 31665 17623 31723 17629
rect 28460 17592 28488 17620
rect 26896 17564 28488 17592
rect 26789 17555 26847 17561
rect 22281 17527 22339 17533
rect 22281 17493 22293 17527
rect 22327 17493 22339 17527
rect 22281 17487 22339 17493
rect 25958 17484 25964 17536
rect 26016 17524 26022 17536
rect 26252 17524 26280 17555
rect 26016 17496 26280 17524
rect 26016 17484 26022 17496
rect 26694 17484 26700 17536
rect 26752 17484 26758 17536
rect 26804 17524 26832 17555
rect 30466 17552 30472 17604
rect 30524 17592 30530 17604
rect 31113 17595 31171 17601
rect 31113 17592 31125 17595
rect 30524 17564 31125 17592
rect 30524 17552 30530 17564
rect 31113 17561 31125 17564
rect 31159 17561 31171 17595
rect 31113 17555 31171 17561
rect 27062 17524 27068 17536
rect 26804 17496 27068 17524
rect 27062 17484 27068 17496
rect 27120 17484 27126 17536
rect 28537 17527 28595 17533
rect 28537 17493 28549 17527
rect 28583 17524 28595 17527
rect 28626 17524 28632 17536
rect 28583 17496 28632 17524
rect 28583 17493 28595 17496
rect 28537 17487 28595 17493
rect 28626 17484 28632 17496
rect 28684 17484 28690 17536
rect 1104 17434 32844 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 32844 17434
rect 1104 17360 32844 17382
rect 3234 17320 3240 17332
rect 2424 17292 3240 17320
rect 2424 17193 2452 17292
rect 3234 17280 3240 17292
rect 3292 17280 3298 17332
rect 5534 17320 5540 17332
rect 4448 17292 5540 17320
rect 2593 17255 2651 17261
rect 2593 17221 2605 17255
rect 2639 17252 2651 17255
rect 3970 17252 3976 17264
rect 2639 17224 3976 17252
rect 2639 17221 2651 17224
rect 2593 17215 2651 17221
rect 3970 17212 3976 17224
rect 4028 17212 4034 17264
rect 4154 17212 4160 17264
rect 4212 17252 4218 17264
rect 4448 17261 4476 17292
rect 4433 17255 4491 17261
rect 4433 17252 4445 17255
rect 4212 17224 4445 17252
rect 4212 17212 4218 17224
rect 4433 17221 4445 17224
rect 4479 17221 4491 17255
rect 4433 17215 4491 17221
rect 4525 17255 4583 17261
rect 4525 17221 4537 17255
rect 4571 17252 4583 17255
rect 4706 17252 4712 17264
rect 4571 17224 4712 17252
rect 4571 17221 4583 17224
rect 4525 17215 4583 17221
rect 4706 17212 4712 17224
rect 4764 17212 4770 17264
rect 5460 17261 5488 17292
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 5813 17323 5871 17329
rect 5813 17289 5825 17323
rect 5859 17320 5871 17323
rect 6546 17320 6552 17332
rect 5859 17292 6552 17320
rect 5859 17289 5871 17292
rect 5813 17283 5871 17289
rect 6546 17280 6552 17292
rect 6604 17280 6610 17332
rect 7101 17323 7159 17329
rect 7101 17289 7113 17323
rect 7147 17320 7159 17323
rect 7190 17320 7196 17332
rect 7147 17292 7196 17320
rect 7147 17289 7159 17292
rect 7101 17283 7159 17289
rect 5445 17255 5503 17261
rect 5445 17221 5457 17255
rect 5491 17221 5503 17255
rect 6454 17252 6460 17264
rect 5445 17215 5503 17221
rect 5552 17224 6460 17252
rect 2409 17187 2467 17193
rect 2409 17153 2421 17187
rect 2455 17153 2467 17187
rect 2409 17147 2467 17153
rect 2682 17144 2688 17196
rect 2740 17144 2746 17196
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17184 2835 17187
rect 3878 17184 3884 17196
rect 2823 17156 3884 17184
rect 2823 17153 2835 17156
rect 2777 17147 2835 17153
rect 3878 17144 3884 17156
rect 3936 17144 3942 17196
rect 4246 17144 4252 17196
rect 4304 17144 4310 17196
rect 4614 17144 4620 17196
rect 4672 17144 4678 17196
rect 4798 17144 4804 17196
rect 4856 17184 4862 17196
rect 5552 17193 5580 17224
rect 6454 17212 6460 17224
rect 6512 17212 6518 17264
rect 7116 17252 7144 17283
rect 7190 17280 7196 17292
rect 7248 17280 7254 17332
rect 7282 17280 7288 17332
rect 7340 17320 7346 17332
rect 7340 17292 7604 17320
rect 7340 17280 7346 17292
rect 6564 17224 7144 17252
rect 5261 17187 5319 17193
rect 5261 17184 5273 17187
rect 4856 17156 5273 17184
rect 4856 17144 4862 17156
rect 5261 17153 5273 17156
rect 5307 17153 5319 17187
rect 5261 17147 5319 17153
rect 5537 17187 5595 17193
rect 5537 17153 5549 17187
rect 5583 17153 5595 17187
rect 5537 17147 5595 17153
rect 5629 17187 5687 17193
rect 5629 17153 5641 17187
rect 5675 17184 5687 17187
rect 5718 17184 5724 17196
rect 5675 17156 5724 17184
rect 5675 17153 5687 17156
rect 5629 17147 5687 17153
rect 4264 17116 4292 17144
rect 2746 17088 4292 17116
rect 4632 17116 4660 17144
rect 5644 17116 5672 17147
rect 5718 17144 5724 17156
rect 5776 17144 5782 17196
rect 6362 17144 6368 17196
rect 6420 17144 6426 17196
rect 6564 17193 6592 17224
rect 7374 17212 7380 17264
rect 7432 17212 7438 17264
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 6638 17144 6644 17196
rect 6696 17144 6702 17196
rect 6914 17144 6920 17196
rect 6972 17144 6978 17196
rect 7576 17193 7604 17292
rect 7650 17280 7656 17332
rect 7708 17320 7714 17332
rect 7708 17292 7972 17320
rect 7708 17280 7714 17292
rect 7193 17187 7251 17193
rect 7193 17153 7205 17187
rect 7239 17153 7251 17187
rect 7193 17147 7251 17153
rect 7469 17187 7527 17193
rect 7469 17153 7481 17187
rect 7515 17153 7527 17187
rect 7469 17147 7527 17153
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 7208 17116 7236 17147
rect 4632 17088 5672 17116
rect 5736 17088 7236 17116
rect 2746 17060 2774 17088
rect 2682 17008 2688 17060
rect 2740 17020 2774 17060
rect 3878 17048 3884 17060
rect 2976 17020 3884 17048
rect 2740 17008 2746 17020
rect 2976 16989 3004 17020
rect 3878 17008 3884 17020
rect 3936 17008 3942 17060
rect 4801 17051 4859 17057
rect 4801 17017 4813 17051
rect 4847 17048 4859 17051
rect 4982 17048 4988 17060
rect 4847 17020 4988 17048
rect 4847 17017 4859 17020
rect 4801 17011 4859 17017
rect 4982 17008 4988 17020
rect 5040 17008 5046 17060
rect 2961 16983 3019 16989
rect 2961 16949 2973 16983
rect 3007 16949 3019 16983
rect 2961 16943 3019 16949
rect 3142 16940 3148 16992
rect 3200 16980 3206 16992
rect 3694 16980 3700 16992
rect 3200 16952 3700 16980
rect 3200 16940 3206 16952
rect 3694 16940 3700 16952
rect 3752 16980 3758 16992
rect 5736 16980 5764 17088
rect 7282 17048 7288 17060
rect 6472 17020 7288 17048
rect 6472 16989 6500 17020
rect 7282 17008 7288 17020
rect 7340 17008 7346 17060
rect 7484 16992 7512 17147
rect 7650 17144 7656 17196
rect 7708 17184 7714 17196
rect 7837 17187 7895 17193
rect 7837 17184 7849 17187
rect 7708 17156 7849 17184
rect 7708 17144 7714 17156
rect 7837 17153 7849 17156
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 7944 17048 7972 17292
rect 8018 17280 8024 17332
rect 8076 17320 8082 17332
rect 10318 17320 10324 17332
rect 8076 17292 9996 17320
rect 8076 17280 8082 17292
rect 9309 17255 9367 17261
rect 9309 17221 9321 17255
rect 9355 17252 9367 17255
rect 9858 17252 9864 17264
rect 9355 17224 9674 17252
rect 9355 17221 9367 17224
rect 9309 17215 9367 17221
rect 8113 17187 8171 17193
rect 8113 17153 8125 17187
rect 8159 17184 8171 17187
rect 8202 17184 8208 17196
rect 8159 17156 8208 17184
rect 8159 17153 8171 17156
rect 8113 17147 8171 17153
rect 8202 17144 8208 17156
rect 8260 17144 8266 17196
rect 9122 17144 9128 17196
rect 9180 17184 9186 17196
rect 9493 17187 9551 17193
rect 9493 17184 9505 17187
rect 9180 17156 9505 17184
rect 9180 17144 9186 17156
rect 9493 17153 9505 17156
rect 9539 17153 9551 17187
rect 9493 17147 9551 17153
rect 8021 17119 8079 17125
rect 8021 17085 8033 17119
rect 8067 17116 8079 17119
rect 8662 17116 8668 17128
rect 8067 17088 8668 17116
rect 8067 17085 8079 17088
rect 8021 17079 8079 17085
rect 8662 17076 8668 17088
rect 8720 17076 8726 17128
rect 9646 17116 9674 17224
rect 9784 17224 9864 17252
rect 9784 17193 9812 17224
rect 9858 17212 9864 17224
rect 9916 17212 9922 17264
rect 9769 17187 9827 17193
rect 9769 17153 9781 17187
rect 9815 17153 9827 17187
rect 9968 17184 9996 17292
rect 10060 17292 10324 17320
rect 10060 17261 10088 17292
rect 10318 17280 10324 17292
rect 10376 17280 10382 17332
rect 10597 17323 10655 17329
rect 10597 17289 10609 17323
rect 10643 17320 10655 17323
rect 11054 17320 11060 17332
rect 10643 17292 11060 17320
rect 10643 17289 10655 17292
rect 10597 17283 10655 17289
rect 11054 17280 11060 17292
rect 11112 17280 11118 17332
rect 11790 17280 11796 17332
rect 11848 17320 11854 17332
rect 12618 17320 12624 17332
rect 11848 17292 12624 17320
rect 11848 17280 11854 17292
rect 12618 17280 12624 17292
rect 12676 17280 12682 17332
rect 12710 17280 12716 17332
rect 12768 17320 12774 17332
rect 15010 17320 15016 17332
rect 12768 17292 15016 17320
rect 12768 17280 12774 17292
rect 15010 17280 15016 17292
rect 15068 17280 15074 17332
rect 15105 17323 15163 17329
rect 15105 17289 15117 17323
rect 15151 17320 15163 17323
rect 15286 17320 15292 17332
rect 15151 17292 15292 17320
rect 15151 17289 15163 17292
rect 15105 17283 15163 17289
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 15654 17280 15660 17332
rect 15712 17320 15718 17332
rect 17770 17320 17776 17332
rect 15712 17292 17776 17320
rect 15712 17280 15718 17292
rect 17770 17280 17776 17292
rect 17828 17280 17834 17332
rect 17862 17280 17868 17332
rect 17920 17320 17926 17332
rect 18141 17323 18199 17329
rect 18141 17320 18153 17323
rect 17920 17292 18153 17320
rect 17920 17280 17926 17292
rect 18141 17289 18153 17292
rect 18187 17320 18199 17323
rect 24394 17320 24400 17332
rect 18187 17292 24400 17320
rect 18187 17289 18199 17292
rect 18141 17283 18199 17289
rect 24394 17280 24400 17292
rect 24452 17280 24458 17332
rect 24673 17323 24731 17329
rect 24673 17289 24685 17323
rect 24719 17320 24731 17323
rect 27246 17320 27252 17332
rect 24719 17292 25636 17320
rect 24719 17289 24731 17292
rect 24673 17283 24731 17289
rect 10045 17255 10103 17261
rect 10045 17221 10057 17255
rect 10091 17221 10103 17255
rect 10045 17215 10103 17221
rect 10134 17212 10140 17264
rect 10192 17212 10198 17264
rect 10336 17252 10364 17280
rect 10336 17224 11376 17252
rect 10321 17187 10379 17193
rect 10321 17184 10333 17187
rect 9968 17156 10333 17184
rect 9769 17147 9827 17153
rect 10321 17153 10333 17156
rect 10367 17153 10379 17187
rect 10321 17147 10379 17153
rect 10410 17144 10416 17196
rect 10468 17144 10474 17196
rect 10502 17144 10508 17196
rect 10560 17184 10566 17196
rect 10873 17187 10931 17193
rect 10873 17184 10885 17187
rect 10560 17156 10885 17184
rect 10560 17144 10566 17156
rect 10873 17153 10885 17156
rect 10919 17153 10931 17187
rect 10873 17147 10931 17153
rect 11054 17144 11060 17196
rect 11112 17144 11118 17196
rect 11149 17187 11207 17193
rect 11149 17153 11161 17187
rect 11195 17184 11207 17187
rect 11238 17184 11244 17196
rect 11195 17156 11244 17184
rect 11195 17153 11207 17156
rect 11149 17147 11207 17153
rect 11238 17144 11244 17156
rect 11296 17144 11302 17196
rect 11348 17184 11376 17224
rect 12158 17212 12164 17264
rect 12216 17252 12222 17264
rect 12253 17255 12311 17261
rect 12253 17252 12265 17255
rect 12216 17224 12265 17252
rect 12216 17212 12222 17224
rect 12253 17221 12265 17224
rect 12299 17221 12311 17255
rect 12253 17215 12311 17221
rect 12342 17212 12348 17264
rect 12400 17252 12406 17264
rect 12400 17224 15884 17252
rect 12400 17212 12406 17224
rect 11348 17156 11560 17184
rect 9858 17116 9864 17128
rect 9646 17088 9864 17116
rect 9858 17076 9864 17088
rect 9916 17076 9922 17128
rect 9953 17119 10011 17125
rect 9953 17085 9965 17119
rect 9999 17116 10011 17119
rect 10226 17116 10232 17128
rect 9999 17088 10232 17116
rect 9999 17085 10011 17088
rect 9953 17079 10011 17085
rect 10226 17076 10232 17088
rect 10284 17116 10290 17128
rect 11532 17116 11560 17156
rect 11698 17144 11704 17196
rect 11756 17144 11762 17196
rect 11974 17144 11980 17196
rect 12032 17184 12038 17196
rect 12529 17187 12587 17193
rect 12529 17184 12541 17187
rect 12032 17156 12541 17184
rect 12032 17144 12038 17156
rect 12529 17153 12541 17156
rect 12575 17153 12587 17187
rect 12529 17147 12587 17153
rect 13814 17144 13820 17196
rect 13872 17184 13878 17196
rect 13909 17187 13967 17193
rect 13909 17184 13921 17187
rect 13872 17156 13921 17184
rect 13872 17144 13878 17156
rect 13909 17153 13921 17156
rect 13955 17153 13967 17187
rect 13909 17147 13967 17153
rect 14458 17144 14464 17196
rect 14516 17184 14522 17196
rect 14737 17187 14795 17193
rect 14737 17184 14749 17187
rect 14516 17156 14749 17184
rect 14516 17144 14522 17156
rect 14737 17153 14749 17156
rect 14783 17153 14795 17187
rect 15856 17184 15884 17224
rect 15930 17212 15936 17264
rect 15988 17252 15994 17264
rect 16390 17252 16396 17264
rect 15988 17224 16396 17252
rect 15988 17212 15994 17224
rect 16390 17212 16396 17224
rect 16448 17212 16454 17264
rect 16669 17255 16727 17261
rect 16669 17221 16681 17255
rect 16715 17252 16727 17255
rect 17954 17252 17960 17264
rect 16715 17224 17960 17252
rect 16715 17221 16727 17224
rect 16669 17215 16727 17221
rect 17954 17212 17960 17224
rect 18012 17212 18018 17264
rect 18046 17212 18052 17264
rect 18104 17252 18110 17264
rect 22002 17252 22008 17264
rect 18104 17224 22008 17252
rect 18104 17212 18110 17224
rect 22002 17212 22008 17224
rect 22060 17212 22066 17264
rect 22554 17252 22560 17264
rect 22112 17224 22560 17252
rect 16574 17184 16580 17196
rect 15856 17156 16580 17184
rect 14737 17147 14795 17153
rect 16574 17144 16580 17156
rect 16632 17184 16638 17196
rect 17586 17184 17592 17196
rect 16632 17156 17592 17184
rect 16632 17144 16638 17156
rect 17586 17144 17592 17156
rect 17644 17144 17650 17196
rect 19610 17144 19616 17196
rect 19668 17184 19674 17196
rect 22112 17193 22140 17224
rect 22554 17212 22560 17224
rect 22612 17212 22618 17264
rect 23842 17212 23848 17264
rect 23900 17252 23906 17264
rect 25608 17261 25636 17292
rect 27172 17292 27252 17320
rect 25593 17255 25651 17261
rect 23900 17224 24532 17252
rect 23900 17212 23906 17224
rect 21913 17187 21971 17193
rect 21913 17184 21925 17187
rect 19668 17156 21925 17184
rect 19668 17144 19674 17156
rect 21913 17153 21925 17156
rect 21959 17153 21971 17187
rect 21913 17147 21971 17153
rect 22097 17187 22155 17193
rect 22097 17153 22109 17187
rect 22143 17153 22155 17187
rect 22097 17147 22155 17153
rect 22189 17187 22247 17193
rect 22189 17153 22201 17187
rect 22235 17153 22247 17187
rect 22189 17147 22247 17153
rect 22741 17187 22799 17193
rect 22741 17153 22753 17187
rect 22787 17184 22799 17187
rect 23198 17184 23204 17196
rect 22787 17156 23204 17184
rect 22787 17153 22799 17156
rect 22741 17147 22799 17153
rect 11885 17119 11943 17125
rect 11885 17116 11897 17119
rect 10284 17088 10640 17116
rect 11532 17088 11897 17116
rect 10284 17076 10290 17088
rect 9585 17051 9643 17057
rect 7944 17020 8156 17048
rect 3752 16952 5764 16980
rect 6457 16983 6515 16989
rect 3752 16940 3758 16952
rect 6457 16949 6469 16983
rect 6503 16949 6515 16983
rect 6457 16943 6515 16949
rect 6546 16940 6552 16992
rect 6604 16980 6610 16992
rect 6825 16983 6883 16989
rect 6825 16980 6837 16983
rect 6604 16952 6837 16980
rect 6604 16940 6610 16952
rect 6825 16949 6837 16952
rect 6871 16949 6883 16983
rect 6825 16943 6883 16949
rect 7466 16940 7472 16992
rect 7524 16940 7530 16992
rect 7650 16940 7656 16992
rect 7708 16980 7714 16992
rect 8128 16989 8156 17020
rect 9585 17017 9597 17051
rect 9631 17048 9643 17051
rect 10612 17048 10640 17088
rect 11885 17085 11897 17088
rect 11931 17116 11943 17119
rect 12158 17116 12164 17128
rect 11931 17088 12164 17116
rect 11931 17085 11943 17088
rect 11885 17079 11943 17085
rect 12158 17076 12164 17088
rect 12216 17076 12222 17128
rect 12345 17119 12403 17125
rect 12345 17085 12357 17119
rect 12391 17085 12403 17119
rect 12345 17079 12403 17085
rect 11333 17051 11391 17057
rect 9631 17020 10180 17048
rect 10612 17020 11008 17048
rect 9631 17017 9643 17020
rect 9585 17011 9643 17017
rect 7745 16983 7803 16989
rect 7745 16980 7757 16983
rect 7708 16952 7757 16980
rect 7708 16940 7714 16952
rect 7745 16949 7757 16952
rect 7791 16949 7803 16983
rect 7745 16943 7803 16949
rect 8113 16983 8171 16989
rect 8113 16949 8125 16983
rect 8159 16980 8171 16983
rect 8202 16980 8208 16992
rect 8159 16952 8208 16980
rect 8159 16949 8171 16952
rect 8113 16943 8171 16949
rect 8202 16940 8208 16952
rect 8260 16940 8266 16992
rect 8297 16983 8355 16989
rect 8297 16949 8309 16983
rect 8343 16980 8355 16983
rect 8386 16980 8392 16992
rect 8343 16952 8392 16980
rect 8343 16949 8355 16952
rect 8297 16943 8355 16949
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 9125 16983 9183 16989
rect 9125 16949 9137 16983
rect 9171 16980 9183 16983
rect 9766 16980 9772 16992
rect 9171 16952 9772 16980
rect 9171 16949 9183 16952
rect 9125 16943 9183 16949
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 10152 16989 10180 17020
rect 10137 16983 10195 16989
rect 10137 16949 10149 16983
rect 10183 16949 10195 16983
rect 10137 16943 10195 16949
rect 10870 16940 10876 16992
rect 10928 16940 10934 16992
rect 10980 16980 11008 17020
rect 11333 17017 11345 17051
rect 11379 17048 11391 17051
rect 12360 17048 12388 17079
rect 14826 17076 14832 17128
rect 14884 17076 14890 17128
rect 14918 17076 14924 17128
rect 14976 17116 14982 17128
rect 17862 17116 17868 17128
rect 14976 17088 17868 17116
rect 14976 17076 14982 17088
rect 17862 17076 17868 17088
rect 17920 17076 17926 17128
rect 18230 17076 18236 17128
rect 18288 17116 18294 17128
rect 20254 17116 20260 17128
rect 18288 17088 20260 17116
rect 18288 17076 18294 17088
rect 20254 17076 20260 17088
rect 20312 17076 20318 17128
rect 20622 17076 20628 17128
rect 20680 17116 20686 17128
rect 22204 17116 22232 17147
rect 23198 17144 23204 17156
rect 23256 17144 23262 17196
rect 24210 17144 24216 17196
rect 24268 17144 24274 17196
rect 24302 17144 24308 17196
rect 24360 17184 24366 17196
rect 24504 17193 24532 17224
rect 25593 17221 25605 17255
rect 25639 17221 25651 17255
rect 25593 17215 25651 17221
rect 24397 17187 24455 17193
rect 24397 17184 24409 17187
rect 24360 17156 24409 17184
rect 24360 17144 24366 17156
rect 24397 17153 24409 17156
rect 24443 17153 24455 17187
rect 24397 17147 24455 17153
rect 24489 17187 24547 17193
rect 24489 17153 24501 17187
rect 24535 17153 24547 17187
rect 24489 17147 24547 17153
rect 25774 17144 25780 17196
rect 25832 17144 25838 17196
rect 26142 17144 26148 17196
rect 26200 17184 26206 17196
rect 26878 17184 26884 17196
rect 26200 17156 26884 17184
rect 26200 17144 26206 17156
rect 26878 17144 26884 17156
rect 26936 17184 26942 17196
rect 27172 17193 27200 17292
rect 27246 17280 27252 17292
rect 27304 17280 27310 17332
rect 27433 17323 27491 17329
rect 27433 17289 27445 17323
rect 27479 17320 27491 17323
rect 28629 17323 28687 17329
rect 27479 17292 28212 17320
rect 27479 17289 27491 17292
rect 27433 17283 27491 17289
rect 28184 17261 28212 17292
rect 28629 17289 28641 17323
rect 28675 17320 28687 17323
rect 30926 17320 30932 17332
rect 28675 17292 30932 17320
rect 28675 17289 28687 17292
rect 28629 17283 28687 17289
rect 30926 17280 30932 17292
rect 30984 17280 30990 17332
rect 28169 17255 28227 17261
rect 27264 17224 27936 17252
rect 27264 17193 27292 17224
rect 26973 17187 27031 17193
rect 26973 17184 26985 17187
rect 26936 17156 26985 17184
rect 26936 17144 26942 17156
rect 26973 17153 26985 17156
rect 27019 17153 27031 17187
rect 26973 17147 27031 17153
rect 27157 17187 27215 17193
rect 27157 17153 27169 17187
rect 27203 17153 27215 17187
rect 27157 17147 27215 17153
rect 27249 17187 27307 17193
rect 27249 17153 27261 17187
rect 27295 17153 27307 17187
rect 27249 17147 27307 17153
rect 22833 17119 22891 17125
rect 22833 17116 22845 17119
rect 20680 17088 22845 17116
rect 20680 17076 20686 17088
rect 22833 17085 22845 17088
rect 22879 17085 22891 17119
rect 22833 17079 22891 17085
rect 23474 17076 23480 17128
rect 23532 17116 23538 17128
rect 27264 17116 27292 17147
rect 27522 17144 27528 17196
rect 27580 17184 27586 17196
rect 27908 17193 27936 17224
rect 28169 17221 28181 17255
rect 28215 17221 28227 17255
rect 28905 17255 28963 17261
rect 28905 17252 28917 17255
rect 28169 17215 28227 17221
rect 28460 17224 28917 17252
rect 28460 17196 28488 17224
rect 28905 17221 28917 17224
rect 28951 17221 28963 17255
rect 28905 17215 28963 17221
rect 27617 17187 27675 17193
rect 27617 17184 27629 17187
rect 27580 17156 27629 17184
rect 27580 17144 27586 17156
rect 27617 17153 27629 17156
rect 27663 17153 27675 17187
rect 27617 17147 27675 17153
rect 27893 17187 27951 17193
rect 27893 17153 27905 17187
rect 27939 17153 27951 17187
rect 27893 17147 27951 17153
rect 28442 17144 28448 17196
rect 28500 17144 28506 17196
rect 28534 17144 28540 17196
rect 28592 17184 28598 17196
rect 28721 17187 28779 17193
rect 28721 17184 28733 17187
rect 28592 17156 28733 17184
rect 28592 17144 28598 17156
rect 28721 17153 28733 17156
rect 28767 17153 28779 17187
rect 28721 17147 28779 17153
rect 30561 17187 30619 17193
rect 30561 17153 30573 17187
rect 30607 17184 30619 17187
rect 30650 17184 30656 17196
rect 30607 17156 30656 17184
rect 30607 17153 30619 17156
rect 30561 17147 30619 17153
rect 30650 17144 30656 17156
rect 30708 17144 30714 17196
rect 30828 17187 30886 17193
rect 30828 17153 30840 17187
rect 30874 17184 30886 17187
rect 31570 17184 31576 17196
rect 30874 17156 31576 17184
rect 30874 17153 30886 17156
rect 30828 17147 30886 17153
rect 31570 17144 31576 17156
rect 31628 17144 31634 17196
rect 32217 17187 32275 17193
rect 32217 17184 32229 17187
rect 31956 17156 32229 17184
rect 23532 17088 27292 17116
rect 23532 17076 23538 17088
rect 27706 17076 27712 17128
rect 27764 17076 27770 17128
rect 27798 17076 27804 17128
rect 27856 17116 27862 17128
rect 28261 17119 28319 17125
rect 28261 17116 28273 17119
rect 27856 17088 28273 17116
rect 27856 17076 27862 17088
rect 28261 17085 28273 17088
rect 28307 17085 28319 17119
rect 28261 17079 28319 17085
rect 11379 17020 12388 17048
rect 11379 17017 11391 17020
rect 11333 17011 11391 17017
rect 13906 17008 13912 17060
rect 13964 17048 13970 17060
rect 14093 17051 14151 17057
rect 14093 17048 14105 17051
rect 13964 17020 14105 17048
rect 13964 17008 13970 17020
rect 14093 17017 14105 17020
rect 14139 17048 14151 17051
rect 16850 17048 16856 17060
rect 14139 17020 16856 17048
rect 14139 17017 14151 17020
rect 14093 17011 14151 17017
rect 16850 17008 16856 17020
rect 16908 17008 16914 17060
rect 18138 17008 18144 17060
rect 18196 17048 18202 17060
rect 22278 17048 22284 17060
rect 18196 17020 22284 17048
rect 18196 17008 18202 17020
rect 22278 17008 22284 17020
rect 22336 17008 22342 17060
rect 22373 17051 22431 17057
rect 22373 17017 22385 17051
rect 22419 17048 22431 17051
rect 24118 17048 24124 17060
rect 22419 17020 24124 17048
rect 22419 17017 22431 17020
rect 22373 17011 22431 17017
rect 24118 17008 24124 17020
rect 24176 17048 24182 17060
rect 31956 17057 31984 17156
rect 32217 17153 32229 17156
rect 32263 17184 32275 17187
rect 32306 17184 32312 17196
rect 32263 17156 32312 17184
rect 32263 17153 32275 17156
rect 32217 17147 32275 17153
rect 32306 17144 32312 17156
rect 32364 17144 32370 17196
rect 25961 17051 26019 17057
rect 24176 17020 25912 17048
rect 24176 17008 24182 17020
rect 11701 16983 11759 16989
rect 11701 16980 11713 16983
rect 10980 16952 11713 16980
rect 11701 16949 11713 16952
rect 11747 16949 11759 16983
rect 11701 16943 11759 16949
rect 12158 16940 12164 16992
rect 12216 16940 12222 16992
rect 12250 16940 12256 16992
rect 12308 16940 12314 16992
rect 12710 16940 12716 16992
rect 12768 16940 12774 16992
rect 12802 16940 12808 16992
rect 12860 16980 12866 16992
rect 13998 16980 14004 16992
rect 12860 16952 14004 16980
rect 12860 16940 12866 16952
rect 13998 16940 14004 16952
rect 14056 16940 14062 16992
rect 14182 16940 14188 16992
rect 14240 16980 14246 16992
rect 14737 16983 14795 16989
rect 14737 16980 14749 16983
rect 14240 16952 14749 16980
rect 14240 16940 14246 16952
rect 14737 16949 14749 16952
rect 14783 16949 14795 16983
rect 14737 16943 14795 16949
rect 16022 16940 16028 16992
rect 16080 16980 16086 16992
rect 16942 16980 16948 16992
rect 16080 16952 16948 16980
rect 16080 16940 16086 16952
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17770 16940 17776 16992
rect 17828 16980 17834 16992
rect 21913 16983 21971 16989
rect 21913 16980 21925 16983
rect 17828 16952 21925 16980
rect 17828 16940 17834 16952
rect 21913 16949 21925 16952
rect 21959 16980 21971 16983
rect 22741 16983 22799 16989
rect 22741 16980 22753 16983
rect 21959 16952 22753 16980
rect 21959 16949 21971 16952
rect 21913 16943 21971 16949
rect 22741 16949 22753 16952
rect 22787 16949 22799 16983
rect 22741 16943 22799 16949
rect 23106 16940 23112 16992
rect 23164 16940 23170 16992
rect 23842 16940 23848 16992
rect 23900 16980 23906 16992
rect 24029 16983 24087 16989
rect 24029 16980 24041 16983
rect 23900 16952 24041 16980
rect 23900 16940 23906 16952
rect 24029 16949 24041 16952
rect 24075 16949 24087 16983
rect 24029 16943 24087 16949
rect 24210 16940 24216 16992
rect 24268 16980 24274 16992
rect 24489 16983 24547 16989
rect 24489 16980 24501 16983
rect 24268 16952 24501 16980
rect 24268 16940 24274 16952
rect 24489 16949 24501 16952
rect 24535 16980 24547 16983
rect 24670 16980 24676 16992
rect 24535 16952 24676 16980
rect 24535 16949 24547 16952
rect 24489 16943 24547 16949
rect 24670 16940 24676 16952
rect 24728 16940 24734 16992
rect 25884 16980 25912 17020
rect 25961 17017 25973 17051
rect 26007 17048 26019 17051
rect 31941 17051 31999 17057
rect 26007 17020 28212 17048
rect 26007 17017 26019 17020
rect 25961 17011 26019 17017
rect 26973 16983 27031 16989
rect 26973 16980 26985 16983
rect 25884 16952 26985 16980
rect 26973 16949 26985 16952
rect 27019 16980 27031 16983
rect 27617 16983 27675 16989
rect 27617 16980 27629 16983
rect 27019 16952 27629 16980
rect 27019 16949 27031 16952
rect 26973 16943 27031 16949
rect 27617 16949 27629 16952
rect 27663 16949 27675 16983
rect 27617 16943 27675 16949
rect 28074 16940 28080 16992
rect 28132 16940 28138 16992
rect 28184 16989 28212 17020
rect 31941 17017 31953 17051
rect 31987 17017 31999 17051
rect 31941 17011 31999 17017
rect 32398 17008 32404 17060
rect 32456 17008 32462 17060
rect 28169 16983 28227 16989
rect 28169 16949 28181 16983
rect 28215 16949 28227 16983
rect 28169 16943 28227 16949
rect 29089 16983 29147 16989
rect 29089 16949 29101 16983
rect 29135 16980 29147 16983
rect 30282 16980 30288 16992
rect 29135 16952 30288 16980
rect 29135 16949 29147 16952
rect 29089 16943 29147 16949
rect 30282 16940 30288 16952
rect 30340 16940 30346 16992
rect 1104 16890 32844 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 32844 16890
rect 1104 16816 32844 16838
rect 3234 16736 3240 16788
rect 3292 16776 3298 16788
rect 3510 16776 3516 16788
rect 3292 16748 3516 16776
rect 3292 16736 3298 16748
rect 3510 16736 3516 16748
rect 3568 16776 3574 16788
rect 7466 16776 7472 16788
rect 3568 16748 7472 16776
rect 3568 16736 3574 16748
rect 7466 16736 7472 16748
rect 7524 16736 7530 16788
rect 8018 16736 8024 16788
rect 8076 16736 8082 16788
rect 8389 16779 8447 16785
rect 8389 16745 8401 16779
rect 8435 16776 8447 16779
rect 8478 16776 8484 16788
rect 8435 16748 8484 16776
rect 8435 16745 8447 16748
rect 8389 16739 8447 16745
rect 8478 16736 8484 16748
rect 8536 16736 8542 16788
rect 9953 16779 10011 16785
rect 9953 16745 9965 16779
rect 9999 16776 10011 16779
rect 10410 16776 10416 16788
rect 9999 16748 10416 16776
rect 9999 16745 10011 16748
rect 9953 16739 10011 16745
rect 10410 16736 10416 16748
rect 10468 16736 10474 16788
rect 10686 16736 10692 16788
rect 10744 16776 10750 16788
rect 11790 16776 11796 16788
rect 10744 16748 11796 16776
rect 10744 16736 10750 16748
rect 11790 16736 11796 16748
rect 11848 16736 11854 16788
rect 12158 16736 12164 16788
rect 12216 16776 12222 16788
rect 12805 16779 12863 16785
rect 12805 16776 12817 16779
rect 12216 16748 12817 16776
rect 12216 16736 12222 16748
rect 12805 16745 12817 16748
rect 12851 16745 12863 16779
rect 12805 16739 12863 16745
rect 13170 16736 13176 16788
rect 13228 16776 13234 16788
rect 13265 16779 13323 16785
rect 13265 16776 13277 16779
rect 13228 16748 13277 16776
rect 13228 16736 13234 16748
rect 13265 16745 13277 16748
rect 13311 16745 13323 16779
rect 13265 16739 13323 16745
rect 13998 16736 14004 16788
rect 14056 16776 14062 16788
rect 15654 16776 15660 16788
rect 14056 16748 15660 16776
rect 14056 16736 14062 16748
rect 15654 16736 15660 16748
rect 15712 16736 15718 16788
rect 15749 16779 15807 16785
rect 15749 16745 15761 16779
rect 15795 16776 15807 16779
rect 15930 16776 15936 16788
rect 15795 16748 15936 16776
rect 15795 16745 15807 16748
rect 15749 16739 15807 16745
rect 15930 16736 15936 16748
rect 15988 16736 15994 16788
rect 16022 16736 16028 16788
rect 16080 16736 16086 16788
rect 16482 16736 16488 16788
rect 16540 16736 16546 16788
rect 16574 16736 16580 16788
rect 16632 16776 16638 16788
rect 16669 16779 16727 16785
rect 16669 16776 16681 16779
rect 16632 16748 16681 16776
rect 16632 16736 16638 16748
rect 16669 16745 16681 16748
rect 16715 16745 16727 16779
rect 16669 16739 16727 16745
rect 17129 16779 17187 16785
rect 17129 16745 17141 16779
rect 17175 16745 17187 16779
rect 17129 16739 17187 16745
rect 474 16668 480 16720
rect 532 16708 538 16720
rect 532 16680 4220 16708
rect 532 16668 538 16680
rect 3602 16640 3608 16652
rect 2976 16612 3608 16640
rect 2976 16584 3004 16612
rect 3602 16600 3608 16612
rect 3660 16600 3666 16652
rect 842 16532 848 16584
rect 900 16572 906 16584
rect 1397 16575 1455 16581
rect 1397 16572 1409 16575
rect 900 16544 1409 16572
rect 900 16532 906 16544
rect 1397 16541 1409 16544
rect 1443 16541 1455 16575
rect 1397 16535 1455 16541
rect 2682 16532 2688 16584
rect 2740 16532 2746 16584
rect 2958 16532 2964 16584
rect 3016 16532 3022 16584
rect 3050 16532 3056 16584
rect 3108 16532 3114 16584
rect 2406 16464 2412 16516
rect 2464 16504 2470 16516
rect 2590 16504 2596 16516
rect 2464 16476 2596 16504
rect 2464 16464 2470 16476
rect 2590 16464 2596 16476
rect 2648 16504 2654 16516
rect 2869 16507 2927 16513
rect 2869 16504 2881 16507
rect 2648 16476 2881 16504
rect 2648 16464 2654 16476
rect 2869 16473 2881 16476
rect 2915 16473 2927 16507
rect 2869 16467 2927 16473
rect 1578 16396 1584 16448
rect 1636 16396 1642 16448
rect 2222 16396 2228 16448
rect 2280 16436 2286 16448
rect 3068 16436 3096 16532
rect 2280 16408 3096 16436
rect 2280 16396 2286 16408
rect 3234 16396 3240 16448
rect 3292 16396 3298 16448
rect 4192 16436 4220 16680
rect 4430 16668 4436 16720
rect 4488 16708 4494 16720
rect 5994 16708 6000 16720
rect 4488 16680 6000 16708
rect 4488 16668 4494 16680
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 9766 16668 9772 16720
rect 9824 16708 9830 16720
rect 11974 16708 11980 16720
rect 9824 16680 11980 16708
rect 9824 16668 9830 16680
rect 11974 16668 11980 16680
rect 12032 16668 12038 16720
rect 14826 16708 14832 16720
rect 12084 16680 14832 16708
rect 4522 16600 4528 16652
rect 4580 16600 4586 16652
rect 4982 16600 4988 16652
rect 5040 16640 5046 16652
rect 5040 16612 8064 16640
rect 5040 16600 5046 16612
rect 4341 16575 4399 16581
rect 4341 16541 4353 16575
rect 4387 16572 4399 16575
rect 4540 16572 4568 16600
rect 4387 16544 4568 16572
rect 4387 16541 4399 16544
rect 4341 16535 4399 16541
rect 4614 16532 4620 16584
rect 4672 16532 4678 16584
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16572 4767 16575
rect 5166 16572 5172 16584
rect 4755 16544 5172 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 5166 16532 5172 16544
rect 5224 16532 5230 16584
rect 5350 16532 5356 16584
rect 5408 16532 5414 16584
rect 5534 16532 5540 16584
rect 5592 16532 5598 16584
rect 5718 16532 5724 16584
rect 5776 16532 5782 16584
rect 6086 16532 6092 16584
rect 6144 16572 6150 16584
rect 7466 16572 7472 16584
rect 6144 16544 7472 16572
rect 6144 16532 6150 16544
rect 7466 16532 7472 16544
rect 7524 16532 7530 16584
rect 4522 16464 4528 16516
rect 4580 16464 4586 16516
rect 5626 16464 5632 16516
rect 5684 16464 5690 16516
rect 8036 16504 8064 16612
rect 8294 16600 8300 16652
rect 8352 16640 8358 16652
rect 8352 16612 9628 16640
rect 8352 16600 8358 16612
rect 8386 16532 8392 16584
rect 8444 16532 8450 16584
rect 9493 16575 9551 16581
rect 9493 16541 9505 16575
rect 9539 16541 9551 16575
rect 9600 16572 9628 16612
rect 9858 16600 9864 16652
rect 9916 16640 9922 16652
rect 12084 16640 12112 16680
rect 14826 16668 14832 16680
rect 14884 16668 14890 16720
rect 14921 16711 14979 16717
rect 14921 16677 14933 16711
rect 14967 16708 14979 16711
rect 15010 16708 15016 16720
rect 14967 16680 15016 16708
rect 14967 16677 14979 16680
rect 14921 16671 14979 16677
rect 15010 16668 15016 16680
rect 15068 16668 15074 16720
rect 15378 16668 15384 16720
rect 15436 16708 15442 16720
rect 16942 16708 16948 16720
rect 15436 16680 15608 16708
rect 15436 16668 15442 16680
rect 15580 16649 15608 16680
rect 15764 16680 16948 16708
rect 9916 16612 12112 16640
rect 15565 16643 15623 16649
rect 9916 16600 9922 16612
rect 15565 16609 15577 16643
rect 15611 16609 15623 16643
rect 15565 16603 15623 16609
rect 9600 16544 11836 16572
rect 9493 16535 9551 16541
rect 9508 16504 9536 16535
rect 8036 16476 9536 16504
rect 9508 16448 9536 16476
rect 9950 16464 9956 16516
rect 10008 16504 10014 16516
rect 10137 16507 10195 16513
rect 10137 16504 10149 16507
rect 10008 16476 10149 16504
rect 10008 16464 10014 16476
rect 10137 16473 10149 16476
rect 10183 16473 10195 16507
rect 10137 16467 10195 16473
rect 10321 16507 10379 16513
rect 10321 16473 10333 16507
rect 10367 16504 10379 16507
rect 11698 16504 11704 16516
rect 10367 16476 11704 16504
rect 10367 16473 10379 16476
rect 10321 16467 10379 16473
rect 11698 16464 11704 16476
rect 11756 16464 11762 16516
rect 11808 16504 11836 16544
rect 11974 16532 11980 16584
rect 12032 16572 12038 16584
rect 12032 16544 12756 16572
rect 12032 16532 12038 16544
rect 12728 16504 12756 16544
rect 12802 16532 12808 16584
rect 12860 16532 12866 16584
rect 12986 16532 12992 16584
rect 13044 16532 13050 16584
rect 13446 16532 13452 16584
rect 13504 16532 13510 16584
rect 14366 16532 14372 16584
rect 14424 16572 14430 16584
rect 14737 16575 14795 16581
rect 14737 16572 14749 16575
rect 14424 16544 14749 16572
rect 14424 16532 14430 16544
rect 14737 16541 14749 16544
rect 14783 16541 14795 16575
rect 15102 16572 15108 16584
rect 14737 16535 14795 16541
rect 14936 16544 15108 16572
rect 13633 16507 13691 16513
rect 13633 16504 13645 16507
rect 11808 16476 12572 16504
rect 12728 16476 13645 16504
rect 4706 16436 4712 16448
rect 4192 16408 4712 16436
rect 4706 16396 4712 16408
rect 4764 16396 4770 16448
rect 4798 16396 4804 16448
rect 4856 16436 4862 16448
rect 4893 16439 4951 16445
rect 4893 16436 4905 16439
rect 4856 16408 4905 16436
rect 4856 16396 4862 16408
rect 4893 16405 4905 16408
rect 4939 16405 4951 16439
rect 4893 16399 4951 16405
rect 5905 16439 5963 16445
rect 5905 16405 5917 16439
rect 5951 16436 5963 16439
rect 6086 16436 6092 16448
rect 5951 16408 6092 16436
rect 5951 16405 5963 16408
rect 5905 16399 5963 16405
rect 6086 16396 6092 16408
rect 6144 16396 6150 16448
rect 9490 16396 9496 16448
rect 9548 16396 9554 16448
rect 9677 16439 9735 16445
rect 9677 16405 9689 16439
rect 9723 16436 9735 16439
rect 9858 16436 9864 16448
rect 9723 16408 9864 16436
rect 9723 16405 9735 16408
rect 9677 16399 9735 16405
rect 9858 16396 9864 16408
rect 9916 16396 9922 16448
rect 11146 16396 11152 16448
rect 11204 16436 11210 16448
rect 12434 16436 12440 16448
rect 11204 16408 12440 16436
rect 11204 16396 11210 16408
rect 12434 16396 12440 16408
rect 12492 16396 12498 16448
rect 12544 16436 12572 16476
rect 13633 16473 13645 16476
rect 13679 16504 13691 16507
rect 14936 16504 14964 16544
rect 15102 16532 15108 16544
rect 15160 16532 15166 16584
rect 15194 16532 15200 16584
rect 15252 16532 15258 16584
rect 15764 16581 15792 16680
rect 16942 16668 16948 16680
rect 17000 16708 17006 16720
rect 17144 16708 17172 16739
rect 17862 16736 17868 16788
rect 17920 16776 17926 16788
rect 17957 16779 18015 16785
rect 17957 16776 17969 16779
rect 17920 16748 17969 16776
rect 17920 16736 17926 16748
rect 17957 16745 17969 16748
rect 18003 16745 18015 16779
rect 17957 16739 18015 16745
rect 18693 16779 18751 16785
rect 18693 16745 18705 16779
rect 18739 16776 18751 16779
rect 18782 16776 18788 16788
rect 18739 16748 18788 16776
rect 18739 16745 18751 16748
rect 18693 16739 18751 16745
rect 18782 16736 18788 16748
rect 18840 16736 18846 16788
rect 20349 16779 20407 16785
rect 20349 16745 20361 16779
rect 20395 16745 20407 16779
rect 20349 16739 20407 16745
rect 17000 16680 17172 16708
rect 17236 16680 18552 16708
rect 17000 16668 17006 16680
rect 16022 16600 16028 16652
rect 16080 16640 16086 16652
rect 16080 16612 16528 16640
rect 16080 16600 16086 16612
rect 15381 16575 15439 16581
rect 15381 16541 15393 16575
rect 15427 16572 15439 16575
rect 15749 16575 15807 16581
rect 15749 16572 15761 16575
rect 15427 16544 15761 16572
rect 15427 16541 15439 16544
rect 15381 16535 15439 16541
rect 15749 16541 15761 16544
rect 15795 16541 15807 16575
rect 15749 16535 15807 16541
rect 13679 16476 14964 16504
rect 13679 16473 13691 16476
rect 13633 16467 13691 16473
rect 15010 16464 15016 16516
rect 15068 16464 15074 16516
rect 15470 16464 15476 16516
rect 15528 16464 15534 16516
rect 16209 16507 16267 16513
rect 16209 16473 16221 16507
rect 16255 16504 16267 16507
rect 16298 16504 16304 16516
rect 16255 16476 16304 16504
rect 16255 16473 16267 16476
rect 16209 16467 16267 16473
rect 16298 16464 16304 16476
rect 16356 16464 16362 16516
rect 16390 16464 16396 16516
rect 16448 16464 16454 16516
rect 16500 16504 16528 16612
rect 16574 16600 16580 16652
rect 16632 16640 16638 16652
rect 16761 16643 16819 16649
rect 16761 16640 16773 16643
rect 16632 16612 16773 16640
rect 16632 16600 16638 16612
rect 16761 16609 16773 16612
rect 16807 16609 16819 16643
rect 17236 16640 17264 16680
rect 16761 16603 16819 16609
rect 16868 16612 17264 16640
rect 16666 16532 16672 16584
rect 16724 16532 16730 16584
rect 16868 16504 16896 16612
rect 17310 16600 17316 16652
rect 17368 16600 17374 16652
rect 18414 16640 18420 16652
rect 18064 16612 18420 16640
rect 18064 16584 18092 16612
rect 18414 16600 18420 16612
rect 18472 16600 18478 16652
rect 18524 16649 18552 16680
rect 20254 16668 20260 16720
rect 20312 16668 20318 16720
rect 18509 16643 18567 16649
rect 18509 16609 18521 16643
rect 18555 16609 18567 16643
rect 18509 16603 18567 16609
rect 20165 16643 20223 16649
rect 20165 16609 20177 16643
rect 20211 16640 20223 16643
rect 20272 16640 20300 16668
rect 20211 16612 20300 16640
rect 20364 16640 20392 16739
rect 22278 16736 22284 16788
rect 22336 16776 22342 16788
rect 23842 16776 23848 16788
rect 22336 16748 23848 16776
rect 22336 16736 22342 16748
rect 23842 16736 23848 16748
rect 23900 16736 23906 16788
rect 25406 16736 25412 16788
rect 25464 16736 25470 16788
rect 25685 16779 25743 16785
rect 25685 16745 25697 16779
rect 25731 16776 25743 16779
rect 25774 16776 25780 16788
rect 25731 16748 25780 16776
rect 25731 16745 25743 16748
rect 25685 16739 25743 16745
rect 25774 16736 25780 16748
rect 25832 16736 25838 16788
rect 27154 16736 27160 16788
rect 27212 16736 27218 16788
rect 28074 16736 28080 16788
rect 28132 16736 28138 16788
rect 28353 16779 28411 16785
rect 28353 16745 28365 16779
rect 28399 16776 28411 16779
rect 28534 16776 28540 16788
rect 28399 16748 28540 16776
rect 28399 16745 28411 16748
rect 28353 16739 28411 16745
rect 28534 16736 28540 16748
rect 28592 16736 28598 16788
rect 28718 16736 28724 16788
rect 28776 16736 28782 16788
rect 28997 16779 29055 16785
rect 28997 16745 29009 16779
rect 29043 16776 29055 16779
rect 29362 16776 29368 16788
rect 29043 16748 29368 16776
rect 29043 16745 29055 16748
rect 28997 16739 29055 16745
rect 21634 16668 21640 16720
rect 21692 16708 21698 16720
rect 24486 16708 24492 16720
rect 21692 16680 24492 16708
rect 21692 16668 21698 16680
rect 24486 16668 24492 16680
rect 24544 16668 24550 16720
rect 27172 16708 27200 16736
rect 25516 16680 27200 16708
rect 22462 16640 22468 16652
rect 20364 16612 22468 16640
rect 20211 16609 20223 16612
rect 20165 16603 20223 16609
rect 22462 16600 22468 16612
rect 22520 16640 22526 16652
rect 23382 16640 23388 16652
rect 22520 16612 23388 16640
rect 22520 16600 22526 16612
rect 23382 16600 23388 16612
rect 23440 16600 23446 16652
rect 23658 16600 23664 16652
rect 23716 16640 23722 16652
rect 25317 16643 25375 16649
rect 25317 16640 25329 16643
rect 23716 16612 25329 16640
rect 23716 16600 23722 16612
rect 25317 16609 25329 16612
rect 25363 16609 25375 16643
rect 25317 16603 25375 16609
rect 17405 16575 17463 16581
rect 17405 16541 17417 16575
rect 17451 16572 17463 16575
rect 17494 16572 17500 16584
rect 17451 16544 17500 16572
rect 17451 16541 17463 16544
rect 17405 16535 17463 16541
rect 17494 16532 17500 16544
rect 17552 16532 17558 16584
rect 17954 16532 17960 16584
rect 18012 16532 18018 16584
rect 18046 16532 18052 16584
rect 18104 16532 18110 16584
rect 18340 16544 18644 16572
rect 16500 16476 16896 16504
rect 16945 16507 17003 16513
rect 16945 16473 16957 16507
rect 16991 16473 17003 16507
rect 16945 16467 17003 16473
rect 12894 16436 12900 16448
rect 12544 16408 12900 16436
rect 12894 16396 12900 16408
rect 12952 16396 12958 16448
rect 13173 16439 13231 16445
rect 13173 16405 13185 16439
rect 13219 16436 13231 16439
rect 15654 16436 15660 16448
rect 13219 16408 15660 16436
rect 13219 16405 13231 16408
rect 13173 16399 13231 16405
rect 15654 16396 15660 16408
rect 15712 16396 15718 16448
rect 15930 16396 15936 16448
rect 15988 16396 15994 16448
rect 16960 16436 16988 16467
rect 17126 16464 17132 16516
rect 17184 16464 17190 16516
rect 18340 16504 18368 16544
rect 17604 16476 18368 16504
rect 17494 16436 17500 16448
rect 16960 16408 17500 16436
rect 17494 16396 17500 16408
rect 17552 16396 17558 16448
rect 17604 16445 17632 16476
rect 18414 16464 18420 16516
rect 18472 16464 18478 16516
rect 18616 16504 18644 16544
rect 18690 16532 18696 16584
rect 18748 16532 18754 16584
rect 20073 16575 20131 16581
rect 20073 16541 20085 16575
rect 20119 16572 20131 16575
rect 20990 16572 20996 16584
rect 20119 16544 20996 16572
rect 20119 16541 20131 16544
rect 20073 16535 20131 16541
rect 20990 16532 20996 16544
rect 21048 16532 21054 16584
rect 23566 16532 23572 16584
rect 23624 16572 23630 16584
rect 25516 16581 25544 16680
rect 27614 16668 27620 16720
rect 27672 16708 27678 16720
rect 29012 16708 29040 16739
rect 29362 16736 29368 16748
rect 29420 16736 29426 16788
rect 31570 16736 31576 16788
rect 31628 16736 31634 16788
rect 27672 16680 29040 16708
rect 27672 16668 27678 16680
rect 26878 16600 26884 16652
rect 26936 16640 26942 16652
rect 27154 16640 27160 16652
rect 26936 16612 27160 16640
rect 26936 16600 26942 16612
rect 27154 16600 27160 16612
rect 27212 16600 27218 16652
rect 27522 16600 27528 16652
rect 27580 16640 27586 16652
rect 27798 16640 27804 16652
rect 27580 16612 27804 16640
rect 27580 16600 27586 16612
rect 27798 16600 27804 16612
rect 27856 16640 27862 16652
rect 27985 16643 28043 16649
rect 27985 16640 27997 16643
rect 27856 16612 27997 16640
rect 27856 16600 27862 16612
rect 27985 16609 27997 16612
rect 28031 16609 28043 16643
rect 27985 16603 28043 16609
rect 28074 16600 28080 16652
rect 28132 16640 28138 16652
rect 28721 16643 28779 16649
rect 28721 16640 28733 16643
rect 28132 16612 28733 16640
rect 28132 16600 28138 16612
rect 28721 16609 28733 16612
rect 28767 16609 28779 16643
rect 28721 16603 28779 16609
rect 28902 16600 28908 16652
rect 28960 16640 28966 16652
rect 29089 16643 29147 16649
rect 29089 16640 29101 16643
rect 28960 16612 29101 16640
rect 28960 16600 28966 16612
rect 29089 16609 29101 16612
rect 29135 16609 29147 16643
rect 29089 16603 29147 16609
rect 32306 16600 32312 16652
rect 32364 16600 32370 16652
rect 25501 16575 25559 16581
rect 25501 16572 25513 16575
rect 23624 16544 25513 16572
rect 23624 16532 23630 16544
rect 25501 16541 25513 16544
rect 25547 16541 25559 16575
rect 25501 16535 25559 16541
rect 26694 16532 26700 16584
rect 26752 16572 26758 16584
rect 27893 16575 27951 16581
rect 27893 16572 27905 16575
rect 26752 16544 27905 16572
rect 26752 16532 26758 16544
rect 27893 16541 27905 16544
rect 27939 16541 27951 16575
rect 27893 16535 27951 16541
rect 28169 16575 28227 16581
rect 28169 16541 28181 16575
rect 28215 16541 28227 16575
rect 28169 16535 28227 16541
rect 20349 16507 20407 16513
rect 18616 16476 20300 16504
rect 17589 16439 17647 16445
rect 17589 16405 17601 16439
rect 17635 16405 17647 16439
rect 17589 16399 17647 16405
rect 18322 16396 18328 16448
rect 18380 16396 18386 16448
rect 18874 16396 18880 16448
rect 18932 16396 18938 16448
rect 19889 16439 19947 16445
rect 19889 16405 19901 16439
rect 19935 16436 19947 16439
rect 19978 16436 19984 16448
rect 19935 16408 19984 16436
rect 19935 16405 19947 16408
rect 19889 16399 19947 16405
rect 19978 16396 19984 16408
rect 20036 16396 20042 16448
rect 20272 16436 20300 16476
rect 20349 16473 20361 16507
rect 20395 16504 20407 16507
rect 20530 16504 20536 16516
rect 20395 16476 20536 16504
rect 20395 16473 20407 16476
rect 20349 16467 20407 16473
rect 20530 16464 20536 16476
rect 20588 16464 20594 16516
rect 22278 16464 22284 16516
rect 22336 16504 22342 16516
rect 24854 16504 24860 16516
rect 22336 16476 24860 16504
rect 22336 16464 22342 16476
rect 24854 16464 24860 16476
rect 24912 16464 24918 16516
rect 25130 16464 25136 16516
rect 25188 16504 25194 16516
rect 25225 16507 25283 16513
rect 25225 16504 25237 16507
rect 25188 16476 25237 16504
rect 25188 16464 25194 16476
rect 25225 16473 25237 16476
rect 25271 16504 25283 16507
rect 25406 16504 25412 16516
rect 25271 16476 25412 16504
rect 25271 16473 25283 16476
rect 25225 16467 25283 16473
rect 25406 16464 25412 16476
rect 25464 16464 25470 16516
rect 28184 16436 28212 16535
rect 28258 16532 28264 16584
rect 28316 16572 28322 16584
rect 28813 16575 28871 16581
rect 28813 16572 28825 16575
rect 28316 16544 28825 16572
rect 28316 16532 28322 16544
rect 28813 16541 28825 16544
rect 28859 16541 28871 16575
rect 28813 16535 28871 16541
rect 28997 16575 29055 16581
rect 28997 16541 29009 16575
rect 29043 16541 29055 16575
rect 28997 16535 29055 16541
rect 29012 16504 29040 16535
rect 30282 16532 30288 16584
rect 30340 16572 30346 16584
rect 31021 16575 31079 16581
rect 31021 16572 31033 16575
rect 30340 16544 31033 16572
rect 30340 16532 30346 16544
rect 31021 16541 31033 16544
rect 31067 16541 31079 16575
rect 31021 16535 31079 16541
rect 31389 16575 31447 16581
rect 31389 16541 31401 16575
rect 31435 16572 31447 16575
rect 31757 16575 31815 16581
rect 31757 16572 31769 16575
rect 31435 16544 31769 16572
rect 31435 16541 31447 16544
rect 31389 16535 31447 16541
rect 31757 16541 31769 16544
rect 31803 16541 31815 16575
rect 31757 16535 31815 16541
rect 29454 16504 29460 16516
rect 29012 16476 29460 16504
rect 29454 16464 29460 16476
rect 29512 16464 29518 16516
rect 30926 16464 30932 16516
rect 30984 16504 30990 16516
rect 31205 16507 31263 16513
rect 31205 16504 31217 16507
rect 30984 16476 31217 16504
rect 30984 16464 30990 16476
rect 31205 16473 31217 16476
rect 31251 16473 31263 16507
rect 31205 16467 31263 16473
rect 31297 16507 31355 16513
rect 31297 16473 31309 16507
rect 31343 16473 31355 16507
rect 31297 16467 31355 16473
rect 28258 16436 28264 16448
rect 20272 16408 28264 16436
rect 28258 16396 28264 16408
rect 28316 16396 28322 16448
rect 28445 16439 28503 16445
rect 28445 16405 28457 16439
rect 28491 16436 28503 16439
rect 28626 16436 28632 16448
rect 28491 16408 28632 16436
rect 28491 16405 28503 16408
rect 28445 16399 28503 16405
rect 28626 16396 28632 16408
rect 28684 16396 28690 16448
rect 29362 16396 29368 16448
rect 29420 16396 29426 16448
rect 30374 16396 30380 16448
rect 30432 16436 30438 16448
rect 31312 16436 31340 16467
rect 30432 16408 31340 16436
rect 30432 16396 30438 16408
rect 1104 16346 32844 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 32844 16346
rect 1104 16272 32844 16294
rect 2958 16232 2964 16244
rect 2884 16204 2964 16232
rect 2884 16173 2912 16204
rect 2958 16192 2964 16204
rect 3016 16192 3022 16244
rect 4157 16235 4215 16241
rect 4157 16201 4169 16235
rect 4203 16232 4215 16235
rect 4430 16232 4436 16244
rect 4203 16204 4436 16232
rect 4203 16201 4215 16204
rect 4157 16195 4215 16201
rect 4430 16192 4436 16204
rect 4488 16192 4494 16244
rect 4522 16192 4528 16244
rect 4580 16232 4586 16244
rect 7006 16232 7012 16244
rect 4580 16204 7012 16232
rect 4580 16192 4586 16204
rect 7006 16192 7012 16204
rect 7064 16192 7070 16244
rect 9122 16192 9128 16244
rect 9180 16232 9186 16244
rect 9858 16232 9864 16244
rect 9180 16204 9864 16232
rect 9180 16192 9186 16204
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 10134 16192 10140 16244
rect 10192 16232 10198 16244
rect 10505 16235 10563 16241
rect 10505 16232 10517 16235
rect 10192 16204 10517 16232
rect 10192 16192 10198 16204
rect 10505 16201 10517 16204
rect 10551 16201 10563 16235
rect 10505 16195 10563 16201
rect 12452 16204 12664 16232
rect 2869 16167 2927 16173
rect 2869 16133 2881 16167
rect 2915 16133 2927 16167
rect 2869 16127 2927 16133
rect 2976 16136 5304 16164
rect 2976 16108 3004 16136
rect 2593 16099 2651 16105
rect 2593 16065 2605 16099
rect 2639 16096 2651 16099
rect 2682 16096 2688 16108
rect 2639 16068 2688 16096
rect 2639 16065 2651 16068
rect 2593 16059 2651 16065
rect 2682 16056 2688 16068
rect 2740 16056 2746 16108
rect 2777 16099 2835 16105
rect 2777 16065 2789 16099
rect 2823 16065 2835 16099
rect 2777 16059 2835 16065
rect 2792 16028 2820 16059
rect 2958 16056 2964 16108
rect 3016 16056 3022 16108
rect 4338 16056 4344 16108
rect 4396 16056 4402 16108
rect 4525 16099 4583 16105
rect 4525 16065 4537 16099
rect 4571 16096 4583 16099
rect 5166 16096 5172 16108
rect 4571 16068 5172 16096
rect 4571 16065 4583 16068
rect 4525 16059 4583 16065
rect 5166 16056 5172 16068
rect 5224 16056 5230 16108
rect 5276 16096 5304 16136
rect 5810 16124 5816 16176
rect 5868 16164 5874 16176
rect 5997 16167 6055 16173
rect 5997 16164 6009 16167
rect 5868 16136 6009 16164
rect 5868 16124 5874 16136
rect 5997 16133 6009 16136
rect 6043 16133 6055 16167
rect 5997 16127 6055 16133
rect 6641 16167 6699 16173
rect 6641 16133 6653 16167
rect 6687 16164 6699 16167
rect 6914 16164 6920 16176
rect 6687 16136 6920 16164
rect 6687 16133 6699 16136
rect 6641 16127 6699 16133
rect 6914 16124 6920 16136
rect 6972 16124 6978 16176
rect 8478 16124 8484 16176
rect 8536 16124 8542 16176
rect 9490 16124 9496 16176
rect 9548 16164 9554 16176
rect 12452 16164 12480 16204
rect 9548 16136 12480 16164
rect 9548 16124 9554 16136
rect 12526 16124 12532 16176
rect 12584 16124 12590 16176
rect 12636 16164 12664 16204
rect 12802 16192 12808 16244
rect 12860 16232 12866 16244
rect 12989 16235 13047 16241
rect 12989 16232 13001 16235
rect 12860 16204 13001 16232
rect 12860 16192 12866 16204
rect 12989 16201 13001 16204
rect 13035 16201 13047 16235
rect 12989 16195 13047 16201
rect 13078 16192 13084 16244
rect 13136 16232 13142 16244
rect 16666 16232 16672 16244
rect 13136 16204 16672 16232
rect 13136 16192 13142 16204
rect 16666 16192 16672 16204
rect 16724 16192 16730 16244
rect 19334 16232 19340 16244
rect 16776 16204 19340 16232
rect 14274 16164 14280 16176
rect 12636 16136 14280 16164
rect 14274 16124 14280 16136
rect 14332 16124 14338 16176
rect 14476 16136 15700 16164
rect 6178 16096 6184 16108
rect 5276 16068 6184 16096
rect 6178 16056 6184 16068
rect 6236 16056 6242 16108
rect 6730 16056 6736 16108
rect 6788 16096 6794 16108
rect 6825 16099 6883 16105
rect 6825 16096 6837 16099
rect 6788 16068 6837 16096
rect 6788 16056 6794 16068
rect 6825 16065 6837 16068
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 3142 16028 3148 16040
rect 2792 16000 3148 16028
rect 3142 15988 3148 16000
rect 3200 16028 3206 16040
rect 5902 16028 5908 16040
rect 3200 16000 5908 16028
rect 3200 15988 3206 16000
rect 5902 15988 5908 16000
rect 5960 15988 5966 16040
rect 6840 16028 6868 16059
rect 7006 16056 7012 16108
rect 7064 16056 7070 16108
rect 8662 16056 8668 16108
rect 8720 16056 8726 16108
rect 8846 16056 8852 16108
rect 8904 16096 8910 16108
rect 9030 16096 9036 16108
rect 8904 16068 9036 16096
rect 8904 16056 8910 16068
rect 9030 16056 9036 16068
rect 9088 16056 9094 16108
rect 10689 16099 10747 16105
rect 10689 16065 10701 16099
rect 10735 16065 10747 16099
rect 10689 16059 10747 16065
rect 7193 16031 7251 16037
rect 7193 16028 7205 16031
rect 6840 16000 7205 16028
rect 7193 15997 7205 16000
rect 7239 15997 7251 16031
rect 10704 16028 10732 16059
rect 10778 16056 10784 16108
rect 10836 16056 10842 16108
rect 10962 16056 10968 16108
rect 11020 16056 11026 16108
rect 11241 16099 11299 16105
rect 11241 16065 11253 16099
rect 11287 16096 11299 16099
rect 12158 16096 12164 16108
rect 11287 16068 12164 16096
rect 11287 16065 11299 16068
rect 11241 16059 11299 16065
rect 12158 16056 12164 16068
rect 12216 16056 12222 16108
rect 12802 16056 12808 16108
rect 12860 16096 12866 16108
rect 14476 16096 14504 16136
rect 12860 16068 14504 16096
rect 12860 16056 12866 16068
rect 15010 16056 15016 16108
rect 15068 16096 15074 16108
rect 15278 16099 15336 16105
rect 15278 16096 15290 16099
rect 15068 16068 15290 16096
rect 15068 16056 15074 16068
rect 15278 16065 15290 16068
rect 15324 16065 15336 16099
rect 15278 16059 15336 16065
rect 15378 16056 15384 16108
rect 15436 16096 15442 16108
rect 15473 16099 15531 16105
rect 15473 16096 15485 16099
rect 15436 16068 15485 16096
rect 15436 16056 15442 16068
rect 15473 16065 15485 16068
rect 15519 16065 15531 16099
rect 15473 16059 15531 16065
rect 15565 16099 15623 16105
rect 15565 16065 15577 16099
rect 15611 16065 15623 16099
rect 15672 16096 15700 16136
rect 16390 16124 16396 16176
rect 16448 16164 16454 16176
rect 16776 16164 16804 16204
rect 19334 16192 19340 16204
rect 19392 16192 19398 16244
rect 20441 16235 20499 16241
rect 20441 16201 20453 16235
rect 20487 16232 20499 16235
rect 20487 16204 23428 16232
rect 20487 16201 20499 16204
rect 20441 16195 20499 16201
rect 16448 16136 16804 16164
rect 16448 16124 16454 16136
rect 16942 16124 16948 16176
rect 17000 16164 17006 16176
rect 19150 16164 19156 16176
rect 17000 16136 19156 16164
rect 17000 16124 17006 16136
rect 19150 16124 19156 16136
rect 19208 16124 19214 16176
rect 19702 16124 19708 16176
rect 19760 16164 19766 16176
rect 19797 16167 19855 16173
rect 19797 16164 19809 16167
rect 19760 16136 19809 16164
rect 19760 16124 19766 16136
rect 19797 16133 19809 16136
rect 19843 16133 19855 16167
rect 19797 16127 19855 16133
rect 19978 16124 19984 16176
rect 20036 16124 20042 16176
rect 22830 16124 22836 16176
rect 22888 16124 22894 16176
rect 23400 16164 23428 16204
rect 23474 16192 23480 16244
rect 23532 16192 23538 16244
rect 25869 16235 25927 16241
rect 25869 16201 25881 16235
rect 25915 16232 25927 16235
rect 27522 16232 27528 16244
rect 25915 16204 27528 16232
rect 25915 16201 25927 16204
rect 25869 16195 25927 16201
rect 27522 16192 27528 16204
rect 27580 16192 27586 16244
rect 30190 16192 30196 16244
rect 30248 16192 30254 16244
rect 30558 16192 30564 16244
rect 30616 16232 30622 16244
rect 31754 16232 31760 16244
rect 30616 16204 31760 16232
rect 30616 16192 30622 16204
rect 31754 16192 31760 16204
rect 31812 16192 31818 16244
rect 23400 16136 30236 16164
rect 30208 16108 30236 16136
rect 30742 16124 30748 16176
rect 30800 16164 30806 16176
rect 30929 16167 30987 16173
rect 30929 16164 30941 16167
rect 30800 16136 30941 16164
rect 30800 16124 30806 16136
rect 30929 16133 30941 16136
rect 30975 16133 30987 16167
rect 30929 16127 30987 16133
rect 17678 16096 17684 16108
rect 15672 16068 17684 16096
rect 15565 16059 15623 16065
rect 11146 16028 11152 16040
rect 10704 16000 11152 16028
rect 7193 15991 7251 15997
rect 11146 15988 11152 16000
rect 11204 15988 11210 16040
rect 11606 15988 11612 16040
rect 11664 16028 11670 16040
rect 12618 16028 12624 16040
rect 11664 16000 12624 16028
rect 11664 15988 11670 16000
rect 12618 15988 12624 16000
rect 12676 15988 12682 16040
rect 12713 16031 12771 16037
rect 12713 15997 12725 16031
rect 12759 16028 12771 16031
rect 13170 16028 13176 16040
rect 12759 16000 13176 16028
rect 12759 15997 12771 16000
rect 12713 15991 12771 15997
rect 13170 15988 13176 16000
rect 13228 15988 13234 16040
rect 15580 16028 15608 16059
rect 17678 16056 17684 16068
rect 17736 16056 17742 16108
rect 18322 16056 18328 16108
rect 18380 16096 18386 16108
rect 20257 16099 20315 16105
rect 20257 16096 20269 16099
rect 18380 16068 20269 16096
rect 18380 16056 18386 16068
rect 20257 16065 20269 16068
rect 20303 16065 20315 16099
rect 20257 16059 20315 16065
rect 20530 16056 20536 16108
rect 20588 16056 20594 16108
rect 20714 16056 20720 16108
rect 20772 16056 20778 16108
rect 20809 16099 20867 16105
rect 20809 16065 20821 16099
rect 20855 16096 20867 16099
rect 20898 16096 20904 16108
rect 20855 16068 20904 16096
rect 20855 16065 20867 16068
rect 20809 16059 20867 16065
rect 20898 16056 20904 16068
rect 20956 16056 20962 16108
rect 23109 16099 23167 16105
rect 23109 16065 23121 16099
rect 23155 16065 23167 16099
rect 23109 16059 23167 16065
rect 23569 16099 23627 16105
rect 23569 16065 23581 16099
rect 23615 16096 23627 16099
rect 24302 16096 24308 16108
rect 23615 16068 24308 16096
rect 23615 16065 23627 16068
rect 23569 16059 23627 16065
rect 15396 16000 15608 16028
rect 1118 15920 1124 15972
rect 1176 15960 1182 15972
rect 1176 15932 4660 15960
rect 1176 15920 1182 15932
rect 3145 15895 3203 15901
rect 3145 15861 3157 15895
rect 3191 15892 3203 15895
rect 3602 15892 3608 15904
rect 3191 15864 3608 15892
rect 3191 15861 3203 15864
rect 3145 15855 3203 15861
rect 3602 15852 3608 15864
rect 3660 15852 3666 15904
rect 4632 15892 4660 15932
rect 4706 15920 4712 15972
rect 4764 15920 4770 15972
rect 5994 15920 6000 15972
rect 6052 15960 6058 15972
rect 6270 15960 6276 15972
rect 6052 15932 6276 15960
rect 6052 15920 6058 15932
rect 6270 15920 6276 15932
rect 6328 15920 6334 15972
rect 6457 15963 6515 15969
rect 6457 15929 6469 15963
rect 6503 15960 6515 15963
rect 8294 15960 8300 15972
rect 6503 15932 8300 15960
rect 6503 15929 6515 15932
rect 6457 15923 6515 15929
rect 8294 15920 8300 15932
rect 8352 15920 8358 15972
rect 12434 15960 12440 15972
rect 8404 15932 12440 15960
rect 5810 15892 5816 15904
rect 4632 15864 5816 15892
rect 5810 15852 5816 15864
rect 5868 15892 5874 15904
rect 6089 15895 6147 15901
rect 6089 15892 6101 15895
rect 5868 15864 6101 15892
rect 5868 15852 5874 15864
rect 6089 15861 6101 15864
rect 6135 15861 6147 15895
rect 6089 15855 6147 15861
rect 6178 15852 6184 15904
rect 6236 15892 6242 15904
rect 8404 15892 8432 15932
rect 12434 15920 12440 15932
rect 12492 15920 12498 15972
rect 12894 15920 12900 15972
rect 12952 15960 12958 15972
rect 13998 15960 14004 15972
rect 12952 15932 14004 15960
rect 12952 15920 12958 15932
rect 13998 15920 14004 15932
rect 14056 15920 14062 15972
rect 15396 15960 15424 16000
rect 16298 15988 16304 16040
rect 16356 16028 16362 16040
rect 18782 16028 18788 16040
rect 16356 16000 18788 16028
rect 16356 15988 16362 16000
rect 18782 15988 18788 16000
rect 18840 15988 18846 16040
rect 19702 15988 19708 16040
rect 19760 16028 19766 16040
rect 20073 16031 20131 16037
rect 20073 16028 20085 16031
rect 19760 16000 20085 16028
rect 19760 15988 19766 16000
rect 20073 15997 20085 16000
rect 20119 15997 20131 16031
rect 20073 15991 20131 15997
rect 22922 15988 22928 16040
rect 22980 15988 22986 16040
rect 15304 15932 15424 15960
rect 6236 15864 8432 15892
rect 6236 15852 6242 15864
rect 8846 15852 8852 15904
rect 8904 15892 8910 15904
rect 10318 15892 10324 15904
rect 8904 15864 10324 15892
rect 8904 15852 8910 15864
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 10686 15852 10692 15904
rect 10744 15852 10750 15904
rect 11146 15852 11152 15904
rect 11204 15852 11210 15904
rect 11790 15852 11796 15904
rect 11848 15892 11854 15904
rect 12529 15895 12587 15901
rect 12529 15892 12541 15895
rect 11848 15864 12541 15892
rect 11848 15852 11854 15864
rect 12529 15861 12541 15864
rect 12575 15861 12587 15895
rect 12529 15855 12587 15861
rect 13906 15852 13912 15904
rect 13964 15892 13970 15904
rect 15304 15892 15332 15932
rect 15746 15920 15752 15972
rect 15804 15920 15810 15972
rect 15930 15920 15936 15972
rect 15988 15960 15994 15972
rect 23124 15960 23152 16059
rect 24302 16056 24308 16068
rect 24360 16096 24366 16108
rect 24360 16068 24808 16096
rect 24360 16056 24366 16068
rect 23382 15988 23388 16040
rect 23440 16028 23446 16040
rect 23661 16031 23719 16037
rect 23661 16028 23673 16031
rect 23440 16000 23673 16028
rect 23440 15988 23446 16000
rect 23661 15997 23673 16000
rect 23707 15997 23719 16031
rect 23661 15991 23719 15997
rect 15988 15932 23152 15960
rect 24780 15960 24808 16068
rect 24854 16056 24860 16108
rect 24912 16096 24918 16108
rect 25501 16099 25559 16105
rect 25501 16096 25513 16099
rect 24912 16068 25513 16096
rect 24912 16056 24918 16068
rect 25501 16065 25513 16068
rect 25547 16065 25559 16099
rect 25501 16059 25559 16065
rect 25685 16099 25743 16105
rect 25685 16065 25697 16099
rect 25731 16096 25743 16099
rect 25774 16096 25780 16108
rect 25731 16068 25780 16096
rect 25731 16065 25743 16068
rect 25685 16059 25743 16065
rect 25774 16056 25780 16068
rect 25832 16056 25838 16108
rect 26418 16056 26424 16108
rect 26476 16056 26482 16108
rect 29638 16056 29644 16108
rect 29696 16096 29702 16108
rect 29733 16099 29791 16105
rect 29733 16096 29745 16099
rect 29696 16068 29745 16096
rect 29696 16056 29702 16068
rect 29733 16065 29745 16068
rect 29779 16065 29791 16099
rect 29733 16059 29791 16065
rect 30006 16056 30012 16108
rect 30064 16056 30070 16108
rect 30190 16056 30196 16108
rect 30248 16056 30254 16108
rect 30558 16056 30564 16108
rect 30616 16056 30622 16108
rect 30653 16099 30711 16105
rect 30653 16065 30665 16099
rect 30699 16065 30711 16099
rect 30653 16059 30711 16065
rect 26326 15988 26332 16040
rect 26384 16028 26390 16040
rect 26513 16031 26571 16037
rect 26513 16028 26525 16031
rect 26384 16000 26525 16028
rect 26384 15988 26390 16000
rect 26513 15997 26525 16000
rect 26559 15997 26571 16031
rect 29270 16028 29276 16040
rect 26513 15991 26571 15997
rect 26620 16000 29276 16028
rect 26620 15960 26648 16000
rect 29270 15988 29276 16000
rect 29328 15988 29334 16040
rect 29822 15988 29828 16040
rect 29880 15988 29886 16040
rect 24780 15932 26648 15960
rect 15988 15920 15994 15932
rect 26786 15920 26792 15972
rect 26844 15920 26850 15972
rect 30558 15920 30564 15972
rect 30616 15960 30622 15972
rect 30668 15960 30696 16059
rect 30834 16056 30840 16108
rect 30892 16056 30898 16108
rect 31021 16099 31079 16105
rect 31021 16065 31033 16099
rect 31067 16096 31079 16099
rect 31297 16099 31355 16105
rect 31297 16096 31309 16099
rect 31067 16068 31309 16096
rect 31067 16065 31079 16068
rect 31021 16059 31079 16065
rect 31297 16065 31309 16068
rect 31343 16065 31355 16099
rect 31297 16059 31355 16065
rect 31941 16099 31999 16105
rect 31941 16065 31953 16099
rect 31987 16096 31999 16099
rect 32214 16096 32220 16108
rect 31987 16068 32220 16096
rect 31987 16065 31999 16068
rect 31941 16059 31999 16065
rect 32214 16056 32220 16068
rect 32272 16056 32278 16108
rect 30616 15932 30696 15960
rect 30616 15920 30622 15932
rect 13964 15864 15332 15892
rect 15565 15895 15623 15901
rect 13964 15852 13970 15864
rect 15565 15861 15577 15895
rect 15611 15892 15623 15895
rect 17034 15892 17040 15904
rect 15611 15864 17040 15892
rect 15611 15861 15623 15864
rect 15565 15855 15623 15861
rect 17034 15852 17040 15864
rect 17092 15852 17098 15904
rect 18138 15852 18144 15904
rect 18196 15892 18202 15904
rect 18690 15892 18696 15904
rect 18196 15864 18696 15892
rect 18196 15852 18202 15864
rect 18690 15852 18696 15864
rect 18748 15852 18754 15904
rect 19886 15852 19892 15904
rect 19944 15892 19950 15904
rect 19981 15895 20039 15901
rect 19981 15892 19993 15895
rect 19944 15864 19993 15892
rect 19944 15852 19950 15864
rect 19981 15861 19993 15864
rect 20027 15861 20039 15895
rect 19981 15855 20039 15861
rect 20438 15852 20444 15904
rect 20496 15892 20502 15904
rect 20533 15895 20591 15901
rect 20533 15892 20545 15895
rect 20496 15864 20545 15892
rect 20496 15852 20502 15864
rect 20533 15861 20545 15864
rect 20579 15861 20591 15895
rect 20533 15855 20591 15861
rect 20993 15895 21051 15901
rect 20993 15861 21005 15895
rect 21039 15892 21051 15895
rect 21174 15892 21180 15904
rect 21039 15864 21180 15892
rect 21039 15861 21051 15864
rect 20993 15855 21051 15861
rect 21174 15852 21180 15864
rect 21232 15852 21238 15904
rect 21266 15852 21272 15904
rect 21324 15892 21330 15904
rect 21910 15892 21916 15904
rect 21324 15864 21916 15892
rect 21324 15852 21330 15864
rect 21910 15852 21916 15864
rect 21968 15852 21974 15904
rect 22462 15852 22468 15904
rect 22520 15892 22526 15904
rect 22833 15895 22891 15901
rect 22833 15892 22845 15895
rect 22520 15864 22845 15892
rect 22520 15852 22526 15864
rect 22833 15861 22845 15864
rect 22879 15861 22891 15895
rect 22833 15855 22891 15861
rect 23290 15852 23296 15904
rect 23348 15852 23354 15904
rect 23474 15852 23480 15904
rect 23532 15892 23538 15904
rect 23569 15895 23627 15901
rect 23569 15892 23581 15895
rect 23532 15864 23581 15892
rect 23532 15852 23538 15864
rect 23569 15861 23581 15864
rect 23615 15861 23627 15895
rect 23569 15855 23627 15861
rect 23842 15852 23848 15904
rect 23900 15892 23906 15904
rect 23937 15895 23995 15901
rect 23937 15892 23949 15895
rect 23900 15864 23949 15892
rect 23900 15852 23906 15864
rect 23937 15861 23949 15864
rect 23983 15861 23995 15895
rect 23937 15855 23995 15861
rect 25498 15852 25504 15904
rect 25556 15852 25562 15904
rect 26329 15895 26387 15901
rect 26329 15861 26341 15895
rect 26375 15892 26387 15895
rect 26421 15895 26479 15901
rect 26421 15892 26433 15895
rect 26375 15864 26433 15892
rect 26375 15861 26387 15864
rect 26329 15855 26387 15861
rect 26421 15861 26433 15864
rect 26467 15892 26479 15895
rect 26694 15892 26700 15904
rect 26467 15864 26700 15892
rect 26467 15861 26479 15864
rect 26421 15855 26479 15861
rect 26694 15852 26700 15864
rect 26752 15852 26758 15904
rect 29454 15852 29460 15904
rect 29512 15892 29518 15904
rect 29733 15895 29791 15901
rect 29733 15892 29745 15895
rect 29512 15864 29745 15892
rect 29512 15852 29518 15864
rect 29733 15861 29745 15864
rect 29779 15861 29791 15895
rect 29733 15855 29791 15861
rect 30377 15895 30435 15901
rect 30377 15861 30389 15895
rect 30423 15892 30435 15895
rect 30466 15892 30472 15904
rect 30423 15864 30472 15892
rect 30423 15861 30435 15864
rect 30377 15855 30435 15861
rect 30466 15852 30472 15864
rect 30524 15852 30530 15904
rect 31202 15852 31208 15904
rect 31260 15852 31266 15904
rect 32398 15852 32404 15904
rect 32456 15852 32462 15904
rect 1104 15802 32844 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 32844 15802
rect 1104 15728 32844 15750
rect 3878 15688 3884 15700
rect 3436 15660 3884 15688
rect 3436 15493 3464 15660
rect 3878 15648 3884 15660
rect 3936 15688 3942 15700
rect 3973 15691 4031 15697
rect 3973 15688 3985 15691
rect 3936 15660 3985 15688
rect 3936 15648 3942 15660
rect 3973 15657 3985 15660
rect 4019 15657 4031 15691
rect 3973 15651 4031 15657
rect 5445 15691 5503 15697
rect 5445 15657 5457 15691
rect 5491 15688 5503 15691
rect 5534 15688 5540 15700
rect 5491 15660 5540 15688
rect 5491 15657 5503 15660
rect 5445 15651 5503 15657
rect 5534 15648 5540 15660
rect 5592 15688 5598 15700
rect 5994 15688 6000 15700
rect 5592 15660 6000 15688
rect 5592 15648 5598 15660
rect 5994 15648 6000 15660
rect 6052 15648 6058 15700
rect 6270 15648 6276 15700
rect 6328 15688 6334 15700
rect 6328 15660 6684 15688
rect 6328 15648 6334 15660
rect 6546 15580 6552 15632
rect 6604 15580 6610 15632
rect 6656 15620 6684 15660
rect 6730 15648 6736 15700
rect 6788 15688 6794 15700
rect 7834 15688 7840 15700
rect 6788 15660 7840 15688
rect 6788 15648 6794 15660
rect 7834 15648 7840 15660
rect 7892 15648 7898 15700
rect 12802 15688 12808 15700
rect 7944 15660 12808 15688
rect 7944 15620 7972 15660
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 13725 15691 13783 15697
rect 13725 15657 13737 15691
rect 13771 15688 13783 15691
rect 14918 15688 14924 15700
rect 13771 15660 14924 15688
rect 13771 15657 13783 15660
rect 13725 15651 13783 15657
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 15013 15691 15071 15697
rect 15013 15657 15025 15691
rect 15059 15688 15071 15691
rect 15102 15688 15108 15700
rect 15059 15660 15108 15688
rect 15059 15657 15071 15660
rect 15013 15651 15071 15657
rect 15102 15648 15108 15660
rect 15160 15648 15166 15700
rect 15194 15648 15200 15700
rect 15252 15648 15258 15700
rect 15286 15648 15292 15700
rect 15344 15688 15350 15700
rect 16393 15691 16451 15697
rect 16393 15688 16405 15691
rect 15344 15660 16405 15688
rect 15344 15648 15350 15660
rect 16393 15657 16405 15660
rect 16439 15657 16451 15691
rect 16393 15651 16451 15657
rect 16758 15648 16764 15700
rect 16816 15648 16822 15700
rect 18138 15648 18144 15700
rect 18196 15688 18202 15700
rect 18506 15688 18512 15700
rect 18196 15660 18512 15688
rect 18196 15648 18202 15660
rect 18506 15648 18512 15660
rect 18564 15688 18570 15700
rect 20438 15688 20444 15700
rect 18564 15660 20444 15688
rect 18564 15648 18570 15660
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 21818 15648 21824 15700
rect 21876 15688 21882 15700
rect 21913 15691 21971 15697
rect 21913 15688 21925 15691
rect 21876 15660 21925 15688
rect 21876 15648 21882 15660
rect 21913 15657 21925 15660
rect 21959 15657 21971 15691
rect 21913 15651 21971 15657
rect 22373 15691 22431 15697
rect 22373 15657 22385 15691
rect 22419 15688 22431 15691
rect 22462 15688 22468 15700
rect 22419 15660 22468 15688
rect 22419 15657 22431 15660
rect 22373 15651 22431 15657
rect 22462 15648 22468 15660
rect 22520 15648 22526 15700
rect 23014 15648 23020 15700
rect 23072 15648 23078 15700
rect 27249 15691 27307 15697
rect 27249 15657 27261 15691
rect 27295 15688 27307 15691
rect 27522 15688 27528 15700
rect 27295 15660 27528 15688
rect 27295 15657 27307 15660
rect 27249 15651 27307 15657
rect 27522 15648 27528 15660
rect 27580 15648 27586 15700
rect 29454 15648 29460 15700
rect 29512 15688 29518 15700
rect 29641 15691 29699 15697
rect 29641 15688 29653 15691
rect 29512 15660 29653 15688
rect 29512 15648 29518 15660
rect 29641 15657 29653 15660
rect 29687 15657 29699 15691
rect 29641 15651 29699 15657
rect 30190 15648 30196 15700
rect 30248 15648 30254 15700
rect 30558 15648 30564 15700
rect 30616 15648 30622 15700
rect 32214 15648 32220 15700
rect 32272 15688 32278 15700
rect 32493 15691 32551 15697
rect 32493 15688 32505 15691
rect 32272 15660 32505 15688
rect 32272 15648 32278 15660
rect 32493 15657 32505 15660
rect 32539 15657 32551 15691
rect 32493 15651 32551 15657
rect 6656 15592 7972 15620
rect 9122 15580 9128 15632
rect 9180 15620 9186 15632
rect 9306 15620 9312 15632
rect 9180 15592 9312 15620
rect 9180 15580 9186 15592
rect 9306 15580 9312 15592
rect 9364 15620 9370 15632
rect 9585 15623 9643 15629
rect 9585 15620 9597 15623
rect 9364 15592 9597 15620
rect 9364 15580 9370 15592
rect 9585 15589 9597 15592
rect 9631 15589 9643 15623
rect 9585 15583 9643 15589
rect 10226 15580 10232 15632
rect 10284 15580 10290 15632
rect 10410 15580 10416 15632
rect 10468 15620 10474 15632
rect 10597 15623 10655 15629
rect 10597 15620 10609 15623
rect 10468 15592 10609 15620
rect 10468 15580 10474 15592
rect 10597 15589 10609 15592
rect 10643 15589 10655 15623
rect 15378 15620 15384 15632
rect 10597 15583 10655 15589
rect 11440 15592 15384 15620
rect 3786 15512 3792 15564
rect 3844 15552 3850 15564
rect 4341 15555 4399 15561
rect 4341 15552 4353 15555
rect 3844 15524 4353 15552
rect 3844 15512 3850 15524
rect 4341 15521 4353 15524
rect 4387 15552 4399 15555
rect 6178 15552 6184 15564
rect 4387 15524 6184 15552
rect 4387 15521 4399 15524
rect 4341 15515 4399 15521
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 6564 15552 6592 15580
rect 6564 15524 6684 15552
rect 3421 15487 3479 15493
rect 3421 15453 3433 15487
rect 3467 15453 3479 15487
rect 3421 15447 3479 15453
rect 3878 15444 3884 15496
rect 3936 15444 3942 15496
rect 4522 15444 4528 15496
rect 4580 15484 4586 15496
rect 4617 15487 4675 15493
rect 4617 15484 4629 15487
rect 4580 15456 4629 15484
rect 4580 15444 4586 15456
rect 4617 15453 4629 15456
rect 4663 15453 4675 15487
rect 4617 15447 4675 15453
rect 5258 15444 5264 15496
rect 5316 15444 5322 15496
rect 5626 15444 5632 15496
rect 5684 15484 5690 15496
rect 6273 15487 6331 15493
rect 6273 15484 6285 15487
rect 5684 15456 6285 15484
rect 5684 15444 5690 15456
rect 6273 15453 6285 15456
rect 6319 15453 6331 15487
rect 6273 15447 6331 15453
rect 6546 15444 6552 15496
rect 6604 15444 6610 15496
rect 6656 15493 6684 15524
rect 7650 15512 7656 15564
rect 7708 15552 7714 15564
rect 10502 15552 10508 15564
rect 7708 15524 10508 15552
rect 7708 15512 7714 15524
rect 10502 15512 10508 15524
rect 10560 15552 10566 15564
rect 10560 15524 10916 15552
rect 10560 15512 10566 15524
rect 6641 15487 6699 15493
rect 6641 15453 6653 15487
rect 6687 15453 6699 15487
rect 6641 15447 6699 15453
rect 6730 15444 6736 15496
rect 6788 15484 6794 15496
rect 6825 15487 6883 15493
rect 6825 15484 6837 15487
rect 6788 15456 6837 15484
rect 6788 15444 6794 15456
rect 6825 15453 6837 15456
rect 6871 15453 6883 15487
rect 6825 15447 6883 15453
rect 6917 15487 6975 15493
rect 6917 15453 6929 15487
rect 6963 15484 6975 15487
rect 8294 15484 8300 15496
rect 6963 15456 8300 15484
rect 6963 15453 6975 15456
rect 6917 15447 6975 15453
rect 8294 15444 8300 15456
rect 8352 15444 8358 15496
rect 9766 15444 9772 15496
rect 9824 15444 9830 15496
rect 10042 15444 10048 15496
rect 10100 15444 10106 15496
rect 10413 15487 10471 15493
rect 10413 15453 10425 15487
rect 10459 15484 10471 15487
rect 10594 15484 10600 15496
rect 10459 15456 10600 15484
rect 10459 15453 10471 15456
rect 10413 15447 10471 15453
rect 10594 15444 10600 15456
rect 10652 15444 10658 15496
rect 10778 15444 10784 15496
rect 10836 15444 10842 15496
rect 10888 15493 10916 15524
rect 10873 15487 10931 15493
rect 10873 15453 10885 15487
rect 10919 15453 10931 15487
rect 10873 15447 10931 15453
rect 2498 15376 2504 15428
rect 2556 15416 2562 15428
rect 7374 15416 7380 15428
rect 2556 15388 7380 15416
rect 2556 15376 2562 15388
rect 7374 15376 7380 15388
rect 7432 15376 7438 15428
rect 7466 15376 7472 15428
rect 7524 15416 7530 15428
rect 11440 15416 11468 15592
rect 15378 15580 15384 15592
rect 15436 15580 15442 15632
rect 15473 15623 15531 15629
rect 15473 15589 15485 15623
rect 15519 15620 15531 15623
rect 16206 15620 16212 15632
rect 15519 15592 16212 15620
rect 15519 15589 15531 15592
rect 15473 15583 15531 15589
rect 12342 15512 12348 15564
rect 12400 15552 12406 15564
rect 13906 15552 13912 15564
rect 12400 15524 13912 15552
rect 12400 15512 12406 15524
rect 13906 15512 13912 15524
rect 13964 15512 13970 15564
rect 13998 15512 14004 15564
rect 14056 15552 14062 15564
rect 14829 15555 14887 15561
rect 14829 15552 14841 15555
rect 14056 15524 14841 15552
rect 14056 15512 14062 15524
rect 14829 15521 14841 15524
rect 14875 15552 14887 15555
rect 15488 15552 15516 15583
rect 16206 15580 16212 15592
rect 16264 15580 16270 15632
rect 18874 15580 18880 15632
rect 18932 15620 18938 15632
rect 21634 15620 21640 15632
rect 18932 15592 21640 15620
rect 18932 15580 18938 15592
rect 21634 15580 21640 15592
rect 21692 15580 21698 15632
rect 22278 15620 22284 15632
rect 22066 15592 22284 15620
rect 14875 15524 15516 15552
rect 14875 15521 14887 15524
rect 14829 15515 14887 15521
rect 15654 15512 15660 15564
rect 15712 15552 15718 15564
rect 16485 15555 16543 15561
rect 16485 15552 16497 15555
rect 15712 15524 16497 15552
rect 15712 15512 15718 15524
rect 16485 15521 16497 15524
rect 16531 15521 16543 15555
rect 16485 15515 16543 15521
rect 17954 15512 17960 15564
rect 18012 15552 18018 15564
rect 22066 15552 22094 15592
rect 22278 15580 22284 15592
rect 22336 15580 22342 15632
rect 27433 15623 27491 15629
rect 27433 15589 27445 15623
rect 27479 15620 27491 15623
rect 30101 15623 30159 15629
rect 27479 15592 30052 15620
rect 27479 15589 27491 15592
rect 27433 15583 27491 15589
rect 18012 15524 22094 15552
rect 18012 15512 18018 15524
rect 22186 15512 22192 15564
rect 22244 15512 22250 15564
rect 22922 15512 22928 15564
rect 22980 15512 22986 15564
rect 23109 15555 23167 15561
rect 23109 15521 23121 15555
rect 23155 15552 23167 15555
rect 23566 15552 23572 15564
rect 23155 15524 23572 15552
rect 23155 15521 23167 15524
rect 23109 15515 23167 15521
rect 23566 15512 23572 15524
rect 23624 15512 23630 15564
rect 27062 15512 27068 15564
rect 27120 15512 27126 15564
rect 27172 15524 29776 15552
rect 12158 15444 12164 15496
rect 12216 15484 12222 15496
rect 12216 15456 12388 15484
rect 12216 15444 12222 15456
rect 7524 15388 11468 15416
rect 12360 15416 12388 15456
rect 12434 15444 12440 15496
rect 12492 15484 12498 15496
rect 12492 15456 14872 15484
rect 12492 15444 12498 15456
rect 12802 15416 12808 15428
rect 12360 15388 12808 15416
rect 7524 15376 7530 15388
rect 12802 15376 12808 15388
rect 12860 15376 12866 15428
rect 13078 15376 13084 15428
rect 13136 15416 13142 15428
rect 13357 15419 13415 15425
rect 13357 15416 13369 15419
rect 13136 15388 13369 15416
rect 13136 15376 13142 15388
rect 13357 15385 13369 15388
rect 13403 15385 13415 15419
rect 13357 15379 13415 15385
rect 13538 15376 13544 15428
rect 13596 15376 13602 15428
rect 14737 15419 14795 15425
rect 14737 15385 14749 15419
rect 14783 15385 14795 15419
rect 14844 15416 14872 15456
rect 15010 15444 15016 15496
rect 15068 15444 15074 15496
rect 15289 15487 15347 15493
rect 15289 15453 15301 15487
rect 15335 15453 15347 15487
rect 15289 15447 15347 15453
rect 15304 15416 15332 15447
rect 15378 15444 15384 15496
rect 15436 15484 15442 15496
rect 15565 15487 15623 15493
rect 15565 15484 15577 15487
rect 15436 15456 15577 15484
rect 15436 15444 15442 15456
rect 15565 15453 15577 15456
rect 15611 15453 15623 15487
rect 15565 15447 15623 15453
rect 16114 15444 16120 15496
rect 16172 15484 16178 15496
rect 16393 15487 16451 15493
rect 16393 15484 16405 15487
rect 16172 15456 16405 15484
rect 16172 15444 16178 15456
rect 16393 15453 16405 15456
rect 16439 15453 16451 15487
rect 16393 15447 16451 15453
rect 18782 15444 18788 15496
rect 18840 15484 18846 15496
rect 20438 15484 20444 15496
rect 18840 15456 20444 15484
rect 18840 15444 18846 15456
rect 20438 15444 20444 15456
rect 20496 15444 20502 15496
rect 22002 15444 22008 15496
rect 22060 15484 22066 15496
rect 22097 15487 22155 15493
rect 22097 15484 22109 15487
rect 22060 15456 22109 15484
rect 22060 15444 22066 15456
rect 22097 15453 22109 15456
rect 22143 15453 22155 15487
rect 22833 15487 22891 15493
rect 22833 15484 22845 15487
rect 22097 15447 22155 15453
rect 22197 15456 22845 15484
rect 14844 15388 15332 15416
rect 14737 15379 14795 15385
rect 3605 15351 3663 15357
rect 3605 15317 3617 15351
rect 3651 15348 3663 15351
rect 4062 15348 4068 15360
rect 3651 15320 4068 15348
rect 3651 15317 3663 15320
rect 3605 15311 3663 15317
rect 4062 15308 4068 15320
rect 4120 15308 4126 15360
rect 7101 15351 7159 15357
rect 7101 15317 7113 15351
rect 7147 15348 7159 15351
rect 8386 15348 8392 15360
rect 7147 15320 8392 15348
rect 7147 15317 7159 15320
rect 7101 15311 7159 15317
rect 8386 15308 8392 15320
rect 8444 15308 8450 15360
rect 8478 15308 8484 15360
rect 8536 15348 8542 15360
rect 9306 15348 9312 15360
rect 8536 15320 9312 15348
rect 8536 15308 8542 15320
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 9766 15308 9772 15360
rect 9824 15348 9830 15360
rect 9861 15351 9919 15357
rect 9861 15348 9873 15351
rect 9824 15320 9873 15348
rect 9824 15308 9830 15320
rect 9861 15317 9873 15320
rect 9907 15317 9919 15351
rect 9861 15311 9919 15317
rect 10318 15308 10324 15360
rect 10376 15348 10382 15360
rect 10778 15348 10784 15360
rect 10376 15320 10784 15348
rect 10376 15308 10382 15320
rect 10778 15308 10784 15320
rect 10836 15308 10842 15360
rect 10870 15308 10876 15360
rect 10928 15348 10934 15360
rect 11057 15351 11115 15357
rect 11057 15348 11069 15351
rect 10928 15320 11069 15348
rect 10928 15308 10934 15320
rect 11057 15317 11069 15320
rect 11103 15348 11115 15351
rect 14182 15348 14188 15360
rect 11103 15320 14188 15348
rect 11103 15317 11115 15320
rect 11057 15311 11115 15317
rect 14182 15308 14188 15320
rect 14240 15308 14246 15360
rect 14752 15348 14780 15379
rect 17218 15376 17224 15428
rect 17276 15416 17282 15428
rect 17276 15388 18644 15416
rect 17276 15376 17282 15388
rect 15749 15351 15807 15357
rect 15749 15348 15761 15351
rect 14752 15320 15761 15348
rect 15749 15317 15761 15320
rect 15795 15348 15807 15351
rect 15838 15348 15844 15360
rect 15795 15320 15844 15348
rect 15795 15317 15807 15320
rect 15749 15311 15807 15317
rect 15838 15308 15844 15320
rect 15896 15308 15902 15360
rect 18616 15348 18644 15388
rect 19334 15376 19340 15428
rect 19392 15416 19398 15428
rect 19610 15416 19616 15428
rect 19392 15388 19616 15416
rect 19392 15376 19398 15388
rect 19610 15376 19616 15388
rect 19668 15416 19674 15428
rect 19981 15419 20039 15425
rect 19981 15416 19993 15419
rect 19668 15388 19993 15416
rect 19668 15376 19674 15388
rect 19981 15385 19993 15388
rect 20027 15385 20039 15419
rect 19981 15379 20039 15385
rect 20165 15419 20223 15425
rect 20165 15385 20177 15419
rect 20211 15385 20223 15419
rect 20165 15379 20223 15385
rect 19702 15348 19708 15360
rect 18616 15320 19708 15348
rect 19702 15308 19708 15320
rect 19760 15348 19766 15360
rect 20180 15348 20208 15379
rect 21818 15376 21824 15428
rect 21876 15416 21882 15428
rect 22197 15416 22225 15456
rect 22833 15453 22845 15456
rect 22879 15484 22891 15487
rect 22940 15484 22968 15512
rect 22879 15456 22968 15484
rect 22879 15453 22891 15456
rect 22833 15447 22891 15453
rect 23198 15444 23204 15496
rect 23256 15484 23262 15496
rect 23293 15487 23351 15493
rect 23293 15484 23305 15487
rect 23256 15456 23305 15484
rect 23256 15444 23262 15456
rect 23293 15453 23305 15456
rect 23339 15453 23351 15487
rect 23293 15447 23351 15453
rect 24946 15444 24952 15496
rect 25004 15484 25010 15496
rect 25498 15484 25504 15496
rect 25004 15456 25504 15484
rect 25004 15444 25010 15456
rect 25498 15444 25504 15456
rect 25556 15444 25562 15496
rect 27172 15484 27200 15524
rect 25884 15456 27200 15484
rect 27249 15487 27307 15493
rect 21876 15388 22225 15416
rect 22373 15419 22431 15425
rect 21876 15376 21882 15388
rect 22373 15385 22385 15419
rect 22419 15416 22431 15419
rect 22462 15416 22468 15428
rect 22419 15388 22468 15416
rect 22419 15385 22431 15388
rect 22373 15379 22431 15385
rect 22462 15376 22468 15388
rect 22520 15376 22526 15428
rect 22646 15376 22652 15428
rect 22704 15376 22710 15428
rect 22922 15376 22928 15428
rect 22980 15416 22986 15428
rect 23017 15419 23075 15425
rect 23017 15416 23029 15419
rect 22980 15388 23029 15416
rect 22980 15376 22986 15388
rect 23017 15385 23029 15388
rect 23063 15385 23075 15419
rect 25317 15419 25375 15425
rect 25317 15416 25329 15419
rect 23017 15379 23075 15385
rect 23400 15388 25329 15416
rect 19760 15320 20208 15348
rect 19760 15308 19766 15320
rect 20254 15308 20260 15360
rect 20312 15348 20318 15360
rect 20349 15351 20407 15357
rect 20349 15348 20361 15351
rect 20312 15320 20361 15348
rect 20312 15308 20318 15320
rect 20349 15317 20361 15320
rect 20395 15348 20407 15351
rect 20530 15348 20536 15360
rect 20395 15320 20536 15348
rect 20395 15317 20407 15320
rect 20349 15311 20407 15317
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 20806 15308 20812 15360
rect 20864 15348 20870 15360
rect 23400 15348 23428 15388
rect 25317 15385 25329 15388
rect 25363 15385 25375 15419
rect 25317 15379 25375 15385
rect 25884 15360 25912 15456
rect 27249 15453 27261 15487
rect 27295 15484 27307 15487
rect 27338 15484 27344 15496
rect 27295 15456 27344 15484
rect 27295 15453 27307 15456
rect 27249 15447 27307 15453
rect 27338 15444 27344 15456
rect 27396 15444 27402 15496
rect 27522 15444 27528 15496
rect 27580 15484 27586 15496
rect 27893 15487 27951 15493
rect 27893 15484 27905 15487
rect 27580 15456 27905 15484
rect 27580 15444 27586 15456
rect 27893 15453 27905 15456
rect 27939 15453 27951 15487
rect 27893 15447 27951 15453
rect 28810 15444 28816 15496
rect 28868 15484 28874 15496
rect 29641 15487 29699 15493
rect 29641 15484 29653 15487
rect 28868 15456 29653 15484
rect 28868 15444 28874 15456
rect 29641 15453 29653 15456
rect 29687 15453 29699 15487
rect 29748 15484 29776 15524
rect 29822 15512 29828 15564
rect 29880 15512 29886 15564
rect 29917 15487 29975 15493
rect 29917 15484 29929 15487
rect 29748 15456 29929 15484
rect 29641 15447 29699 15453
rect 29917 15453 29929 15456
rect 29963 15453 29975 15487
rect 30024 15484 30052 15592
rect 30101 15589 30113 15623
rect 30147 15620 30159 15623
rect 30147 15592 30328 15620
rect 30147 15589 30159 15592
rect 30101 15583 30159 15589
rect 30300 15561 30328 15592
rect 30285 15555 30343 15561
rect 30285 15521 30297 15555
rect 30331 15521 30343 15555
rect 30285 15515 30343 15521
rect 30650 15512 30656 15564
rect 30708 15552 30714 15564
rect 31113 15555 31171 15561
rect 31113 15552 31125 15555
rect 30708 15524 31125 15552
rect 30708 15512 30714 15524
rect 31113 15521 31125 15524
rect 31159 15521 31171 15555
rect 31113 15515 31171 15521
rect 30193 15487 30251 15493
rect 30193 15484 30205 15487
rect 30024 15456 30205 15484
rect 29917 15447 29975 15453
rect 30193 15453 30205 15456
rect 30239 15453 30251 15487
rect 30193 15447 30251 15453
rect 26970 15376 26976 15428
rect 27028 15376 27034 15428
rect 27430 15376 27436 15428
rect 27488 15416 27494 15428
rect 28077 15419 28135 15425
rect 28077 15416 28089 15419
rect 27488 15388 28089 15416
rect 27488 15376 27494 15388
rect 28077 15385 28089 15388
rect 28123 15416 28135 15419
rect 28534 15416 28540 15428
rect 28123 15388 28540 15416
rect 28123 15385 28135 15388
rect 28077 15379 28135 15385
rect 28534 15376 28540 15388
rect 28592 15376 28598 15428
rect 29270 15376 29276 15428
rect 29328 15416 29334 15428
rect 29454 15416 29460 15428
rect 29328 15388 29460 15416
rect 29328 15376 29334 15388
rect 29454 15376 29460 15388
rect 29512 15416 29518 15428
rect 29730 15416 29736 15428
rect 29512 15388 29736 15416
rect 29512 15376 29518 15388
rect 29730 15376 29736 15388
rect 29788 15376 29794 15428
rect 29932 15416 29960 15447
rect 31202 15444 31208 15496
rect 31260 15484 31266 15496
rect 31369 15487 31427 15493
rect 31369 15484 31381 15487
rect 31260 15456 31381 15484
rect 31260 15444 31266 15456
rect 31369 15453 31381 15456
rect 31415 15453 31427 15487
rect 31369 15447 31427 15453
rect 30006 15416 30012 15428
rect 29932 15388 30012 15416
rect 30006 15376 30012 15388
rect 30064 15376 30070 15428
rect 20864 15320 23428 15348
rect 20864 15308 20870 15320
rect 23474 15308 23480 15360
rect 23532 15308 23538 15360
rect 25685 15351 25743 15357
rect 25685 15317 25697 15351
rect 25731 15348 25743 15351
rect 25866 15348 25872 15360
rect 25731 15320 25872 15348
rect 25731 15317 25743 15320
rect 25685 15311 25743 15317
rect 25866 15308 25872 15320
rect 25924 15308 25930 15360
rect 28166 15308 28172 15360
rect 28224 15348 28230 15360
rect 28261 15351 28319 15357
rect 28261 15348 28273 15351
rect 28224 15320 28273 15348
rect 28224 15308 28230 15320
rect 28261 15317 28273 15320
rect 28307 15348 28319 15351
rect 28442 15348 28448 15360
rect 28307 15320 28448 15348
rect 28307 15317 28319 15320
rect 28261 15311 28319 15317
rect 28442 15308 28448 15320
rect 28500 15308 28506 15360
rect 30558 15308 30564 15360
rect 30616 15348 30622 15360
rect 30926 15348 30932 15360
rect 30616 15320 30932 15348
rect 30616 15308 30622 15320
rect 30926 15308 30932 15320
rect 30984 15308 30990 15360
rect 1104 15258 32844 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 32844 15258
rect 1104 15184 32844 15206
rect 2869 15147 2927 15153
rect 2869 15113 2881 15147
rect 2915 15144 2927 15147
rect 3050 15144 3056 15156
rect 2915 15116 3056 15144
rect 2915 15113 2927 15116
rect 2869 15107 2927 15113
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 3878 15104 3884 15156
rect 3936 15144 3942 15156
rect 6730 15144 6736 15156
rect 3936 15116 6736 15144
rect 3936 15104 3942 15116
rect 6730 15104 6736 15116
rect 6788 15104 6794 15156
rect 7006 15104 7012 15156
rect 7064 15144 7070 15156
rect 8113 15147 8171 15153
rect 8113 15144 8125 15147
rect 7064 15116 8125 15144
rect 7064 15104 7070 15116
rect 8113 15113 8125 15116
rect 8159 15113 8171 15147
rect 8846 15144 8852 15156
rect 8113 15107 8171 15113
rect 8220 15116 8852 15144
rect 4706 15076 4712 15088
rect 4356 15048 4712 15076
rect 2222 14968 2228 15020
rect 2280 14968 2286 15020
rect 2406 14968 2412 15020
rect 2464 14968 2470 15020
rect 2685 15011 2743 15017
rect 2685 14977 2697 15011
rect 2731 14977 2743 15011
rect 2685 14971 2743 14977
rect 2700 14940 2728 14971
rect 2958 14968 2964 15020
rect 3016 14968 3022 15020
rect 3142 14968 3148 15020
rect 3200 14968 3206 15020
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 3697 15011 3755 15017
rect 3697 14977 3709 15011
rect 3743 15008 3755 15011
rect 3786 15008 3792 15020
rect 3743 14980 3792 15008
rect 3743 14977 3755 14980
rect 3697 14971 3755 14977
rect 3436 14940 3464 14971
rect 3786 14968 3792 14980
rect 3844 14968 3850 15020
rect 4356 15017 4384 15048
rect 4706 15036 4712 15048
rect 4764 15036 4770 15088
rect 5442 15076 5448 15088
rect 5184 15048 5448 15076
rect 4341 15011 4399 15017
rect 4341 14977 4353 15011
rect 4387 14977 4399 15011
rect 4341 14971 4399 14977
rect 4614 14968 4620 15020
rect 4672 14968 4678 15020
rect 4798 14968 4804 15020
rect 4856 15008 4862 15020
rect 5184 15017 5212 15048
rect 5442 15036 5448 15048
rect 5500 15036 5506 15088
rect 7374 15036 7380 15088
rect 7432 15076 7438 15088
rect 8220 15076 8248 15116
rect 8846 15104 8852 15116
rect 8904 15104 8910 15156
rect 9125 15147 9183 15153
rect 9125 15113 9137 15147
rect 9171 15144 9183 15147
rect 10597 15147 10655 15153
rect 9171 15116 10088 15144
rect 9171 15113 9183 15116
rect 9125 15107 9183 15113
rect 10060 15088 10088 15116
rect 10597 15113 10609 15147
rect 10643 15144 10655 15147
rect 10962 15144 10968 15156
rect 10643 15116 10968 15144
rect 10643 15113 10655 15116
rect 10597 15107 10655 15113
rect 10962 15104 10968 15116
rect 11020 15104 11026 15156
rect 12158 15104 12164 15156
rect 12216 15144 12222 15156
rect 12216 15116 14596 15144
rect 12216 15104 12222 15116
rect 7432 15048 8248 15076
rect 7432 15036 7438 15048
rect 8754 15036 8760 15088
rect 8812 15076 8818 15088
rect 8812 15048 9444 15076
rect 8812 15036 8818 15048
rect 4893 15011 4951 15017
rect 4893 15008 4905 15011
rect 4856 14980 4905 15008
rect 4856 14968 4862 14980
rect 4893 14977 4905 14980
rect 4939 14977 4951 15011
rect 4893 14971 4951 14977
rect 5169 15011 5227 15017
rect 5169 14977 5181 15011
rect 5215 14977 5227 15011
rect 7466 15008 7472 15020
rect 5169 14971 5227 14977
rect 5276 14980 7472 15008
rect 2700 14912 3464 14940
rect 3436 14872 3464 14912
rect 3970 14900 3976 14952
rect 4028 14900 4034 14952
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14940 4583 14943
rect 4706 14940 4712 14952
rect 4571 14912 4712 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 4706 14900 4712 14912
rect 4764 14900 4770 14952
rect 4982 14900 4988 14952
rect 5040 14940 5046 14952
rect 5276 14940 5304 14980
rect 7466 14968 7472 14980
rect 7524 14968 7530 15020
rect 7929 15011 7987 15017
rect 7929 14977 7941 15011
rect 7975 15008 7987 15011
rect 8110 15008 8116 15020
rect 7975 14980 8116 15008
rect 7975 14977 7987 14980
rect 7929 14971 7987 14977
rect 8110 14968 8116 14980
rect 8168 14968 8174 15020
rect 8294 14968 8300 15020
rect 8352 14968 8358 15020
rect 8386 14968 8392 15020
rect 8444 14968 8450 15020
rect 8478 14968 8484 15020
rect 8536 15008 8542 15020
rect 8573 15011 8631 15017
rect 8573 15008 8585 15011
rect 8536 14980 8585 15008
rect 8536 14968 8542 14980
rect 8573 14977 8585 14980
rect 8619 14977 8631 15011
rect 8573 14971 8631 14977
rect 8665 15011 8723 15017
rect 8665 14977 8677 15011
rect 8711 15008 8723 15011
rect 8846 15008 8852 15020
rect 8711 14980 8852 15008
rect 8711 14977 8723 14980
rect 8665 14971 8723 14977
rect 8846 14968 8852 14980
rect 8904 14968 8910 15020
rect 8941 15012 8999 15017
rect 9217 15014 9275 15017
rect 9306 15014 9312 15020
rect 8941 15011 9076 15012
rect 8941 14977 8953 15011
rect 8987 15008 9076 15011
rect 9217 15011 9312 15014
rect 8987 14984 9175 15008
rect 8987 14977 8999 14984
rect 9048 14980 9175 14984
rect 8941 14971 8999 14977
rect 5040 14912 5304 14940
rect 5445 14943 5503 14949
rect 5040 14900 5046 14912
rect 5445 14909 5457 14943
rect 5491 14940 5503 14943
rect 5534 14940 5540 14952
rect 5491 14912 5540 14940
rect 5491 14909 5503 14912
rect 5445 14903 5503 14909
rect 5534 14900 5540 14912
rect 5592 14940 5598 14952
rect 5718 14940 5724 14952
rect 5592 14912 5724 14940
rect 5592 14900 5598 14912
rect 5718 14900 5724 14912
rect 5776 14900 5782 14952
rect 6362 14900 6368 14952
rect 6420 14900 6426 14952
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14940 6699 14943
rect 7006 14940 7012 14952
rect 6687 14912 7012 14940
rect 6687 14909 6699 14912
rect 6641 14903 6699 14909
rect 7006 14900 7012 14912
rect 7064 14940 7070 14952
rect 8018 14940 8024 14952
rect 7064 14912 8024 14940
rect 7064 14900 7070 14912
rect 8018 14900 8024 14912
rect 8076 14900 8082 14952
rect 9147 14940 9175 14980
rect 9217 14977 9229 15011
rect 9263 14986 9312 15011
rect 9263 14977 9275 14986
rect 9217 14971 9275 14977
rect 9306 14968 9312 14986
rect 9364 14968 9370 15020
rect 9416 15017 9444 15048
rect 10042 15036 10048 15088
rect 10100 15036 10106 15088
rect 11238 15036 11244 15088
rect 11296 15076 11302 15088
rect 13538 15076 13544 15088
rect 11296 15048 13544 15076
rect 11296 15036 11302 15048
rect 13538 15036 13544 15048
rect 13596 15036 13602 15088
rect 14001 15079 14059 15085
rect 14001 15045 14013 15079
rect 14047 15076 14059 15079
rect 14090 15076 14096 15088
rect 14047 15048 14096 15076
rect 14047 15045 14059 15048
rect 14001 15039 14059 15045
rect 14090 15036 14096 15048
rect 14148 15076 14154 15088
rect 14366 15076 14372 15088
rect 14148 15048 14372 15076
rect 14148 15036 14154 15048
rect 14366 15036 14372 15048
rect 14424 15036 14430 15088
rect 9401 15011 9459 15017
rect 9401 14977 9413 15011
rect 9447 14977 9459 15011
rect 9401 14971 9459 14977
rect 9582 14968 9588 15020
rect 9640 15008 9646 15020
rect 9677 15011 9735 15017
rect 9677 15008 9689 15011
rect 9640 14980 9689 15008
rect 9640 14968 9646 14980
rect 9677 14977 9689 14980
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 10318 14968 10324 15020
rect 10376 14968 10382 15020
rect 10778 14968 10784 15020
rect 10836 14968 10842 15020
rect 10873 15011 10931 15017
rect 10873 14977 10885 15011
rect 10919 15008 10931 15011
rect 10962 15008 10968 15020
rect 10919 14980 10968 15008
rect 10919 14977 10931 14980
rect 10873 14971 10931 14977
rect 10962 14968 10968 14980
rect 11020 14968 11026 15020
rect 11057 15011 11115 15017
rect 11057 14977 11069 15011
rect 11103 15008 11115 15011
rect 11146 15008 11152 15020
rect 11103 14980 11152 15008
rect 11103 14977 11115 14980
rect 11057 14971 11115 14977
rect 11146 14968 11152 14980
rect 11204 15008 11210 15020
rect 11790 15008 11796 15020
rect 11204 14980 11796 15008
rect 11204 14968 11210 14980
rect 11790 14968 11796 14980
rect 11848 14968 11854 15020
rect 11882 14968 11888 15020
rect 11940 15008 11946 15020
rect 12069 15011 12127 15017
rect 12069 15008 12081 15011
rect 11940 14980 12081 15008
rect 11940 14968 11946 14980
rect 12069 14977 12081 14980
rect 12115 14977 12127 15011
rect 13722 15008 13728 15020
rect 12069 14971 12127 14977
rect 12360 14980 13728 15008
rect 10137 14943 10195 14949
rect 8128 14912 8892 14940
rect 9147 14912 9904 14940
rect 3988 14872 4016 14900
rect 8128 14872 8156 14912
rect 3436 14844 8156 14872
rect 8662 14832 8668 14884
rect 8720 14832 8726 14884
rect 8864 14872 8892 14912
rect 8864 14844 8984 14872
rect 3605 14807 3663 14813
rect 3605 14773 3617 14807
rect 3651 14804 3663 14807
rect 3786 14804 3792 14816
rect 3651 14776 3792 14804
rect 3651 14773 3663 14776
rect 3605 14767 3663 14773
rect 3786 14764 3792 14776
rect 3844 14764 3850 14816
rect 3970 14764 3976 14816
rect 4028 14804 4034 14816
rect 4157 14807 4215 14813
rect 4157 14804 4169 14807
rect 4028 14776 4169 14804
rect 4028 14764 4034 14776
rect 4157 14773 4169 14776
rect 4203 14773 4215 14807
rect 4157 14767 4215 14773
rect 4522 14764 4528 14816
rect 4580 14804 4586 14816
rect 4617 14807 4675 14813
rect 4617 14804 4629 14807
rect 4580 14776 4629 14804
rect 4580 14764 4586 14776
rect 4617 14773 4629 14776
rect 4663 14804 4675 14807
rect 4890 14804 4896 14816
rect 4663 14776 4896 14804
rect 4663 14773 4675 14776
rect 4617 14767 4675 14773
rect 4890 14764 4896 14776
rect 4948 14764 4954 14816
rect 5074 14764 5080 14816
rect 5132 14804 5138 14816
rect 7650 14804 7656 14816
rect 5132 14776 7656 14804
rect 5132 14764 5138 14776
rect 7650 14764 7656 14776
rect 7708 14764 7714 14816
rect 7742 14764 7748 14816
rect 7800 14804 7806 14816
rect 8018 14804 8024 14816
rect 7800 14776 8024 14804
rect 7800 14764 7806 14776
rect 8018 14764 8024 14776
rect 8076 14764 8082 14816
rect 8573 14807 8631 14813
rect 8573 14773 8585 14807
rect 8619 14804 8631 14807
rect 8680 14804 8708 14832
rect 8619 14776 8708 14804
rect 8619 14773 8631 14776
rect 8573 14767 8631 14773
rect 8846 14764 8852 14816
rect 8904 14764 8910 14816
rect 8956 14804 8984 14844
rect 9876 14816 9904 14912
rect 10137 14909 10149 14943
rect 10183 14940 10195 14943
rect 11977 14943 12035 14949
rect 10183 14912 11928 14940
rect 10183 14909 10195 14912
rect 10137 14903 10195 14909
rect 11054 14832 11060 14884
rect 11112 14872 11118 14884
rect 11900 14872 11928 14912
rect 11977 14909 11989 14943
rect 12023 14940 12035 14943
rect 12250 14940 12256 14952
rect 12023 14912 12256 14940
rect 12023 14909 12035 14912
rect 11977 14903 12035 14909
rect 12250 14900 12256 14912
rect 12308 14900 12314 14952
rect 12360 14872 12388 14980
rect 13722 14968 13728 14980
rect 13780 14968 13786 15020
rect 14274 14968 14280 15020
rect 14332 14968 14338 15020
rect 14568 15017 14596 15116
rect 15838 15104 15844 15156
rect 15896 15144 15902 15156
rect 16390 15144 16396 15156
rect 15896 15116 16396 15144
rect 15896 15104 15902 15116
rect 16390 15104 16396 15116
rect 16448 15104 16454 15156
rect 16758 15104 16764 15156
rect 16816 15144 16822 15156
rect 17770 15144 17776 15156
rect 16816 15116 17776 15144
rect 16816 15104 16822 15116
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 17957 15147 18015 15153
rect 17957 15113 17969 15147
rect 18003 15144 18015 15147
rect 20622 15144 20628 15156
rect 18003 15116 20628 15144
rect 18003 15113 18015 15116
rect 17957 15107 18015 15113
rect 17972 15076 18000 15107
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 22462 15104 22468 15156
rect 22520 15144 22526 15156
rect 22520 15116 23704 15144
rect 22520 15104 22526 15116
rect 17328 15048 18000 15076
rect 18064 15048 19840 15076
rect 17328 15017 17356 15048
rect 14553 15011 14611 15017
rect 14553 14977 14565 15011
rect 14599 14977 14611 15011
rect 14553 14971 14611 14977
rect 17313 15011 17371 15017
rect 17313 14977 17325 15011
rect 17359 14977 17371 15011
rect 17313 14971 17371 14977
rect 17405 15011 17463 15017
rect 17405 14977 17417 15011
rect 17451 15008 17463 15011
rect 17451 14980 17632 15008
rect 17451 14977 17463 14980
rect 17405 14971 17463 14977
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 13262 14940 13268 14952
rect 12492 14912 13268 14940
rect 12492 14900 12498 14912
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 14093 14943 14151 14949
rect 14093 14940 14105 14943
rect 13556 14912 14105 14940
rect 11112 14844 11744 14872
rect 11900 14844 12388 14872
rect 11112 14832 11118 14844
rect 9582 14804 9588 14816
rect 8956 14776 9588 14804
rect 9582 14764 9588 14776
rect 9640 14764 9646 14816
rect 9858 14764 9864 14816
rect 9916 14764 9922 14816
rect 10042 14764 10048 14816
rect 10100 14764 10106 14816
rect 10505 14807 10563 14813
rect 10505 14773 10517 14807
rect 10551 14804 10563 14807
rect 10686 14804 10692 14816
rect 10551 14776 10692 14804
rect 10551 14773 10563 14776
rect 10505 14767 10563 14773
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 10870 14764 10876 14816
rect 10928 14764 10934 14816
rect 11716 14813 11744 14844
rect 13170 14832 13176 14884
rect 13228 14872 13234 14884
rect 13446 14872 13452 14884
rect 13228 14844 13452 14872
rect 13228 14832 13234 14844
rect 13446 14832 13452 14844
rect 13504 14832 13510 14884
rect 13556 14816 13584 14912
rect 14093 14909 14105 14912
rect 14139 14909 14151 14943
rect 17126 14940 17132 14952
rect 14093 14903 14151 14909
rect 14200 14912 17132 14940
rect 13630 14832 13636 14884
rect 13688 14872 13694 14884
rect 14200 14872 14228 14912
rect 17126 14900 17132 14912
rect 17184 14900 17190 14952
rect 14918 14872 14924 14884
rect 13688 14844 14228 14872
rect 14292 14844 14924 14872
rect 13688 14832 13694 14844
rect 11701 14807 11759 14813
rect 11701 14773 11713 14807
rect 11747 14773 11759 14807
rect 11701 14767 11759 14773
rect 12066 14764 12072 14816
rect 12124 14764 12130 14816
rect 13262 14764 13268 14816
rect 13320 14804 13326 14816
rect 13538 14804 13544 14816
rect 13320 14776 13544 14804
rect 13320 14764 13326 14776
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 14292 14813 14320 14844
rect 14918 14832 14924 14844
rect 14976 14832 14982 14884
rect 17604 14872 17632 14980
rect 17678 14968 17684 15020
rect 17736 14968 17742 15020
rect 17770 14968 17776 15020
rect 17828 14968 17834 15020
rect 18064 14940 18092 15048
rect 18230 14968 18236 15020
rect 18288 15008 18294 15020
rect 18414 15008 18420 15020
rect 18288 14980 18420 15008
rect 18288 14968 18294 14980
rect 18414 14968 18420 14980
rect 18472 14968 18478 15020
rect 18874 14968 18880 15020
rect 18932 14968 18938 15020
rect 19337 15011 19395 15017
rect 19610 15012 19616 15020
rect 19337 14977 19349 15011
rect 19383 15008 19395 15011
rect 19536 15008 19616 15012
rect 19383 14984 19616 15008
rect 19383 14980 19564 14984
rect 19383 14977 19395 14980
rect 19337 14971 19395 14977
rect 19610 14968 19616 14984
rect 19668 14968 19674 15020
rect 19705 15011 19763 15017
rect 19705 14977 19717 15011
rect 19751 14998 19763 15011
rect 19812 14998 19840 15048
rect 20438 15036 20444 15088
rect 20496 15076 20502 15088
rect 20993 15079 21051 15085
rect 20496 15048 20760 15076
rect 20496 15036 20502 15048
rect 19751 14977 19840 14998
rect 20732 15008 20760 15048
rect 20993 15045 21005 15079
rect 21039 15076 21051 15079
rect 21634 15076 21640 15088
rect 21039 15048 21640 15076
rect 21039 15045 21051 15048
rect 20993 15039 21051 15045
rect 21634 15036 21640 15048
rect 21692 15036 21698 15088
rect 23382 15036 23388 15088
rect 23440 15036 23446 15088
rect 23676 15076 23704 15116
rect 23750 15104 23756 15156
rect 23808 15144 23814 15156
rect 23845 15147 23903 15153
rect 23845 15144 23857 15147
rect 23808 15116 23857 15144
rect 23808 15104 23814 15116
rect 23845 15113 23857 15116
rect 23891 15113 23903 15147
rect 23845 15107 23903 15113
rect 26050 15104 26056 15156
rect 26108 15104 26114 15156
rect 29546 15104 29552 15156
rect 29604 15144 29610 15156
rect 30190 15144 30196 15156
rect 29604 15116 30196 15144
rect 29604 15104 29610 15116
rect 30190 15104 30196 15116
rect 30248 15104 30254 15156
rect 32398 15104 32404 15156
rect 32456 15104 32462 15156
rect 27893 15079 27951 15085
rect 27893 15076 27905 15079
rect 23676 15048 27905 15076
rect 23768 15020 23796 15048
rect 27893 15045 27905 15048
rect 27939 15045 27951 15079
rect 27893 15039 27951 15045
rect 30374 15036 30380 15088
rect 30432 15076 30438 15088
rect 31202 15076 31208 15088
rect 30432 15048 31208 15076
rect 30432 15036 30438 15048
rect 31202 15036 31208 15048
rect 31260 15036 31266 15088
rect 21177 15011 21235 15017
rect 21177 15008 21189 15011
rect 20732 14980 21189 15008
rect 19705 14971 19840 14977
rect 21177 14977 21189 14980
rect 21223 14977 21235 15011
rect 21177 14971 21235 14977
rect 21361 15011 21419 15017
rect 21361 14977 21373 15011
rect 21407 15008 21419 15011
rect 22094 15008 22100 15020
rect 21407 14980 22100 15008
rect 21407 14977 21419 14980
rect 21361 14971 21419 14977
rect 19720 14970 19840 14971
rect 22094 14968 22100 14980
rect 22152 15008 22158 15020
rect 23566 15008 23572 15020
rect 22152 14980 23572 15008
rect 22152 14968 22158 14980
rect 23566 14968 23572 14980
rect 23624 14968 23630 15020
rect 23658 14968 23664 15020
rect 23716 14968 23722 15020
rect 23750 14968 23756 15020
rect 23808 14968 23814 15020
rect 24670 14968 24676 15020
rect 24728 15008 24734 15020
rect 25685 15011 25743 15017
rect 25685 15008 25697 15011
rect 24728 14980 25697 15008
rect 24728 14968 24734 14980
rect 25685 14977 25697 14980
rect 25731 14977 25743 15011
rect 25685 14971 25743 14977
rect 28074 14968 28080 15020
rect 28132 14968 28138 15020
rect 30561 15011 30619 15017
rect 30561 14977 30573 15011
rect 30607 15008 30619 15011
rect 30834 15008 30840 15020
rect 30607 14980 30840 15008
rect 30607 14977 30619 14980
rect 30561 14971 30619 14977
rect 30834 14968 30840 14980
rect 30892 14968 30898 15020
rect 31018 14968 31024 15020
rect 31076 15008 31082 15020
rect 31389 15011 31447 15017
rect 31389 15008 31401 15011
rect 31076 14980 31401 15008
rect 31076 14968 31082 14980
rect 31389 14977 31401 14980
rect 31435 14977 31447 15011
rect 31389 14971 31447 14977
rect 32214 14968 32220 15020
rect 32272 14968 32278 15020
rect 17696 14912 18092 14940
rect 18509 14943 18567 14949
rect 17696 14884 17724 14912
rect 18509 14909 18521 14943
rect 18555 14909 18567 14943
rect 22922 14940 22928 14952
rect 18509 14903 18567 14909
rect 19076 14912 22928 14940
rect 16080 14844 17632 14872
rect 13909 14807 13967 14813
rect 13909 14773 13921 14807
rect 13955 14804 13967 14807
rect 14277 14807 14335 14813
rect 14277 14804 14289 14807
rect 13955 14776 14289 14804
rect 13955 14773 13967 14776
rect 13909 14767 13967 14773
rect 14277 14773 14289 14776
rect 14323 14773 14335 14807
rect 14277 14767 14335 14773
rect 14461 14807 14519 14813
rect 14461 14773 14473 14807
rect 14507 14804 14519 14807
rect 14642 14804 14648 14816
rect 14507 14776 14648 14804
rect 14507 14773 14519 14776
rect 14461 14767 14519 14773
rect 14642 14764 14648 14776
rect 14700 14764 14706 14816
rect 14737 14807 14795 14813
rect 14737 14773 14749 14807
rect 14783 14804 14795 14807
rect 15286 14804 15292 14816
rect 14783 14776 15292 14804
rect 14783 14773 14795 14776
rect 14737 14767 14795 14773
rect 15286 14764 15292 14776
rect 15344 14804 15350 14816
rect 16080 14804 16108 14844
rect 15344 14776 16108 14804
rect 15344 14764 15350 14776
rect 16206 14764 16212 14816
rect 16264 14804 16270 14816
rect 16666 14804 16672 14816
rect 16264 14776 16672 14804
rect 16264 14764 16270 14776
rect 16666 14764 16672 14776
rect 16724 14804 16730 14816
rect 16942 14804 16948 14816
rect 16724 14776 16948 14804
rect 16724 14764 16730 14776
rect 16942 14764 16948 14776
rect 17000 14764 17006 14816
rect 17034 14764 17040 14816
rect 17092 14764 17098 14816
rect 17126 14764 17132 14816
rect 17184 14804 17190 14816
rect 17405 14807 17463 14813
rect 17405 14804 17417 14807
rect 17184 14776 17417 14804
rect 17184 14764 17190 14776
rect 17405 14773 17417 14776
rect 17451 14804 17463 14807
rect 17497 14807 17555 14813
rect 17497 14804 17509 14807
rect 17451 14776 17509 14804
rect 17451 14773 17463 14776
rect 17405 14767 17463 14773
rect 17497 14773 17509 14776
rect 17543 14773 17555 14807
rect 17604 14804 17632 14844
rect 17678 14832 17684 14884
rect 17736 14832 17742 14884
rect 17770 14832 17776 14884
rect 17828 14872 17834 14884
rect 18524 14872 18552 14903
rect 17828 14844 18552 14872
rect 17828 14832 17834 14844
rect 18782 14832 18788 14884
rect 18840 14832 18846 14884
rect 18874 14832 18880 14884
rect 18932 14872 18938 14884
rect 19076 14881 19104 14912
rect 22922 14900 22928 14912
rect 22980 14900 22986 14952
rect 23290 14900 23296 14952
rect 23348 14940 23354 14952
rect 23477 14943 23535 14949
rect 23477 14940 23489 14943
rect 23348 14912 23489 14940
rect 23348 14900 23354 14912
rect 23477 14909 23489 14912
rect 23523 14909 23535 14943
rect 23477 14903 23535 14909
rect 24946 14900 24952 14952
rect 25004 14940 25010 14952
rect 25777 14943 25835 14949
rect 25777 14940 25789 14943
rect 25004 14912 25789 14940
rect 25004 14900 25010 14912
rect 25777 14909 25789 14912
rect 25823 14940 25835 14943
rect 26050 14940 26056 14952
rect 25823 14912 26056 14940
rect 25823 14909 25835 14912
rect 25777 14903 25835 14909
rect 26050 14900 26056 14912
rect 26108 14900 26114 14952
rect 30374 14900 30380 14952
rect 30432 14940 30438 14952
rect 31113 14943 31171 14949
rect 31113 14940 31125 14943
rect 30432 14912 31125 14940
rect 30432 14900 30438 14912
rect 31113 14909 31125 14912
rect 31159 14909 31171 14943
rect 31113 14903 31171 14909
rect 19061 14875 19119 14881
rect 19061 14872 19073 14875
rect 18932 14844 19073 14872
rect 18932 14832 18938 14844
rect 19061 14841 19073 14844
rect 19107 14841 19119 14875
rect 19061 14835 19119 14841
rect 19150 14832 19156 14884
rect 19208 14832 19214 14884
rect 24670 14872 24676 14884
rect 19306 14844 24676 14872
rect 18414 14804 18420 14816
rect 17604 14776 18420 14804
rect 17497 14767 17555 14773
rect 18414 14764 18420 14776
rect 18472 14764 18478 14816
rect 18506 14764 18512 14816
rect 18564 14804 18570 14816
rect 19306 14804 19334 14844
rect 24670 14832 24676 14844
rect 24728 14832 24734 14884
rect 30745 14875 30803 14881
rect 30745 14841 30757 14875
rect 30791 14872 30803 14875
rect 30791 14844 31432 14872
rect 30791 14841 30803 14844
rect 30745 14835 30803 14841
rect 31404 14816 31432 14844
rect 18564 14776 19334 14804
rect 18564 14764 18570 14776
rect 19610 14764 19616 14816
rect 19668 14804 19674 14816
rect 19889 14807 19947 14813
rect 19889 14804 19901 14807
rect 19668 14776 19901 14804
rect 19668 14764 19674 14776
rect 19889 14773 19901 14776
rect 19935 14804 19947 14807
rect 20070 14804 20076 14816
rect 19935 14776 20076 14804
rect 19935 14773 19947 14776
rect 19889 14767 19947 14773
rect 20070 14764 20076 14776
rect 20128 14764 20134 14816
rect 21266 14764 21272 14816
rect 21324 14804 21330 14816
rect 23198 14804 23204 14816
rect 21324 14776 23204 14804
rect 21324 14764 21330 14776
rect 23198 14764 23204 14776
rect 23256 14764 23262 14816
rect 23661 14807 23719 14813
rect 23661 14773 23673 14807
rect 23707 14804 23719 14807
rect 23842 14804 23848 14816
rect 23707 14776 23848 14804
rect 23707 14773 23719 14776
rect 23661 14767 23719 14773
rect 23842 14764 23848 14776
rect 23900 14764 23906 14816
rect 24486 14764 24492 14816
rect 24544 14804 24550 14816
rect 24854 14804 24860 14816
rect 24544 14776 24860 14804
rect 24544 14764 24550 14776
rect 24854 14764 24860 14776
rect 24912 14764 24918 14816
rect 25590 14764 25596 14816
rect 25648 14804 25654 14816
rect 25685 14807 25743 14813
rect 25685 14804 25697 14807
rect 25648 14776 25697 14804
rect 25648 14764 25654 14776
rect 25685 14773 25697 14776
rect 25731 14773 25743 14807
rect 25685 14767 25743 14773
rect 28261 14807 28319 14813
rect 28261 14773 28273 14807
rect 28307 14804 28319 14807
rect 28994 14804 29000 14816
rect 28307 14776 29000 14804
rect 28307 14773 28319 14776
rect 28261 14767 28319 14773
rect 28994 14764 29000 14776
rect 29052 14764 29058 14816
rect 29730 14764 29736 14816
rect 29788 14804 29794 14816
rect 30466 14804 30472 14816
rect 29788 14776 30472 14804
rect 29788 14764 29794 14776
rect 30466 14764 30472 14776
rect 30524 14804 30530 14816
rect 30650 14804 30656 14816
rect 30524 14776 30656 14804
rect 30524 14764 30530 14776
rect 30650 14764 30656 14776
rect 30708 14764 30714 14816
rect 30834 14764 30840 14816
rect 30892 14764 30898 14816
rect 31386 14764 31392 14816
rect 31444 14764 31450 14816
rect 1104 14714 32844 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 32844 14714
rect 1104 14640 32844 14662
rect 1486 14560 1492 14612
rect 1544 14600 1550 14612
rect 1581 14603 1639 14609
rect 1581 14600 1593 14603
rect 1544 14572 1593 14600
rect 1544 14560 1550 14572
rect 1581 14569 1593 14572
rect 1627 14569 1639 14603
rect 1581 14563 1639 14569
rect 3878 14560 3884 14612
rect 3936 14560 3942 14612
rect 4062 14560 4068 14612
rect 4120 14560 4126 14612
rect 4249 14603 4307 14609
rect 4249 14569 4261 14603
rect 4295 14600 4307 14603
rect 4706 14600 4712 14612
rect 4295 14572 4712 14600
rect 4295 14569 4307 14572
rect 4249 14563 4307 14569
rect 4706 14560 4712 14572
rect 4764 14560 4770 14612
rect 5445 14603 5503 14609
rect 5445 14569 5457 14603
rect 5491 14600 5503 14603
rect 5534 14600 5540 14612
rect 5491 14572 5540 14600
rect 5491 14569 5503 14572
rect 5445 14563 5503 14569
rect 5534 14560 5540 14572
rect 5592 14560 5598 14612
rect 5718 14560 5724 14612
rect 5776 14560 5782 14612
rect 6089 14603 6147 14609
rect 6089 14600 6101 14603
rect 5828 14572 6101 14600
rect 3896 14532 3924 14560
rect 4985 14535 5043 14541
rect 3896 14504 4108 14532
rect 3234 14424 3240 14476
rect 3292 14464 3298 14476
rect 3881 14467 3939 14473
rect 3881 14464 3893 14467
rect 3292 14436 3893 14464
rect 3292 14424 3298 14436
rect 3881 14433 3893 14436
rect 3927 14433 3939 14467
rect 3881 14427 3939 14433
rect 842 14356 848 14408
rect 900 14396 906 14408
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 900 14368 1409 14396
rect 900 14356 906 14368
rect 1397 14365 1409 14368
rect 1443 14365 1455 14399
rect 1397 14359 1455 14365
rect 3789 14399 3847 14405
rect 3789 14365 3801 14399
rect 3835 14396 3847 14399
rect 3970 14396 3976 14408
rect 3835 14368 3976 14396
rect 3835 14365 3847 14368
rect 3789 14359 3847 14365
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 4080 14405 4108 14504
rect 4985 14501 4997 14535
rect 5031 14532 5043 14535
rect 5828 14532 5856 14572
rect 6089 14569 6101 14572
rect 6135 14569 6147 14603
rect 6089 14563 6147 14569
rect 6549 14603 6607 14609
rect 6549 14569 6561 14603
rect 6595 14600 6607 14603
rect 6638 14600 6644 14612
rect 6595 14572 6644 14600
rect 6595 14569 6607 14572
rect 6549 14563 6607 14569
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 7374 14560 7380 14612
rect 7432 14560 7438 14612
rect 7837 14603 7895 14609
rect 7837 14569 7849 14603
rect 7883 14600 7895 14603
rect 8294 14600 8300 14612
rect 7883 14572 8300 14600
rect 7883 14569 7895 14572
rect 7837 14563 7895 14569
rect 8294 14560 8300 14572
rect 8352 14560 8358 14612
rect 9122 14560 9128 14612
rect 9180 14600 9186 14612
rect 9401 14603 9459 14609
rect 9401 14600 9413 14603
rect 9180 14572 9413 14600
rect 9180 14560 9186 14572
rect 9401 14569 9413 14572
rect 9447 14569 9459 14603
rect 9401 14563 9459 14569
rect 9861 14603 9919 14609
rect 9861 14569 9873 14603
rect 9907 14600 9919 14603
rect 9953 14603 10011 14609
rect 9953 14600 9965 14603
rect 9907 14572 9965 14600
rect 9907 14569 9919 14572
rect 9861 14563 9919 14569
rect 9953 14569 9965 14572
rect 9999 14569 10011 14603
rect 9953 14563 10011 14569
rect 11238 14560 11244 14612
rect 11296 14560 11302 14612
rect 11606 14560 11612 14612
rect 11664 14560 11670 14612
rect 11698 14560 11704 14612
rect 11756 14560 11762 14612
rect 12434 14600 12440 14612
rect 11808 14572 12440 14600
rect 5031 14504 5856 14532
rect 5997 14535 6055 14541
rect 5031 14501 5043 14504
rect 4985 14495 5043 14501
rect 5997 14501 6009 14535
rect 6043 14532 6055 14535
rect 6043 14504 6224 14532
rect 6043 14501 6055 14504
rect 5997 14495 6055 14501
rect 4614 14424 4620 14476
rect 4672 14464 4678 14476
rect 5629 14467 5687 14473
rect 4672 14436 5414 14464
rect 4672 14424 4678 14436
rect 4065 14399 4123 14405
rect 4065 14365 4077 14399
rect 4111 14365 4123 14399
rect 4065 14359 4123 14365
rect 4709 14399 4767 14405
rect 4709 14365 4721 14399
rect 4755 14365 4767 14399
rect 4709 14359 4767 14365
rect 4724 14328 4752 14359
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 5169 14399 5227 14405
rect 5169 14396 5181 14399
rect 4856 14368 5181 14396
rect 4856 14356 4862 14368
rect 5169 14365 5181 14368
rect 5215 14365 5227 14399
rect 5169 14359 5227 14365
rect 5261 14399 5319 14405
rect 5261 14365 5273 14399
rect 5307 14365 5319 14399
rect 5386 14396 5414 14436
rect 5629 14433 5641 14467
rect 5675 14464 5687 14467
rect 5902 14464 5908 14476
rect 5675 14436 5908 14464
rect 5675 14433 5687 14436
rect 5629 14427 5687 14433
rect 5902 14424 5908 14436
rect 5960 14424 5966 14476
rect 6196 14473 6224 14504
rect 6822 14492 6828 14544
rect 6880 14532 6886 14544
rect 7009 14535 7067 14541
rect 7009 14532 7021 14535
rect 6880 14504 7021 14532
rect 6880 14492 6886 14504
rect 7009 14501 7021 14504
rect 7055 14532 7067 14535
rect 8938 14532 8944 14544
rect 7055 14504 8944 14532
rect 7055 14501 7067 14504
rect 7009 14495 7067 14501
rect 8938 14492 8944 14504
rect 8996 14492 9002 14544
rect 9309 14535 9367 14541
rect 9309 14501 9321 14535
rect 9355 14532 9367 14535
rect 9490 14532 9496 14544
rect 9355 14504 9496 14532
rect 9355 14501 9367 14504
rect 9309 14495 9367 14501
rect 9490 14492 9496 14504
rect 9548 14492 9554 14544
rect 9674 14492 9680 14544
rect 9732 14532 9738 14544
rect 9732 14504 10088 14532
rect 9732 14492 9738 14504
rect 6181 14467 6239 14473
rect 6181 14433 6193 14467
rect 6227 14433 6239 14467
rect 6917 14467 6975 14473
rect 6917 14464 6929 14467
rect 6181 14427 6239 14433
rect 6564 14436 6929 14464
rect 6564 14408 6592 14436
rect 6917 14433 6929 14436
rect 6963 14464 6975 14467
rect 7282 14464 7288 14476
rect 6963 14436 7288 14464
rect 6963 14433 6975 14436
rect 6917 14427 6975 14433
rect 7282 14424 7288 14436
rect 7340 14424 7346 14476
rect 7561 14467 7619 14473
rect 7561 14433 7573 14467
rect 7607 14464 7619 14467
rect 7742 14464 7748 14476
rect 7607 14436 7748 14464
rect 7607 14433 7619 14436
rect 7561 14427 7619 14433
rect 7742 14424 7748 14436
rect 7800 14424 7806 14476
rect 7926 14424 7932 14476
rect 7984 14424 7990 14476
rect 8386 14424 8392 14476
rect 8444 14464 8450 14476
rect 9585 14467 9643 14473
rect 8444 14436 9352 14464
rect 8444 14424 8450 14436
rect 9324 14408 9352 14436
rect 9585 14433 9597 14467
rect 9631 14464 9643 14467
rect 9950 14464 9956 14476
rect 9631 14436 9956 14464
rect 9631 14433 9643 14436
rect 9585 14427 9643 14433
rect 9950 14424 9956 14436
rect 10008 14424 10014 14476
rect 10060 14473 10088 14504
rect 10594 14492 10600 14544
rect 10652 14532 10658 14544
rect 10689 14535 10747 14541
rect 10689 14532 10701 14535
rect 10652 14504 10701 14532
rect 10652 14492 10658 14504
rect 10689 14501 10701 14504
rect 10735 14501 10747 14535
rect 10689 14495 10747 14501
rect 11146 14492 11152 14544
rect 11204 14532 11210 14544
rect 11330 14532 11336 14544
rect 11204 14504 11336 14532
rect 11204 14492 11210 14504
rect 10045 14467 10103 14473
rect 10045 14433 10057 14467
rect 10091 14433 10103 14467
rect 10870 14464 10876 14476
rect 10045 14427 10103 14433
rect 10152 14436 10876 14464
rect 5537 14399 5595 14405
rect 5537 14396 5549 14399
rect 5386 14368 5549 14396
rect 5261 14359 5319 14365
rect 5537 14365 5549 14368
rect 5583 14365 5595 14399
rect 5537 14359 5595 14365
rect 4982 14328 4988 14340
rect 4724 14300 4988 14328
rect 4982 14288 4988 14300
rect 5040 14288 5046 14340
rect 5074 14288 5080 14340
rect 5132 14328 5138 14340
rect 5276 14328 5304 14359
rect 5810 14356 5816 14408
rect 5868 14356 5874 14408
rect 6365 14399 6423 14405
rect 6365 14365 6377 14399
rect 6411 14396 6423 14399
rect 6454 14396 6460 14408
rect 6411 14368 6460 14396
rect 6411 14365 6423 14368
rect 6365 14359 6423 14365
rect 6454 14356 6460 14368
rect 6512 14356 6518 14408
rect 6546 14356 6552 14408
rect 6604 14356 6610 14408
rect 6730 14356 6736 14408
rect 6788 14356 6794 14408
rect 7006 14356 7012 14408
rect 7064 14396 7070 14408
rect 7193 14399 7251 14405
rect 7193 14396 7205 14399
rect 7064 14368 7205 14396
rect 7064 14356 7070 14368
rect 7193 14365 7205 14368
rect 7239 14365 7251 14399
rect 7193 14359 7251 14365
rect 7650 14356 7656 14408
rect 7708 14396 7714 14408
rect 8205 14399 8263 14405
rect 8205 14396 8217 14399
rect 7708 14368 8217 14396
rect 7708 14356 7714 14368
rect 8205 14365 8217 14368
rect 8251 14365 8263 14399
rect 8205 14359 8263 14365
rect 8294 14356 8300 14408
rect 8352 14396 8358 14408
rect 9125 14399 9183 14405
rect 9125 14396 9137 14399
rect 8352 14368 9137 14396
rect 8352 14356 8358 14368
rect 9125 14365 9137 14368
rect 9171 14365 9183 14399
rect 9125 14359 9183 14365
rect 9306 14356 9312 14408
rect 9364 14356 9370 14408
rect 9677 14399 9735 14405
rect 9677 14365 9689 14399
rect 9723 14396 9735 14399
rect 9766 14396 9772 14408
rect 9723 14368 9772 14396
rect 9723 14365 9735 14368
rect 9677 14359 9735 14365
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 10152 14396 10180 14436
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 11256 14473 11284 14504
rect 11330 14492 11336 14504
rect 11388 14492 11394 14544
rect 11517 14535 11575 14541
rect 11517 14501 11529 14535
rect 11563 14532 11575 14535
rect 11716 14532 11744 14560
rect 11563 14504 11744 14532
rect 11563 14501 11575 14504
rect 11517 14495 11575 14501
rect 11241 14467 11299 14473
rect 11241 14433 11253 14467
rect 11287 14433 11299 14467
rect 11241 14427 11299 14433
rect 11698 14424 11704 14476
rect 11756 14424 11762 14476
rect 11808 14408 11836 14572
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 13078 14560 13084 14612
rect 13136 14600 13142 14612
rect 13357 14603 13415 14609
rect 13357 14600 13369 14603
rect 13136 14572 13369 14600
rect 13136 14560 13142 14572
rect 13357 14569 13369 14572
rect 13403 14569 13415 14603
rect 13357 14563 13415 14569
rect 15010 14560 15016 14612
rect 15068 14600 15074 14612
rect 15841 14603 15899 14609
rect 15841 14600 15853 14603
rect 15068 14572 15853 14600
rect 15068 14560 15074 14572
rect 15841 14569 15853 14572
rect 15887 14569 15899 14603
rect 15841 14563 15899 14569
rect 15948 14572 16436 14600
rect 11974 14492 11980 14544
rect 12032 14532 12038 14544
rect 12069 14535 12127 14541
rect 12069 14532 12081 14535
rect 12032 14504 12081 14532
rect 12032 14492 12038 14504
rect 12069 14501 12081 14504
rect 12115 14501 12127 14535
rect 12069 14495 12127 14501
rect 12161 14535 12219 14541
rect 12161 14501 12173 14535
rect 12207 14532 12219 14535
rect 12618 14532 12624 14544
rect 12207 14504 12624 14532
rect 12207 14501 12219 14504
rect 12161 14495 12219 14501
rect 12176 14464 12204 14495
rect 12618 14492 12624 14504
rect 12676 14492 12682 14544
rect 14642 14492 14648 14544
rect 14700 14532 14706 14544
rect 15948 14532 15976 14572
rect 14700 14504 15976 14532
rect 14700 14492 14706 14504
rect 16114 14492 16120 14544
rect 16172 14492 16178 14544
rect 16301 14535 16359 14541
rect 16301 14501 16313 14535
rect 16347 14501 16359 14535
rect 16408 14532 16436 14572
rect 16482 14560 16488 14612
rect 16540 14600 16546 14612
rect 16666 14600 16672 14612
rect 16540 14572 16672 14600
rect 16540 14560 16546 14572
rect 16666 14560 16672 14572
rect 16724 14560 16730 14612
rect 16758 14560 16764 14612
rect 16816 14560 16822 14612
rect 17497 14603 17555 14609
rect 17497 14569 17509 14603
rect 17543 14600 17555 14603
rect 17586 14600 17592 14612
rect 17543 14572 17592 14600
rect 17543 14569 17555 14572
rect 17497 14563 17555 14569
rect 17586 14560 17592 14572
rect 17644 14600 17650 14612
rect 18506 14600 18512 14612
rect 17644 14572 18512 14600
rect 17644 14560 17650 14572
rect 18506 14560 18512 14572
rect 18564 14560 18570 14612
rect 18601 14603 18659 14609
rect 18601 14569 18613 14603
rect 18647 14600 18659 14603
rect 18874 14600 18880 14612
rect 18647 14572 18880 14600
rect 18647 14569 18659 14572
rect 18601 14563 18659 14569
rect 18874 14560 18880 14572
rect 18932 14560 18938 14612
rect 19518 14560 19524 14612
rect 19576 14600 19582 14612
rect 19613 14603 19671 14609
rect 19613 14600 19625 14603
rect 19576 14572 19625 14600
rect 19576 14560 19582 14572
rect 19613 14569 19625 14572
rect 19659 14569 19671 14603
rect 19613 14563 19671 14569
rect 19904 14572 20116 14600
rect 19904 14532 19932 14572
rect 16408 14504 19932 14532
rect 16301 14495 16359 14501
rect 11992 14436 12204 14464
rect 9876 14368 10180 14396
rect 5132 14300 5304 14328
rect 5445 14331 5503 14337
rect 5132 14288 5138 14300
rect 5445 14297 5457 14331
rect 5491 14328 5503 14331
rect 5994 14328 6000 14340
rect 5491 14300 6000 14328
rect 5491 14297 5503 14300
rect 5445 14291 5503 14297
rect 5994 14288 6000 14300
rect 6052 14288 6058 14340
rect 6089 14331 6147 14337
rect 6089 14297 6101 14331
rect 6135 14328 6147 14331
rect 6178 14328 6184 14340
rect 6135 14300 6184 14328
rect 6135 14297 6147 14300
rect 6089 14291 6147 14297
rect 6178 14288 6184 14300
rect 6236 14288 6242 14340
rect 7282 14288 7288 14340
rect 7340 14328 7346 14340
rect 7377 14331 7435 14337
rect 7377 14328 7389 14331
rect 7340 14300 7389 14328
rect 7340 14288 7346 14300
rect 7377 14297 7389 14300
rect 7423 14297 7435 14331
rect 7377 14291 7435 14297
rect 8846 14288 8852 14340
rect 8904 14328 8910 14340
rect 9401 14331 9459 14337
rect 9401 14328 9413 14331
rect 8904 14300 9413 14328
rect 8904 14288 8910 14300
rect 9401 14297 9413 14300
rect 9447 14328 9459 14331
rect 9876 14328 9904 14368
rect 10226 14356 10232 14408
rect 10284 14356 10290 14408
rect 11149 14399 11207 14405
rect 11149 14396 11161 14399
rect 10336 14368 11161 14396
rect 9447 14300 9904 14328
rect 9447 14297 9459 14300
rect 9401 14291 9459 14297
rect 9950 14288 9956 14340
rect 10008 14288 10014 14340
rect 4893 14263 4951 14269
rect 4893 14229 4905 14263
rect 4939 14260 4951 14263
rect 5534 14260 5540 14272
rect 4939 14232 5540 14260
rect 4939 14229 4951 14232
rect 4893 14223 4951 14229
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 5810 14220 5816 14272
rect 5868 14260 5874 14272
rect 6822 14260 6828 14272
rect 5868 14232 6828 14260
rect 5868 14220 5874 14232
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 7466 14220 7472 14272
rect 7524 14260 7530 14272
rect 10336 14260 10364 14368
rect 11149 14365 11161 14368
rect 11195 14396 11207 14399
rect 11790 14396 11796 14408
rect 11195 14368 11796 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 11882 14356 11888 14408
rect 11940 14356 11946 14408
rect 10594 14288 10600 14340
rect 10652 14328 10658 14340
rect 10873 14331 10931 14337
rect 10873 14328 10885 14331
rect 10652 14300 10885 14328
rect 10652 14288 10658 14300
rect 10873 14297 10885 14300
rect 10919 14328 10931 14331
rect 10962 14328 10968 14340
rect 10919 14300 10968 14328
rect 10919 14297 10931 14300
rect 10873 14291 10931 14297
rect 10962 14288 10968 14300
rect 11020 14288 11026 14340
rect 11057 14331 11115 14337
rect 11057 14297 11069 14331
rect 11103 14297 11115 14331
rect 11057 14291 11115 14297
rect 7524 14232 10364 14260
rect 7524 14220 7530 14232
rect 10410 14220 10416 14272
rect 10468 14220 10474 14272
rect 11072 14260 11100 14291
rect 11514 14288 11520 14340
rect 11572 14328 11578 14340
rect 11609 14331 11667 14337
rect 11609 14328 11621 14331
rect 11572 14300 11621 14328
rect 11572 14288 11578 14300
rect 11609 14297 11621 14300
rect 11655 14297 11667 14331
rect 11609 14291 11667 14297
rect 11698 14288 11704 14340
rect 11756 14328 11762 14340
rect 11992 14328 12020 14436
rect 12250 14424 12256 14476
rect 12308 14464 12314 14476
rect 13449 14467 13507 14473
rect 13449 14464 13461 14467
rect 12308 14436 13461 14464
rect 12308 14424 12314 14436
rect 13449 14433 13461 14436
rect 13495 14433 13507 14467
rect 16132 14464 16160 14492
rect 13449 14427 13507 14433
rect 14016 14436 16160 14464
rect 12066 14356 12072 14408
rect 12124 14396 12130 14408
rect 12345 14399 12403 14405
rect 12345 14396 12357 14399
rect 12124 14368 12357 14396
rect 12124 14356 12130 14368
rect 12345 14365 12357 14368
rect 12391 14365 12403 14399
rect 13078 14396 13084 14408
rect 12345 14359 12403 14365
rect 12544 14368 13084 14396
rect 11756 14300 12020 14328
rect 11756 14288 11762 14300
rect 12250 14288 12256 14340
rect 12308 14328 12314 14340
rect 12544 14328 12572 14368
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 13262 14356 13268 14408
rect 13320 14396 13326 14408
rect 13357 14399 13415 14405
rect 13357 14396 13369 14399
rect 13320 14368 13369 14396
rect 13320 14356 13326 14368
rect 13357 14365 13369 14368
rect 13403 14365 13415 14399
rect 14016 14396 14044 14436
rect 13357 14359 13415 14365
rect 13556 14368 14044 14396
rect 12308 14300 12572 14328
rect 12308 14288 12314 14300
rect 12618 14288 12624 14340
rect 12676 14328 12682 14340
rect 13556 14328 13584 14368
rect 14090 14356 14096 14408
rect 14148 14396 14154 14408
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 14148 14368 15853 14396
rect 14148 14356 14154 14368
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 16025 14399 16083 14405
rect 16025 14365 16037 14399
rect 16071 14365 16083 14399
rect 16025 14359 16083 14365
rect 16117 14399 16175 14405
rect 16117 14365 16129 14399
rect 16163 14396 16175 14399
rect 16206 14396 16212 14408
rect 16163 14368 16212 14396
rect 16163 14365 16175 14368
rect 16117 14359 16175 14365
rect 14642 14328 14648 14340
rect 12676 14300 13584 14328
rect 13648 14300 14648 14328
rect 12676 14288 12682 14300
rect 11330 14260 11336 14272
rect 11072 14232 11336 14260
rect 11330 14220 11336 14232
rect 11388 14260 11394 14272
rect 13648 14260 13676 14300
rect 14642 14288 14648 14300
rect 14700 14288 14706 14340
rect 15378 14288 15384 14340
rect 15436 14288 15442 14340
rect 15562 14288 15568 14340
rect 15620 14288 15626 14340
rect 16040 14328 16068 14359
rect 16206 14356 16212 14368
rect 16264 14356 16270 14408
rect 16316 14328 16344 14495
rect 19978 14492 19984 14544
rect 20036 14492 20042 14544
rect 20088 14532 20116 14572
rect 20806 14560 20812 14612
rect 20864 14600 20870 14612
rect 22097 14603 22155 14609
rect 22097 14600 22109 14603
rect 20864 14572 22109 14600
rect 20864 14560 20870 14572
rect 22097 14569 22109 14572
rect 22143 14569 22155 14603
rect 22097 14563 22155 14569
rect 23569 14603 23627 14609
rect 23569 14569 23581 14603
rect 23615 14569 23627 14603
rect 23569 14563 23627 14569
rect 20088 14504 20300 14532
rect 17034 14424 17040 14476
rect 17092 14464 17098 14476
rect 17313 14467 17371 14473
rect 17313 14464 17325 14467
rect 17092 14436 17325 14464
rect 17092 14424 17098 14436
rect 17313 14433 17325 14436
rect 17359 14433 17371 14467
rect 17770 14464 17776 14476
rect 17313 14427 17371 14433
rect 17420 14436 17776 14464
rect 16390 14356 16396 14408
rect 16448 14356 16454 14408
rect 16482 14356 16488 14408
rect 16540 14356 16546 14408
rect 16942 14356 16948 14408
rect 17000 14396 17006 14408
rect 17420 14396 17448 14436
rect 17770 14424 17776 14436
rect 17828 14464 17834 14476
rect 18417 14467 18475 14473
rect 18417 14464 18429 14467
rect 17828 14436 18429 14464
rect 17828 14424 17834 14436
rect 18417 14433 18429 14436
rect 18463 14433 18475 14467
rect 18417 14427 18475 14433
rect 18524 14436 19564 14464
rect 17000 14368 17448 14396
rect 17497 14399 17555 14405
rect 17000 14356 17006 14368
rect 17497 14365 17509 14399
rect 17543 14396 17555 14399
rect 18524 14396 18552 14436
rect 17543 14368 18552 14396
rect 18601 14399 18659 14405
rect 17543 14365 17555 14368
rect 17497 14359 17555 14365
rect 18601 14365 18613 14399
rect 18647 14396 18659 14399
rect 18782 14396 18788 14408
rect 18647 14368 18788 14396
rect 18647 14365 18659 14368
rect 18601 14359 18659 14365
rect 18782 14356 18788 14368
rect 18840 14356 18846 14408
rect 17221 14331 17279 14337
rect 17221 14328 17233 14331
rect 16040 14300 16160 14328
rect 16316 14300 17233 14328
rect 11388 14232 13676 14260
rect 13725 14263 13783 14269
rect 11388 14220 11394 14232
rect 13725 14229 13737 14263
rect 13771 14260 13783 14263
rect 15194 14260 15200 14272
rect 13771 14232 15200 14260
rect 13771 14229 13783 14232
rect 13725 14223 13783 14229
rect 15194 14220 15200 14232
rect 15252 14220 15258 14272
rect 15749 14263 15807 14269
rect 15749 14229 15761 14263
rect 15795 14260 15807 14263
rect 16022 14260 16028 14272
rect 15795 14232 16028 14260
rect 15795 14229 15807 14232
rect 15749 14223 15807 14229
rect 16022 14220 16028 14232
rect 16080 14220 16086 14272
rect 16132 14260 16160 14300
rect 17221 14297 17233 14300
rect 17267 14297 17279 14331
rect 17221 14291 17279 14297
rect 17328 14300 17816 14328
rect 17328 14260 17356 14300
rect 16132 14232 17356 14260
rect 17678 14220 17684 14272
rect 17736 14220 17742 14272
rect 17788 14260 17816 14300
rect 18230 14288 18236 14340
rect 18288 14328 18294 14340
rect 18325 14331 18383 14337
rect 18325 14328 18337 14331
rect 18288 14300 18337 14328
rect 18288 14288 18294 14300
rect 18325 14297 18337 14300
rect 18371 14297 18383 14331
rect 19334 14328 19340 14340
rect 18325 14291 18383 14297
rect 18432 14300 19340 14328
rect 18432 14260 18460 14300
rect 19334 14288 19340 14300
rect 19392 14288 19398 14340
rect 19536 14328 19564 14436
rect 19613 14399 19671 14405
rect 19613 14365 19625 14399
rect 19659 14396 19671 14399
rect 19702 14396 19708 14408
rect 19659 14368 19708 14396
rect 19659 14365 19671 14368
rect 19613 14359 19671 14365
rect 19702 14356 19708 14368
rect 19760 14356 19766 14408
rect 19794 14356 19800 14408
rect 19852 14356 19858 14408
rect 20070 14356 20076 14408
rect 20128 14356 20134 14408
rect 20272 14405 20300 14504
rect 20714 14492 20720 14544
rect 20772 14532 20778 14544
rect 22005 14535 22063 14541
rect 22005 14532 22017 14535
rect 20772 14504 22017 14532
rect 20772 14492 20778 14504
rect 22005 14501 22017 14504
rect 22051 14532 22063 14535
rect 23584 14532 23612 14563
rect 24302 14560 24308 14612
rect 24360 14600 24366 14612
rect 24673 14603 24731 14609
rect 24673 14600 24685 14603
rect 24360 14572 24685 14600
rect 24360 14560 24366 14572
rect 24673 14569 24685 14572
rect 24719 14569 24731 14603
rect 24673 14563 24731 14569
rect 24762 14560 24768 14612
rect 24820 14600 24826 14612
rect 25041 14603 25099 14609
rect 25041 14600 25053 14603
rect 24820 14572 25053 14600
rect 24820 14560 24826 14572
rect 25041 14569 25053 14572
rect 25087 14569 25099 14603
rect 27062 14600 27068 14612
rect 25041 14563 25099 14569
rect 25608 14572 27068 14600
rect 22051 14504 23612 14532
rect 23937 14535 23995 14541
rect 22051 14501 22063 14504
rect 22005 14495 22063 14501
rect 23937 14501 23949 14535
rect 23983 14532 23995 14535
rect 25608 14532 25636 14572
rect 27062 14560 27068 14572
rect 27120 14560 27126 14612
rect 27522 14560 27528 14612
rect 27580 14600 27586 14612
rect 28813 14603 28871 14609
rect 28813 14600 28825 14603
rect 27580 14572 28825 14600
rect 27580 14560 27586 14572
rect 28813 14569 28825 14572
rect 28859 14569 28871 14603
rect 28813 14563 28871 14569
rect 30282 14560 30288 14612
rect 30340 14560 30346 14612
rect 30377 14603 30435 14609
rect 30377 14569 30389 14603
rect 30423 14600 30435 14603
rect 30558 14600 30564 14612
rect 30423 14572 30564 14600
rect 30423 14569 30435 14572
rect 30377 14563 30435 14569
rect 30558 14560 30564 14572
rect 30616 14560 30622 14612
rect 30653 14603 30711 14609
rect 30653 14569 30665 14603
rect 30699 14600 30711 14603
rect 30742 14600 30748 14612
rect 30699 14572 30748 14600
rect 30699 14569 30711 14572
rect 30653 14563 30711 14569
rect 23983 14504 25636 14532
rect 25685 14535 25743 14541
rect 23983 14501 23995 14504
rect 23937 14495 23995 14501
rect 25685 14501 25697 14535
rect 25731 14532 25743 14535
rect 27798 14532 27804 14544
rect 25731 14504 27804 14532
rect 25731 14501 25743 14504
rect 25685 14495 25743 14501
rect 27798 14492 27804 14504
rect 27856 14492 27862 14544
rect 28537 14535 28595 14541
rect 28537 14501 28549 14535
rect 28583 14532 28595 14535
rect 30006 14532 30012 14544
rect 28583 14504 30012 14532
rect 28583 14501 28595 14504
rect 28537 14495 28595 14501
rect 30006 14492 30012 14504
rect 30064 14492 30070 14544
rect 30668 14532 30696 14563
rect 30742 14560 30748 14572
rect 30800 14560 30806 14612
rect 30926 14560 30932 14612
rect 30984 14600 30990 14612
rect 31205 14603 31263 14609
rect 31205 14600 31217 14603
rect 30984 14572 31217 14600
rect 30984 14560 30990 14572
rect 31205 14569 31217 14572
rect 31251 14569 31263 14603
rect 31205 14563 31263 14569
rect 30116 14504 30696 14532
rect 20441 14467 20499 14473
rect 20441 14433 20453 14467
rect 20487 14464 20499 14467
rect 24486 14464 24492 14476
rect 20487 14436 24492 14464
rect 20487 14433 20499 14436
rect 20441 14427 20499 14433
rect 20257 14399 20315 14405
rect 20257 14365 20269 14399
rect 20303 14365 20315 14399
rect 20257 14359 20315 14365
rect 20346 14356 20352 14408
rect 20404 14396 20410 14408
rect 20456 14396 20484 14427
rect 23290 14396 23296 14408
rect 20404 14368 20484 14396
rect 21376 14368 23296 14396
rect 20404 14356 20410 14368
rect 21376 14328 21404 14368
rect 23290 14356 23296 14368
rect 23348 14396 23354 14408
rect 23584 14405 23612 14436
rect 24486 14424 24492 14436
rect 24544 14424 24550 14476
rect 25222 14464 25228 14476
rect 24688 14436 25228 14464
rect 24688 14405 24716 14436
rect 25222 14424 25228 14436
rect 25280 14424 25286 14476
rect 26252 14436 27568 14464
rect 23569 14399 23627 14405
rect 23348 14368 23520 14396
rect 23348 14356 23354 14368
rect 19536 14300 20024 14328
rect 17788 14232 18460 14260
rect 18785 14263 18843 14269
rect 18785 14229 18797 14263
rect 18831 14260 18843 14263
rect 19242 14260 19248 14272
rect 18831 14232 19248 14260
rect 18831 14229 18843 14232
rect 18785 14223 18843 14229
rect 19242 14220 19248 14232
rect 19300 14220 19306 14272
rect 19996 14260 20024 14300
rect 20456 14300 21404 14328
rect 20456 14260 20484 14300
rect 21450 14288 21456 14340
rect 21508 14288 21514 14340
rect 21634 14288 21640 14340
rect 21692 14288 21698 14340
rect 21913 14331 21971 14337
rect 21913 14328 21925 14331
rect 21744 14300 21925 14328
rect 19996 14232 20484 14260
rect 20530 14220 20536 14272
rect 20588 14260 20594 14272
rect 21744 14260 21772 14300
rect 21913 14297 21925 14300
rect 21959 14297 21971 14331
rect 22281 14331 22339 14337
rect 22281 14328 22293 14331
rect 21913 14291 21971 14297
rect 22066 14300 22293 14328
rect 20588 14232 21772 14260
rect 21821 14263 21879 14269
rect 20588 14220 20594 14232
rect 21821 14229 21833 14263
rect 21867 14260 21879 14263
rect 22066 14260 22094 14300
rect 22281 14297 22293 14300
rect 22327 14328 22339 14331
rect 22554 14328 22560 14340
rect 22327 14300 22560 14328
rect 22327 14297 22339 14300
rect 22281 14291 22339 14297
rect 22554 14288 22560 14300
rect 22612 14288 22618 14340
rect 22922 14288 22928 14340
rect 22980 14328 22986 14340
rect 23198 14328 23204 14340
rect 22980 14300 23204 14328
rect 22980 14288 22986 14300
rect 23198 14288 23204 14300
rect 23256 14288 23262 14340
rect 23492 14328 23520 14368
rect 23569 14365 23581 14399
rect 23615 14365 23627 14399
rect 23569 14359 23627 14365
rect 23661 14399 23719 14405
rect 23661 14365 23673 14399
rect 23707 14365 23719 14399
rect 23661 14359 23719 14365
rect 24673 14399 24731 14405
rect 24673 14365 24685 14399
rect 24719 14365 24731 14399
rect 24673 14359 24731 14365
rect 23676 14328 23704 14359
rect 24762 14356 24768 14408
rect 24820 14356 24826 14408
rect 25501 14399 25559 14405
rect 25501 14396 25513 14399
rect 24872 14368 25513 14396
rect 24872 14328 24900 14368
rect 25501 14365 25513 14368
rect 25547 14365 25559 14399
rect 25501 14359 25559 14365
rect 26252 14340 26280 14436
rect 26970 14396 26976 14408
rect 26528 14368 26976 14396
rect 23492 14300 23704 14328
rect 23860 14300 24900 14328
rect 24949 14331 25007 14337
rect 21867 14232 22094 14260
rect 22189 14263 22247 14269
rect 21867 14229 21879 14232
rect 21821 14223 21879 14229
rect 22189 14229 22201 14263
rect 22235 14260 22247 14263
rect 23860 14260 23888 14300
rect 24949 14297 24961 14331
rect 24995 14297 25007 14331
rect 24949 14291 25007 14297
rect 22235 14232 23888 14260
rect 22235 14229 22247 14232
rect 22189 14223 22247 14229
rect 24486 14220 24492 14272
rect 24544 14220 24550 14272
rect 24964 14260 24992 14291
rect 25222 14288 25228 14340
rect 25280 14288 25286 14340
rect 25409 14331 25467 14337
rect 25409 14297 25421 14331
rect 25455 14328 25467 14331
rect 25590 14328 25596 14340
rect 25455 14300 25596 14328
rect 25455 14297 25467 14300
rect 25409 14291 25467 14297
rect 25590 14288 25596 14300
rect 25648 14328 25654 14340
rect 25958 14328 25964 14340
rect 25648 14300 25964 14328
rect 25648 14288 25654 14300
rect 25958 14288 25964 14300
rect 26016 14288 26022 14340
rect 26234 14288 26240 14340
rect 26292 14288 26298 14340
rect 26528 14260 26556 14368
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 27062 14356 27068 14408
rect 27120 14396 27126 14408
rect 27430 14396 27436 14408
rect 27120 14368 27436 14396
rect 27120 14356 27126 14368
rect 27430 14356 27436 14368
rect 27488 14356 27494 14408
rect 27540 14328 27568 14436
rect 27614 14424 27620 14476
rect 27672 14464 27678 14476
rect 28629 14467 28687 14473
rect 28629 14464 28641 14467
rect 27672 14436 28641 14464
rect 27672 14424 27678 14436
rect 28629 14433 28641 14436
rect 28675 14433 28687 14467
rect 28629 14427 28687 14433
rect 27982 14356 27988 14408
rect 28040 14396 28046 14408
rect 28169 14399 28227 14405
rect 28169 14396 28181 14399
rect 28040 14368 28181 14396
rect 28040 14356 28046 14368
rect 28169 14365 28181 14368
rect 28215 14365 28227 14399
rect 28644 14396 28672 14427
rect 28994 14424 29000 14476
rect 29052 14464 29058 14476
rect 29822 14464 29828 14476
rect 29052 14436 29828 14464
rect 29052 14424 29058 14436
rect 29822 14424 29828 14436
rect 29880 14424 29886 14476
rect 29089 14399 29147 14405
rect 29089 14396 29101 14399
rect 28644 14368 29101 14396
rect 28169 14359 28227 14365
rect 29089 14365 29101 14368
rect 29135 14365 29147 14399
rect 29089 14359 29147 14365
rect 29178 14356 29184 14408
rect 29236 14396 29242 14408
rect 30116 14405 30144 14504
rect 30944 14464 30972 14560
rect 30576 14436 30972 14464
rect 30576 14405 30604 14436
rect 31754 14424 31760 14476
rect 31812 14464 31818 14476
rect 31941 14467 31999 14473
rect 31941 14464 31953 14467
rect 31812 14436 31953 14464
rect 31812 14424 31818 14436
rect 31941 14433 31953 14436
rect 31987 14433 31999 14467
rect 31941 14427 31999 14433
rect 30101 14399 30159 14405
rect 29236 14368 30052 14396
rect 29236 14356 29242 14368
rect 27614 14328 27620 14340
rect 27540 14300 27620 14328
rect 27614 14288 27620 14300
rect 27672 14288 27678 14340
rect 27706 14288 27712 14340
rect 27764 14328 27770 14340
rect 28353 14331 28411 14337
rect 28353 14328 28365 14331
rect 27764 14300 28365 14328
rect 27764 14288 27770 14300
rect 28353 14297 28365 14300
rect 28399 14297 28411 14331
rect 28353 14291 28411 14297
rect 28810 14288 28816 14340
rect 28868 14288 28874 14340
rect 24964 14232 26556 14260
rect 26602 14220 26608 14272
rect 26660 14260 26666 14272
rect 27430 14260 27436 14272
rect 26660 14232 27436 14260
rect 26660 14220 26666 14232
rect 27430 14220 27436 14232
rect 27488 14220 27494 14272
rect 29273 14263 29331 14269
rect 29273 14229 29285 14263
rect 29319 14260 29331 14263
rect 29822 14260 29828 14272
rect 29319 14232 29828 14260
rect 29319 14229 29331 14232
rect 29273 14223 29331 14229
rect 29822 14220 29828 14232
rect 29880 14220 29886 14272
rect 30024 14260 30052 14368
rect 30101 14365 30113 14399
rect 30147 14365 30159 14399
rect 30101 14359 30159 14365
rect 30561 14399 30619 14405
rect 30561 14365 30573 14399
rect 30607 14365 30619 14399
rect 30561 14359 30619 14365
rect 30837 14399 30895 14405
rect 30837 14365 30849 14399
rect 30883 14365 30895 14399
rect 30837 14359 30895 14365
rect 30852 14328 30880 14359
rect 30926 14356 30932 14408
rect 30984 14356 30990 14408
rect 31386 14356 31392 14408
rect 31444 14356 31450 14408
rect 31662 14356 31668 14408
rect 31720 14356 31726 14408
rect 30852 14300 31064 14328
rect 31036 14272 31064 14300
rect 30282 14260 30288 14272
rect 30024 14232 30288 14260
rect 30282 14220 30288 14232
rect 30340 14220 30346 14272
rect 31018 14220 31024 14272
rect 31076 14260 31082 14272
rect 31113 14263 31171 14269
rect 31113 14260 31125 14263
rect 31076 14232 31125 14260
rect 31076 14220 31082 14232
rect 31113 14229 31125 14232
rect 31159 14229 31171 14263
rect 31113 14223 31171 14229
rect 31846 14220 31852 14272
rect 31904 14260 31910 14272
rect 32122 14260 32128 14272
rect 31904 14232 32128 14260
rect 31904 14220 31910 14232
rect 32122 14220 32128 14232
rect 32180 14220 32186 14272
rect 1104 14170 32844 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 32844 14170
rect 1104 14096 32844 14118
rect 3697 14059 3755 14065
rect 3697 14025 3709 14059
rect 3743 14025 3755 14059
rect 3697 14019 3755 14025
rect 3973 14059 4031 14065
rect 3973 14025 3985 14059
rect 4019 14056 4031 14059
rect 4614 14056 4620 14068
rect 4019 14028 4620 14056
rect 4019 14025 4031 14028
rect 3973 14019 4031 14025
rect 3712 13988 3740 14019
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 4706 14016 4712 14068
rect 4764 14056 4770 14068
rect 5718 14056 5724 14068
rect 4764 14028 5724 14056
rect 4764 14016 4770 14028
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 5994 14016 6000 14068
rect 6052 14016 6058 14068
rect 7282 14016 7288 14068
rect 7340 14016 7346 14068
rect 8202 14056 8208 14068
rect 7668 14028 8208 14056
rect 3712 13960 4568 13988
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 3142 13920 3148 13932
rect 2731 13892 3148 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 3142 13880 3148 13892
rect 3200 13880 3206 13932
rect 3510 13880 3516 13932
rect 3568 13880 3574 13932
rect 3694 13880 3700 13932
rect 3752 13920 3758 13932
rect 3789 13923 3847 13929
rect 3789 13920 3801 13923
rect 3752 13892 3801 13920
rect 3752 13880 3758 13892
rect 3789 13889 3801 13892
rect 3835 13889 3847 13923
rect 3789 13883 3847 13889
rect 3878 13880 3884 13932
rect 3936 13920 3942 13932
rect 4540 13929 4568 13960
rect 5534 13948 5540 14000
rect 5592 13948 5598 14000
rect 7668 13988 7696 14028
rect 8202 14016 8208 14028
rect 8260 14056 8266 14068
rect 8260 14028 9175 14056
rect 8260 14016 8266 14028
rect 5828 13960 7696 13988
rect 4065 13923 4123 13929
rect 4065 13920 4077 13923
rect 3936 13892 4077 13920
rect 3936 13880 3942 13892
rect 4065 13889 4077 13892
rect 4111 13889 4123 13923
rect 4065 13883 4123 13889
rect 4525 13923 4583 13929
rect 4525 13889 4537 13923
rect 4571 13920 4583 13923
rect 4982 13920 4988 13932
rect 4571 13892 4988 13920
rect 4571 13889 4583 13892
rect 4525 13883 4583 13889
rect 4982 13880 4988 13892
rect 5040 13880 5046 13932
rect 5350 13880 5356 13932
rect 5408 13920 5414 13932
rect 5718 13920 5724 13932
rect 5408 13892 5724 13920
rect 5408 13880 5414 13892
rect 5718 13880 5724 13892
rect 5776 13880 5782 13932
rect 5828 13929 5856 13960
rect 7742 13948 7748 14000
rect 7800 13948 7806 14000
rect 8386 13948 8392 14000
rect 8444 13988 8450 14000
rect 9033 13991 9091 13997
rect 9033 13988 9045 13991
rect 8444 13960 9045 13988
rect 8444 13948 8450 13960
rect 9033 13957 9045 13960
rect 9079 13957 9091 13991
rect 9033 13951 9091 13957
rect 5813 13923 5871 13929
rect 5813 13889 5825 13923
rect 5859 13889 5871 13923
rect 5813 13883 5871 13889
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 8570 13920 8576 13932
rect 7515 13892 8576 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 8570 13880 8576 13892
rect 8628 13880 8634 13932
rect 8662 13880 8668 13932
rect 8720 13880 8726 13932
rect 8757 13923 8815 13929
rect 8757 13889 8769 13923
rect 8803 13889 8815 13923
rect 8757 13883 8815 13889
rect 3970 13812 3976 13864
rect 4028 13852 4034 13864
rect 4890 13852 4896 13864
rect 4028 13824 4896 13852
rect 4028 13812 4034 13824
rect 4890 13812 4896 13824
rect 4948 13812 4954 13864
rect 5626 13812 5632 13864
rect 5684 13812 5690 13864
rect 5994 13812 6000 13864
rect 6052 13852 6058 13864
rect 6362 13852 6368 13864
rect 6052 13824 6368 13852
rect 6052 13812 6058 13824
rect 6362 13812 6368 13824
rect 6420 13812 6426 13864
rect 6917 13855 6975 13861
rect 6917 13821 6929 13855
rect 6963 13821 6975 13855
rect 6917 13815 6975 13821
rect 2682 13744 2688 13796
rect 2740 13784 2746 13796
rect 6932 13784 6960 13815
rect 7190 13812 7196 13864
rect 7248 13812 7254 13864
rect 7374 13812 7380 13864
rect 7432 13852 7438 13864
rect 7561 13855 7619 13861
rect 7561 13852 7573 13855
rect 7432 13824 7573 13852
rect 7432 13812 7438 13824
rect 7561 13821 7573 13824
rect 7607 13821 7619 13855
rect 7561 13815 7619 13821
rect 7650 13812 7656 13864
rect 7708 13852 7714 13864
rect 8772 13852 8800 13883
rect 7708 13824 8800 13852
rect 7708 13812 7714 13824
rect 7006 13784 7012 13796
rect 2740 13756 7012 13784
rect 2740 13744 2746 13756
rect 7006 13744 7012 13756
rect 7064 13744 7070 13796
rect 8662 13744 8668 13796
rect 8720 13784 8726 13796
rect 8720 13756 9076 13784
rect 8720 13744 8726 13756
rect 9048 13728 9076 13756
rect 2498 13676 2504 13728
rect 2556 13676 2562 13728
rect 3694 13676 3700 13728
rect 3752 13716 3758 13728
rect 4246 13716 4252 13728
rect 3752 13688 4252 13716
rect 3752 13676 3758 13688
rect 4246 13676 4252 13688
rect 4304 13676 4310 13728
rect 4341 13719 4399 13725
rect 4341 13685 4353 13719
rect 4387 13716 4399 13719
rect 4706 13716 4712 13728
rect 4387 13688 4712 13716
rect 4387 13685 4399 13688
rect 4341 13679 4399 13685
rect 4706 13676 4712 13688
rect 4764 13676 4770 13728
rect 5813 13719 5871 13725
rect 5813 13685 5825 13719
rect 5859 13716 5871 13719
rect 6638 13716 6644 13728
rect 5859 13688 6644 13716
rect 5859 13685 5871 13688
rect 5813 13679 5871 13685
rect 6638 13676 6644 13688
rect 6696 13676 6702 13728
rect 7466 13676 7472 13728
rect 7524 13676 7530 13728
rect 8478 13676 8484 13728
rect 8536 13676 8542 13728
rect 8846 13676 8852 13728
rect 8904 13716 8910 13728
rect 8941 13719 8999 13725
rect 8941 13716 8953 13719
rect 8904 13688 8953 13716
rect 8904 13676 8910 13688
rect 8941 13685 8953 13688
rect 8987 13685 8999 13719
rect 8941 13679 8999 13685
rect 9030 13676 9036 13728
rect 9088 13676 9094 13728
rect 9147 13716 9175 14028
rect 9306 14016 9312 14068
rect 9364 14016 9370 14068
rect 9493 14059 9551 14065
rect 9493 14025 9505 14059
rect 9539 14056 9551 14059
rect 10226 14056 10232 14068
rect 9539 14028 10232 14056
rect 9539 14025 9551 14028
rect 9493 14019 9551 14025
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 10410 14016 10416 14068
rect 10468 14056 10474 14068
rect 11238 14056 11244 14068
rect 10468 14028 11244 14056
rect 10468 14016 10474 14028
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 11330 14016 11336 14068
rect 11388 14016 11394 14068
rect 11514 14016 11520 14068
rect 11572 14056 11578 14068
rect 12250 14056 12256 14068
rect 11572 14028 12256 14056
rect 11572 14016 11578 14028
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 12437 14059 12495 14065
rect 12437 14025 12449 14059
rect 12483 14056 12495 14059
rect 12526 14056 12532 14068
rect 12483 14028 12532 14056
rect 12483 14025 12495 14028
rect 12437 14019 12495 14025
rect 12526 14016 12532 14028
rect 12584 14016 12590 14068
rect 13170 14016 13176 14068
rect 13228 14016 13234 14068
rect 13446 14016 13452 14068
rect 13504 14016 13510 14068
rect 13541 14059 13599 14065
rect 13541 14025 13553 14059
rect 13587 14056 13599 14059
rect 13630 14056 13636 14068
rect 13587 14028 13636 14056
rect 13587 14025 13599 14028
rect 13541 14019 13599 14025
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 14645 14059 14703 14065
rect 14645 14025 14657 14059
rect 14691 14025 14703 14059
rect 14645 14019 14703 14025
rect 9324 13988 9352 14016
rect 9324 13960 11928 13988
rect 9306 13880 9312 13932
rect 9364 13880 9370 13932
rect 9582 13880 9588 13932
rect 9640 13920 9646 13932
rect 9769 13923 9827 13929
rect 9769 13920 9781 13923
rect 9640 13892 9781 13920
rect 9640 13880 9646 13892
rect 9769 13889 9781 13892
rect 9815 13889 9827 13923
rect 9769 13883 9827 13889
rect 9858 13880 9864 13932
rect 9916 13880 9922 13932
rect 10134 13880 10140 13932
rect 10192 13920 10198 13932
rect 10321 13923 10379 13929
rect 10321 13920 10333 13923
rect 10192 13892 10333 13920
rect 10192 13880 10198 13892
rect 10321 13889 10333 13892
rect 10367 13889 10379 13923
rect 10321 13883 10379 13889
rect 10870 13880 10876 13932
rect 10928 13920 10934 13932
rect 11149 13923 11207 13929
rect 11149 13920 11161 13923
rect 10928 13892 11161 13920
rect 10928 13880 10934 13892
rect 11149 13889 11161 13892
rect 11195 13889 11207 13923
rect 11149 13883 11207 13889
rect 11698 13880 11704 13932
rect 11756 13880 11762 13932
rect 11900 13920 11928 13960
rect 11974 13948 11980 14000
rect 12032 13948 12038 14000
rect 14660 13988 14688 14019
rect 14918 14016 14924 14068
rect 14976 14056 14982 14068
rect 20806 14056 20812 14068
rect 14976 14028 20812 14056
rect 14976 14016 14982 14028
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 21082 14016 21088 14068
rect 21140 14016 21146 14068
rect 21177 14059 21235 14065
rect 21177 14025 21189 14059
rect 21223 14056 21235 14059
rect 24305 14059 24363 14065
rect 21223 14028 24164 14056
rect 21223 14025 21235 14028
rect 21177 14019 21235 14025
rect 15105 13991 15163 13997
rect 15105 13988 15117 13991
rect 12084 13960 14688 13988
rect 14752 13960 15117 13988
rect 12084 13920 12112 13960
rect 11900 13892 12112 13920
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13920 12311 13923
rect 12434 13920 12440 13932
rect 12299 13892 12440 13920
rect 12299 13889 12311 13892
rect 12253 13883 12311 13889
rect 12434 13880 12440 13892
rect 12492 13880 12498 13932
rect 12526 13880 12532 13932
rect 12584 13920 12590 13932
rect 12713 13923 12771 13929
rect 12713 13920 12725 13923
rect 12584 13892 12725 13920
rect 12584 13880 12590 13892
rect 12713 13889 12725 13892
rect 12759 13889 12771 13923
rect 12713 13883 12771 13889
rect 12802 13880 12808 13932
rect 12860 13920 12866 13932
rect 12897 13923 12955 13929
rect 12897 13920 12909 13923
rect 12860 13892 12909 13920
rect 12860 13880 12866 13892
rect 12897 13889 12909 13892
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 12989 13923 13047 13929
rect 12989 13889 13001 13923
rect 13035 13889 13047 13923
rect 12989 13883 13047 13889
rect 9217 13855 9275 13861
rect 9217 13821 9229 13855
rect 9263 13852 9275 13855
rect 9490 13852 9496 13864
rect 9263 13824 9496 13852
rect 9263 13821 9275 13824
rect 9217 13815 9275 13821
rect 9490 13812 9496 13824
rect 9548 13852 9554 13864
rect 9548 13824 9628 13852
rect 9548 13812 9554 13824
rect 9600 13793 9628 13824
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 11514 13852 11520 13864
rect 11112 13824 11520 13852
rect 11112 13812 11118 13824
rect 11514 13812 11520 13824
rect 11572 13812 11578 13864
rect 12158 13852 12164 13864
rect 11900 13824 12164 13852
rect 9585 13787 9643 13793
rect 9585 13753 9597 13787
rect 9631 13753 9643 13787
rect 11330 13784 11336 13796
rect 9585 13747 9643 13753
rect 9692 13756 11336 13784
rect 9692 13716 9720 13756
rect 11330 13744 11336 13756
rect 11388 13744 11394 13796
rect 11422 13744 11428 13796
rect 11480 13784 11486 13796
rect 11698 13784 11704 13796
rect 11480 13756 11704 13784
rect 11480 13744 11486 13756
rect 11698 13744 11704 13756
rect 11756 13744 11762 13796
rect 11900 13793 11928 13824
rect 12158 13812 12164 13824
rect 12216 13812 12222 13864
rect 13004 13852 13032 13883
rect 13170 13880 13176 13932
rect 13228 13920 13234 13932
rect 13265 13923 13323 13929
rect 13265 13920 13277 13923
rect 13228 13892 13277 13920
rect 13228 13880 13234 13892
rect 13265 13889 13277 13892
rect 13311 13889 13323 13923
rect 13265 13883 13323 13889
rect 13722 13880 13728 13932
rect 13780 13880 13786 13932
rect 14550 13880 14556 13932
rect 14608 13920 14614 13932
rect 14752 13920 14780 13960
rect 15105 13957 15117 13960
rect 15151 13957 15163 13991
rect 16298 13988 16304 14000
rect 15105 13951 15163 13957
rect 15304 13960 16304 13988
rect 14608 13892 14780 13920
rect 14829 13923 14887 13929
rect 14608 13880 14614 13892
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 15304 13920 15332 13960
rect 16298 13948 16304 13960
rect 16356 13948 16362 14000
rect 19886 13988 19892 14000
rect 18616 13960 19892 13988
rect 14875 13892 15332 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 13446 13852 13452 13864
rect 13004 13824 13452 13852
rect 13446 13812 13452 13824
rect 13504 13852 13510 13864
rect 13504 13824 14412 13852
rect 13504 13812 13510 13824
rect 11885 13787 11943 13793
rect 11885 13753 11897 13787
rect 11931 13753 11943 13787
rect 11885 13747 11943 13753
rect 12802 13744 12808 13796
rect 12860 13784 12866 13796
rect 14274 13784 14280 13796
rect 12860 13756 14280 13784
rect 12860 13744 12866 13756
rect 14274 13744 14280 13756
rect 14332 13744 14338 13796
rect 14384 13784 14412 13824
rect 15010 13812 15016 13864
rect 15068 13812 15074 13864
rect 15304 13852 15332 13892
rect 15381 13923 15439 13929
rect 15381 13889 15393 13923
rect 15427 13920 15439 13923
rect 15930 13920 15936 13932
rect 15427 13892 15936 13920
rect 15427 13889 15439 13892
rect 15381 13883 15439 13889
rect 15930 13880 15936 13892
rect 15988 13880 15994 13932
rect 16206 13880 16212 13932
rect 16264 13920 16270 13932
rect 16666 13920 16672 13932
rect 16264 13892 16672 13920
rect 16264 13880 16270 13892
rect 16666 13880 16672 13892
rect 16724 13880 16730 13932
rect 18616 13929 18644 13960
rect 19886 13948 19892 13960
rect 19944 13948 19950 14000
rect 20530 13948 20536 14000
rect 20588 13988 20594 14000
rect 21192 13988 21220 14019
rect 22370 13988 22376 14000
rect 20588 13960 21220 13988
rect 22204 13960 22376 13988
rect 20588 13948 20594 13960
rect 18601 13923 18659 13929
rect 18601 13889 18613 13923
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 18690 13880 18696 13932
rect 18748 13880 18754 13932
rect 18782 13880 18788 13932
rect 18840 13920 18846 13932
rect 18877 13923 18935 13929
rect 18877 13920 18889 13923
rect 18840 13892 18889 13920
rect 18840 13880 18846 13892
rect 18877 13889 18889 13892
rect 18923 13889 18935 13923
rect 18877 13883 18935 13889
rect 18966 13880 18972 13932
rect 19024 13920 19030 13932
rect 19061 13923 19119 13929
rect 19061 13920 19073 13923
rect 19024 13892 19073 13920
rect 19024 13880 19030 13892
rect 19061 13889 19073 13892
rect 19107 13889 19119 13923
rect 19061 13883 19119 13889
rect 20438 13880 20444 13932
rect 20496 13920 20502 13932
rect 20625 13923 20683 13929
rect 20625 13920 20637 13923
rect 20496 13892 20637 13920
rect 20496 13880 20502 13892
rect 20625 13889 20637 13892
rect 20671 13889 20683 13923
rect 20625 13883 20683 13889
rect 20901 13923 20959 13929
rect 20901 13889 20913 13923
rect 20947 13920 20959 13923
rect 21082 13920 21088 13932
rect 20947 13892 21088 13920
rect 20947 13889 20959 13892
rect 20901 13883 20959 13889
rect 21082 13880 21088 13892
rect 21140 13920 21146 13932
rect 21266 13920 21272 13932
rect 21140 13892 21272 13920
rect 21140 13880 21146 13892
rect 21266 13880 21272 13892
rect 21324 13880 21330 13932
rect 21358 13880 21364 13932
rect 21416 13880 21422 13932
rect 21450 13880 21456 13932
rect 21508 13880 21514 13932
rect 21726 13880 21732 13932
rect 21784 13920 21790 13932
rect 22204 13929 22232 13960
rect 22370 13948 22376 13960
rect 22428 13948 22434 14000
rect 23198 13948 23204 14000
rect 23256 13988 23262 14000
rect 23566 13988 23572 14000
rect 23256 13960 23572 13988
rect 23256 13948 23262 13960
rect 23566 13948 23572 13960
rect 23624 13988 23630 14000
rect 23845 13991 23903 13997
rect 23845 13988 23857 13991
rect 23624 13960 23857 13988
rect 23624 13948 23630 13960
rect 23845 13957 23857 13960
rect 23891 13957 23903 13991
rect 23845 13951 23903 13957
rect 23934 13948 23940 14000
rect 23992 13988 23998 14000
rect 23992 13960 24072 13988
rect 23992 13948 23998 13960
rect 22005 13923 22063 13929
rect 22005 13920 22017 13923
rect 21784 13892 22017 13920
rect 21784 13880 21790 13892
rect 22005 13889 22017 13892
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 22189 13923 22247 13929
rect 22189 13889 22201 13923
rect 22235 13889 22247 13923
rect 22189 13883 22247 13889
rect 22281 13923 22339 13929
rect 22281 13889 22293 13923
rect 22327 13889 22339 13923
rect 22281 13883 22339 13889
rect 15304 13824 15424 13852
rect 15286 13784 15292 13796
rect 14384 13756 15292 13784
rect 15286 13744 15292 13756
rect 15344 13744 15350 13796
rect 9147 13688 9720 13716
rect 10042 13676 10048 13728
rect 10100 13676 10106 13728
rect 10134 13676 10140 13728
rect 10192 13676 10198 13728
rect 10594 13676 10600 13728
rect 10652 13716 10658 13728
rect 11977 13719 12035 13725
rect 11977 13716 11989 13719
rect 10652 13688 11989 13716
rect 10652 13676 10658 13688
rect 11977 13685 11989 13688
rect 12023 13685 12035 13719
rect 11977 13679 12035 13685
rect 12989 13719 13047 13725
rect 12989 13685 13001 13719
rect 13035 13716 13047 13719
rect 14734 13716 14740 13728
rect 13035 13688 14740 13716
rect 13035 13685 13047 13688
rect 12989 13679 13047 13685
rect 14734 13676 14740 13688
rect 14792 13676 14798 13728
rect 14918 13676 14924 13728
rect 14976 13676 14982 13728
rect 15197 13719 15255 13725
rect 15197 13685 15209 13719
rect 15243 13716 15255 13719
rect 15396 13716 15424 13824
rect 16022 13812 16028 13864
rect 16080 13852 16086 13864
rect 20714 13852 20720 13864
rect 16080 13824 20720 13852
rect 16080 13812 16086 13824
rect 20714 13812 20720 13824
rect 20772 13812 20778 13864
rect 20809 13855 20867 13861
rect 20809 13821 20821 13855
rect 20855 13852 20867 13855
rect 22094 13852 22100 13864
rect 20855 13824 22100 13852
rect 20855 13821 20867 13824
rect 20809 13815 20867 13821
rect 22094 13812 22100 13824
rect 22152 13812 22158 13864
rect 15838 13744 15844 13796
rect 15896 13784 15902 13796
rect 16298 13784 16304 13796
rect 15896 13756 16304 13784
rect 15896 13744 15902 13756
rect 16298 13744 16304 13756
rect 16356 13744 16362 13796
rect 18230 13744 18236 13796
rect 18288 13784 18294 13796
rect 18288 13756 18552 13784
rect 18288 13744 18294 13756
rect 15243 13688 15424 13716
rect 15243 13685 15255 13688
rect 15197 13679 15255 13685
rect 18322 13676 18328 13728
rect 18380 13676 18386 13728
rect 18524 13725 18552 13756
rect 20346 13744 20352 13796
rect 20404 13784 20410 13796
rect 21634 13784 21640 13796
rect 20404 13756 21640 13784
rect 20404 13744 20410 13756
rect 21634 13744 21640 13756
rect 21692 13744 21698 13796
rect 22289 13784 22317 13883
rect 22462 13880 22468 13932
rect 22520 13920 22526 13932
rect 22557 13923 22615 13929
rect 22557 13920 22569 13923
rect 22520 13892 22569 13920
rect 22520 13880 22526 13892
rect 22557 13889 22569 13892
rect 22603 13889 22615 13923
rect 22557 13883 22615 13889
rect 22646 13812 22652 13864
rect 22704 13852 22710 13864
rect 23106 13852 23112 13864
rect 22704 13824 23112 13852
rect 22704 13812 22710 13824
rect 23106 13812 23112 13824
rect 23164 13812 23170 13864
rect 23934 13812 23940 13864
rect 23992 13812 23998 13864
rect 24044 13852 24072 13960
rect 24136 13929 24164 14028
rect 24305 14025 24317 14059
rect 24351 14056 24363 14059
rect 25222 14056 25228 14068
rect 24351 14028 25228 14056
rect 24351 14025 24363 14028
rect 24305 14019 24363 14025
rect 25222 14016 25228 14028
rect 25280 14056 25286 14068
rect 25280 14028 26924 14056
rect 25280 14016 25286 14028
rect 26418 13948 26424 14000
rect 26476 13988 26482 14000
rect 26786 13988 26792 14000
rect 26476 13960 26792 13988
rect 26476 13948 26482 13960
rect 26786 13948 26792 13960
rect 26844 13948 26850 14000
rect 26896 13988 26924 14028
rect 26970 14016 26976 14068
rect 27028 14056 27034 14068
rect 27893 14059 27951 14065
rect 27893 14056 27905 14059
rect 27028 14028 27905 14056
rect 27028 14016 27034 14028
rect 27893 14025 27905 14028
rect 27939 14056 27951 14059
rect 28810 14056 28816 14068
rect 27939 14028 28816 14056
rect 27939 14025 27951 14028
rect 27893 14019 27951 14025
rect 28810 14016 28816 14028
rect 28868 14016 28874 14068
rect 30101 14059 30159 14065
rect 30101 14025 30113 14059
rect 30147 14056 30159 14059
rect 30926 14056 30932 14068
rect 30147 14028 30932 14056
rect 30147 14025 30159 14028
rect 30101 14019 30159 14025
rect 30926 14016 30932 14028
rect 30984 14016 30990 14068
rect 31941 14059 31999 14065
rect 31941 14025 31953 14059
rect 31987 14056 31999 14059
rect 32214 14056 32220 14068
rect 31987 14028 32220 14056
rect 31987 14025 31999 14028
rect 31941 14019 31999 14025
rect 32214 14016 32220 14028
rect 32272 14016 32278 14068
rect 32398 14016 32404 14068
rect 32456 14016 32462 14068
rect 26896 13960 27200 13988
rect 24121 13923 24179 13929
rect 24121 13889 24133 13923
rect 24167 13920 24179 13923
rect 24210 13920 24216 13932
rect 24167 13892 24216 13920
rect 24167 13889 24179 13892
rect 24121 13883 24179 13889
rect 24210 13880 24216 13892
rect 24268 13880 24274 13932
rect 26234 13880 26240 13932
rect 26292 13920 26298 13932
rect 26329 13923 26387 13929
rect 26329 13920 26341 13923
rect 26292 13892 26341 13920
rect 26292 13880 26298 13892
rect 26329 13889 26341 13892
rect 26375 13889 26387 13923
rect 26329 13883 26387 13889
rect 26602 13880 26608 13932
rect 26660 13880 26666 13932
rect 26878 13920 26884 13932
rect 26804 13892 26884 13920
rect 24044 13824 24624 13852
rect 24596 13796 24624 13824
rect 26510 13812 26516 13864
rect 26568 13812 26574 13864
rect 21836 13756 22317 13784
rect 21836 13728 21864 13756
rect 22922 13744 22928 13796
rect 22980 13744 22986 13796
rect 24578 13744 24584 13796
rect 24636 13744 24642 13796
rect 18509 13719 18567 13725
rect 18509 13685 18521 13719
rect 18555 13685 18567 13719
rect 18509 13679 18567 13685
rect 20070 13676 20076 13728
rect 20128 13716 20134 13728
rect 20530 13716 20536 13728
rect 20128 13688 20536 13716
rect 20128 13676 20134 13688
rect 20530 13676 20536 13688
rect 20588 13676 20594 13728
rect 20714 13676 20720 13728
rect 20772 13676 20778 13728
rect 21818 13676 21824 13728
rect 21876 13676 21882 13728
rect 22278 13676 22284 13728
rect 22336 13676 22342 13728
rect 22462 13676 22468 13728
rect 22520 13676 22526 13728
rect 22554 13676 22560 13728
rect 22612 13676 22618 13728
rect 24118 13676 24124 13728
rect 24176 13676 24182 13728
rect 26234 13676 26240 13728
rect 26292 13716 26298 13728
rect 26329 13719 26387 13725
rect 26329 13716 26341 13719
rect 26292 13688 26341 13716
rect 26292 13676 26298 13688
rect 26329 13685 26341 13688
rect 26375 13716 26387 13719
rect 26694 13716 26700 13728
rect 26375 13688 26700 13716
rect 26375 13685 26387 13688
rect 26329 13679 26387 13685
rect 26694 13676 26700 13688
rect 26752 13676 26758 13728
rect 26804 13725 26832 13892
rect 26878 13880 26884 13892
rect 26936 13920 26942 13932
rect 27172 13929 27200 13960
rect 27430 13948 27436 14000
rect 27488 13988 27494 14000
rect 27488 13960 27660 13988
rect 27488 13948 27494 13960
rect 26973 13923 27031 13929
rect 26973 13920 26985 13923
rect 26936 13892 26985 13920
rect 26936 13880 26942 13892
rect 26973 13889 26985 13892
rect 27019 13889 27031 13923
rect 26973 13883 27031 13889
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13889 27215 13923
rect 27157 13883 27215 13889
rect 27246 13880 27252 13932
rect 27304 13880 27310 13932
rect 27632 13929 27660 13960
rect 27798 13948 27804 14000
rect 27856 13988 27862 14000
rect 27856 13960 30236 13988
rect 27856 13948 27862 13960
rect 27525 13923 27583 13929
rect 27525 13889 27537 13923
rect 27571 13889 27583 13923
rect 27525 13883 27583 13889
rect 27617 13923 27675 13929
rect 27617 13889 27629 13923
rect 27663 13889 27675 13923
rect 29641 13923 29699 13929
rect 29641 13920 29653 13923
rect 27617 13883 27675 13889
rect 29472 13892 29653 13920
rect 27264 13852 27292 13880
rect 26988 13824 27292 13852
rect 26988 13796 27016 13824
rect 27430 13812 27436 13864
rect 27488 13852 27494 13864
rect 27540 13852 27568 13883
rect 27488 13824 27568 13852
rect 27488 13812 27494 13824
rect 29270 13812 29276 13864
rect 29328 13852 29334 13864
rect 29472 13861 29500 13892
rect 29641 13889 29653 13892
rect 29687 13889 29699 13923
rect 29641 13883 29699 13889
rect 29822 13880 29828 13932
rect 29880 13880 29886 13932
rect 30208 13929 30236 13960
rect 29917 13923 29975 13929
rect 29917 13889 29929 13923
rect 29963 13889 29975 13923
rect 29917 13883 29975 13889
rect 30193 13923 30251 13929
rect 30193 13889 30205 13923
rect 30239 13889 30251 13923
rect 30193 13883 30251 13889
rect 29457 13855 29515 13861
rect 29457 13852 29469 13855
rect 29328 13824 29469 13852
rect 29328 13812 29334 13824
rect 29457 13821 29469 13824
rect 29503 13821 29515 13855
rect 29932 13852 29960 13883
rect 30282 13880 30288 13932
rect 30340 13920 30346 13932
rect 30377 13923 30435 13929
rect 30377 13920 30389 13923
rect 30340 13892 30389 13920
rect 30340 13880 30346 13892
rect 30377 13889 30389 13892
rect 30423 13889 30435 13923
rect 30377 13883 30435 13889
rect 30828 13923 30886 13929
rect 30828 13889 30840 13923
rect 30874 13920 30886 13923
rect 31754 13920 31760 13932
rect 30874 13892 31760 13920
rect 30874 13889 30886 13892
rect 30828 13883 30886 13889
rect 31754 13880 31760 13892
rect 31812 13880 31818 13932
rect 32122 13880 32128 13932
rect 32180 13920 32186 13932
rect 32217 13923 32275 13929
rect 32217 13920 32229 13923
rect 32180 13892 32229 13920
rect 32180 13880 32186 13892
rect 32217 13889 32229 13892
rect 32263 13889 32275 13923
rect 32217 13883 32275 13889
rect 30006 13852 30012 13864
rect 29457 13815 29515 13821
rect 29564 13824 30012 13852
rect 26970 13744 26976 13796
rect 27028 13744 27034 13796
rect 28258 13744 28264 13796
rect 28316 13784 28322 13796
rect 28442 13784 28448 13796
rect 28316 13756 28448 13784
rect 28316 13744 28322 13756
rect 28442 13744 28448 13756
rect 28500 13744 28506 13796
rect 29178 13744 29184 13796
rect 29236 13784 29242 13796
rect 29564 13784 29592 13824
rect 30006 13812 30012 13824
rect 30064 13812 30070 13864
rect 30558 13812 30564 13864
rect 30616 13812 30622 13864
rect 30285 13787 30343 13793
rect 30285 13784 30297 13787
rect 29236 13756 29592 13784
rect 29932 13756 30297 13784
rect 29236 13744 29242 13756
rect 26789 13719 26847 13725
rect 26789 13685 26801 13719
rect 26835 13685 26847 13719
rect 26789 13679 26847 13685
rect 26878 13676 26884 13728
rect 26936 13716 26942 13728
rect 27154 13716 27160 13728
rect 26936 13688 27160 13716
rect 26936 13676 26942 13688
rect 27154 13676 27160 13688
rect 27212 13676 27218 13728
rect 27430 13676 27436 13728
rect 27488 13676 27494 13728
rect 27706 13676 27712 13728
rect 27764 13676 27770 13728
rect 29932 13725 29960 13756
rect 30285 13753 30297 13756
rect 30331 13753 30343 13787
rect 30285 13747 30343 13753
rect 29917 13719 29975 13725
rect 29917 13685 29929 13719
rect 29963 13685 29975 13719
rect 29917 13679 29975 13685
rect 1104 13626 32844 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 32844 13626
rect 1104 13552 32844 13574
rect 2317 13515 2375 13521
rect 2317 13481 2329 13515
rect 2363 13512 2375 13515
rect 3234 13512 3240 13524
rect 2363 13484 3240 13512
rect 2363 13481 2375 13484
rect 2317 13475 2375 13481
rect 3234 13472 3240 13484
rect 3292 13472 3298 13524
rect 3605 13515 3663 13521
rect 3605 13481 3617 13515
rect 3651 13512 3663 13515
rect 3970 13512 3976 13524
rect 3651 13484 3976 13512
rect 3651 13481 3663 13484
rect 3605 13475 3663 13481
rect 3970 13472 3976 13484
rect 4028 13472 4034 13524
rect 4522 13472 4528 13524
rect 4580 13512 4586 13524
rect 4580 13484 6500 13512
rect 4580 13472 4586 13484
rect 566 13404 572 13456
rect 624 13444 630 13456
rect 3418 13444 3424 13456
rect 624 13416 3424 13444
rect 624 13404 630 13416
rect 3418 13404 3424 13416
rect 3476 13404 3482 13456
rect 4706 13444 4712 13456
rect 3804 13416 4712 13444
rect 2774 13336 2780 13388
rect 2832 13376 2838 13388
rect 3804 13376 3832 13416
rect 4706 13404 4712 13416
rect 4764 13404 4770 13456
rect 4982 13404 4988 13456
rect 5040 13444 5046 13456
rect 6362 13444 6368 13456
rect 5040 13416 6368 13444
rect 5040 13404 5046 13416
rect 6362 13404 6368 13416
rect 6420 13404 6426 13456
rect 2832 13348 3832 13376
rect 2832 13336 2838 13348
rect 2498 13268 2504 13320
rect 2556 13268 2562 13320
rect 2866 13268 2872 13320
rect 2924 13308 2930 13320
rect 3421 13311 3479 13317
rect 3421 13308 3433 13311
rect 2924 13280 3433 13308
rect 2924 13268 2930 13280
rect 3421 13277 3433 13280
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 3694 13268 3700 13320
rect 3752 13268 3758 13320
rect 3804 13317 3832 13348
rect 3896 13348 4200 13376
rect 3789 13311 3847 13317
rect 3789 13277 3801 13311
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 2685 13243 2743 13249
rect 2685 13209 2697 13243
rect 2731 13240 2743 13243
rect 2958 13240 2964 13252
rect 2731 13212 2964 13240
rect 2731 13209 2743 13212
rect 2685 13203 2743 13209
rect 2958 13200 2964 13212
rect 3016 13200 3022 13252
rect 3712 13240 3740 13268
rect 3896 13240 3924 13348
rect 3970 13268 3976 13320
rect 4028 13268 4034 13320
rect 4172 13317 4200 13348
rect 4430 13336 4436 13388
rect 4488 13376 4494 13388
rect 6181 13379 6239 13385
rect 6181 13376 6193 13379
rect 4488 13348 6193 13376
rect 4488 13336 4494 13348
rect 6181 13345 6193 13348
rect 6227 13345 6239 13379
rect 6472 13376 6500 13484
rect 7834 13472 7840 13524
rect 7892 13512 7898 13524
rect 8113 13515 8171 13521
rect 8113 13512 8125 13515
rect 7892 13484 8125 13512
rect 7892 13472 7898 13484
rect 8113 13481 8125 13484
rect 8159 13481 8171 13515
rect 8113 13475 8171 13481
rect 8754 13472 8760 13524
rect 8812 13512 8818 13524
rect 9582 13512 9588 13524
rect 8812 13484 9588 13512
rect 8812 13472 8818 13484
rect 9582 13472 9588 13484
rect 9640 13472 9646 13524
rect 9766 13472 9772 13524
rect 9824 13512 9830 13524
rect 10226 13512 10232 13524
rect 9824 13484 10232 13512
rect 9824 13472 9830 13484
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 11238 13472 11244 13524
rect 11296 13472 11302 13524
rect 11422 13472 11428 13524
rect 11480 13512 11486 13524
rect 12066 13512 12072 13524
rect 11480 13484 12072 13512
rect 11480 13472 11486 13484
rect 12066 13472 12072 13484
rect 12124 13472 12130 13524
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 13265 13515 13323 13521
rect 12492 13484 12756 13512
rect 12492 13472 12498 13484
rect 7282 13453 7288 13456
rect 7266 13447 7288 13453
rect 7266 13413 7278 13447
rect 7266 13407 7288 13413
rect 7282 13404 7288 13407
rect 7340 13404 7346 13456
rect 7377 13447 7435 13453
rect 7377 13413 7389 13447
rect 7423 13444 7435 13447
rect 7742 13444 7748 13456
rect 7423 13416 7748 13444
rect 7423 13413 7435 13416
rect 7377 13407 7435 13413
rect 7742 13404 7748 13416
rect 7800 13404 7806 13456
rect 12526 13444 12532 13456
rect 7852 13416 12532 13444
rect 7466 13376 7472 13388
rect 6472 13348 7472 13376
rect 6181 13339 6239 13345
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 7650 13336 7656 13388
rect 7708 13376 7714 13388
rect 7852 13376 7880 13416
rect 12526 13404 12532 13416
rect 12584 13404 12590 13456
rect 12728 13453 12756 13484
rect 13265 13481 13277 13515
rect 13311 13512 13323 13515
rect 13630 13512 13636 13524
rect 13311 13484 13636 13512
rect 13311 13481 13323 13484
rect 13265 13475 13323 13481
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 14461 13515 14519 13521
rect 14461 13481 14473 13515
rect 14507 13512 14519 13515
rect 14550 13512 14556 13524
rect 14507 13484 14556 13512
rect 14507 13481 14519 13484
rect 14461 13475 14519 13481
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 17770 13472 17776 13524
rect 17828 13512 17834 13524
rect 18141 13515 18199 13521
rect 17828 13484 18000 13512
rect 17828 13472 17834 13484
rect 12713 13447 12771 13453
rect 12713 13413 12725 13447
rect 12759 13444 12771 13447
rect 12759 13416 17908 13444
rect 12759 13413 12771 13416
rect 12713 13407 12771 13413
rect 10134 13376 10140 13388
rect 7708 13348 7880 13376
rect 8404 13348 10140 13376
rect 7708 13336 7714 13348
rect 4157 13311 4215 13317
rect 4157 13277 4169 13311
rect 4203 13277 4215 13311
rect 4157 13271 4215 13277
rect 4338 13268 4344 13320
rect 4396 13308 4402 13320
rect 4396 13280 4568 13308
rect 4396 13268 4402 13280
rect 3712 13212 3924 13240
rect 4065 13243 4123 13249
rect 4065 13209 4077 13243
rect 4111 13240 4123 13243
rect 4540 13240 4568 13280
rect 4614 13268 4620 13320
rect 4672 13308 4678 13320
rect 4672 13280 5580 13308
rect 4672 13268 4678 13280
rect 4890 13240 4896 13252
rect 4111 13212 4476 13240
rect 4540 13212 4896 13240
rect 4111 13209 4123 13212
rect 4065 13203 4123 13209
rect 3694 13132 3700 13184
rect 3752 13172 3758 13184
rect 4264 13172 4292 13212
rect 3752 13144 4292 13172
rect 3752 13132 3758 13144
rect 4338 13132 4344 13184
rect 4396 13132 4402 13184
rect 4448 13181 4476 13212
rect 4890 13200 4896 13212
rect 4948 13200 4954 13252
rect 4433 13175 4491 13181
rect 4433 13141 4445 13175
rect 4479 13141 4491 13175
rect 4433 13135 4491 13141
rect 4614 13132 4620 13184
rect 4672 13172 4678 13184
rect 5442 13172 5448 13184
rect 4672 13144 5448 13172
rect 4672 13132 4678 13144
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 5552 13172 5580 13280
rect 5810 13268 5816 13320
rect 5868 13268 5874 13320
rect 5902 13268 5908 13320
rect 5960 13308 5966 13320
rect 6089 13311 6147 13317
rect 6089 13308 6101 13311
rect 5960 13280 6101 13308
rect 5960 13268 5966 13280
rect 6089 13277 6101 13280
rect 6135 13277 6147 13311
rect 6089 13271 6147 13277
rect 6270 13268 6276 13320
rect 6328 13308 6334 13320
rect 6457 13311 6515 13317
rect 6457 13308 6469 13311
rect 6328 13280 6469 13308
rect 6328 13268 6334 13280
rect 6457 13277 6469 13280
rect 6503 13277 6515 13311
rect 8404 13308 8432 13348
rect 6457 13271 6515 13277
rect 6886 13280 8432 13308
rect 5626 13200 5632 13252
rect 5684 13240 5690 13252
rect 6886 13240 6914 13280
rect 8478 13268 8484 13320
rect 8536 13308 8542 13320
rect 9324 13317 9352 13348
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 12802 13376 12808 13388
rect 11348 13348 12808 13376
rect 9033 13311 9091 13317
rect 9033 13308 9045 13311
rect 8536 13280 9045 13308
rect 8536 13268 8542 13280
rect 9033 13277 9045 13280
rect 9079 13277 9091 13311
rect 9033 13271 9091 13277
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13277 9367 13311
rect 9309 13271 9367 13277
rect 9401 13311 9459 13317
rect 9401 13277 9413 13311
rect 9447 13308 9459 13311
rect 9447 13280 9674 13308
rect 9447 13277 9459 13280
rect 9401 13271 9459 13277
rect 5684 13212 6914 13240
rect 7101 13243 7159 13249
rect 5684 13200 5690 13212
rect 7101 13209 7113 13243
rect 7147 13240 7159 13243
rect 7374 13240 7380 13252
rect 7147 13212 7380 13240
rect 7147 13209 7159 13212
rect 7101 13203 7159 13209
rect 7374 13200 7380 13212
rect 7432 13240 7438 13252
rect 7650 13240 7656 13252
rect 7432 13212 7656 13240
rect 7432 13200 7438 13212
rect 7650 13200 7656 13212
rect 7708 13200 7714 13252
rect 7834 13200 7840 13252
rect 7892 13200 7898 13252
rect 8021 13243 8079 13249
rect 8021 13209 8033 13243
rect 8067 13209 8079 13243
rect 8021 13203 8079 13209
rect 6178 13172 6184 13184
rect 5552 13144 6184 13172
rect 6178 13132 6184 13144
rect 6236 13132 6242 13184
rect 6730 13132 6736 13184
rect 6788 13172 6794 13184
rect 8036 13172 8064 13203
rect 8846 13200 8852 13252
rect 8904 13240 8910 13252
rect 9217 13243 9275 13249
rect 9217 13240 9229 13243
rect 8904 13212 9229 13240
rect 8904 13200 8910 13212
rect 9217 13209 9229 13212
rect 9263 13209 9275 13243
rect 9646 13240 9674 13280
rect 9858 13268 9864 13320
rect 9916 13308 9922 13320
rect 11348 13308 11376 13348
rect 12802 13336 12808 13348
rect 12860 13336 12866 13388
rect 12986 13336 12992 13388
rect 13044 13336 13050 13388
rect 13078 13336 13084 13388
rect 13136 13336 13142 13388
rect 13538 13376 13544 13388
rect 13188 13348 13544 13376
rect 9916 13280 11376 13308
rect 11425 13311 11483 13317
rect 9916 13268 9922 13280
rect 11425 13277 11437 13311
rect 11471 13308 11483 13311
rect 11698 13308 11704 13320
rect 11471 13280 11704 13308
rect 11471 13277 11483 13280
rect 11425 13271 11483 13277
rect 11698 13268 11704 13280
rect 11756 13268 11762 13320
rect 11882 13268 11888 13320
rect 11940 13308 11946 13320
rect 12250 13308 12256 13320
rect 11940 13280 12256 13308
rect 11940 13268 11946 13280
rect 12250 13268 12256 13280
rect 12308 13268 12314 13320
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13308 12955 13311
rect 13004 13308 13032 13336
rect 12943 13280 13032 13308
rect 12943 13277 12955 13280
rect 12897 13271 12955 13277
rect 10134 13240 10140 13252
rect 9646 13212 10140 13240
rect 9217 13203 9275 13209
rect 10134 13200 10140 13212
rect 10192 13200 10198 13252
rect 10962 13200 10968 13252
rect 11020 13240 11026 13252
rect 12989 13243 13047 13249
rect 11020 13212 11192 13240
rect 11020 13200 11026 13212
rect 6788 13144 8064 13172
rect 6788 13132 6794 13144
rect 8202 13132 8208 13184
rect 8260 13172 8266 13184
rect 10870 13172 10876 13184
rect 8260 13144 10876 13172
rect 8260 13132 8266 13144
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 11164 13172 11192 13212
rect 12989 13209 13001 13243
rect 13035 13240 13047 13243
rect 13078 13240 13084 13252
rect 13035 13212 13084 13240
rect 13035 13209 13047 13212
rect 12989 13203 13047 13209
rect 13078 13200 13084 13212
rect 13136 13240 13142 13252
rect 13188 13240 13216 13348
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 13262 13268 13268 13320
rect 13320 13268 13326 13320
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 13372 13280 14289 13308
rect 13136 13212 13216 13240
rect 13136 13200 13142 13212
rect 13372 13172 13400 13280
rect 14277 13277 14289 13280
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 14734 13268 14740 13320
rect 14792 13308 14798 13320
rect 15105 13311 15163 13317
rect 15105 13308 15117 13311
rect 14792 13280 15117 13308
rect 14792 13268 14798 13280
rect 15105 13277 15117 13280
rect 15151 13277 15163 13311
rect 15105 13271 15163 13277
rect 15286 13268 15292 13320
rect 15344 13268 15350 13320
rect 15838 13268 15844 13320
rect 15896 13308 15902 13320
rect 17218 13308 17224 13320
rect 15896 13280 17224 13308
rect 15896 13268 15902 13280
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 14090 13200 14096 13252
rect 14148 13200 14154 13252
rect 15473 13243 15531 13249
rect 15473 13209 15485 13243
rect 15519 13240 15531 13243
rect 15930 13240 15936 13252
rect 15519 13212 15936 13240
rect 15519 13209 15531 13212
rect 15473 13203 15531 13209
rect 15930 13200 15936 13212
rect 15988 13200 15994 13252
rect 16666 13200 16672 13252
rect 16724 13240 16730 13252
rect 17586 13240 17592 13252
rect 16724 13212 17592 13240
rect 16724 13200 16730 13212
rect 17586 13200 17592 13212
rect 17644 13200 17650 13252
rect 17880 13249 17908 13416
rect 17972 13385 18000 13484
rect 18141 13481 18153 13515
rect 18187 13481 18199 13515
rect 18141 13475 18199 13481
rect 18325 13515 18383 13521
rect 18325 13481 18337 13515
rect 18371 13512 18383 13515
rect 18690 13512 18696 13524
rect 18371 13484 18696 13512
rect 18371 13481 18383 13484
rect 18325 13475 18383 13481
rect 18156 13444 18184 13475
rect 18690 13472 18696 13484
rect 18748 13472 18754 13524
rect 20070 13472 20076 13524
rect 20128 13512 20134 13524
rect 20441 13515 20499 13521
rect 20441 13512 20453 13515
rect 20128 13484 20453 13512
rect 20128 13472 20134 13484
rect 20441 13481 20453 13484
rect 20487 13481 20499 13515
rect 20993 13515 21051 13521
rect 20993 13512 21005 13515
rect 20441 13475 20499 13481
rect 20548 13484 21005 13512
rect 18598 13444 18604 13456
rect 18156 13416 18604 13444
rect 18598 13404 18604 13416
rect 18656 13404 18662 13456
rect 20548 13444 20576 13484
rect 20993 13481 21005 13484
rect 21039 13481 21051 13515
rect 20993 13475 21051 13481
rect 22554 13472 22560 13524
rect 22612 13512 22618 13524
rect 22922 13512 22928 13524
rect 22612 13484 22928 13512
rect 22612 13472 22618 13484
rect 22922 13472 22928 13484
rect 22980 13472 22986 13524
rect 28261 13515 28319 13521
rect 28261 13481 28273 13515
rect 28307 13512 28319 13515
rect 28350 13512 28356 13524
rect 28307 13484 28356 13512
rect 28307 13481 28319 13484
rect 28261 13475 28319 13481
rect 28350 13472 28356 13484
rect 28408 13472 28414 13524
rect 28626 13472 28632 13524
rect 28684 13512 28690 13524
rect 28721 13515 28779 13521
rect 28721 13512 28733 13515
rect 28684 13484 28733 13512
rect 28684 13472 28690 13484
rect 28721 13481 28733 13484
rect 28767 13481 28779 13515
rect 28721 13475 28779 13481
rect 29273 13515 29331 13521
rect 29273 13481 29285 13515
rect 29319 13512 29331 13515
rect 30374 13512 30380 13524
rect 29319 13484 30380 13512
rect 29319 13481 29331 13484
rect 29273 13475 29331 13481
rect 30374 13472 30380 13484
rect 30432 13472 30438 13524
rect 31481 13515 31539 13521
rect 31481 13481 31493 13515
rect 31527 13512 31539 13515
rect 31754 13512 31760 13524
rect 31527 13484 31760 13512
rect 31527 13481 31539 13484
rect 31481 13475 31539 13481
rect 31754 13472 31760 13484
rect 31812 13472 31818 13524
rect 20088 13416 20576 13444
rect 20901 13447 20959 13453
rect 17957 13379 18015 13385
rect 17957 13345 17969 13379
rect 18003 13345 18015 13379
rect 17957 13339 18015 13345
rect 18141 13311 18199 13317
rect 18141 13277 18153 13311
rect 18187 13308 18199 13311
rect 18966 13308 18972 13320
rect 18187 13280 18972 13308
rect 18187 13277 18199 13280
rect 18141 13271 18199 13277
rect 18966 13268 18972 13280
rect 19024 13268 19030 13320
rect 19518 13268 19524 13320
rect 19576 13308 19582 13320
rect 19794 13308 19800 13320
rect 19576 13280 19800 13308
rect 19576 13268 19582 13280
rect 19794 13268 19800 13280
rect 19852 13268 19858 13320
rect 17865 13243 17923 13249
rect 17865 13209 17877 13243
rect 17911 13240 17923 13243
rect 20088 13240 20116 13416
rect 20901 13413 20913 13447
rect 20947 13444 20959 13447
rect 21266 13444 21272 13456
rect 20947 13416 21272 13444
rect 20947 13413 20959 13416
rect 20901 13407 20959 13413
rect 21266 13404 21272 13416
rect 21324 13404 21330 13456
rect 21634 13404 21640 13456
rect 21692 13444 21698 13456
rect 22370 13444 22376 13456
rect 21692 13416 22376 13444
rect 21692 13404 21698 13416
rect 22370 13404 22376 13416
rect 22428 13444 22434 13456
rect 25774 13444 25780 13456
rect 22428 13416 25780 13444
rect 22428 13404 22434 13416
rect 25774 13404 25780 13416
rect 25832 13404 25838 13456
rect 26421 13447 26479 13453
rect 26421 13413 26433 13447
rect 26467 13444 26479 13447
rect 28445 13447 28503 13453
rect 26467 13416 27936 13444
rect 26467 13413 26479 13416
rect 26421 13407 26479 13413
rect 20346 13336 20352 13388
rect 20404 13376 20410 13388
rect 20533 13379 20591 13385
rect 20533 13376 20545 13379
rect 20404 13348 20545 13376
rect 20404 13336 20410 13348
rect 20533 13345 20545 13348
rect 20579 13345 20591 13379
rect 20533 13339 20591 13345
rect 20640 13348 21680 13376
rect 20165 13311 20223 13317
rect 20165 13277 20177 13311
rect 20211 13308 20223 13311
rect 20640 13308 20668 13348
rect 20211 13280 20668 13308
rect 20717 13311 20775 13317
rect 20211 13277 20223 13280
rect 20165 13271 20223 13277
rect 20717 13277 20729 13311
rect 20763 13277 20775 13311
rect 20717 13271 20775 13277
rect 20441 13243 20499 13249
rect 20441 13240 20453 13243
rect 17911 13212 20453 13240
rect 17911 13209 17923 13212
rect 17865 13203 17923 13209
rect 20441 13209 20453 13212
rect 20487 13209 20499 13243
rect 20441 13203 20499 13209
rect 20530 13200 20536 13252
rect 20588 13240 20594 13252
rect 20732 13240 20760 13271
rect 20806 13268 20812 13320
rect 20864 13308 20870 13320
rect 20993 13311 21051 13317
rect 20993 13308 21005 13311
rect 20864 13280 21005 13308
rect 20864 13268 20870 13280
rect 20993 13277 21005 13280
rect 21039 13277 21051 13311
rect 20993 13271 21051 13277
rect 21177 13311 21235 13317
rect 21177 13277 21189 13311
rect 21223 13308 21235 13311
rect 21358 13308 21364 13320
rect 21223 13280 21364 13308
rect 21223 13277 21235 13280
rect 21177 13271 21235 13277
rect 20588 13212 20760 13240
rect 20588 13200 20594 13212
rect 11164 13144 13400 13172
rect 13446 13132 13452 13184
rect 13504 13132 13510 13184
rect 13906 13132 13912 13184
rect 13964 13172 13970 13184
rect 14366 13172 14372 13184
rect 13964 13144 14372 13172
rect 13964 13132 13970 13144
rect 14366 13132 14372 13144
rect 14424 13132 14430 13184
rect 14918 13132 14924 13184
rect 14976 13172 14982 13184
rect 18690 13172 18696 13184
rect 14976 13144 18696 13172
rect 14976 13132 14982 13144
rect 18690 13132 18696 13144
rect 18748 13132 18754 13184
rect 20349 13175 20407 13181
rect 20349 13141 20361 13175
rect 20395 13172 20407 13175
rect 21192 13172 21220 13271
rect 21358 13268 21364 13280
rect 21416 13268 21422 13320
rect 21652 13308 21680 13348
rect 21726 13336 21732 13388
rect 21784 13376 21790 13388
rect 24854 13376 24860 13388
rect 21784 13348 24860 13376
rect 21784 13336 21790 13348
rect 24854 13336 24860 13348
rect 24912 13336 24918 13388
rect 24118 13308 24124 13320
rect 21652 13280 24124 13308
rect 24118 13268 24124 13280
rect 24176 13268 24182 13320
rect 24394 13268 24400 13320
rect 24452 13268 24458 13320
rect 25792 13308 25820 13404
rect 26145 13379 26203 13385
rect 26145 13345 26157 13379
rect 26191 13376 26203 13379
rect 26191 13348 27752 13376
rect 26191 13345 26203 13348
rect 26145 13339 26203 13345
rect 26237 13311 26295 13317
rect 26237 13308 26249 13311
rect 25792 13280 26249 13308
rect 26237 13277 26249 13280
rect 26283 13277 26295 13311
rect 26237 13271 26295 13277
rect 26421 13311 26479 13317
rect 26421 13277 26433 13311
rect 26467 13277 26479 13311
rect 26421 13271 26479 13277
rect 21266 13200 21272 13252
rect 21324 13240 21330 13252
rect 21324 13212 22317 13240
rect 21324 13200 21330 13212
rect 20395 13144 21220 13172
rect 21361 13175 21419 13181
rect 20395 13141 20407 13144
rect 20349 13135 20407 13141
rect 21361 13141 21373 13175
rect 21407 13172 21419 13175
rect 21542 13172 21548 13184
rect 21407 13144 21548 13172
rect 21407 13141 21419 13144
rect 21361 13135 21419 13141
rect 21542 13132 21548 13144
rect 21600 13132 21606 13184
rect 22289 13172 22317 13212
rect 22370 13200 22376 13252
rect 22428 13240 22434 13252
rect 26050 13240 26056 13252
rect 22428 13212 26056 13240
rect 22428 13200 22434 13212
rect 26050 13200 26056 13212
rect 26108 13200 26114 13252
rect 23106 13172 23112 13184
rect 22289 13144 23112 13172
rect 23106 13132 23112 13144
rect 23164 13132 23170 13184
rect 24578 13132 24584 13184
rect 24636 13172 24642 13184
rect 26436 13172 26464 13271
rect 27724 13240 27752 13348
rect 27798 13268 27804 13320
rect 27856 13268 27862 13320
rect 27908 13317 27936 13416
rect 28445 13413 28457 13447
rect 28491 13444 28503 13447
rect 28813 13447 28871 13453
rect 28813 13444 28825 13447
rect 28491 13416 28825 13444
rect 28491 13413 28503 13416
rect 28445 13407 28503 13413
rect 28813 13413 28825 13416
rect 28859 13413 28871 13447
rect 28813 13407 28871 13413
rect 29454 13404 29460 13456
rect 29512 13444 29518 13456
rect 29914 13444 29920 13456
rect 29512 13416 29920 13444
rect 29512 13404 29518 13416
rect 29914 13404 29920 13416
rect 29972 13404 29978 13456
rect 30558 13376 30564 13388
rect 28828 13348 30564 13376
rect 27893 13311 27951 13317
rect 27893 13277 27905 13311
rect 27939 13277 27951 13311
rect 27893 13271 27951 13277
rect 28261 13311 28319 13317
rect 28261 13277 28273 13311
rect 28307 13308 28319 13311
rect 28442 13308 28448 13320
rect 28307 13280 28448 13308
rect 28307 13277 28319 13280
rect 28261 13271 28319 13277
rect 28442 13268 28448 13280
rect 28500 13268 28506 13320
rect 28534 13268 28540 13320
rect 28592 13268 28598 13320
rect 28828 13240 28856 13348
rect 30558 13336 30564 13348
rect 30616 13336 30622 13388
rect 32214 13336 32220 13388
rect 32272 13336 32278 13388
rect 28902 13268 28908 13320
rect 28960 13268 28966 13320
rect 28997 13311 29055 13317
rect 28997 13277 29009 13311
rect 29043 13308 29055 13311
rect 30282 13308 30288 13320
rect 29043 13280 30288 13308
rect 29043 13277 29055 13280
rect 28997 13271 29055 13277
rect 30282 13268 30288 13280
rect 30340 13268 30346 13320
rect 30926 13268 30932 13320
rect 30984 13268 30990 13320
rect 31202 13268 31208 13320
rect 31260 13268 31266 13320
rect 31297 13311 31355 13317
rect 31297 13277 31309 13311
rect 31343 13308 31355 13311
rect 31665 13311 31723 13317
rect 31665 13308 31677 13311
rect 31343 13280 31677 13308
rect 31343 13277 31355 13280
rect 31297 13271 31355 13277
rect 31665 13277 31677 13280
rect 31711 13277 31723 13311
rect 31665 13271 31723 13277
rect 27724 13212 28856 13240
rect 29730 13200 29736 13252
rect 29788 13240 29794 13252
rect 30098 13240 30104 13252
rect 29788 13212 30104 13240
rect 29788 13200 29794 13212
rect 30098 13200 30104 13212
rect 30156 13200 30162 13252
rect 30650 13200 30656 13252
rect 30708 13240 30714 13252
rect 30834 13240 30840 13252
rect 30708 13212 30840 13240
rect 30708 13200 30714 13212
rect 30834 13200 30840 13212
rect 30892 13240 30898 13252
rect 31113 13243 31171 13249
rect 31113 13240 31125 13243
rect 30892 13212 31125 13240
rect 30892 13200 30898 13212
rect 31113 13209 31125 13212
rect 31159 13209 31171 13243
rect 31113 13203 31171 13209
rect 24636 13144 26464 13172
rect 27617 13175 27675 13181
rect 24636 13132 24642 13144
rect 27617 13141 27629 13175
rect 27663 13172 27675 13175
rect 27706 13172 27712 13184
rect 27663 13144 27712 13172
rect 27663 13141 27675 13144
rect 27617 13135 27675 13141
rect 27706 13132 27712 13144
rect 27764 13172 27770 13184
rect 28442 13172 28448 13184
rect 27764 13144 28448 13172
rect 27764 13132 27770 13144
rect 28442 13132 28448 13144
rect 28500 13132 28506 13184
rect 1104 13082 32844 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 32844 13082
rect 1104 13008 32844 13030
rect 2498 12928 2504 12980
rect 2556 12968 2562 12980
rect 6086 12968 6092 12980
rect 2556 12940 6092 12968
rect 2556 12928 2562 12940
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 6365 12971 6423 12977
rect 6365 12937 6377 12971
rect 6411 12968 6423 12971
rect 6454 12968 6460 12980
rect 6411 12940 6460 12968
rect 6411 12937 6423 12940
rect 6365 12931 6423 12937
rect 6454 12928 6460 12940
rect 6512 12968 6518 12980
rect 6730 12968 6736 12980
rect 6512 12940 6736 12968
rect 6512 12928 6518 12940
rect 6730 12928 6736 12940
rect 6788 12928 6794 12980
rect 8202 12968 8208 12980
rect 6886 12940 8208 12968
rect 3513 12903 3571 12909
rect 3513 12900 3525 12903
rect 3160 12872 3525 12900
rect 3160 12764 3188 12872
rect 3513 12869 3525 12872
rect 3559 12900 3571 12903
rect 4617 12903 4675 12909
rect 4617 12900 4629 12903
rect 3559 12872 4629 12900
rect 3559 12869 3571 12872
rect 3513 12863 3571 12869
rect 4617 12869 4629 12872
rect 4663 12869 4675 12903
rect 4617 12863 4675 12869
rect 4715 12872 5479 12900
rect 3234 12792 3240 12844
rect 3292 12792 3298 12844
rect 3329 12835 3387 12841
rect 3329 12801 3341 12835
rect 3375 12832 3387 12835
rect 3602 12832 3608 12844
rect 3375 12804 3608 12832
rect 3375 12801 3387 12804
rect 3329 12795 3387 12801
rect 3602 12792 3608 12804
rect 3660 12792 3666 12844
rect 3786 12792 3792 12844
rect 3844 12792 3850 12844
rect 3878 12792 3884 12844
rect 3936 12832 3942 12844
rect 3973 12835 4031 12841
rect 3973 12832 3985 12835
rect 3936 12804 3985 12832
rect 3936 12792 3942 12804
rect 3973 12801 3985 12804
rect 4019 12832 4031 12835
rect 4522 12832 4528 12844
rect 4019 12804 4528 12832
rect 4019 12801 4031 12804
rect 3973 12795 4031 12801
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 3160 12736 3280 12764
rect 3252 12708 3280 12736
rect 3053 12699 3111 12705
rect 3053 12665 3065 12699
rect 3099 12696 3111 12699
rect 3142 12696 3148 12708
rect 3099 12668 3148 12696
rect 3099 12665 3111 12668
rect 3053 12659 3111 12665
rect 3142 12656 3148 12668
rect 3200 12656 3206 12708
rect 3234 12656 3240 12708
rect 3292 12656 3298 12708
rect 4715 12696 4743 12872
rect 4801 12835 4859 12841
rect 4801 12801 4813 12835
rect 4847 12801 4859 12835
rect 4801 12795 4859 12801
rect 4985 12835 5043 12841
rect 4985 12801 4997 12835
rect 5031 12832 5043 12835
rect 5031 12804 5212 12832
rect 5031 12801 5043 12804
rect 4985 12795 5043 12801
rect 4816 12764 4844 12795
rect 5184 12764 5212 12804
rect 5258 12792 5264 12844
rect 5316 12792 5322 12844
rect 4816 12736 5120 12764
rect 5184 12736 5396 12764
rect 5092 12708 5120 12736
rect 3528 12668 4743 12696
rect 3528 12637 3556 12668
rect 5074 12656 5080 12708
rect 5132 12656 5138 12708
rect 3513 12631 3571 12637
rect 3513 12597 3525 12631
rect 3559 12597 3571 12631
rect 3513 12591 3571 12597
rect 3786 12588 3792 12640
rect 3844 12628 3850 12640
rect 5258 12628 5264 12640
rect 3844 12600 5264 12628
rect 3844 12588 3850 12600
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 5368 12637 5396 12736
rect 5451 12696 5479 12872
rect 5718 12860 5724 12912
rect 5776 12860 5782 12912
rect 6886 12900 6914 12940
rect 8202 12928 8208 12940
rect 8260 12928 8266 12980
rect 14090 12968 14096 12980
rect 8680 12940 14096 12968
rect 6472 12872 6914 12900
rect 5537 12835 5595 12841
rect 5537 12801 5549 12835
rect 5583 12801 5595 12835
rect 5736 12832 5764 12860
rect 5902 12832 5908 12844
rect 5736 12804 5908 12832
rect 5537 12795 5595 12801
rect 5552 12764 5580 12795
rect 5902 12792 5908 12804
rect 5960 12792 5966 12844
rect 6089 12835 6147 12841
rect 6089 12801 6101 12835
rect 6135 12832 6147 12835
rect 6472 12832 6500 12872
rect 7650 12860 7656 12912
rect 7708 12900 7714 12912
rect 8680 12909 8708 12940
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 15381 12971 15439 12977
rect 15381 12937 15393 12971
rect 15427 12968 15439 12971
rect 15470 12968 15476 12980
rect 15427 12940 15476 12968
rect 15427 12937 15439 12940
rect 15381 12931 15439 12937
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 15580 12940 19932 12968
rect 8665 12903 8723 12909
rect 8665 12900 8677 12903
rect 7708 12872 8677 12900
rect 7708 12860 7714 12872
rect 8665 12869 8677 12872
rect 8711 12869 8723 12903
rect 10410 12900 10416 12912
rect 8665 12863 8723 12869
rect 8864 12872 10416 12900
rect 6135 12804 6500 12832
rect 6135 12801 6147 12804
rect 6089 12795 6147 12801
rect 6546 12792 6552 12844
rect 6604 12792 6610 12844
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12832 6883 12835
rect 7006 12832 7012 12844
rect 6871 12804 7012 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 7006 12792 7012 12804
rect 7064 12792 7070 12844
rect 7282 12792 7288 12844
rect 7340 12832 7346 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 7340 12804 7389 12832
rect 7340 12792 7346 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 8389 12835 8447 12841
rect 8389 12801 8401 12835
rect 8435 12832 8447 12835
rect 8570 12832 8576 12844
rect 8435 12804 8576 12832
rect 8435 12801 8447 12804
rect 8389 12795 8447 12801
rect 8570 12792 8576 12804
rect 8628 12792 8634 12844
rect 8754 12792 8760 12844
rect 8812 12832 8818 12844
rect 8864 12841 8892 12872
rect 10410 12860 10416 12872
rect 10468 12860 10474 12912
rect 11517 12903 11575 12909
rect 11517 12869 11529 12903
rect 11563 12900 11575 12903
rect 11563 12872 11928 12900
rect 11563 12869 11575 12872
rect 11517 12863 11575 12869
rect 11900 12844 11928 12872
rect 12526 12860 12532 12912
rect 12584 12900 12590 12912
rect 14921 12903 14979 12909
rect 14921 12900 14933 12903
rect 12584 12872 14933 12900
rect 12584 12860 12590 12872
rect 14921 12869 14933 12872
rect 14967 12900 14979 12903
rect 15580 12900 15608 12940
rect 14967 12872 15608 12900
rect 14967 12869 14979 12872
rect 14921 12863 14979 12869
rect 15654 12860 15660 12912
rect 15712 12860 15718 12912
rect 16758 12900 16764 12912
rect 15856 12872 16764 12900
rect 8849 12835 8907 12841
rect 8849 12832 8861 12835
rect 8812 12804 8861 12832
rect 8812 12792 8818 12804
rect 8849 12801 8861 12804
rect 8895 12801 8907 12835
rect 8849 12795 8907 12801
rect 8938 12792 8944 12844
rect 8996 12792 9002 12844
rect 9490 12792 9496 12844
rect 9548 12792 9554 12844
rect 9769 12835 9827 12841
rect 9769 12801 9781 12835
rect 9815 12832 9827 12835
rect 9858 12832 9864 12844
rect 9815 12804 9864 12832
rect 9815 12801 9827 12804
rect 9769 12795 9827 12801
rect 9858 12792 9864 12804
rect 9916 12792 9922 12844
rect 10042 12792 10048 12844
rect 10100 12832 10106 12844
rect 11040 12835 11098 12841
rect 11040 12832 11052 12835
rect 10100 12804 11052 12832
rect 10100 12792 10106 12804
rect 11040 12801 11052 12804
rect 11086 12801 11098 12835
rect 11040 12795 11098 12801
rect 11333 12835 11391 12841
rect 11333 12801 11345 12835
rect 11379 12822 11391 12835
rect 11422 12822 11428 12844
rect 11379 12801 11428 12822
rect 11333 12795 11428 12801
rect 11348 12794 11428 12795
rect 11422 12792 11428 12794
rect 11480 12792 11486 12844
rect 11790 12792 11796 12844
rect 11848 12792 11854 12844
rect 11882 12792 11888 12844
rect 11940 12792 11946 12844
rect 11974 12792 11980 12844
rect 12032 12792 12038 12844
rect 12342 12792 12348 12844
rect 12400 12792 12406 12844
rect 15102 12792 15108 12844
rect 15160 12792 15166 12844
rect 15197 12835 15255 12841
rect 15197 12801 15209 12835
rect 15243 12832 15255 12835
rect 15286 12832 15292 12844
rect 15243 12804 15292 12832
rect 15243 12801 15255 12804
rect 15197 12795 15255 12801
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 15378 12792 15384 12844
rect 15436 12832 15442 12844
rect 15473 12835 15531 12841
rect 15473 12832 15485 12835
rect 15436 12804 15485 12832
rect 15436 12792 15442 12804
rect 15473 12801 15485 12804
rect 15519 12801 15531 12835
rect 15473 12795 15531 12801
rect 6178 12764 6184 12776
rect 5552 12736 6184 12764
rect 6178 12724 6184 12736
rect 6236 12724 6242 12776
rect 6270 12724 6276 12776
rect 6328 12764 6334 12776
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 6328 12736 6653 12764
rect 6328 12724 6334 12736
rect 6641 12733 6653 12736
rect 6687 12733 6699 12767
rect 6641 12727 6699 12733
rect 6748 12736 6960 12764
rect 5721 12699 5779 12705
rect 5721 12696 5733 12699
rect 5451 12668 5733 12696
rect 5721 12665 5733 12668
rect 5767 12696 5779 12699
rect 6546 12696 6552 12708
rect 5767 12668 6552 12696
rect 5767 12665 5779 12668
rect 5721 12659 5779 12665
rect 6546 12656 6552 12668
rect 6604 12656 6610 12708
rect 6748 12696 6776 12736
rect 6656 12668 6776 12696
rect 5353 12631 5411 12637
rect 5353 12597 5365 12631
rect 5399 12628 5411 12631
rect 6656 12628 6684 12668
rect 6822 12656 6828 12708
rect 6880 12656 6886 12708
rect 6932 12696 6960 12736
rect 7098 12724 7104 12776
rect 7156 12724 7162 12776
rect 9306 12764 9312 12776
rect 7208 12736 9312 12764
rect 7208 12696 7236 12736
rect 9306 12724 9312 12736
rect 9364 12724 9370 12776
rect 10870 12724 10876 12776
rect 10928 12724 10934 12776
rect 11238 12724 11244 12776
rect 11296 12724 11302 12776
rect 11701 12767 11759 12773
rect 11701 12733 11713 12767
rect 11747 12764 11759 12767
rect 11992 12764 12020 12792
rect 12434 12764 12440 12776
rect 11747 12736 12440 12764
rect 11747 12733 11759 12736
rect 11701 12727 11759 12733
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 12526 12724 12532 12776
rect 12584 12764 12590 12776
rect 12986 12764 12992 12776
rect 12584 12736 12992 12764
rect 12584 12724 12590 12736
rect 12986 12724 12992 12736
rect 13044 12764 13050 12776
rect 14918 12764 14924 12776
rect 13044 12736 14924 12764
rect 13044 12724 13050 12736
rect 14918 12724 14924 12736
rect 14976 12764 14982 12776
rect 15013 12767 15071 12773
rect 15013 12764 15025 12767
rect 14976 12736 15025 12764
rect 14976 12724 14982 12736
rect 15013 12733 15025 12736
rect 15059 12733 15071 12767
rect 15120 12764 15148 12792
rect 15856 12773 15884 12872
rect 16758 12860 16764 12872
rect 16816 12860 16822 12912
rect 19904 12909 19932 12940
rect 20530 12928 20536 12980
rect 20588 12968 20594 12980
rect 22738 12968 22744 12980
rect 20588 12940 22744 12968
rect 20588 12928 20594 12940
rect 22738 12928 22744 12940
rect 22796 12928 22802 12980
rect 23750 12928 23756 12980
rect 23808 12968 23814 12980
rect 23845 12971 23903 12977
rect 23845 12968 23857 12971
rect 23808 12940 23857 12968
rect 23808 12928 23814 12940
rect 23845 12937 23857 12940
rect 23891 12937 23903 12971
rect 23845 12931 23903 12937
rect 23934 12928 23940 12980
rect 23992 12968 23998 12980
rect 24394 12968 24400 12980
rect 23992 12940 24164 12968
rect 23992 12928 23998 12940
rect 19889 12903 19947 12909
rect 17144 12872 19334 12900
rect 15930 12792 15936 12844
rect 15988 12792 15994 12844
rect 16022 12792 16028 12844
rect 16080 12832 16086 12844
rect 16209 12835 16267 12841
rect 16209 12832 16221 12835
rect 16080 12804 16221 12832
rect 16080 12792 16086 12804
rect 16209 12801 16221 12804
rect 16255 12832 16267 12835
rect 16482 12832 16488 12844
rect 16255 12804 16488 12832
rect 16255 12801 16267 12804
rect 16209 12795 16267 12801
rect 16482 12792 16488 12804
rect 16540 12792 16546 12844
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 15841 12767 15899 12773
rect 15841 12764 15853 12767
rect 15120 12736 15853 12764
rect 15013 12727 15071 12733
rect 15841 12733 15853 12736
rect 15887 12733 15899 12767
rect 15841 12727 15899 12733
rect 16117 12767 16175 12773
rect 16117 12733 16129 12767
rect 16163 12764 16175 12767
rect 16390 12764 16396 12776
rect 16163 12736 16396 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 16390 12724 16396 12736
rect 16448 12724 16454 12776
rect 16853 12767 16911 12773
rect 16853 12733 16865 12767
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 6932 12668 7236 12696
rect 8573 12699 8631 12705
rect 8573 12665 8585 12699
rect 8619 12696 8631 12699
rect 8754 12696 8760 12708
rect 8619 12668 8760 12696
rect 8619 12665 8631 12668
rect 8573 12659 8631 12665
rect 8754 12656 8760 12668
rect 8812 12656 8818 12708
rect 8956 12668 9720 12696
rect 5399 12600 6684 12628
rect 6733 12631 6791 12637
rect 5399 12597 5411 12600
rect 5353 12591 5411 12597
rect 6733 12597 6745 12631
rect 6779 12628 6791 12631
rect 6840 12628 6868 12656
rect 6779 12600 6868 12628
rect 6779 12597 6791 12600
rect 6733 12591 6791 12597
rect 7006 12588 7012 12640
rect 7064 12628 7070 12640
rect 7926 12628 7932 12640
rect 7064 12600 7932 12628
rect 7064 12588 7070 12600
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 8956 12637 8984 12668
rect 8941 12631 8999 12637
rect 8941 12597 8953 12631
rect 8987 12597 8999 12631
rect 8941 12591 8999 12597
rect 9122 12588 9128 12640
rect 9180 12588 9186 12640
rect 9306 12588 9312 12640
rect 9364 12588 9370 12640
rect 9490 12588 9496 12640
rect 9548 12628 9554 12640
rect 9585 12631 9643 12637
rect 9585 12628 9597 12631
rect 9548 12600 9597 12628
rect 9548 12588 9554 12600
rect 9585 12597 9597 12600
rect 9631 12597 9643 12631
rect 9692 12628 9720 12668
rect 9766 12656 9772 12708
rect 9824 12696 9830 12708
rect 10594 12696 10600 12708
rect 9824 12668 10600 12696
rect 9824 12656 9830 12668
rect 10594 12656 10600 12668
rect 10652 12656 10658 12708
rect 10888 12696 10916 12724
rect 11977 12699 12035 12705
rect 10888 12668 11560 12696
rect 10042 12628 10048 12640
rect 9692 12600 10048 12628
rect 9585 12591 9643 12597
rect 10042 12588 10048 12600
rect 10100 12588 10106 12640
rect 10870 12588 10876 12640
rect 10928 12588 10934 12640
rect 11146 12588 11152 12640
rect 11204 12588 11210 12640
rect 11532 12637 11560 12668
rect 11977 12665 11989 12699
rect 12023 12696 12035 12699
rect 12023 12668 12940 12696
rect 12023 12665 12035 12668
rect 11977 12659 12035 12665
rect 11517 12631 11575 12637
rect 11517 12597 11529 12631
rect 11563 12597 11575 12631
rect 11517 12591 11575 12597
rect 12066 12588 12072 12640
rect 12124 12628 12130 12640
rect 12161 12631 12219 12637
rect 12161 12628 12173 12631
rect 12124 12600 12173 12628
rect 12124 12588 12130 12600
rect 12161 12597 12173 12600
rect 12207 12628 12219 12631
rect 12526 12628 12532 12640
rect 12207 12600 12532 12628
rect 12207 12597 12219 12600
rect 12161 12591 12219 12597
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 12912 12628 12940 12668
rect 14826 12656 14832 12708
rect 14884 12696 14890 12708
rect 16868 12696 16896 12727
rect 16942 12724 16948 12776
rect 17000 12764 17006 12776
rect 17052 12764 17080 12795
rect 17000 12736 17080 12764
rect 17000 12724 17006 12736
rect 14884 12668 16896 12696
rect 14884 12656 14890 12668
rect 13722 12628 13728 12640
rect 12912 12600 13728 12628
rect 13722 12588 13728 12600
rect 13780 12588 13786 12640
rect 15105 12631 15163 12637
rect 15105 12597 15117 12631
rect 15151 12628 15163 12631
rect 15194 12628 15200 12640
rect 15151 12600 15200 12628
rect 15151 12597 15163 12600
rect 15105 12591 15163 12597
rect 15194 12588 15200 12600
rect 15252 12588 15258 12640
rect 15470 12588 15476 12640
rect 15528 12628 15534 12640
rect 15654 12628 15660 12640
rect 15528 12600 15660 12628
rect 15528 12588 15534 12600
rect 15654 12588 15660 12600
rect 15712 12588 15718 12640
rect 16206 12588 16212 12640
rect 16264 12588 16270 12640
rect 16298 12588 16304 12640
rect 16356 12628 16362 12640
rect 16393 12631 16451 12637
rect 16393 12628 16405 12631
rect 16356 12600 16405 12628
rect 16356 12588 16362 12600
rect 16393 12597 16405 12600
rect 16439 12597 16451 12631
rect 16393 12591 16451 12597
rect 16853 12631 16911 12637
rect 16853 12597 16865 12631
rect 16899 12628 16911 12631
rect 17144 12628 17172 12872
rect 17310 12792 17316 12844
rect 17368 12792 17374 12844
rect 18506 12792 18512 12844
rect 18564 12832 18570 12844
rect 18601 12835 18659 12841
rect 18601 12832 18613 12835
rect 18564 12804 18613 12832
rect 18564 12792 18570 12804
rect 18601 12801 18613 12804
rect 18647 12801 18659 12835
rect 18601 12795 18659 12801
rect 18690 12792 18696 12844
rect 18748 12792 18754 12844
rect 19306 12832 19334 12872
rect 19889 12869 19901 12903
rect 19935 12869 19947 12903
rect 20257 12903 20315 12909
rect 19889 12863 19947 12869
rect 19996 12872 20208 12900
rect 19996 12832 20024 12872
rect 19306 12804 20024 12832
rect 20070 12792 20076 12844
rect 20128 12792 20134 12844
rect 20180 12832 20208 12872
rect 20257 12869 20269 12903
rect 20303 12900 20315 12903
rect 21082 12900 21088 12912
rect 20303 12872 21088 12900
rect 20303 12869 20315 12872
rect 20257 12863 20315 12869
rect 21082 12860 21088 12872
rect 21140 12860 21146 12912
rect 22005 12835 22063 12841
rect 20180 12804 21772 12832
rect 17954 12764 17960 12776
rect 17236 12736 17960 12764
rect 17236 12637 17264 12736
rect 17954 12724 17960 12736
rect 18012 12724 18018 12776
rect 18782 12724 18788 12776
rect 18840 12764 18846 12776
rect 21634 12764 21640 12776
rect 18840 12736 21640 12764
rect 18840 12724 18846 12736
rect 21634 12724 21640 12736
rect 21692 12724 21698 12776
rect 21744 12764 21772 12804
rect 22005 12801 22017 12835
rect 22051 12832 22063 12835
rect 22094 12832 22100 12844
rect 22051 12804 22100 12832
rect 22051 12801 22063 12804
rect 22005 12795 22063 12801
rect 22094 12792 22100 12804
rect 22152 12792 22158 12844
rect 22186 12792 22192 12844
rect 22244 12792 22250 12844
rect 22462 12792 22468 12844
rect 22520 12832 22526 12844
rect 23385 12835 23443 12841
rect 23385 12832 23397 12835
rect 22520 12804 23397 12832
rect 22520 12792 22526 12804
rect 23385 12801 23397 12804
rect 23431 12801 23443 12835
rect 23385 12795 23443 12801
rect 23934 12792 23940 12844
rect 23992 12832 23998 12844
rect 24029 12835 24087 12841
rect 24029 12832 24041 12835
rect 23992 12804 24041 12832
rect 23992 12792 23998 12804
rect 24029 12801 24041 12804
rect 24075 12801 24087 12835
rect 24136 12832 24164 12940
rect 24228 12940 24400 12968
rect 24228 12909 24256 12940
rect 24394 12928 24400 12940
rect 24452 12928 24458 12980
rect 24670 12928 24676 12980
rect 24728 12968 24734 12980
rect 27617 12971 27675 12977
rect 24728 12940 26280 12968
rect 24728 12928 24734 12940
rect 24213 12903 24271 12909
rect 24213 12869 24225 12903
rect 24259 12869 24271 12903
rect 25777 12903 25835 12909
rect 25777 12900 25789 12903
rect 24213 12863 24271 12869
rect 24412 12872 25789 12900
rect 24305 12835 24363 12841
rect 24305 12832 24317 12835
rect 24136 12804 24317 12832
rect 24029 12795 24087 12801
rect 24305 12801 24317 12804
rect 24351 12801 24363 12835
rect 24305 12795 24363 12801
rect 21910 12764 21916 12776
rect 21744 12736 21916 12764
rect 21910 12724 21916 12736
rect 21968 12764 21974 12776
rect 22646 12764 22652 12776
rect 21968 12736 22652 12764
rect 21968 12724 21974 12736
rect 22646 12724 22652 12736
rect 22704 12724 22710 12776
rect 23198 12724 23204 12776
rect 23256 12764 23262 12776
rect 23477 12767 23535 12773
rect 23256 12736 23428 12764
rect 23256 12724 23262 12736
rect 17497 12699 17555 12705
rect 17497 12665 17509 12699
rect 17543 12696 17555 12699
rect 17586 12696 17592 12708
rect 17543 12668 17592 12696
rect 17543 12665 17555 12668
rect 17497 12659 17555 12665
rect 17586 12656 17592 12668
rect 17644 12696 17650 12708
rect 17770 12696 17776 12708
rect 17644 12668 17776 12696
rect 17644 12656 17650 12668
rect 17770 12656 17776 12668
rect 17828 12696 17834 12708
rect 22462 12696 22468 12708
rect 17828 12668 22468 12696
rect 17828 12656 17834 12668
rect 22462 12656 22468 12668
rect 22520 12656 22526 12708
rect 16899 12600 17172 12628
rect 17221 12631 17279 12637
rect 16899 12597 16911 12600
rect 16853 12591 16911 12597
rect 17221 12597 17233 12631
rect 17267 12597 17279 12631
rect 17221 12591 17279 12597
rect 17310 12588 17316 12640
rect 17368 12628 17374 12640
rect 18601 12631 18659 12637
rect 18601 12628 18613 12631
rect 17368 12600 18613 12628
rect 17368 12588 17374 12600
rect 18601 12597 18613 12600
rect 18647 12628 18659 12631
rect 18782 12628 18788 12640
rect 18647 12600 18788 12628
rect 18647 12597 18659 12600
rect 18601 12591 18659 12597
rect 18782 12588 18788 12600
rect 18840 12588 18846 12640
rect 18874 12588 18880 12640
rect 18932 12628 18938 12640
rect 18969 12631 19027 12637
rect 18969 12628 18981 12631
rect 18932 12600 18981 12628
rect 18932 12588 18938 12600
rect 18969 12597 18981 12600
rect 19015 12597 19027 12631
rect 18969 12591 19027 12597
rect 21634 12588 21640 12640
rect 21692 12628 21698 12640
rect 22097 12631 22155 12637
rect 22097 12628 22109 12631
rect 21692 12600 22109 12628
rect 21692 12588 21698 12600
rect 22097 12597 22109 12600
rect 22143 12597 22155 12631
rect 22097 12591 22155 12597
rect 22373 12631 22431 12637
rect 22373 12597 22385 12631
rect 22419 12628 22431 12631
rect 22830 12628 22836 12640
rect 22419 12600 22836 12628
rect 22419 12597 22431 12600
rect 22373 12591 22431 12597
rect 22830 12588 22836 12600
rect 22888 12588 22894 12640
rect 23400 12628 23428 12736
rect 23477 12733 23489 12767
rect 23523 12764 23535 12767
rect 23658 12764 23664 12776
rect 23523 12736 23664 12764
rect 23523 12733 23535 12736
rect 23477 12727 23535 12733
rect 23658 12724 23664 12736
rect 23716 12764 23722 12776
rect 24412 12764 24440 12872
rect 25777 12869 25789 12872
rect 25823 12900 25835 12903
rect 26142 12900 26148 12912
rect 25823 12872 26148 12900
rect 25823 12869 25835 12872
rect 25777 12863 25835 12869
rect 26142 12860 26148 12872
rect 26200 12860 26206 12912
rect 26252 12900 26280 12940
rect 27617 12937 27629 12971
rect 27663 12968 27675 12971
rect 28902 12968 28908 12980
rect 27663 12940 28908 12968
rect 27663 12937 27675 12940
rect 27617 12931 27675 12937
rect 28902 12928 28908 12940
rect 28960 12928 28966 12980
rect 29546 12928 29552 12980
rect 29604 12968 29610 12980
rect 30098 12968 30104 12980
rect 29604 12940 30104 12968
rect 29604 12928 29610 12940
rect 30098 12928 30104 12940
rect 30156 12928 30162 12980
rect 30377 12971 30435 12977
rect 30377 12937 30389 12971
rect 30423 12968 30435 12971
rect 31662 12968 31668 12980
rect 30423 12940 31668 12968
rect 30423 12937 30435 12940
rect 30377 12931 30435 12937
rect 31662 12928 31668 12940
rect 31720 12928 31726 12980
rect 28074 12900 28080 12912
rect 26252 12872 28080 12900
rect 28074 12860 28080 12872
rect 28132 12860 28138 12912
rect 28166 12860 28172 12912
rect 28224 12860 28230 12912
rect 30558 12860 30564 12912
rect 30616 12900 30622 12912
rect 30616 12872 31984 12900
rect 30616 12860 30622 12872
rect 24762 12792 24768 12844
rect 24820 12792 24826 12844
rect 24854 12792 24860 12844
rect 24912 12792 24918 12844
rect 26050 12792 26056 12844
rect 26108 12792 26114 12844
rect 27154 12792 27160 12844
rect 27212 12792 27218 12844
rect 27430 12792 27436 12844
rect 27488 12792 27494 12844
rect 28445 12835 28503 12841
rect 28445 12832 28457 12835
rect 28368 12804 28457 12832
rect 25869 12767 25927 12773
rect 25869 12764 25881 12767
rect 23716 12736 24440 12764
rect 25056 12736 25881 12764
rect 23716 12724 23722 12736
rect 24489 12699 24547 12705
rect 24489 12665 24501 12699
rect 24535 12696 24547 12699
rect 24670 12696 24676 12708
rect 24535 12668 24676 12696
rect 24535 12665 24547 12668
rect 24489 12659 24547 12665
rect 24670 12656 24676 12668
rect 24728 12656 24734 12708
rect 25056 12640 25084 12736
rect 25869 12733 25881 12736
rect 25915 12764 25927 12767
rect 26878 12764 26884 12776
rect 25915 12736 26884 12764
rect 25915 12733 25927 12736
rect 25869 12727 25927 12733
rect 26878 12724 26884 12736
rect 26936 12724 26942 12776
rect 27246 12724 27252 12776
rect 27304 12724 27310 12776
rect 27448 12764 27476 12792
rect 28261 12767 28319 12773
rect 28261 12764 28273 12767
rect 27448 12736 28273 12764
rect 28261 12733 28273 12736
rect 28307 12733 28319 12767
rect 28261 12727 28319 12733
rect 26237 12699 26295 12705
rect 26237 12665 26249 12699
rect 26283 12696 26295 12699
rect 28368 12696 28396 12804
rect 28445 12801 28457 12804
rect 28491 12801 28503 12835
rect 28445 12795 28503 12801
rect 30282 12792 30288 12844
rect 30340 12792 30346 12844
rect 30650 12792 30656 12844
rect 30708 12832 30714 12844
rect 31202 12832 31208 12844
rect 30708 12804 31208 12832
rect 30708 12792 30714 12804
rect 31202 12792 31208 12804
rect 31260 12792 31266 12844
rect 31956 12841 31984 12872
rect 31685 12835 31743 12841
rect 31685 12801 31697 12835
rect 31731 12832 31743 12835
rect 31941 12835 31999 12841
rect 31731 12804 31892 12832
rect 31731 12801 31743 12804
rect 31685 12795 31743 12801
rect 28626 12724 28632 12776
rect 28684 12724 28690 12776
rect 28644 12696 28672 12724
rect 26283 12668 28396 12696
rect 28460 12668 28672 12696
rect 30300 12696 30328 12792
rect 31864 12764 31892 12804
rect 31941 12801 31953 12835
rect 31987 12801 31999 12835
rect 31941 12795 31999 12801
rect 32490 12792 32496 12844
rect 32548 12792 32554 12844
rect 31864 12736 32352 12764
rect 32324 12705 32352 12736
rect 30561 12699 30619 12705
rect 30561 12696 30573 12699
rect 30300 12668 30573 12696
rect 26283 12665 26295 12668
rect 26237 12659 26295 12665
rect 23477 12631 23535 12637
rect 23477 12628 23489 12631
rect 23400 12600 23489 12628
rect 23477 12597 23489 12600
rect 23523 12597 23535 12631
rect 23477 12591 23535 12597
rect 23750 12588 23756 12640
rect 23808 12588 23814 12640
rect 24118 12588 24124 12640
rect 24176 12628 24182 12640
rect 24394 12628 24400 12640
rect 24176 12600 24400 12628
rect 24176 12588 24182 12600
rect 24394 12588 24400 12600
rect 24452 12628 24458 12640
rect 24581 12631 24639 12637
rect 24581 12628 24593 12631
rect 24452 12600 24593 12628
rect 24452 12588 24458 12600
rect 24581 12597 24593 12600
rect 24627 12597 24639 12631
rect 24581 12591 24639 12597
rect 25038 12588 25044 12640
rect 25096 12588 25102 12640
rect 25774 12588 25780 12640
rect 25832 12588 25838 12640
rect 26602 12588 26608 12640
rect 26660 12628 26666 12640
rect 28460 12637 28488 12668
rect 30561 12665 30573 12668
rect 30607 12665 30619 12699
rect 30561 12659 30619 12665
rect 32309 12699 32367 12705
rect 32309 12665 32321 12699
rect 32355 12665 32367 12699
rect 32309 12659 32367 12665
rect 27157 12631 27215 12637
rect 27157 12628 27169 12631
rect 26660 12600 27169 12628
rect 26660 12588 26666 12600
rect 27157 12597 27169 12600
rect 27203 12597 27215 12631
rect 27157 12591 27215 12597
rect 28445 12631 28503 12637
rect 28445 12597 28457 12631
rect 28491 12597 28503 12631
rect 28445 12591 28503 12597
rect 28629 12631 28687 12637
rect 28629 12597 28641 12631
rect 28675 12628 28687 12631
rect 30926 12628 30932 12640
rect 28675 12600 30932 12628
rect 28675 12597 28687 12600
rect 28629 12591 28687 12597
rect 30926 12588 30932 12600
rect 30984 12588 30990 12640
rect 1104 12538 32844 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 32844 12538
rect 1104 12464 32844 12486
rect 3050 12384 3056 12436
rect 3108 12384 3114 12436
rect 3145 12427 3203 12433
rect 3145 12393 3157 12427
rect 3191 12424 3203 12427
rect 3191 12396 4936 12424
rect 3191 12393 3203 12396
rect 3145 12387 3203 12393
rect 3160 12356 3188 12387
rect 2884 12328 3188 12356
rect 2774 12288 2780 12300
rect 2424 12260 2780 12288
rect 2424 12229 2452 12260
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 2884 12232 2912 12328
rect 3786 12316 3792 12368
rect 3844 12356 3850 12368
rect 4908 12356 4936 12396
rect 4982 12384 4988 12436
rect 5040 12424 5046 12436
rect 6089 12427 6147 12433
rect 6089 12424 6101 12427
rect 5040 12396 6101 12424
rect 5040 12384 5046 12396
rect 6089 12393 6101 12396
rect 6135 12393 6147 12427
rect 6089 12387 6147 12393
rect 6362 12384 6368 12436
rect 6420 12424 6426 12436
rect 6822 12424 6828 12436
rect 6420 12396 6828 12424
rect 6420 12384 6426 12396
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 7926 12424 7932 12436
rect 6972 12396 7932 12424
rect 6972 12384 6978 12396
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 9306 12384 9312 12436
rect 9364 12424 9370 12436
rect 9401 12427 9459 12433
rect 9401 12424 9413 12427
rect 9364 12396 9413 12424
rect 9364 12384 9370 12396
rect 9401 12393 9413 12396
rect 9447 12424 9459 12427
rect 11333 12427 11391 12433
rect 9447 12396 11284 12424
rect 9447 12393 9459 12396
rect 9401 12387 9459 12393
rect 5074 12356 5080 12368
rect 3844 12328 4844 12356
rect 4908 12328 5080 12356
rect 3844 12316 3850 12328
rect 3050 12248 3056 12300
rect 3108 12288 3114 12300
rect 3108 12260 3832 12288
rect 3108 12248 3114 12260
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12189 2467 12223
rect 2409 12183 2467 12189
rect 2501 12223 2559 12229
rect 2501 12189 2513 12223
rect 2547 12189 2559 12223
rect 2501 12183 2559 12189
rect 2516 12152 2544 12183
rect 2866 12180 2872 12232
rect 2924 12180 2930 12232
rect 3329 12223 3387 12229
rect 3329 12189 3341 12223
rect 3375 12220 3387 12223
rect 3418 12220 3424 12232
rect 3375 12192 3424 12220
rect 3375 12189 3387 12192
rect 3329 12183 3387 12189
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3605 12223 3663 12229
rect 3605 12189 3617 12223
rect 3651 12220 3663 12223
rect 3694 12220 3700 12232
rect 3651 12192 3700 12220
rect 3651 12189 3663 12192
rect 3605 12183 3663 12189
rect 3694 12180 3700 12192
rect 3752 12180 3758 12232
rect 2240 12124 2544 12152
rect 2685 12155 2743 12161
rect 2240 12096 2268 12124
rect 2685 12121 2697 12155
rect 2731 12121 2743 12155
rect 2685 12115 2743 12121
rect 2222 12044 2228 12096
rect 2280 12044 2286 12096
rect 2700 12084 2728 12115
rect 2774 12112 2780 12164
rect 2832 12152 2838 12164
rect 3804 12152 3832 12260
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4709 12223 4767 12229
rect 4709 12220 4721 12223
rect 4120 12192 4721 12220
rect 4120 12180 4126 12192
rect 4709 12189 4721 12192
rect 4755 12189 4767 12223
rect 4816 12220 4844 12328
rect 5074 12316 5080 12328
rect 5132 12316 5138 12368
rect 5261 12359 5319 12365
rect 5261 12325 5273 12359
rect 5307 12356 5319 12359
rect 5307 12328 5672 12356
rect 5307 12325 5319 12328
rect 5261 12319 5319 12325
rect 5276 12260 5580 12288
rect 4982 12220 4988 12232
rect 4816 12192 4988 12220
rect 4709 12183 4767 12189
rect 4982 12180 4988 12192
rect 5040 12180 5046 12232
rect 5074 12180 5080 12232
rect 5132 12229 5138 12232
rect 5132 12223 5159 12229
rect 5147 12189 5159 12223
rect 5132 12183 5159 12189
rect 5132 12180 5138 12183
rect 4893 12155 4951 12161
rect 4893 12152 4905 12155
rect 2832 12124 3464 12152
rect 3804 12124 4905 12152
rect 2832 12112 2838 12124
rect 2958 12084 2964 12096
rect 2700 12056 2964 12084
rect 2958 12044 2964 12056
rect 3016 12044 3022 12096
rect 3436 12093 3464 12124
rect 4893 12121 4905 12124
rect 4939 12152 4951 12155
rect 5276 12152 5304 12260
rect 5552 12229 5580 12260
rect 5353 12223 5411 12229
rect 5353 12189 5365 12223
rect 5399 12189 5411 12223
rect 5353 12183 5411 12189
rect 5537 12223 5595 12229
rect 5537 12189 5549 12223
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 4939 12124 5304 12152
rect 4939 12121 4951 12124
rect 4893 12115 4951 12121
rect 3421 12087 3479 12093
rect 3421 12053 3433 12087
rect 3467 12053 3479 12087
rect 3421 12047 3479 12053
rect 3510 12044 3516 12096
rect 3568 12084 3574 12096
rect 5368 12084 5396 12183
rect 3568 12056 5396 12084
rect 5644 12084 5672 12328
rect 5810 12316 5816 12368
rect 5868 12316 5874 12368
rect 11256 12356 11284 12396
rect 11333 12393 11345 12427
rect 11379 12424 11391 12427
rect 11422 12424 11428 12436
rect 11379 12396 11428 12424
rect 11379 12393 11391 12396
rect 11333 12387 11391 12393
rect 11422 12384 11428 12396
rect 11480 12384 11486 12436
rect 11885 12427 11943 12433
rect 11885 12424 11897 12427
rect 11532 12396 11897 12424
rect 11532 12356 11560 12396
rect 11885 12393 11897 12396
rect 11931 12424 11943 12427
rect 15838 12424 15844 12436
rect 11931 12396 15844 12424
rect 11931 12393 11943 12396
rect 11885 12387 11943 12393
rect 15838 12384 15844 12396
rect 15896 12384 15902 12436
rect 16390 12384 16396 12436
rect 16448 12384 16454 12436
rect 16666 12384 16672 12436
rect 16724 12424 16730 12436
rect 16761 12427 16819 12433
rect 16761 12424 16773 12427
rect 16724 12396 16773 12424
rect 16724 12384 16730 12396
rect 16761 12393 16773 12396
rect 16807 12393 16819 12427
rect 20070 12424 20076 12436
rect 16761 12387 16819 12393
rect 16868 12396 20076 12424
rect 6472 12328 9076 12356
rect 11256 12328 11560 12356
rect 5828 12288 5856 12316
rect 6086 12288 6092 12300
rect 5828 12260 6092 12288
rect 6086 12248 6092 12260
rect 6144 12288 6150 12300
rect 6144 12260 6316 12288
rect 6144 12248 6150 12260
rect 5718 12180 5724 12232
rect 5776 12220 5782 12232
rect 6288 12229 6316 12260
rect 5813 12223 5871 12229
rect 5813 12220 5825 12223
rect 5776 12192 5825 12220
rect 5776 12180 5782 12192
rect 5813 12189 5825 12192
rect 5859 12189 5871 12223
rect 5813 12183 5871 12189
rect 6273 12223 6331 12229
rect 6273 12189 6285 12223
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 5997 12155 6055 12161
rect 5997 12121 6009 12155
rect 6043 12152 6055 12155
rect 6472 12152 6500 12328
rect 6546 12248 6552 12300
rect 6604 12288 6610 12300
rect 8570 12288 8576 12300
rect 6604 12260 8576 12288
rect 6604 12248 6610 12260
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 9048 12288 9076 12328
rect 11790 12316 11796 12368
rect 11848 12356 11854 12368
rect 12526 12356 12532 12368
rect 11848 12328 12532 12356
rect 11848 12316 11854 12328
rect 12526 12316 12532 12328
rect 12584 12316 12590 12368
rect 13078 12316 13084 12368
rect 13136 12356 13142 12368
rect 16868 12356 16896 12396
rect 20070 12384 20076 12396
rect 20128 12384 20134 12436
rect 20530 12384 20536 12436
rect 20588 12424 20594 12436
rect 21450 12424 21456 12436
rect 20588 12396 21456 12424
rect 20588 12384 20594 12396
rect 21450 12384 21456 12396
rect 21508 12384 21514 12436
rect 21910 12384 21916 12436
rect 21968 12384 21974 12436
rect 22094 12384 22100 12436
rect 22152 12424 22158 12436
rect 22649 12427 22707 12433
rect 22649 12424 22661 12427
rect 22152 12396 22661 12424
rect 22152 12384 22158 12396
rect 22649 12393 22661 12396
rect 22695 12424 22707 12427
rect 23290 12424 23296 12436
rect 22695 12396 23296 12424
rect 22695 12393 22707 12396
rect 22649 12387 22707 12393
rect 23290 12384 23296 12396
rect 23348 12384 23354 12436
rect 23658 12384 23664 12436
rect 23716 12384 23722 12436
rect 24394 12384 24400 12436
rect 24452 12384 24458 12436
rect 24946 12384 24952 12436
rect 25004 12384 25010 12436
rect 25409 12427 25467 12433
rect 25409 12393 25421 12427
rect 25455 12393 25467 12427
rect 25409 12387 25467 12393
rect 13136 12328 16896 12356
rect 13136 12316 13142 12328
rect 17218 12316 17224 12368
rect 17276 12316 17282 12368
rect 18782 12316 18788 12368
rect 18840 12356 18846 12368
rect 18840 12328 22876 12356
rect 18840 12316 18846 12328
rect 10226 12288 10232 12300
rect 9048 12260 10232 12288
rect 10226 12248 10232 12260
rect 10284 12248 10290 12300
rect 10428 12260 11652 12288
rect 6638 12180 6644 12232
rect 6696 12220 6702 12232
rect 6733 12223 6791 12229
rect 6733 12220 6745 12223
rect 6696 12192 6745 12220
rect 6696 12180 6702 12192
rect 6733 12189 6745 12192
rect 6779 12189 6791 12223
rect 6733 12183 6791 12189
rect 6917 12223 6975 12229
rect 6917 12189 6929 12223
rect 6963 12220 6975 12223
rect 7006 12220 7012 12232
rect 6963 12192 7012 12220
rect 6963 12189 6975 12192
rect 6917 12183 6975 12189
rect 7006 12180 7012 12192
rect 7064 12180 7070 12232
rect 7193 12223 7251 12229
rect 7193 12189 7205 12223
rect 7239 12220 7251 12223
rect 7282 12220 7288 12232
rect 7239 12192 7288 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 7282 12180 7288 12192
rect 7340 12180 7346 12232
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 8021 12223 8079 12229
rect 8021 12220 8033 12223
rect 7524 12192 8033 12220
rect 7524 12180 7530 12192
rect 8021 12189 8033 12192
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 9122 12180 9128 12232
rect 9180 12229 9186 12232
rect 9180 12220 9190 12229
rect 9180 12192 9225 12220
rect 9180 12183 9190 12192
rect 9180 12180 9186 12183
rect 9306 12180 9312 12232
rect 9364 12180 9370 12232
rect 9401 12223 9459 12229
rect 9401 12189 9413 12223
rect 9447 12220 9459 12223
rect 9674 12220 9680 12232
rect 9447 12192 9680 12220
rect 9447 12189 9459 12192
rect 9401 12183 9459 12189
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 6043 12124 6500 12152
rect 6043 12121 6055 12124
rect 5997 12115 6055 12121
rect 6546 12112 6552 12164
rect 6604 12112 6610 12164
rect 7834 12112 7840 12164
rect 7892 12112 7898 12164
rect 7926 12112 7932 12164
rect 7984 12152 7990 12164
rect 10428 12152 10456 12260
rect 11149 12223 11207 12229
rect 11149 12189 11161 12223
rect 11195 12220 11207 12223
rect 11422 12220 11428 12232
rect 11195 12192 11428 12220
rect 11195 12189 11207 12192
rect 11149 12183 11207 12189
rect 11422 12180 11428 12192
rect 11480 12180 11486 12232
rect 11624 12220 11652 12260
rect 11698 12248 11704 12300
rect 11756 12248 11762 12300
rect 12066 12288 12072 12300
rect 11808 12260 12072 12288
rect 11808 12230 11836 12260
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 12802 12248 12808 12300
rect 12860 12288 12866 12300
rect 16022 12288 16028 12300
rect 12860 12260 16028 12288
rect 12860 12248 12866 12260
rect 16022 12248 16028 12260
rect 16080 12248 16086 12300
rect 16758 12248 16764 12300
rect 16816 12288 16822 12300
rect 16853 12291 16911 12297
rect 16853 12288 16865 12291
rect 16816 12260 16865 12288
rect 16816 12248 16822 12260
rect 16853 12257 16865 12260
rect 16899 12257 16911 12291
rect 16853 12251 16911 12257
rect 16960 12260 19288 12288
rect 11808 12229 11928 12230
rect 11808 12223 11943 12229
rect 11624 12192 11744 12220
rect 11808 12202 11897 12223
rect 7984 12124 10456 12152
rect 7984 12112 7990 12124
rect 10502 12112 10508 12164
rect 10560 12152 10566 12164
rect 10778 12152 10784 12164
rect 10560 12124 10784 12152
rect 10560 12112 10566 12124
rect 10778 12112 10784 12124
rect 10836 12112 10842 12164
rect 10870 12112 10876 12164
rect 10928 12152 10934 12164
rect 11609 12155 11667 12161
rect 11609 12152 11621 12155
rect 10928 12124 11621 12152
rect 10928 12112 10934 12124
rect 11609 12121 11621 12124
rect 11655 12121 11667 12155
rect 11716 12152 11744 12192
rect 11885 12189 11897 12202
rect 11931 12189 11943 12223
rect 11885 12183 11943 12189
rect 13078 12180 13084 12232
rect 13136 12220 13142 12232
rect 13136 12192 13768 12220
rect 13136 12180 13142 12192
rect 13740 12152 13768 12192
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 16209 12223 16267 12229
rect 16209 12220 16221 12223
rect 13872 12192 16221 12220
rect 13872 12180 13878 12192
rect 16209 12189 16221 12192
rect 16255 12189 16267 12223
rect 16960 12220 16988 12260
rect 16209 12183 16267 12189
rect 16316 12192 16988 12220
rect 17037 12223 17095 12229
rect 16316 12152 16344 12192
rect 17037 12189 17049 12223
rect 17083 12220 17095 12223
rect 17586 12220 17592 12232
rect 17083 12192 17592 12220
rect 17083 12189 17095 12192
rect 17037 12183 17095 12189
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 19260 12229 19288 12260
rect 21266 12248 21272 12300
rect 21324 12288 21330 12300
rect 21324 12260 21588 12288
rect 21324 12248 21330 12260
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12189 18015 12223
rect 17957 12183 18015 12189
rect 18233 12223 18291 12229
rect 18233 12189 18245 12223
rect 18279 12189 18291 12223
rect 18233 12183 18291 12189
rect 19245 12223 19303 12229
rect 19245 12189 19257 12223
rect 19291 12220 19303 12223
rect 21450 12220 21456 12232
rect 19291 12192 21456 12220
rect 19291 12189 19303 12192
rect 19245 12183 19303 12189
rect 11716 12124 13676 12152
rect 13740 12124 16344 12152
rect 16761 12155 16819 12161
rect 11609 12115 11667 12121
rect 6914 12084 6920 12096
rect 5644 12056 6920 12084
rect 3568 12044 3574 12056
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 8205 12087 8263 12093
rect 8205 12053 8217 12087
rect 8251 12084 8263 12087
rect 8754 12084 8760 12096
rect 8251 12056 8760 12084
rect 8251 12053 8263 12056
rect 8205 12047 8263 12053
rect 8754 12044 8760 12056
rect 8812 12044 8818 12096
rect 9398 12044 9404 12096
rect 9456 12084 9462 12096
rect 9585 12087 9643 12093
rect 9585 12084 9597 12087
rect 9456 12056 9597 12084
rect 9456 12044 9462 12056
rect 9585 12053 9597 12056
rect 9631 12053 9643 12087
rect 9585 12047 9643 12053
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 11882 12084 11888 12096
rect 9732 12056 11888 12084
rect 9732 12044 9738 12056
rect 11882 12044 11888 12056
rect 11940 12044 11946 12096
rect 12069 12087 12127 12093
rect 12069 12053 12081 12087
rect 12115 12084 12127 12087
rect 12158 12084 12164 12096
rect 12115 12056 12164 12084
rect 12115 12053 12127 12056
rect 12069 12047 12127 12053
rect 12158 12044 12164 12056
rect 12216 12044 12222 12096
rect 13648 12084 13676 12124
rect 16761 12121 16773 12155
rect 16807 12152 16819 12155
rect 17126 12152 17132 12164
rect 16807 12124 17132 12152
rect 16807 12121 16819 12124
rect 16761 12115 16819 12121
rect 17126 12112 17132 12124
rect 17184 12112 17190 12164
rect 17972 12152 18000 12183
rect 17926 12124 18000 12152
rect 18248 12152 18276 12183
rect 21450 12180 21456 12192
rect 21508 12180 21514 12232
rect 21560 12220 21588 12260
rect 21634 12248 21640 12300
rect 21692 12288 21698 12300
rect 21913 12291 21971 12297
rect 21913 12288 21925 12291
rect 21692 12260 21925 12288
rect 21692 12248 21698 12260
rect 21913 12257 21925 12260
rect 21959 12257 21971 12291
rect 22465 12291 22523 12297
rect 22465 12288 22477 12291
rect 21913 12251 21971 12257
rect 22009 12260 22477 12288
rect 22009 12220 22037 12260
rect 22465 12257 22477 12260
rect 22511 12257 22523 12291
rect 22465 12251 22523 12257
rect 21560 12192 22037 12220
rect 22094 12180 22100 12232
rect 22152 12180 22158 12232
rect 22649 12223 22707 12229
rect 22649 12189 22661 12223
rect 22695 12220 22707 12223
rect 22738 12220 22744 12232
rect 22695 12192 22744 12220
rect 22695 12189 22707 12192
rect 22649 12183 22707 12189
rect 22738 12180 22744 12192
rect 22796 12180 22802 12232
rect 22848 12220 22876 12328
rect 23934 12316 23940 12368
rect 23992 12356 23998 12368
rect 23992 12328 24624 12356
rect 23992 12316 23998 12328
rect 23014 12248 23020 12300
rect 23072 12288 23078 12300
rect 23198 12288 23204 12300
rect 23072 12260 23204 12288
rect 23072 12248 23078 12260
rect 23198 12248 23204 12260
rect 23256 12248 23262 12300
rect 23750 12248 23756 12300
rect 23808 12288 23814 12300
rect 24489 12291 24547 12297
rect 24489 12288 24501 12291
rect 23808 12260 24501 12288
rect 23808 12248 23814 12260
rect 24489 12257 24501 12260
rect 24535 12257 24547 12291
rect 24596 12288 24624 12328
rect 24762 12316 24768 12368
rect 24820 12356 24826 12368
rect 24857 12359 24915 12365
rect 24857 12356 24869 12359
rect 24820 12328 24869 12356
rect 24820 12316 24826 12328
rect 24857 12325 24869 12328
rect 24903 12325 24915 12359
rect 24857 12319 24915 12325
rect 25314 12316 25320 12368
rect 25372 12356 25378 12368
rect 25424 12356 25452 12387
rect 25590 12384 25596 12436
rect 25648 12384 25654 12436
rect 25961 12427 26019 12433
rect 25961 12393 25973 12427
rect 26007 12424 26019 12427
rect 26602 12424 26608 12436
rect 26007 12396 26608 12424
rect 26007 12393 26019 12396
rect 25961 12387 26019 12393
rect 26602 12384 26608 12396
rect 26660 12384 26666 12436
rect 26878 12384 26884 12436
rect 26936 12384 26942 12436
rect 27065 12427 27123 12433
rect 27065 12393 27077 12427
rect 27111 12424 27123 12427
rect 27154 12424 27160 12436
rect 27111 12396 27160 12424
rect 27111 12393 27123 12396
rect 27065 12387 27123 12393
rect 27154 12384 27160 12396
rect 27212 12384 27218 12436
rect 27798 12384 27804 12436
rect 27856 12384 27862 12436
rect 27985 12427 28043 12433
rect 27985 12393 27997 12427
rect 28031 12424 28043 12427
rect 28074 12424 28080 12436
rect 28031 12396 28080 12424
rect 28031 12393 28043 12396
rect 27985 12387 28043 12393
rect 28074 12384 28080 12396
rect 28132 12384 28138 12436
rect 29454 12384 29460 12436
rect 29512 12424 29518 12436
rect 30101 12427 30159 12433
rect 30101 12424 30113 12427
rect 29512 12396 30113 12424
rect 29512 12384 29518 12396
rect 30101 12393 30113 12396
rect 30147 12393 30159 12427
rect 30101 12387 30159 12393
rect 25372 12328 25452 12356
rect 25372 12316 25378 12328
rect 25498 12316 25504 12368
rect 25556 12316 25562 12368
rect 25774 12316 25780 12368
rect 25832 12316 25838 12368
rect 25041 12291 25099 12297
rect 25041 12288 25053 12291
rect 24596 12260 25053 12288
rect 24489 12251 24547 12257
rect 25041 12257 25053 12260
rect 25087 12257 25099 12291
rect 25041 12251 25099 12257
rect 23845 12223 23903 12229
rect 23845 12220 23857 12223
rect 22848 12192 23857 12220
rect 23845 12189 23857 12192
rect 23891 12189 23903 12223
rect 23845 12183 23903 12189
rect 24029 12223 24087 12229
rect 24029 12189 24041 12223
rect 24075 12220 24087 12223
rect 24578 12220 24584 12232
rect 24075 12192 24584 12220
rect 24075 12189 24087 12192
rect 24029 12183 24087 12189
rect 24578 12180 24584 12192
rect 24636 12180 24642 12232
rect 24673 12223 24731 12229
rect 24673 12189 24685 12223
rect 24719 12220 24731 12223
rect 24854 12220 24860 12232
rect 24719 12192 24860 12220
rect 24719 12189 24731 12192
rect 24673 12183 24731 12189
rect 24854 12180 24860 12192
rect 24912 12180 24918 12232
rect 25225 12223 25283 12229
rect 25225 12189 25237 12223
rect 25271 12220 25283 12223
rect 25516 12220 25544 12316
rect 25792 12288 25820 12316
rect 25271 12192 25544 12220
rect 25608 12260 25820 12288
rect 25271 12189 25283 12192
rect 25225 12183 25283 12189
rect 19334 12152 19340 12164
rect 18248 12124 19340 12152
rect 16574 12084 16580 12096
rect 13648 12056 16580 12084
rect 16574 12044 16580 12056
rect 16632 12084 16638 12096
rect 17926 12084 17954 12124
rect 19334 12112 19340 12124
rect 19392 12112 19398 12164
rect 19426 12112 19432 12164
rect 19484 12112 19490 12164
rect 19610 12112 19616 12164
rect 19668 12112 19674 12164
rect 20990 12112 20996 12164
rect 21048 12152 21054 12164
rect 21634 12152 21640 12164
rect 21048 12124 21640 12152
rect 21048 12112 21054 12124
rect 21634 12112 21640 12124
rect 21692 12112 21698 12164
rect 21818 12112 21824 12164
rect 21876 12112 21882 12164
rect 22370 12112 22376 12164
rect 22428 12112 22434 12164
rect 23474 12112 23480 12164
rect 23532 12152 23538 12164
rect 24397 12155 24455 12161
rect 24397 12152 24409 12155
rect 23532 12124 24409 12152
rect 23532 12112 23538 12124
rect 24397 12121 24409 12124
rect 24443 12121 24455 12155
rect 24596 12152 24624 12180
rect 24949 12155 25007 12161
rect 24949 12152 24961 12155
rect 24596 12124 24961 12152
rect 24397 12115 24455 12121
rect 24949 12121 24961 12124
rect 24995 12121 25007 12155
rect 24949 12115 25007 12121
rect 25501 12155 25559 12161
rect 25501 12121 25513 12155
rect 25547 12152 25559 12155
rect 25608 12152 25636 12260
rect 25958 12248 25964 12300
rect 26016 12248 26022 12300
rect 25685 12223 25743 12229
rect 25685 12189 25697 12223
rect 25731 12189 25743 12223
rect 25685 12183 25743 12189
rect 25777 12223 25835 12229
rect 25777 12189 25789 12223
rect 25823 12220 25835 12223
rect 25976 12220 26004 12248
rect 25823 12192 26004 12220
rect 25823 12189 25835 12192
rect 25777 12183 25835 12189
rect 25547 12124 25636 12152
rect 25700 12152 25728 12183
rect 26142 12180 26148 12232
rect 26200 12220 26206 12232
rect 26697 12223 26755 12229
rect 26697 12220 26709 12223
rect 26200 12192 26709 12220
rect 26200 12180 26206 12192
rect 26697 12189 26709 12192
rect 26743 12189 26755 12223
rect 26697 12183 26755 12189
rect 26789 12223 26847 12229
rect 26789 12189 26801 12223
rect 26835 12189 26847 12223
rect 26896 12220 26924 12384
rect 27816 12356 27844 12384
rect 28902 12356 28908 12368
rect 27816 12328 28908 12356
rect 28902 12316 28908 12328
rect 28960 12316 28966 12368
rect 27154 12248 27160 12300
rect 27212 12288 27218 12300
rect 27801 12291 27859 12297
rect 27801 12288 27813 12291
rect 27212 12260 27813 12288
rect 27212 12248 27218 12260
rect 27801 12257 27813 12260
rect 27847 12257 27859 12291
rect 27801 12251 27859 12257
rect 28258 12248 28264 12300
rect 28316 12288 28322 12300
rect 28534 12288 28540 12300
rect 28316 12260 28540 12288
rect 28316 12248 28322 12260
rect 28534 12248 28540 12260
rect 28592 12248 28598 12300
rect 29914 12248 29920 12300
rect 29972 12288 29978 12300
rect 30193 12291 30251 12297
rect 30193 12288 30205 12291
rect 29972 12260 30205 12288
rect 29972 12248 29978 12260
rect 30193 12257 30205 12260
rect 30239 12257 30251 12291
rect 30193 12251 30251 12257
rect 27985 12223 28043 12229
rect 27985 12220 27997 12223
rect 26896 12192 27997 12220
rect 26789 12183 26847 12189
rect 27985 12189 27997 12192
rect 28031 12189 28043 12223
rect 30101 12223 30159 12229
rect 30101 12220 30113 12223
rect 27985 12183 28043 12189
rect 28092 12192 30113 12220
rect 25958 12152 25964 12164
rect 25700 12124 25964 12152
rect 25547 12121 25559 12124
rect 25501 12115 25559 12121
rect 25958 12112 25964 12124
rect 26016 12112 26022 12164
rect 26602 12112 26608 12164
rect 26660 12152 26666 12164
rect 26804 12152 26832 12183
rect 26660 12124 26832 12152
rect 27709 12155 27767 12161
rect 26660 12112 26666 12124
rect 27709 12121 27721 12155
rect 27755 12152 27767 12155
rect 27798 12152 27804 12164
rect 27755 12124 27804 12152
rect 27755 12121 27767 12124
rect 27709 12115 27767 12121
rect 27798 12112 27804 12124
rect 27856 12112 27862 12164
rect 16632 12056 17954 12084
rect 16632 12044 16638 12056
rect 18506 12044 18512 12096
rect 18564 12084 18570 12096
rect 19058 12084 19064 12096
rect 18564 12056 19064 12084
rect 18564 12044 18570 12056
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 19518 12044 19524 12096
rect 19576 12084 19582 12096
rect 22186 12084 22192 12096
rect 19576 12056 22192 12084
rect 19576 12044 19582 12056
rect 22186 12044 22192 12056
rect 22244 12044 22250 12096
rect 22281 12087 22339 12093
rect 22281 12053 22293 12087
rect 22327 12084 22339 12087
rect 22738 12084 22744 12096
rect 22327 12056 22744 12084
rect 22327 12053 22339 12056
rect 22281 12047 22339 12053
rect 22738 12044 22744 12056
rect 22796 12044 22802 12096
rect 22833 12087 22891 12093
rect 22833 12053 22845 12087
rect 22879 12084 22891 12087
rect 28092 12084 28120 12192
rect 30101 12189 30113 12192
rect 30147 12189 30159 12223
rect 30101 12183 30159 12189
rect 30926 12180 30932 12232
rect 30984 12180 30990 12232
rect 31297 12223 31355 12229
rect 31297 12189 31309 12223
rect 31343 12220 31355 12223
rect 31665 12223 31723 12229
rect 31665 12220 31677 12223
rect 31343 12192 31677 12220
rect 31343 12189 31355 12192
rect 31297 12183 31355 12189
rect 31665 12189 31677 12192
rect 31711 12189 31723 12223
rect 31665 12183 31723 12189
rect 32214 12180 32220 12232
rect 32272 12180 32278 12232
rect 30374 12112 30380 12164
rect 30432 12152 30438 12164
rect 30834 12152 30840 12164
rect 30432 12124 30840 12152
rect 30432 12112 30438 12124
rect 30834 12112 30840 12124
rect 30892 12152 30898 12164
rect 31113 12155 31171 12161
rect 31113 12152 31125 12155
rect 30892 12124 31125 12152
rect 30892 12112 30898 12124
rect 31113 12121 31125 12124
rect 31159 12121 31171 12155
rect 31113 12115 31171 12121
rect 31202 12112 31208 12164
rect 31260 12112 31266 12164
rect 22879 12056 28120 12084
rect 28169 12087 28227 12093
rect 22879 12053 22891 12056
rect 22833 12047 22891 12053
rect 28169 12053 28181 12087
rect 28215 12084 28227 12087
rect 28442 12084 28448 12096
rect 28215 12056 28448 12084
rect 28215 12053 28227 12056
rect 28169 12047 28227 12053
rect 28442 12044 28448 12056
rect 28500 12044 28506 12096
rect 30466 12044 30472 12096
rect 30524 12044 30530 12096
rect 30650 12044 30656 12096
rect 30708 12084 30714 12096
rect 31220 12084 31248 12112
rect 30708 12056 31248 12084
rect 30708 12044 30714 12056
rect 31478 12044 31484 12096
rect 31536 12044 31542 12096
rect 1104 11994 32844 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 32844 11994
rect 1104 11920 32844 11942
rect 3237 11883 3295 11889
rect 3237 11849 3249 11883
rect 3283 11880 3295 11883
rect 3510 11880 3516 11892
rect 3283 11852 3516 11880
rect 3283 11849 3295 11852
rect 3237 11843 3295 11849
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 4249 11883 4307 11889
rect 4249 11849 4261 11883
rect 4295 11880 4307 11883
rect 4338 11880 4344 11892
rect 4295 11852 4344 11880
rect 4295 11849 4307 11852
rect 4249 11843 4307 11849
rect 2130 11704 2136 11756
rect 2188 11744 2194 11756
rect 2777 11747 2835 11753
rect 2777 11744 2789 11747
rect 2188 11716 2789 11744
rect 2188 11704 2194 11716
rect 2777 11713 2789 11716
rect 2823 11713 2835 11747
rect 2777 11707 2835 11713
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11744 3111 11747
rect 3326 11744 3332 11756
rect 3099 11716 3332 11744
rect 3099 11713 3111 11716
rect 3053 11707 3111 11713
rect 3326 11704 3332 11716
rect 3384 11704 3390 11756
rect 3510 11704 3516 11756
rect 3568 11704 3574 11756
rect 3602 11704 3608 11756
rect 3660 11744 3666 11756
rect 3789 11747 3847 11753
rect 3789 11744 3801 11747
rect 3660 11716 3801 11744
rect 3660 11704 3666 11716
rect 3789 11713 3801 11716
rect 3835 11713 3847 11747
rect 3789 11707 3847 11713
rect 4157 11747 4215 11753
rect 4157 11713 4169 11747
rect 4203 11744 4215 11747
rect 4264 11744 4292 11843
rect 4338 11840 4344 11852
rect 4396 11840 4402 11892
rect 5350 11880 5356 11892
rect 4632 11852 5356 11880
rect 4203 11716 4292 11744
rect 4203 11713 4215 11716
rect 4157 11707 4215 11713
rect 4430 11704 4436 11756
rect 4488 11704 4494 11756
rect 4632 11753 4660 11852
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 5626 11840 5632 11892
rect 5684 11840 5690 11892
rect 5718 11840 5724 11892
rect 5776 11880 5782 11892
rect 7006 11880 7012 11892
rect 5776 11852 6684 11880
rect 5776 11840 5782 11852
rect 5644 11812 5672 11840
rect 6454 11812 6460 11824
rect 4715 11784 5396 11812
rect 5644 11784 6460 11812
rect 4617 11747 4675 11753
rect 4617 11713 4629 11747
rect 4663 11713 4675 11747
rect 4617 11707 4675 11713
rect 3418 11636 3424 11688
rect 3476 11676 3482 11688
rect 4715 11676 4743 11784
rect 5368 11756 5396 11784
rect 6454 11772 6460 11784
rect 6512 11772 6518 11824
rect 6656 11812 6684 11852
rect 6840 11852 7012 11880
rect 6840 11812 6868 11852
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 7469 11883 7527 11889
rect 7469 11849 7481 11883
rect 7515 11880 7527 11883
rect 7834 11880 7840 11892
rect 7515 11852 7840 11880
rect 7515 11849 7527 11852
rect 7469 11843 7527 11849
rect 7834 11840 7840 11852
rect 7892 11880 7898 11892
rect 9217 11883 9275 11889
rect 7892 11852 8984 11880
rect 7892 11840 7898 11852
rect 6656 11784 6868 11812
rect 6917 11815 6975 11821
rect 6917 11781 6929 11815
rect 6963 11812 6975 11815
rect 7190 11812 7196 11824
rect 6963 11784 7196 11812
rect 6963 11781 6975 11784
rect 6917 11775 6975 11781
rect 7190 11772 7196 11784
rect 7248 11772 7254 11824
rect 7650 11772 7656 11824
rect 7708 11812 7714 11824
rect 8205 11815 8263 11821
rect 8205 11812 8217 11815
rect 7708 11784 8217 11812
rect 7708 11772 7714 11784
rect 8205 11781 8217 11784
rect 8251 11781 8263 11815
rect 8205 11775 8263 11781
rect 4798 11704 4804 11756
rect 4856 11744 4862 11756
rect 5169 11747 5227 11753
rect 5169 11744 5181 11747
rect 4856 11716 5181 11744
rect 4856 11704 4862 11716
rect 5169 11713 5181 11716
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 5350 11704 5356 11756
rect 5408 11744 5414 11756
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 5408 11716 5457 11744
rect 5408 11704 5414 11716
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 5626 11704 5632 11756
rect 5684 11744 5690 11756
rect 6157 11747 6215 11753
rect 6157 11744 6169 11747
rect 5684 11716 6169 11744
rect 5684 11704 5690 11716
rect 6157 11713 6169 11716
rect 6203 11713 6215 11747
rect 6157 11707 6215 11713
rect 6270 11704 6276 11756
rect 6328 11744 6334 11756
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 6328 11716 6561 11744
rect 6328 11704 6334 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 7006 11704 7012 11756
rect 7064 11744 7070 11756
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 7064 11716 7297 11744
rect 7064 11704 7070 11716
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 8757 11747 8815 11753
rect 8757 11713 8769 11747
rect 8803 11713 8815 11747
rect 8757 11707 8815 11713
rect 3476 11648 4743 11676
rect 6380 11648 8524 11676
rect 3476 11636 3482 11648
rect 1854 11568 1860 11620
rect 1912 11608 1918 11620
rect 3050 11608 3056 11620
rect 1912 11580 3056 11608
rect 1912 11568 1918 11580
rect 3050 11568 3056 11580
rect 3108 11568 3114 11620
rect 3142 11568 3148 11620
rect 3200 11608 3206 11620
rect 3200 11580 3464 11608
rect 3200 11568 3206 11580
rect 2498 11500 2504 11552
rect 2556 11540 2562 11552
rect 2774 11540 2780 11552
rect 2556 11512 2780 11540
rect 2556 11500 2562 11512
rect 2774 11500 2780 11512
rect 2832 11500 2838 11552
rect 2958 11500 2964 11552
rect 3016 11500 3022 11552
rect 3326 11500 3332 11552
rect 3384 11500 3390 11552
rect 3436 11540 3464 11580
rect 3510 11568 3516 11620
rect 3568 11608 3574 11620
rect 3605 11611 3663 11617
rect 3605 11608 3617 11611
rect 3568 11580 3617 11608
rect 3568 11568 3574 11580
rect 3605 11577 3617 11580
rect 3651 11577 3663 11611
rect 3605 11571 3663 11577
rect 4801 11611 4859 11617
rect 4801 11577 4813 11611
rect 4847 11608 4859 11611
rect 5902 11608 5908 11620
rect 4847 11580 5908 11608
rect 4847 11577 4859 11580
rect 4801 11571 4859 11577
rect 5902 11568 5908 11580
rect 5960 11608 5966 11620
rect 6380 11608 6408 11648
rect 5960 11580 6408 11608
rect 5960 11568 5966 11580
rect 3973 11543 4031 11549
rect 3973 11540 3985 11543
rect 3436 11512 3985 11540
rect 3973 11509 3985 11512
rect 4019 11509 4031 11543
rect 3973 11503 4031 11509
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 4985 11543 5043 11549
rect 4985 11540 4997 11543
rect 4120 11512 4997 11540
rect 4120 11500 4126 11512
rect 4985 11509 4997 11512
rect 5031 11509 5043 11543
rect 4985 11503 5043 11509
rect 5074 11500 5080 11552
rect 5132 11540 5138 11552
rect 5261 11543 5319 11549
rect 5261 11540 5273 11543
rect 5132 11512 5273 11540
rect 5132 11500 5138 11512
rect 5261 11509 5273 11512
rect 5307 11509 5319 11543
rect 5261 11503 5319 11509
rect 5994 11500 6000 11552
rect 6052 11500 6058 11552
rect 6380 11540 6408 11580
rect 6454 11568 6460 11620
rect 6512 11608 6518 11620
rect 7190 11608 7196 11620
rect 6512 11580 7196 11608
rect 6512 11568 6518 11580
rect 7190 11568 7196 11580
rect 7248 11568 7254 11620
rect 8496 11617 8524 11648
rect 8481 11611 8539 11617
rect 8481 11577 8493 11611
rect 8527 11577 8539 11611
rect 8772 11608 8800 11707
rect 8956 11685 8984 11852
rect 9217 11849 9229 11883
rect 9263 11880 9275 11883
rect 9950 11880 9956 11892
rect 9263 11852 9956 11880
rect 9263 11849 9275 11852
rect 9217 11843 9275 11849
rect 9950 11840 9956 11852
rect 10008 11840 10014 11892
rect 10226 11840 10232 11892
rect 10284 11880 10290 11892
rect 10873 11883 10931 11889
rect 10284 11852 10824 11880
rect 10284 11840 10290 11852
rect 10502 11812 10508 11824
rect 9048 11784 10508 11812
rect 9048 11753 9076 11784
rect 10502 11772 10508 11784
rect 10560 11772 10566 11824
rect 9033 11747 9091 11753
rect 9033 11713 9045 11747
rect 9079 11713 9091 11747
rect 9033 11707 9091 11713
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 10042 11744 10048 11756
rect 9640 11716 10048 11744
rect 9640 11704 9646 11716
rect 10042 11704 10048 11716
rect 10100 11704 10106 11756
rect 10410 11704 10416 11756
rect 10468 11744 10474 11756
rect 10597 11747 10655 11753
rect 10597 11744 10609 11747
rect 10468 11716 10609 11744
rect 10468 11704 10474 11716
rect 10597 11713 10609 11716
rect 10643 11713 10655 11747
rect 10597 11707 10655 11713
rect 10689 11747 10747 11753
rect 10689 11713 10701 11747
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 8941 11679 8999 11685
rect 8941 11645 8953 11679
rect 8987 11676 8999 11679
rect 9674 11676 9680 11688
rect 8987 11648 9680 11676
rect 8987 11645 8999 11648
rect 8941 11639 8999 11645
rect 9674 11636 9680 11648
rect 9732 11636 9738 11688
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 10704 11676 10732 11707
rect 10008 11648 10732 11676
rect 10796 11676 10824 11852
rect 10873 11849 10885 11883
rect 10919 11880 10931 11883
rect 10962 11880 10968 11892
rect 10919 11852 10968 11880
rect 10919 11849 10931 11852
rect 10873 11843 10931 11849
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 11146 11840 11152 11892
rect 11204 11880 11210 11892
rect 12802 11880 12808 11892
rect 11204 11852 12808 11880
rect 11204 11840 11210 11852
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 13722 11840 13728 11892
rect 13780 11880 13786 11892
rect 13780 11852 14872 11880
rect 13780 11840 13786 11852
rect 10980 11753 11008 11840
rect 11072 11784 12480 11812
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 11072 11676 11100 11784
rect 11422 11704 11428 11756
rect 11480 11744 11486 11756
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 11480 11716 11529 11744
rect 11480 11704 11486 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11790 11704 11796 11756
rect 11848 11704 11854 11756
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11744 12219 11747
rect 12250 11744 12256 11756
rect 12207 11716 12256 11744
rect 12207 11713 12219 11716
rect 12161 11707 12219 11713
rect 12250 11704 12256 11716
rect 12308 11704 12314 11756
rect 12342 11704 12348 11756
rect 12400 11704 12406 11756
rect 12452 11744 12480 11784
rect 12618 11772 12624 11824
rect 12676 11812 12682 11824
rect 12676 11784 13216 11812
rect 12676 11772 12682 11784
rect 12897 11747 12955 11753
rect 12897 11744 12909 11747
rect 12452 11716 12909 11744
rect 12897 11713 12909 11716
rect 12943 11744 12955 11747
rect 13078 11744 13084 11756
rect 12943 11716 13084 11744
rect 12943 11713 12955 11716
rect 12897 11707 12955 11713
rect 13078 11704 13084 11716
rect 13136 11704 13142 11756
rect 13188 11753 13216 11784
rect 14090 11772 14096 11824
rect 14148 11812 14154 11824
rect 14550 11812 14556 11824
rect 14148 11784 14556 11812
rect 14148 11772 14154 11784
rect 14550 11772 14556 11784
rect 14608 11812 14614 11824
rect 14737 11815 14795 11821
rect 14737 11812 14749 11815
rect 14608 11784 14749 11812
rect 14608 11772 14614 11784
rect 14737 11781 14749 11784
rect 14783 11781 14795 11815
rect 14844 11812 14872 11852
rect 15102 11840 15108 11892
rect 15160 11880 15166 11892
rect 15160 11852 17080 11880
rect 15160 11840 15166 11852
rect 15197 11815 15255 11821
rect 14844 11784 15148 11812
rect 14737 11775 14795 11781
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 13354 11704 13360 11756
rect 13412 11744 13418 11756
rect 14461 11747 14519 11753
rect 14461 11744 14473 11747
rect 13412 11716 14473 11744
rect 13412 11704 13418 11716
rect 14461 11713 14473 11716
rect 14507 11713 14519 11747
rect 14461 11707 14519 11713
rect 14826 11704 14832 11756
rect 14884 11704 14890 11756
rect 15010 11704 15016 11756
rect 15068 11704 15074 11756
rect 15120 11744 15148 11784
rect 15197 11781 15209 11815
rect 15243 11812 15255 11815
rect 15470 11812 15476 11824
rect 15243 11784 15476 11812
rect 15243 11781 15255 11784
rect 15197 11775 15255 11781
rect 15470 11772 15476 11784
rect 15528 11772 15534 11824
rect 16114 11772 16120 11824
rect 16172 11812 16178 11824
rect 17052 11812 17080 11852
rect 17126 11840 17132 11892
rect 17184 11840 17190 11892
rect 17494 11840 17500 11892
rect 17552 11840 17558 11892
rect 17954 11840 17960 11892
rect 18012 11840 18018 11892
rect 18064 11852 18828 11880
rect 16172 11784 16988 11812
rect 17052 11784 17724 11812
rect 16172 11772 16178 11784
rect 16390 11744 16396 11756
rect 15120 11716 16396 11744
rect 16390 11704 16396 11716
rect 16448 11704 16454 11756
rect 16960 11753 16988 11784
rect 16669 11747 16727 11753
rect 16669 11713 16681 11747
rect 16715 11713 16727 11747
rect 16669 11707 16727 11713
rect 16945 11747 17003 11753
rect 16945 11713 16957 11747
rect 16991 11713 17003 11747
rect 16945 11707 17003 11713
rect 10796 11648 11100 11676
rect 10008 11636 10014 11648
rect 11606 11636 11612 11688
rect 11664 11676 11670 11688
rect 12066 11676 12072 11688
rect 11664 11648 12072 11676
rect 11664 11636 11670 11648
rect 12066 11636 12072 11648
rect 12124 11636 12130 11688
rect 12986 11636 12992 11688
rect 13044 11636 13050 11688
rect 14645 11679 14703 11685
rect 14645 11645 14657 11679
rect 14691 11676 14703 11679
rect 15470 11676 15476 11688
rect 14691 11648 15476 11676
rect 14691 11645 14703 11648
rect 14645 11639 14703 11645
rect 15470 11636 15476 11648
rect 15528 11636 15534 11688
rect 16298 11636 16304 11688
rect 16356 11676 16362 11688
rect 16684 11676 16712 11707
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 17696 11753 17724 11784
rect 17862 11772 17868 11824
rect 17920 11812 17926 11824
rect 18064 11812 18092 11852
rect 17920 11784 18092 11812
rect 18141 11815 18199 11821
rect 17920 11772 17926 11784
rect 18141 11781 18153 11815
rect 18187 11812 18199 11815
rect 18322 11812 18328 11824
rect 18187 11784 18328 11812
rect 18187 11781 18199 11784
rect 18141 11775 18199 11781
rect 18322 11772 18328 11784
rect 18380 11772 18386 11824
rect 17681 11747 17739 11753
rect 17092 11716 17356 11744
rect 17092 11704 17098 11716
rect 16356 11648 16712 11676
rect 16853 11679 16911 11685
rect 16356 11636 16362 11648
rect 16853 11645 16865 11679
rect 16899 11676 16911 11679
rect 17218 11676 17224 11688
rect 16899 11648 17224 11676
rect 16899 11645 16911 11648
rect 16853 11639 16911 11645
rect 17218 11636 17224 11648
rect 17276 11636 17282 11688
rect 17328 11676 17356 11716
rect 17681 11713 17693 11747
rect 17727 11713 17739 11747
rect 17681 11707 17739 11713
rect 18417 11747 18475 11753
rect 18417 11713 18429 11747
rect 18463 11744 18475 11747
rect 18506 11744 18512 11756
rect 18463 11716 18512 11744
rect 18463 11713 18475 11716
rect 18417 11707 18475 11713
rect 18506 11704 18512 11716
rect 18564 11704 18570 11756
rect 18693 11747 18751 11753
rect 18693 11713 18705 11747
rect 18739 11713 18751 11747
rect 18800 11744 18828 11852
rect 19058 11840 19064 11892
rect 19116 11840 19122 11892
rect 20714 11840 20720 11892
rect 20772 11840 20778 11892
rect 20993 11883 21051 11889
rect 20993 11849 21005 11883
rect 21039 11880 21051 11883
rect 21358 11880 21364 11892
rect 21039 11852 21364 11880
rect 21039 11849 21051 11852
rect 20993 11843 21051 11849
rect 19889 11815 19947 11821
rect 19889 11781 19901 11815
rect 19935 11812 19947 11815
rect 21008 11812 21036 11843
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 21542 11840 21548 11892
rect 21600 11880 21606 11892
rect 21600 11852 24256 11880
rect 21600 11840 21606 11852
rect 19935 11784 21036 11812
rect 19935 11781 19947 11784
rect 19889 11775 19947 11781
rect 24118 11772 24124 11824
rect 24176 11772 24182 11824
rect 24228 11812 24256 11852
rect 24854 11840 24860 11892
rect 24912 11880 24918 11892
rect 29178 11880 29184 11892
rect 24912 11852 29184 11880
rect 24912 11840 24918 11852
rect 29178 11840 29184 11852
rect 29236 11840 29242 11892
rect 31941 11883 31999 11889
rect 31941 11849 31953 11883
rect 31987 11880 31999 11883
rect 32214 11880 32220 11892
rect 31987 11852 32220 11880
rect 31987 11849 31999 11852
rect 31941 11843 31999 11849
rect 32214 11840 32220 11852
rect 32272 11840 32278 11892
rect 25590 11812 25596 11824
rect 24228 11784 25596 11812
rect 25590 11772 25596 11784
rect 25648 11812 25654 11824
rect 27154 11812 27160 11824
rect 25648 11784 27160 11812
rect 25648 11772 25654 11784
rect 27154 11772 27160 11784
rect 27212 11772 27218 11824
rect 28534 11772 28540 11824
rect 28592 11812 28598 11824
rect 28592 11784 29132 11812
rect 28592 11772 28598 11784
rect 19705 11747 19763 11753
rect 19705 11744 19717 11747
rect 18800 11716 19717 11744
rect 18693 11707 18751 11713
rect 19705 11713 19717 11716
rect 19751 11713 19763 11747
rect 19705 11707 19763 11713
rect 17862 11676 17868 11688
rect 17328 11648 17868 11676
rect 17862 11636 17868 11648
rect 17920 11636 17926 11688
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 18233 11679 18291 11685
rect 18233 11676 18245 11679
rect 18012 11648 18245 11676
rect 18012 11636 18018 11648
rect 18233 11645 18245 11648
rect 18279 11645 18291 11679
rect 18233 11639 18291 11645
rect 10686 11608 10692 11620
rect 8772 11580 10692 11608
rect 8481 11571 8539 11577
rect 10686 11568 10692 11580
rect 10744 11568 10750 11620
rect 12250 11608 12256 11620
rect 12084 11580 12256 11608
rect 6546 11540 6552 11552
rect 6380 11512 6552 11540
rect 6546 11500 6552 11512
rect 6604 11500 6610 11552
rect 6730 11500 6736 11552
rect 6788 11500 6794 11552
rect 7282 11500 7288 11552
rect 7340 11540 7346 11552
rect 7834 11540 7840 11552
rect 7340 11512 7840 11540
rect 7340 11500 7346 11512
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 8018 11500 8024 11552
rect 8076 11540 8082 11552
rect 8202 11540 8208 11552
rect 8076 11512 8208 11540
rect 8076 11500 8082 11512
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8662 11500 8668 11552
rect 8720 11500 8726 11552
rect 9033 11543 9091 11549
rect 9033 11509 9045 11543
rect 9079 11540 9091 11543
rect 9122 11540 9128 11552
rect 9079 11512 9128 11540
rect 9079 11509 9091 11512
rect 9033 11503 9091 11509
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 9674 11500 9680 11552
rect 9732 11540 9738 11552
rect 9950 11540 9956 11552
rect 9732 11512 9956 11540
rect 9732 11500 9738 11512
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 10410 11500 10416 11552
rect 10468 11500 10474 11552
rect 10502 11500 10508 11552
rect 10560 11540 10566 11552
rect 11146 11540 11152 11552
rect 10560 11512 11152 11540
rect 10560 11500 10566 11512
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 11238 11500 11244 11552
rect 11296 11540 11302 11552
rect 11517 11543 11575 11549
rect 11517 11540 11529 11543
rect 11296 11512 11529 11540
rect 11296 11500 11302 11512
rect 11517 11509 11529 11512
rect 11563 11540 11575 11543
rect 11882 11540 11888 11552
rect 11563 11512 11888 11540
rect 11563 11509 11575 11512
rect 11517 11503 11575 11509
rect 11882 11500 11888 11512
rect 11940 11500 11946 11552
rect 11977 11543 12035 11549
rect 11977 11509 11989 11543
rect 12023 11540 12035 11543
rect 12084 11540 12112 11580
rect 12250 11568 12256 11580
rect 12308 11568 12314 11620
rect 12529 11611 12587 11617
rect 12529 11577 12541 11611
rect 12575 11608 12587 11611
rect 17310 11608 17316 11620
rect 12575 11580 17316 11608
rect 12575 11577 12587 11580
rect 12529 11571 12587 11577
rect 17310 11568 17316 11580
rect 17368 11568 17374 11620
rect 17402 11568 17408 11620
rect 17460 11608 17466 11620
rect 18708 11608 18736 11707
rect 20346 11704 20352 11756
rect 20404 11704 20410 11756
rect 20530 11704 20536 11756
rect 20588 11704 20594 11756
rect 20622 11704 20628 11756
rect 20680 11744 20686 11756
rect 20809 11747 20867 11753
rect 20809 11744 20821 11747
rect 20680 11716 20821 11744
rect 20680 11704 20686 11716
rect 20809 11713 20821 11716
rect 20855 11713 20867 11747
rect 20809 11707 20867 11713
rect 23937 11747 23995 11753
rect 23937 11713 23949 11747
rect 23983 11744 23995 11747
rect 25038 11744 25044 11756
rect 23983 11716 25044 11744
rect 23983 11713 23995 11716
rect 23937 11707 23995 11713
rect 25038 11704 25044 11716
rect 25096 11704 25102 11756
rect 25314 11704 25320 11756
rect 25372 11744 25378 11756
rect 25774 11744 25780 11756
rect 25372 11716 25780 11744
rect 25372 11704 25378 11716
rect 25774 11704 25780 11716
rect 25832 11704 25838 11756
rect 28074 11704 28080 11756
rect 28132 11744 28138 11756
rect 28445 11747 28503 11753
rect 28445 11744 28457 11747
rect 28132 11716 28457 11744
rect 28132 11704 28138 11716
rect 28445 11713 28457 11716
rect 28491 11713 28503 11747
rect 28445 11707 28503 11713
rect 28626 11704 28632 11756
rect 28684 11704 28690 11756
rect 28718 11704 28724 11756
rect 28776 11704 28782 11756
rect 29104 11744 29132 11784
rect 29362 11772 29368 11824
rect 29420 11812 29426 11824
rect 29549 11815 29607 11821
rect 29549 11812 29561 11815
rect 29420 11784 29561 11812
rect 29420 11772 29426 11784
rect 29549 11781 29561 11784
rect 29595 11781 29607 11815
rect 29549 11775 29607 11781
rect 30828 11815 30886 11821
rect 30828 11781 30840 11815
rect 30874 11812 30886 11815
rect 31478 11812 31484 11824
rect 30874 11784 31484 11812
rect 30874 11781 30886 11784
rect 30828 11775 30886 11781
rect 31478 11772 31484 11784
rect 31536 11772 31542 11824
rect 29825 11747 29883 11753
rect 29825 11744 29837 11747
rect 29104 11716 29837 11744
rect 29825 11713 29837 11716
rect 29871 11713 29883 11747
rect 29825 11707 29883 11713
rect 32214 11704 32220 11756
rect 32272 11704 32278 11756
rect 18785 11679 18843 11685
rect 18785 11645 18797 11679
rect 18831 11676 18843 11679
rect 19334 11676 19340 11688
rect 18831 11648 19340 11676
rect 18831 11645 18843 11648
rect 18785 11639 18843 11645
rect 19334 11636 19340 11648
rect 19392 11636 19398 11688
rect 20548 11608 20576 11704
rect 21634 11636 21640 11688
rect 21692 11676 21698 11688
rect 22370 11676 22376 11688
rect 21692 11648 22376 11676
rect 21692 11636 21698 11648
rect 22370 11636 22376 11648
rect 22428 11636 22434 11688
rect 22738 11636 22744 11688
rect 22796 11676 22802 11688
rect 29641 11679 29699 11685
rect 29641 11676 29653 11679
rect 22796 11648 29653 11676
rect 22796 11636 22802 11648
rect 29641 11645 29653 11648
rect 29687 11645 29699 11679
rect 29641 11639 29699 11645
rect 30558 11636 30564 11688
rect 30616 11636 30622 11688
rect 22002 11608 22008 11620
rect 17460 11580 18736 11608
rect 18800 11580 20576 11608
rect 21284 11580 22008 11608
rect 17460 11568 17466 11580
rect 18800 11552 18828 11580
rect 12023 11512 12112 11540
rect 12023 11509 12035 11512
rect 11977 11503 12035 11509
rect 12158 11500 12164 11552
rect 12216 11500 12222 11552
rect 12894 11500 12900 11552
rect 12952 11500 12958 11552
rect 13354 11500 13360 11552
rect 13412 11500 13418 11552
rect 14274 11500 14280 11552
rect 14332 11500 14338 11552
rect 14734 11500 14740 11552
rect 14792 11500 14798 11552
rect 15470 11500 15476 11552
rect 15528 11540 15534 11552
rect 16482 11540 16488 11552
rect 15528 11512 16488 11540
rect 15528 11500 15534 11512
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 16758 11500 16764 11552
rect 16816 11500 16822 11552
rect 16850 11500 16856 11552
rect 16908 11540 16914 11552
rect 18141 11543 18199 11549
rect 18141 11540 18153 11543
rect 16908 11512 18153 11540
rect 16908 11500 16914 11512
rect 18141 11509 18153 11512
rect 18187 11509 18199 11543
rect 18141 11503 18199 11509
rect 18598 11500 18604 11552
rect 18656 11500 18662 11552
rect 18690 11500 18696 11552
rect 18748 11500 18754 11552
rect 18782 11500 18788 11552
rect 18840 11500 18846 11552
rect 20073 11543 20131 11549
rect 20073 11509 20085 11543
rect 20119 11540 20131 11543
rect 20530 11540 20536 11552
rect 20119 11512 20536 11540
rect 20119 11509 20131 11512
rect 20073 11503 20131 11509
rect 20530 11500 20536 11512
rect 20588 11540 20594 11552
rect 21284 11540 21312 11580
rect 22002 11568 22008 11580
rect 22060 11568 22066 11620
rect 23290 11568 23296 11620
rect 23348 11608 23354 11620
rect 25958 11608 25964 11620
rect 23348 11580 25964 11608
rect 23348 11568 23354 11580
rect 25958 11568 25964 11580
rect 26016 11568 26022 11620
rect 30466 11608 30472 11620
rect 29840 11580 30472 11608
rect 20588 11512 21312 11540
rect 20588 11500 20594 11512
rect 21358 11500 21364 11552
rect 21416 11540 21422 11552
rect 23474 11540 23480 11552
rect 21416 11512 23480 11540
rect 21416 11500 21422 11512
rect 23474 11500 23480 11512
rect 23532 11500 23538 11552
rect 23753 11543 23811 11549
rect 23753 11509 23765 11543
rect 23799 11540 23811 11543
rect 24026 11540 24032 11552
rect 23799 11512 24032 11540
rect 23799 11509 23811 11512
rect 23753 11503 23811 11509
rect 24026 11500 24032 11512
rect 24084 11540 24090 11552
rect 24486 11540 24492 11552
rect 24084 11512 24492 11540
rect 24084 11500 24090 11512
rect 24486 11500 24492 11512
rect 24544 11500 24550 11552
rect 24762 11500 24768 11552
rect 24820 11540 24826 11552
rect 26786 11540 26792 11552
rect 24820 11512 26792 11540
rect 24820 11500 24826 11512
rect 26786 11500 26792 11512
rect 26844 11500 26850 11552
rect 28442 11500 28448 11552
rect 28500 11500 28506 11552
rect 28905 11543 28963 11549
rect 28905 11509 28917 11543
rect 28951 11540 28963 11543
rect 29086 11540 29092 11552
rect 28951 11512 29092 11540
rect 28951 11509 28963 11512
rect 28905 11503 28963 11509
rect 29086 11500 29092 11512
rect 29144 11500 29150 11552
rect 29840 11549 29868 11580
rect 30466 11568 30472 11580
rect 30524 11568 30530 11620
rect 29825 11543 29883 11549
rect 29825 11509 29837 11543
rect 29871 11509 29883 11543
rect 29825 11503 29883 11509
rect 30006 11500 30012 11552
rect 30064 11500 30070 11552
rect 30576 11540 30604 11636
rect 32398 11568 32404 11620
rect 32456 11568 32462 11620
rect 30834 11540 30840 11552
rect 30576 11512 30840 11540
rect 30834 11500 30840 11512
rect 30892 11500 30898 11552
rect 1104 11450 32844 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 32844 11450
rect 1104 11376 32844 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 1670 11336 1676 11348
rect 1627 11308 1676 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 3602 11336 3608 11348
rect 2792 11308 3608 11336
rect 2498 11200 2504 11212
rect 1964 11172 2504 11200
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 1964 11141 1992 11172
rect 2498 11160 2504 11172
rect 2556 11200 2562 11212
rect 2792 11200 2820 11308
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 4709 11339 4767 11345
rect 4172 11308 4476 11336
rect 2866 11228 2872 11280
rect 2924 11268 2930 11280
rect 3145 11271 3203 11277
rect 3145 11268 3157 11271
rect 2924 11240 3157 11268
rect 2924 11228 2930 11240
rect 3145 11237 3157 11240
rect 3191 11237 3203 11271
rect 3145 11231 3203 11237
rect 3418 11228 3424 11280
rect 3476 11268 3482 11280
rect 4065 11271 4123 11277
rect 4065 11268 4077 11271
rect 3476 11240 4077 11268
rect 3476 11228 3482 11240
rect 4065 11237 4077 11240
rect 4111 11237 4123 11271
rect 4065 11231 4123 11237
rect 4172 11200 4200 11308
rect 4448 11268 4476 11308
rect 4709 11305 4721 11339
rect 4755 11336 4767 11339
rect 6270 11336 6276 11348
rect 4755 11308 6276 11336
rect 4755 11305 4767 11308
rect 4709 11299 4767 11305
rect 6270 11296 6276 11308
rect 6328 11296 6334 11348
rect 6362 11296 6368 11348
rect 6420 11296 6426 11348
rect 6822 11296 6828 11348
rect 6880 11336 6886 11348
rect 6880 11308 6960 11336
rect 6880 11296 6886 11308
rect 4448 11240 5396 11268
rect 2556 11172 2820 11200
rect 2556 11160 2562 11172
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11101 2007 11135
rect 1949 11095 2007 11101
rect 2130 11092 2136 11144
rect 2188 11092 2194 11144
rect 2222 11092 2228 11144
rect 2280 11092 2286 11144
rect 2317 11135 2375 11141
rect 2317 11101 2329 11135
rect 2363 11101 2375 11135
rect 2317 11095 2375 11101
rect 2593 11135 2651 11141
rect 2593 11101 2605 11135
rect 2639 11132 2651 11135
rect 2792 11132 2820 11172
rect 2884 11172 4200 11200
rect 2884 11144 2912 11172
rect 4246 11160 4252 11212
rect 4304 11200 4310 11212
rect 4304 11172 5120 11200
rect 4304 11160 4310 11172
rect 2639 11104 2820 11132
rect 2639 11101 2651 11104
rect 2593 11095 2651 11101
rect 2332 11064 2360 11095
rect 2866 11092 2872 11144
rect 2924 11092 2930 11144
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11132 3019 11135
rect 3326 11132 3332 11144
rect 3007 11104 3332 11132
rect 3007 11101 3019 11104
rect 2961 11095 3019 11101
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11132 3479 11135
rect 3510 11132 3516 11144
rect 3467 11104 3516 11132
rect 3467 11101 3479 11104
rect 3421 11095 3479 11101
rect 2682 11064 2688 11076
rect 2332 11036 2688 11064
rect 2682 11024 2688 11036
rect 2740 11024 2746 11076
rect 2777 11067 2835 11073
rect 2777 11033 2789 11067
rect 2823 11064 2835 11067
rect 3436 11064 3464 11095
rect 3510 11092 3516 11104
rect 3568 11092 3574 11144
rect 3881 11135 3939 11141
rect 3881 11132 3893 11135
rect 3620 11104 3893 11132
rect 3620 11064 3648 11104
rect 3881 11101 3893 11104
rect 3927 11101 3939 11135
rect 3881 11095 3939 11101
rect 4154 11092 4160 11144
rect 4212 11092 4218 11144
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11132 4583 11135
rect 4614 11132 4620 11144
rect 4571 11104 4620 11132
rect 4571 11101 4583 11104
rect 4525 11095 4583 11101
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 5092 11141 5120 11172
rect 5368 11141 5396 11240
rect 6380 11200 6408 11296
rect 6546 11228 6552 11280
rect 6604 11268 6610 11280
rect 6604 11240 6776 11268
rect 6604 11228 6610 11240
rect 6380 11172 6592 11200
rect 4985 11135 5043 11141
rect 4985 11132 4997 11135
rect 4816 11104 4997 11132
rect 2823 11036 3464 11064
rect 3528 11036 3648 11064
rect 2823 11033 2835 11036
rect 2777 11027 2835 11033
rect 2498 10956 2504 11008
rect 2556 10956 2562 11008
rect 3050 10956 3056 11008
rect 3108 10996 3114 11008
rect 3528 10996 3556 11036
rect 3694 11024 3700 11076
rect 3752 11064 3758 11076
rect 4246 11064 4252 11076
rect 3752 11036 4252 11064
rect 3752 11024 3758 11036
rect 4246 11024 4252 11036
rect 4304 11024 4310 11076
rect 4341 11067 4399 11073
rect 4341 11033 4353 11067
rect 4387 11033 4399 11067
rect 4341 11027 4399 11033
rect 3108 10968 3556 10996
rect 3605 10999 3663 11005
rect 3108 10956 3114 10968
rect 3605 10965 3617 10999
rect 3651 10996 3663 10999
rect 3970 10996 3976 11008
rect 3651 10968 3976 10996
rect 3651 10965 3663 10968
rect 3605 10959 3663 10965
rect 3970 10956 3976 10968
rect 4028 10956 4034 11008
rect 4356 10996 4384 11027
rect 4430 11024 4436 11076
rect 4488 11024 4494 11076
rect 4816 11064 4844 11104
rect 4985 11101 4997 11104
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11101 5135 11135
rect 5077 11095 5135 11101
rect 5353 11135 5411 11141
rect 5353 11101 5365 11135
rect 5399 11101 5411 11135
rect 5353 11095 5411 11101
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11132 5503 11135
rect 5626 11132 5632 11144
rect 5491 11104 5632 11132
rect 5491 11101 5503 11104
rect 5445 11095 5503 11101
rect 5626 11092 5632 11104
rect 5684 11092 5690 11144
rect 5905 11135 5963 11141
rect 5905 11101 5917 11135
rect 5951 11101 5963 11135
rect 5905 11095 5963 11101
rect 4724 11036 4844 11064
rect 4724 11008 4752 11036
rect 5258 11024 5264 11076
rect 5316 11024 5322 11076
rect 5810 11064 5816 11076
rect 5644 11036 5816 11064
rect 4522 10996 4528 11008
rect 4356 10968 4528 10996
rect 4522 10956 4528 10968
rect 4580 10956 4586 11008
rect 4706 10956 4712 11008
rect 4764 10956 4770 11008
rect 4801 10999 4859 11005
rect 4801 10965 4813 10999
rect 4847 10996 4859 10999
rect 4890 10996 4896 11008
rect 4847 10968 4896 10996
rect 4847 10965 4859 10968
rect 4801 10959 4859 10965
rect 4890 10956 4896 10968
rect 4948 10996 4954 11008
rect 5166 10996 5172 11008
rect 4948 10968 5172 10996
rect 4948 10956 4954 10968
rect 5166 10956 5172 10968
rect 5224 10956 5230 11008
rect 5644 11005 5672 11036
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 5629 10999 5687 11005
rect 5629 10965 5641 10999
rect 5675 10965 5687 10999
rect 5629 10959 5687 10965
rect 5718 10956 5724 11008
rect 5776 10996 5782 11008
rect 5920 10996 5948 11095
rect 6362 11092 6368 11144
rect 6420 11092 6426 11144
rect 6564 11141 6592 11172
rect 6549 11135 6607 11141
rect 6549 11101 6561 11135
rect 6595 11101 6607 11135
rect 6549 11095 6607 11101
rect 6638 11064 6644 11076
rect 6104 11036 6644 11064
rect 6104 11005 6132 11036
rect 6638 11024 6644 11036
rect 6696 11024 6702 11076
rect 6748 11073 6776 11240
rect 6932 11200 6960 11308
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 7653 11339 7711 11345
rect 7653 11336 7665 11339
rect 7248 11308 7665 11336
rect 7248 11296 7254 11308
rect 7653 11305 7665 11308
rect 7699 11336 7711 11339
rect 9674 11336 9680 11348
rect 7699 11308 9680 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 10060 11308 10364 11336
rect 7101 11271 7159 11277
rect 7101 11237 7113 11271
rect 7147 11268 7159 11271
rect 7742 11268 7748 11280
rect 7147 11240 7748 11268
rect 7147 11237 7159 11240
rect 7101 11231 7159 11237
rect 7742 11228 7748 11240
rect 7800 11228 7806 11280
rect 10060 11277 10088 11308
rect 7929 11271 7987 11277
rect 7929 11237 7941 11271
rect 7975 11268 7987 11271
rect 10045 11271 10103 11277
rect 7975 11240 8064 11268
rect 7975 11237 7987 11240
rect 7929 11231 7987 11237
rect 7282 11200 7288 11212
rect 6840 11172 6960 11200
rect 7116 11172 7288 11200
rect 6840 11141 6868 11172
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11101 6883 11135
rect 6825 11095 6883 11101
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11132 6975 11135
rect 7006 11132 7012 11144
rect 6963 11104 7012 11132
rect 6963 11101 6975 11104
rect 6917 11095 6975 11101
rect 7006 11092 7012 11104
rect 7064 11092 7070 11144
rect 6733 11067 6791 11073
rect 6733 11033 6745 11067
rect 6779 11033 6791 11067
rect 6733 11027 6791 11033
rect 5776 10968 5948 10996
rect 6089 10999 6147 11005
rect 5776 10956 5782 10968
rect 6089 10965 6101 10999
rect 6135 10965 6147 10999
rect 6089 10959 6147 10965
rect 6273 10999 6331 11005
rect 6273 10965 6285 10999
rect 6319 10996 6331 10999
rect 7116 10996 7144 11172
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 7466 11160 7472 11212
rect 7524 11200 7530 11212
rect 7561 11203 7619 11209
rect 7561 11200 7573 11203
rect 7524 11172 7573 11200
rect 7524 11160 7530 11172
rect 7561 11169 7573 11172
rect 7607 11169 7619 11203
rect 7760 11200 7788 11228
rect 8036 11200 8064 11240
rect 10045 11237 10057 11271
rect 10091 11237 10103 11271
rect 10336 11268 10364 11308
rect 10410 11296 10416 11348
rect 10468 11336 10474 11348
rect 10505 11339 10563 11345
rect 10505 11336 10517 11339
rect 10468 11308 10517 11336
rect 10468 11296 10474 11308
rect 10505 11305 10517 11308
rect 10551 11336 10563 11339
rect 10873 11339 10931 11345
rect 10873 11336 10885 11339
rect 10551 11308 10885 11336
rect 10551 11305 10563 11308
rect 10505 11299 10563 11305
rect 10873 11305 10885 11308
rect 10919 11336 10931 11339
rect 11057 11339 11115 11345
rect 10919 11308 11008 11336
rect 10919 11305 10931 11308
rect 10873 11299 10931 11305
rect 10980 11268 11008 11308
rect 11057 11305 11069 11339
rect 11103 11336 11115 11339
rect 11422 11336 11428 11348
rect 11103 11308 11428 11336
rect 11103 11305 11115 11308
rect 11057 11299 11115 11305
rect 11422 11296 11428 11308
rect 11480 11296 11486 11348
rect 11882 11296 11888 11348
rect 11940 11336 11946 11348
rect 12894 11336 12900 11348
rect 11940 11308 12900 11336
rect 11940 11296 11946 11308
rect 12894 11296 12900 11308
rect 12952 11296 12958 11348
rect 13538 11296 13544 11348
rect 13596 11336 13602 11348
rect 14461 11339 14519 11345
rect 14461 11336 14473 11339
rect 13596 11308 14473 11336
rect 13596 11296 13602 11308
rect 14461 11305 14473 11308
rect 14507 11305 14519 11339
rect 14461 11299 14519 11305
rect 14921 11339 14979 11345
rect 14921 11305 14933 11339
rect 14967 11336 14979 11339
rect 15289 11339 15347 11345
rect 15289 11336 15301 11339
rect 14967 11308 15301 11336
rect 14967 11305 14979 11308
rect 14921 11299 14979 11305
rect 15289 11305 15301 11308
rect 15335 11305 15347 11339
rect 15289 11299 15347 11305
rect 15562 11296 15568 11348
rect 15620 11336 15626 11348
rect 16025 11339 16083 11345
rect 16025 11336 16037 11339
rect 15620 11308 16037 11336
rect 15620 11296 15626 11308
rect 16025 11305 16037 11308
rect 16071 11305 16083 11339
rect 16025 11299 16083 11305
rect 16390 11296 16396 11348
rect 16448 11336 16454 11348
rect 19518 11336 19524 11348
rect 16448 11308 19524 11336
rect 16448 11296 16454 11308
rect 19518 11296 19524 11308
rect 19576 11296 19582 11348
rect 19978 11296 19984 11348
rect 20036 11336 20042 11348
rect 20438 11336 20444 11348
rect 20036 11308 20444 11336
rect 20036 11296 20042 11308
rect 20438 11296 20444 11308
rect 20496 11296 20502 11348
rect 20806 11296 20812 11348
rect 20864 11336 20870 11348
rect 20993 11339 21051 11345
rect 20993 11336 21005 11339
rect 20864 11308 21005 11336
rect 20864 11296 20870 11308
rect 20993 11305 21005 11308
rect 21039 11305 21051 11339
rect 20993 11299 21051 11305
rect 21177 11339 21235 11345
rect 21177 11305 21189 11339
rect 21223 11305 21235 11339
rect 22189 11339 22247 11345
rect 22189 11336 22201 11339
rect 21177 11299 21235 11305
rect 22066 11308 22201 11336
rect 14826 11268 14832 11280
rect 10336 11240 10916 11268
rect 10980 11240 14832 11268
rect 10045 11231 10103 11237
rect 8938 11200 8944 11212
rect 7760 11172 7972 11200
rect 8036 11172 8944 11200
rect 7561 11163 7619 11169
rect 7190 11092 7196 11144
rect 7248 11092 7254 11144
rect 7466 11024 7472 11076
rect 7524 11024 7530 11076
rect 7576 11064 7604 11163
rect 7742 11092 7748 11144
rect 7800 11092 7806 11144
rect 7944 11132 7972 11172
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 10321 11203 10379 11209
rect 10321 11200 10333 11203
rect 9508 11172 10333 11200
rect 8297 11135 8355 11141
rect 7944 11104 8248 11132
rect 7576 11036 8064 11064
rect 6319 10968 7144 10996
rect 6319 10965 6331 10968
rect 6273 10959 6331 10965
rect 7282 10956 7288 11008
rect 7340 10996 7346 11008
rect 7377 10999 7435 11005
rect 7377 10996 7389 10999
rect 7340 10968 7389 10996
rect 7340 10956 7346 10968
rect 7377 10965 7389 10968
rect 7423 10996 7435 10999
rect 7926 10996 7932 11008
rect 7423 10968 7932 10996
rect 7423 10965 7435 10968
rect 7377 10959 7435 10965
rect 7926 10956 7932 10968
rect 7984 10956 7990 11008
rect 8036 10996 8064 11036
rect 8110 11024 8116 11076
rect 8168 11024 8174 11076
rect 8220 11064 8248 11104
rect 8297 11101 8309 11135
rect 8343 11132 8355 11135
rect 8570 11132 8576 11144
rect 8343 11104 8576 11132
rect 8343 11101 8355 11104
rect 8297 11095 8355 11101
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 8754 11092 8760 11144
rect 8812 11132 8818 11144
rect 9306 11132 9312 11144
rect 8812 11104 9312 11132
rect 8812 11092 8818 11104
rect 9306 11092 9312 11104
rect 9364 11132 9370 11144
rect 9508 11132 9536 11172
rect 10321 11169 10333 11172
rect 10367 11169 10379 11203
rect 10321 11163 10379 11169
rect 10686 11160 10692 11212
rect 10744 11160 10750 11212
rect 10888 11200 10916 11240
rect 14826 11228 14832 11240
rect 14884 11228 14890 11280
rect 15470 11268 15476 11280
rect 14936 11240 15476 11268
rect 14090 11200 14096 11212
rect 10888 11172 14096 11200
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 14274 11160 14280 11212
rect 14332 11200 14338 11212
rect 14553 11203 14611 11209
rect 14553 11200 14565 11203
rect 14332 11172 14565 11200
rect 14332 11160 14338 11172
rect 14553 11169 14565 11172
rect 14599 11169 14611 11203
rect 14553 11163 14611 11169
rect 9364 11104 9536 11132
rect 9364 11092 9370 11104
rect 10226 11092 10232 11144
rect 10284 11092 10290 11144
rect 10502 11092 10508 11144
rect 10560 11092 10566 11144
rect 10594 11092 10600 11144
rect 10652 11092 10658 11144
rect 10870 11092 10876 11144
rect 10928 11092 10934 11144
rect 14458 11092 14464 11144
rect 14516 11092 14522 11144
rect 14737 11135 14795 11141
rect 14737 11101 14749 11135
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 11793 11067 11851 11073
rect 8220 11036 10272 11064
rect 8386 10996 8392 11008
rect 8036 10968 8392 10996
rect 8386 10956 8392 10968
rect 8444 10996 8450 11008
rect 9122 10996 9128 11008
rect 8444 10968 9128 10996
rect 8444 10956 8450 10968
rect 9122 10956 9128 10968
rect 9180 10956 9186 11008
rect 10244 10996 10272 11036
rect 11793 11033 11805 11067
rect 11839 11064 11851 11067
rect 12158 11064 12164 11076
rect 11839 11036 12164 11064
rect 11839 11033 11851 11036
rect 11793 11027 11851 11033
rect 12158 11024 12164 11036
rect 12216 11024 12222 11076
rect 14745 11064 14773 11095
rect 14826 11092 14832 11144
rect 14884 11132 14890 11144
rect 14936 11132 14964 11240
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 15930 11228 15936 11280
rect 15988 11268 15994 11280
rect 16301 11271 16359 11277
rect 16301 11268 16313 11271
rect 15988 11240 16313 11268
rect 15988 11228 15994 11240
rect 16301 11237 16313 11240
rect 16347 11237 16359 11271
rect 16301 11231 16359 11237
rect 17310 11228 17316 11280
rect 17368 11268 17374 11280
rect 20901 11271 20959 11277
rect 17368 11240 20852 11268
rect 17368 11228 17374 11240
rect 20438 11200 20444 11212
rect 15304 11172 20444 11200
rect 15304 11141 15332 11172
rect 20438 11160 20444 11172
rect 20496 11160 20502 11212
rect 20530 11160 20536 11212
rect 20588 11160 20594 11212
rect 14884 11104 14964 11132
rect 15289 11135 15347 11141
rect 14884 11092 14890 11104
rect 15289 11101 15301 11135
rect 15335 11101 15347 11135
rect 15289 11095 15347 11101
rect 15473 11135 15531 11141
rect 15473 11101 15485 11135
rect 15519 11132 15531 11135
rect 15746 11132 15752 11144
rect 15519 11104 15752 11132
rect 15519 11101 15531 11104
rect 15473 11095 15531 11101
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 15838 11092 15844 11144
rect 15896 11132 15902 11144
rect 16209 11135 16267 11141
rect 16209 11132 16221 11135
rect 15896 11104 16221 11132
rect 15896 11092 15902 11104
rect 16209 11101 16221 11104
rect 16255 11101 16267 11135
rect 16209 11095 16267 11101
rect 16482 11092 16488 11144
rect 16540 11092 16546 11144
rect 16942 11092 16948 11144
rect 17000 11132 17006 11144
rect 17221 11135 17279 11141
rect 17221 11132 17233 11135
rect 17000 11104 17233 11132
rect 17000 11092 17006 11104
rect 17221 11101 17233 11104
rect 17267 11101 17279 11135
rect 17221 11095 17279 11101
rect 17405 11135 17463 11141
rect 17405 11101 17417 11135
rect 17451 11132 17463 11135
rect 17494 11132 17500 11144
rect 17451 11104 17500 11132
rect 17451 11101 17463 11104
rect 17405 11095 17463 11101
rect 17494 11092 17500 11104
rect 17552 11092 17558 11144
rect 18598 11092 18604 11144
rect 18656 11132 18662 11144
rect 18656 11104 20576 11132
rect 18656 11092 18662 11104
rect 14745 11036 15792 11064
rect 15488 11008 15516 11036
rect 11974 10996 11980 11008
rect 10244 10968 11980 10996
rect 11974 10956 11980 10968
rect 12032 10956 12038 11008
rect 12066 10956 12072 11008
rect 12124 10996 12130 11008
rect 15010 10996 15016 11008
rect 12124 10968 15016 10996
rect 12124 10956 12130 10968
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 15470 10956 15476 11008
rect 15528 10956 15534 11008
rect 15654 10956 15660 11008
rect 15712 10956 15718 11008
rect 15764 10996 15792 11036
rect 17310 11024 17316 11076
rect 17368 11064 17374 11076
rect 17589 11067 17647 11073
rect 17589 11064 17601 11067
rect 17368 11036 17601 11064
rect 17368 11024 17374 11036
rect 17589 11033 17601 11036
rect 17635 11064 17647 11067
rect 18690 11064 18696 11076
rect 17635 11036 18696 11064
rect 17635 11033 17647 11036
rect 17589 11027 17647 11033
rect 18690 11024 18696 11036
rect 18748 11024 18754 11076
rect 19886 11024 19892 11076
rect 19944 11064 19950 11076
rect 20441 11067 20499 11073
rect 20441 11064 20453 11067
rect 19944 11036 20453 11064
rect 19944 11024 19950 11036
rect 20441 11033 20453 11036
rect 20487 11033 20499 11067
rect 20548 11064 20576 11104
rect 20714 11092 20720 11144
rect 20772 11092 20778 11144
rect 20824 11132 20852 11240
rect 20901 11237 20913 11271
rect 20947 11237 20959 11271
rect 21192 11268 21220 11299
rect 22066 11280 22094 11308
rect 22189 11305 22201 11308
rect 22235 11336 22247 11339
rect 22922 11336 22928 11348
rect 22235 11308 22928 11336
rect 22235 11305 22247 11308
rect 22189 11299 22247 11305
rect 22922 11296 22928 11308
rect 22980 11296 22986 11348
rect 23658 11296 23664 11348
rect 23716 11336 23722 11348
rect 23845 11339 23903 11345
rect 23845 11336 23857 11339
rect 23716 11308 23857 11336
rect 23716 11296 23722 11308
rect 23845 11305 23857 11308
rect 23891 11336 23903 11339
rect 23934 11336 23940 11348
rect 23891 11308 23940 11336
rect 23891 11305 23903 11308
rect 23845 11299 23903 11305
rect 23934 11296 23940 11308
rect 23992 11296 23998 11348
rect 25498 11296 25504 11348
rect 25556 11336 25562 11348
rect 25685 11339 25743 11345
rect 25685 11336 25697 11339
rect 25556 11308 25697 11336
rect 25556 11296 25562 11308
rect 25685 11305 25697 11308
rect 25731 11305 25743 11339
rect 25685 11299 25743 11305
rect 26234 11296 26240 11348
rect 26292 11296 26298 11348
rect 26786 11296 26792 11348
rect 26844 11296 26850 11348
rect 28074 11296 28080 11348
rect 28132 11296 28138 11348
rect 32122 11296 32128 11348
rect 32180 11336 32186 11348
rect 32217 11339 32275 11345
rect 32217 11336 32229 11339
rect 32180 11308 32229 11336
rect 32180 11296 32186 11308
rect 32217 11305 32229 11308
rect 32263 11305 32275 11339
rect 32217 11299 32275 11305
rect 20901 11231 20959 11237
rect 21100 11240 21220 11268
rect 20916 11200 20944 11231
rect 21100 11200 21128 11240
rect 22002 11228 22008 11280
rect 22060 11240 22094 11280
rect 22373 11271 22431 11277
rect 22060 11228 22066 11240
rect 22373 11237 22385 11271
rect 22419 11268 22431 11271
rect 22462 11268 22468 11280
rect 22419 11240 22468 11268
rect 22419 11237 22431 11240
rect 22373 11231 22431 11237
rect 22462 11228 22468 11240
rect 22520 11228 22526 11280
rect 25958 11268 25964 11280
rect 23584 11240 25964 11268
rect 20916 11172 21128 11200
rect 21174 11160 21180 11212
rect 21232 11200 21238 11212
rect 23584 11200 23612 11240
rect 25958 11228 25964 11240
rect 26016 11228 26022 11280
rect 26053 11271 26111 11277
rect 26053 11237 26065 11271
rect 26099 11237 26111 11271
rect 26053 11231 26111 11237
rect 21232 11172 21404 11200
rect 21232 11160 21238 11172
rect 21376 11141 21404 11172
rect 22020 11172 23612 11200
rect 23661 11203 23719 11209
rect 22020 11141 22048 11172
rect 23661 11169 23673 11203
rect 23707 11169 23719 11203
rect 23661 11163 23719 11169
rect 21269 11135 21327 11141
rect 21269 11132 21281 11135
rect 20824 11104 21281 11132
rect 21269 11101 21281 11104
rect 21315 11101 21327 11135
rect 21269 11095 21327 11101
rect 21361 11135 21419 11141
rect 21361 11101 21373 11135
rect 21407 11101 21419 11135
rect 21361 11095 21419 11101
rect 22005 11135 22063 11141
rect 22005 11101 22017 11135
rect 22051 11101 22063 11135
rect 22005 11095 22063 11101
rect 22186 11092 22192 11144
rect 22244 11092 22250 11144
rect 22646 11092 22652 11144
rect 22704 11092 22710 11144
rect 23106 11092 23112 11144
rect 23164 11132 23170 11144
rect 23569 11135 23627 11141
rect 23569 11132 23581 11135
rect 23164 11104 23581 11132
rect 23164 11092 23170 11104
rect 23569 11101 23581 11104
rect 23615 11101 23627 11135
rect 23569 11095 23627 11101
rect 22278 11064 22284 11076
rect 20548 11036 22284 11064
rect 20441 11027 20499 11033
rect 22278 11024 22284 11036
rect 22336 11024 22342 11076
rect 22388 11036 23244 11064
rect 22388 10996 22416 11036
rect 15764 10968 22416 10996
rect 22465 10999 22523 11005
rect 22465 10965 22477 10999
rect 22511 10996 22523 10999
rect 22554 10996 22560 11008
rect 22511 10968 22560 10996
rect 22511 10965 22523 10968
rect 22465 10959 22523 10965
rect 22554 10956 22560 10968
rect 22612 10956 22618 11008
rect 23216 10996 23244 11036
rect 23290 11024 23296 11076
rect 23348 11064 23354 11076
rect 23676 11064 23704 11163
rect 23845 11135 23903 11141
rect 23845 11101 23857 11135
rect 23891 11132 23903 11135
rect 24210 11132 24216 11144
rect 23891 11104 24216 11132
rect 23891 11101 23903 11104
rect 23845 11095 23903 11101
rect 24210 11092 24216 11104
rect 24268 11092 24274 11144
rect 25682 11092 25688 11144
rect 25740 11092 25746 11144
rect 25777 11135 25835 11141
rect 25777 11101 25789 11135
rect 25823 11101 25835 11135
rect 26068 11132 26096 11231
rect 26326 11228 26332 11280
rect 26384 11268 26390 11280
rect 26697 11271 26755 11277
rect 26697 11268 26709 11271
rect 26384 11240 26709 11268
rect 26384 11228 26390 11240
rect 26697 11237 26709 11240
rect 26743 11237 26755 11271
rect 26697 11231 26755 11237
rect 27157 11271 27215 11277
rect 27157 11237 27169 11271
rect 27203 11268 27215 11271
rect 28626 11268 28632 11280
rect 27203 11240 28632 11268
rect 27203 11237 27215 11240
rect 27157 11231 27215 11237
rect 28626 11228 28632 11240
rect 28684 11228 28690 11280
rect 30745 11271 30803 11277
rect 30745 11237 30757 11271
rect 30791 11237 30803 11271
rect 30745 11231 30803 11237
rect 26421 11203 26479 11209
rect 26421 11169 26433 11203
rect 26467 11200 26479 11203
rect 27338 11200 27344 11212
rect 26467 11172 27344 11200
rect 26467 11169 26479 11172
rect 26421 11163 26479 11169
rect 27338 11160 27344 11172
rect 27396 11160 27402 11212
rect 28258 11160 28264 11212
rect 28316 11200 28322 11212
rect 28442 11200 28448 11212
rect 28316 11172 28448 11200
rect 28316 11160 28322 11172
rect 28442 11160 28448 11172
rect 28500 11160 28506 11212
rect 30760 11200 30788 11231
rect 30760 11172 30972 11200
rect 26237 11135 26295 11141
rect 26237 11132 26249 11135
rect 26068 11104 26249 11132
rect 25777 11095 25835 11101
rect 26237 11101 26249 11104
rect 26283 11101 26295 11135
rect 26237 11095 26295 11101
rect 26513 11135 26571 11141
rect 26513 11101 26525 11135
rect 26559 11132 26571 11135
rect 26602 11132 26608 11144
rect 26559 11104 26608 11132
rect 26559 11101 26571 11104
rect 26513 11095 26571 11101
rect 23348 11036 23704 11064
rect 23952 11036 25360 11064
rect 23348 11024 23354 11036
rect 23952 10996 23980 11036
rect 23216 10968 23980 10996
rect 24026 10956 24032 11008
rect 24084 10956 24090 11008
rect 25332 10996 25360 11036
rect 25406 11024 25412 11076
rect 25464 11064 25470 11076
rect 25792 11064 25820 11095
rect 26602 11092 26608 11104
rect 26660 11092 26666 11144
rect 26786 11092 26792 11144
rect 26844 11092 26850 11144
rect 26881 11135 26939 11141
rect 26881 11101 26893 11135
rect 26927 11132 26939 11135
rect 28534 11132 28540 11144
rect 26927 11104 28540 11132
rect 26927 11101 26939 11104
rect 26881 11095 26939 11101
rect 28534 11092 28540 11104
rect 28592 11092 28598 11144
rect 30190 11092 30196 11144
rect 30248 11092 30254 11144
rect 30374 11092 30380 11144
rect 30432 11092 30438 11144
rect 30558 11092 30564 11144
rect 30616 11092 30622 11144
rect 30834 11092 30840 11144
rect 30892 11092 30898 11144
rect 30944 11132 30972 11172
rect 31093 11135 31151 11141
rect 31093 11132 31105 11135
rect 30944 11104 31105 11132
rect 31093 11101 31105 11104
rect 31139 11101 31151 11135
rect 31093 11095 31151 11101
rect 25464 11036 25820 11064
rect 26620 11064 26648 11092
rect 26970 11064 26976 11076
rect 26620 11036 26976 11064
rect 25464 11024 25470 11036
rect 26970 11024 26976 11036
rect 27028 11024 27034 11076
rect 27709 11067 27767 11073
rect 27709 11033 27721 11067
rect 27755 11033 27767 11067
rect 27709 11027 27767 11033
rect 26602 10996 26608 11008
rect 25332 10968 26608 10996
rect 26602 10956 26608 10968
rect 26660 10956 26666 11008
rect 27430 10956 27436 11008
rect 27488 10996 27494 11008
rect 27724 10996 27752 11027
rect 27798 11024 27804 11076
rect 27856 11064 27862 11076
rect 27893 11067 27951 11073
rect 27893 11064 27905 11067
rect 27856 11036 27905 11064
rect 27856 11024 27862 11036
rect 27893 11033 27905 11036
rect 27939 11033 27951 11067
rect 27893 11027 27951 11033
rect 30469 11067 30527 11073
rect 30469 11033 30481 11067
rect 30515 11064 30527 11067
rect 31202 11064 31208 11076
rect 30515 11036 31208 11064
rect 30515 11033 30527 11036
rect 30469 11027 30527 11033
rect 31202 11024 31208 11036
rect 31260 11024 31266 11076
rect 28258 10996 28264 11008
rect 27488 10968 28264 10996
rect 27488 10956 27494 10968
rect 28258 10956 28264 10968
rect 28316 10956 28322 11008
rect 1104 10906 32844 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 32844 10906
rect 1104 10832 32844 10854
rect 3602 10752 3608 10804
rect 3660 10792 3666 10804
rect 4430 10792 4436 10804
rect 3660 10764 4436 10792
rect 3660 10752 3666 10764
rect 4430 10752 4436 10764
rect 4488 10752 4494 10804
rect 4614 10752 4620 10804
rect 4672 10792 4678 10804
rect 4709 10795 4767 10801
rect 4709 10792 4721 10795
rect 4672 10764 4721 10792
rect 4672 10752 4678 10764
rect 4709 10761 4721 10764
rect 4755 10761 4767 10795
rect 4709 10755 4767 10761
rect 3970 10684 3976 10736
rect 4028 10724 4034 10736
rect 4249 10727 4307 10733
rect 4249 10724 4261 10727
rect 4028 10696 4261 10724
rect 4028 10684 4034 10696
rect 4249 10693 4261 10696
rect 4295 10693 4307 10727
rect 4724 10724 4752 10755
rect 4982 10752 4988 10804
rect 5040 10792 5046 10804
rect 5718 10792 5724 10804
rect 5040 10764 5724 10792
rect 5040 10752 5046 10764
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 5902 10792 5908 10804
rect 5828 10764 5908 10792
rect 5626 10724 5632 10736
rect 4724 10696 5632 10724
rect 4249 10687 4307 10693
rect 5626 10684 5632 10696
rect 5684 10684 5690 10736
rect 5828 10680 5856 10764
rect 5902 10752 5908 10764
rect 5960 10752 5966 10804
rect 6914 10752 6920 10804
rect 6972 10752 6978 10804
rect 7466 10752 7472 10804
rect 7524 10752 7530 10804
rect 9030 10752 9036 10804
rect 9088 10792 9094 10804
rect 11885 10795 11943 10801
rect 9088 10764 11744 10792
rect 9088 10752 9094 10764
rect 6549 10727 6607 10733
rect 6549 10693 6561 10727
rect 6595 10693 6607 10727
rect 6549 10687 6607 10693
rect 7009 10727 7067 10733
rect 7009 10693 7021 10727
rect 7055 10724 7067 10727
rect 7055 10696 7236 10724
rect 7055 10693 7067 10696
rect 7009 10687 7067 10693
rect 5828 10669 5922 10680
rect 3142 10616 3148 10668
rect 3200 10656 3206 10668
rect 3694 10656 3700 10668
rect 3200 10628 3700 10656
rect 3200 10616 3206 10628
rect 3694 10616 3700 10628
rect 3752 10656 3758 10668
rect 4065 10659 4123 10665
rect 4065 10656 4077 10659
rect 3752 10628 4077 10656
rect 3752 10616 3758 10628
rect 4065 10625 4077 10628
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 4338 10616 4344 10668
rect 4396 10616 4402 10668
rect 4433 10659 4491 10665
rect 4433 10625 4445 10659
rect 4479 10656 4491 10659
rect 4614 10656 4620 10668
rect 4479 10628 4620 10656
rect 4479 10625 4491 10628
rect 4433 10619 4491 10625
rect 4614 10616 4620 10628
rect 4672 10656 4678 10668
rect 4672 10628 4752 10656
rect 4672 10616 4678 10628
rect 4356 10588 4384 10616
rect 3160 10560 4384 10588
rect 4448 10560 4660 10588
rect 3160 10532 3188 10560
rect 4448 10532 4476 10560
rect 3142 10480 3148 10532
rect 3200 10480 3206 10532
rect 4430 10480 4436 10532
rect 4488 10480 4494 10532
rect 4632 10529 4660 10560
rect 4617 10523 4675 10529
rect 4617 10489 4629 10523
rect 4663 10489 4675 10523
rect 4724 10520 4752 10628
rect 4890 10616 4896 10668
rect 4948 10616 4954 10668
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10656 5043 10659
rect 5350 10656 5356 10668
rect 5031 10628 5356 10656
rect 5031 10625 5043 10628
rect 4985 10619 5043 10625
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 5445 10659 5503 10665
rect 5445 10625 5457 10659
rect 5491 10625 5503 10659
rect 5828 10663 5937 10669
rect 5997 10668 6055 10669
rect 5828 10652 5891 10663
rect 5445 10619 5503 10625
rect 5879 10629 5891 10652
rect 5925 10629 5937 10663
rect 5879 10623 5937 10629
rect 5074 10548 5080 10600
rect 5132 10588 5138 10600
rect 5460 10588 5488 10619
rect 5994 10616 6000 10668
rect 6052 10616 6058 10668
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 6196 10628 6377 10656
rect 5132 10560 5488 10588
rect 5132 10548 5138 10560
rect 5261 10523 5319 10529
rect 5261 10520 5273 10523
rect 4724 10492 5273 10520
rect 4617 10483 4675 10489
rect 5261 10489 5273 10492
rect 5307 10489 5319 10523
rect 6196 10520 6224 10628
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 6564 10600 6592 10687
rect 6638 10616 6644 10668
rect 6696 10616 6702 10668
rect 6730 10616 6736 10668
rect 6788 10665 6794 10668
rect 6788 10659 6815 10665
rect 6803 10625 6815 10659
rect 6788 10619 6815 10625
rect 6788 10616 6794 10619
rect 6546 10548 6552 10600
rect 6604 10548 6610 10600
rect 7098 10548 7104 10600
rect 7156 10548 7162 10600
rect 5261 10483 5319 10489
rect 5736 10492 6224 10520
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 5166 10452 5172 10464
rect 4580 10424 5172 10452
rect 4580 10412 4586 10424
rect 5166 10412 5172 10424
rect 5224 10412 5230 10464
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 5736 10461 5764 10492
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 7208 10520 7236 10696
rect 7558 10684 7564 10736
rect 7616 10684 7622 10736
rect 9217 10727 9275 10733
rect 9217 10693 9229 10727
rect 9263 10724 9275 10727
rect 9306 10724 9312 10736
rect 9263 10696 9312 10724
rect 9263 10693 9275 10696
rect 9217 10687 9275 10693
rect 9306 10684 9312 10696
rect 9364 10684 9370 10736
rect 9401 10727 9459 10733
rect 9401 10693 9413 10727
rect 9447 10724 9459 10727
rect 11606 10724 11612 10736
rect 9447 10696 11612 10724
rect 9447 10693 9459 10696
rect 9401 10687 9459 10693
rect 11606 10684 11612 10696
rect 11664 10684 11670 10736
rect 11716 10724 11744 10764
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 12710 10792 12716 10804
rect 11931 10764 12716 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 13081 10795 13139 10801
rect 13081 10761 13093 10795
rect 13127 10792 13139 10795
rect 18049 10795 18107 10801
rect 13127 10764 17724 10792
rect 13127 10761 13139 10764
rect 13081 10755 13139 10761
rect 12250 10724 12256 10736
rect 11716 10696 12256 10724
rect 12250 10684 12256 10696
rect 12308 10684 12314 10736
rect 12621 10727 12679 10733
rect 12621 10693 12633 10727
rect 12667 10724 12679 10727
rect 13998 10724 14004 10736
rect 12667 10696 14004 10724
rect 12667 10693 12679 10696
rect 12621 10687 12679 10693
rect 13998 10684 14004 10696
rect 14056 10684 14062 10736
rect 15841 10727 15899 10733
rect 14200 10696 15148 10724
rect 7282 10616 7288 10668
rect 7340 10616 7346 10668
rect 7742 10616 7748 10668
rect 7800 10616 7806 10668
rect 9677 10659 9735 10665
rect 9677 10625 9689 10659
rect 9723 10656 9735 10659
rect 9950 10656 9956 10668
rect 9723 10628 9956 10656
rect 9723 10625 9735 10628
rect 9677 10619 9735 10625
rect 9950 10616 9956 10628
rect 10008 10616 10014 10668
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10962 10656 10968 10668
rect 10192 10628 10968 10656
rect 10192 10616 10198 10628
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 11422 10616 11428 10668
rect 11480 10656 11486 10668
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 11480 10628 11529 10656
rect 11480 10616 11486 10628
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 11698 10616 11704 10668
rect 11756 10616 11762 10668
rect 11974 10616 11980 10668
rect 12032 10616 12038 10668
rect 12897 10659 12955 10665
rect 12406 10628 12848 10656
rect 7650 10548 7656 10600
rect 7708 10588 7714 10600
rect 8386 10588 8392 10600
rect 7708 10560 8392 10588
rect 7708 10548 7714 10560
rect 8386 10548 8392 10560
rect 8444 10548 8450 10600
rect 9033 10591 9091 10597
rect 9033 10557 9045 10591
rect 9079 10588 9091 10591
rect 9582 10588 9588 10600
rect 9079 10560 9588 10588
rect 9079 10557 9091 10560
rect 9033 10551 9091 10557
rect 9582 10548 9588 10560
rect 9640 10588 9646 10600
rect 12406 10588 12434 10628
rect 9640 10560 12434 10588
rect 9640 10548 9646 10560
rect 12710 10548 12716 10600
rect 12768 10548 12774 10600
rect 12820 10588 12848 10628
rect 12897 10625 12909 10659
rect 12943 10656 12955 10659
rect 13078 10656 13084 10668
rect 12943 10628 13084 10656
rect 12943 10625 12955 10628
rect 12897 10619 12955 10625
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 14200 10588 14228 10696
rect 14277 10659 14335 10665
rect 14277 10625 14289 10659
rect 14323 10625 14335 10659
rect 14277 10619 14335 10625
rect 12820 10560 14228 10588
rect 12802 10520 12808 10532
rect 6972 10492 12808 10520
rect 6972 10480 6978 10492
rect 12802 10480 12808 10492
rect 12860 10480 12866 10532
rect 14292 10520 14320 10619
rect 14550 10616 14556 10668
rect 14608 10616 14614 10668
rect 14366 10548 14372 10600
rect 14424 10548 14430 10600
rect 12912 10492 14320 10520
rect 14737 10523 14795 10529
rect 5721 10455 5779 10461
rect 5721 10452 5733 10455
rect 5592 10424 5733 10452
rect 5592 10412 5598 10424
rect 5721 10421 5733 10424
rect 5767 10421 5779 10455
rect 5721 10415 5779 10421
rect 5810 10412 5816 10464
rect 5868 10452 5874 10464
rect 6086 10452 6092 10464
rect 5868 10424 6092 10452
rect 5868 10412 5874 10424
rect 6086 10412 6092 10424
rect 6144 10412 6150 10464
rect 6181 10455 6239 10461
rect 6181 10421 6193 10455
rect 6227 10452 6239 10455
rect 6270 10452 6276 10464
rect 6227 10424 6276 10452
rect 6227 10421 6239 10424
rect 6181 10415 6239 10421
rect 6270 10412 6276 10424
rect 6328 10412 6334 10464
rect 7285 10455 7343 10461
rect 7285 10421 7297 10455
rect 7331 10452 7343 10455
rect 7374 10452 7380 10464
rect 7331 10424 7380 10452
rect 7331 10421 7343 10424
rect 7285 10415 7343 10421
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 7929 10455 7987 10461
rect 7929 10421 7941 10455
rect 7975 10452 7987 10455
rect 9398 10452 9404 10464
rect 7975 10424 9404 10452
rect 7975 10421 7987 10424
rect 7929 10415 7987 10421
rect 9398 10412 9404 10424
rect 9456 10412 9462 10464
rect 9493 10455 9551 10461
rect 9493 10421 9505 10455
rect 9539 10452 9551 10455
rect 9674 10452 9680 10464
rect 9539 10424 9680 10452
rect 9539 10421 9551 10424
rect 9493 10415 9551 10421
rect 9674 10412 9680 10424
rect 9732 10452 9738 10464
rect 11422 10452 11428 10464
rect 9732 10424 11428 10452
rect 9732 10412 9738 10424
rect 11422 10412 11428 10424
rect 11480 10412 11486 10464
rect 11698 10412 11704 10464
rect 11756 10452 11762 10464
rect 12158 10452 12164 10464
rect 11756 10424 12164 10452
rect 11756 10412 11762 10424
rect 12158 10412 12164 10424
rect 12216 10412 12222 10464
rect 12250 10412 12256 10464
rect 12308 10452 12314 10464
rect 12912 10461 12940 10492
rect 14737 10489 14749 10523
rect 14783 10489 14795 10523
rect 15120 10520 15148 10696
rect 15841 10693 15853 10727
rect 15887 10724 15899 10727
rect 15930 10724 15936 10736
rect 15887 10696 15936 10724
rect 15887 10693 15899 10696
rect 15841 10687 15899 10693
rect 15930 10684 15936 10696
rect 15988 10684 15994 10736
rect 15194 10616 15200 10668
rect 15252 10656 15258 10668
rect 16117 10659 16175 10665
rect 16117 10656 16129 10659
rect 15252 10628 16129 10656
rect 15252 10616 15258 10628
rect 16117 10625 16129 10628
rect 16163 10656 16175 10659
rect 16206 10656 16212 10668
rect 16163 10628 16212 10656
rect 16163 10625 16175 10628
rect 16117 10619 16175 10625
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 16758 10616 16764 10668
rect 16816 10656 16822 10668
rect 16945 10659 17003 10665
rect 16945 10656 16957 10659
rect 16816 10628 16957 10656
rect 16816 10616 16822 10628
rect 16945 10625 16957 10628
rect 16991 10625 17003 10659
rect 16945 10619 17003 10625
rect 17129 10659 17187 10665
rect 17129 10625 17141 10659
rect 17175 10656 17187 10659
rect 17402 10656 17408 10668
rect 17175 10628 17408 10656
rect 17175 10625 17187 10628
rect 17129 10619 17187 10625
rect 17402 10616 17408 10628
rect 17460 10616 17466 10668
rect 17586 10616 17592 10668
rect 17644 10616 17650 10668
rect 17696 10665 17724 10764
rect 18049 10761 18061 10795
rect 18095 10792 18107 10795
rect 18095 10764 19012 10792
rect 18095 10761 18107 10764
rect 18049 10755 18107 10761
rect 18414 10684 18420 10736
rect 18472 10724 18478 10736
rect 18874 10724 18880 10736
rect 18472 10696 18880 10724
rect 18472 10684 18478 10696
rect 18874 10684 18880 10696
rect 18932 10684 18938 10736
rect 18984 10733 19012 10764
rect 19426 10752 19432 10804
rect 19484 10752 19490 10804
rect 20346 10792 20352 10804
rect 19996 10764 20352 10792
rect 19996 10733 20024 10764
rect 20346 10752 20352 10764
rect 20404 10752 20410 10804
rect 20530 10752 20536 10804
rect 20588 10752 20594 10804
rect 20625 10795 20683 10801
rect 20625 10761 20637 10795
rect 20671 10792 20683 10795
rect 20714 10792 20720 10804
rect 20671 10764 20720 10792
rect 20671 10761 20683 10764
rect 20625 10755 20683 10761
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 22094 10792 22100 10804
rect 22066 10752 22100 10792
rect 22152 10752 22158 10804
rect 22186 10752 22192 10804
rect 22244 10752 22250 10804
rect 22833 10795 22891 10801
rect 22833 10761 22845 10795
rect 22879 10792 22891 10795
rect 24397 10795 24455 10801
rect 22879 10764 24348 10792
rect 22879 10761 22891 10764
rect 22833 10755 22891 10761
rect 18969 10727 19027 10733
rect 18969 10693 18981 10727
rect 19015 10693 19027 10727
rect 18969 10687 19027 10693
rect 19974 10727 20032 10733
rect 19974 10693 19986 10727
rect 20020 10693 20032 10727
rect 20548 10724 20576 10752
rect 19974 10687 20032 10693
rect 20456 10696 20576 10724
rect 17681 10659 17739 10665
rect 17681 10625 17693 10659
rect 17727 10625 17739 10659
rect 17681 10619 17739 10625
rect 18782 10616 18788 10668
rect 18840 10656 18846 10668
rect 19245 10659 19303 10665
rect 18840 10628 19196 10656
rect 18840 10616 18846 10628
rect 16025 10591 16083 10597
rect 16025 10557 16037 10591
rect 16071 10557 16083 10591
rect 17773 10591 17831 10597
rect 17773 10588 17785 10591
rect 16025 10551 16083 10557
rect 16224 10560 17785 10588
rect 16040 10520 16068 10551
rect 16114 10520 16120 10532
rect 15120 10492 15976 10520
rect 16040 10492 16120 10520
rect 14737 10483 14795 10489
rect 12897 10455 12955 10461
rect 12897 10452 12909 10455
rect 12308 10424 12909 10452
rect 12308 10412 12314 10424
rect 12897 10421 12909 10424
rect 12943 10421 12955 10455
rect 12897 10415 12955 10421
rect 13078 10412 13084 10464
rect 13136 10452 13142 10464
rect 14277 10455 14335 10461
rect 14277 10452 14289 10455
rect 13136 10424 14289 10452
rect 13136 10412 13142 10424
rect 14277 10421 14289 10424
rect 14323 10421 14335 10455
rect 14752 10452 14780 10483
rect 15470 10452 15476 10464
rect 14752 10424 15476 10452
rect 14277 10415 14335 10421
rect 15470 10412 15476 10424
rect 15528 10412 15534 10464
rect 15562 10412 15568 10464
rect 15620 10452 15626 10464
rect 15841 10455 15899 10461
rect 15841 10452 15853 10455
rect 15620 10424 15853 10452
rect 15620 10412 15626 10424
rect 15841 10421 15853 10424
rect 15887 10421 15899 10455
rect 15948 10452 15976 10492
rect 16114 10480 16120 10492
rect 16172 10480 16178 10532
rect 16224 10452 16252 10560
rect 17773 10557 17785 10560
rect 17819 10588 17831 10591
rect 18138 10588 18144 10600
rect 17819 10560 18144 10588
rect 17819 10557 17831 10560
rect 17773 10551 17831 10557
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 19058 10548 19064 10600
rect 19116 10548 19122 10600
rect 19168 10588 19196 10628
rect 19245 10625 19257 10659
rect 19291 10656 19303 10659
rect 19334 10656 19340 10668
rect 19291 10628 19340 10656
rect 19291 10625 19303 10628
rect 19245 10619 19303 10625
rect 19334 10616 19340 10628
rect 19392 10616 19398 10668
rect 19705 10659 19763 10665
rect 19705 10625 19717 10659
rect 19751 10625 19763 10659
rect 20073 10659 20131 10665
rect 20073 10656 20085 10659
rect 19705 10619 19763 10625
rect 19812 10628 20085 10656
rect 19720 10588 19748 10619
rect 19168 10560 19748 10588
rect 17313 10523 17371 10529
rect 17313 10489 17325 10523
rect 17359 10520 17371 10523
rect 18046 10520 18052 10532
rect 17359 10492 18052 10520
rect 17359 10489 17371 10492
rect 17313 10483 17371 10489
rect 18046 10480 18052 10492
rect 18104 10480 18110 10532
rect 18414 10480 18420 10532
rect 18472 10520 18478 10532
rect 19812 10520 19840 10628
rect 20073 10625 20085 10628
rect 20119 10625 20131 10659
rect 20456 10656 20484 10696
rect 21082 10684 21088 10736
rect 21140 10684 21146 10736
rect 22066 10724 22094 10752
rect 22554 10724 22560 10736
rect 21468 10696 22560 10724
rect 20073 10619 20131 10625
rect 20297 10628 20484 10656
rect 19889 10591 19947 10597
rect 19889 10557 19901 10591
rect 19935 10588 19947 10591
rect 20297 10588 20325 10628
rect 20530 10616 20536 10668
rect 20588 10616 20594 10668
rect 20809 10659 20867 10665
rect 20809 10625 20821 10659
rect 20855 10656 20867 10659
rect 21269 10659 21327 10665
rect 20855 10628 21036 10656
rect 20855 10625 20867 10628
rect 20809 10619 20867 10625
rect 19935 10560 20325 10588
rect 19935 10557 19947 10560
rect 19889 10551 19947 10557
rect 20898 10548 20904 10600
rect 20956 10548 20962 10600
rect 21008 10588 21036 10628
rect 21269 10625 21281 10659
rect 21315 10656 21327 10659
rect 21358 10656 21364 10668
rect 21315 10628 21364 10656
rect 21315 10625 21327 10628
rect 21269 10619 21327 10625
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 21468 10665 21496 10696
rect 22554 10684 22560 10696
rect 22612 10684 22618 10736
rect 23566 10684 23572 10736
rect 23624 10684 23630 10736
rect 23934 10684 23940 10736
rect 23992 10684 23998 10736
rect 24320 10724 24348 10764
rect 24397 10761 24409 10795
rect 24443 10792 24455 10795
rect 25133 10795 25191 10801
rect 24443 10764 24716 10792
rect 24443 10761 24455 10764
rect 24397 10755 24455 10761
rect 24688 10733 24716 10764
rect 25133 10761 25145 10795
rect 25179 10792 25191 10795
rect 25961 10795 26019 10801
rect 25179 10764 25544 10792
rect 25179 10761 25191 10764
rect 25133 10755 25191 10761
rect 25516 10733 25544 10764
rect 25961 10761 25973 10795
rect 26007 10792 26019 10795
rect 26786 10792 26792 10804
rect 26007 10764 26792 10792
rect 26007 10761 26019 10764
rect 25961 10755 26019 10761
rect 26786 10752 26792 10764
rect 26844 10752 26850 10804
rect 27062 10752 27068 10804
rect 27120 10792 27126 10804
rect 27525 10795 27583 10801
rect 27525 10792 27537 10795
rect 27120 10764 27537 10792
rect 27120 10752 27126 10764
rect 27525 10761 27537 10764
rect 27571 10761 27583 10795
rect 27525 10755 27583 10761
rect 27982 10752 27988 10804
rect 28040 10752 28046 10804
rect 28350 10752 28356 10804
rect 28408 10792 28414 10804
rect 28445 10795 28503 10801
rect 28445 10792 28457 10795
rect 28408 10764 28457 10792
rect 28408 10752 28414 10764
rect 28445 10761 28457 10764
rect 28491 10761 28503 10795
rect 28445 10755 28503 10761
rect 30558 10752 30564 10804
rect 30616 10792 30622 10804
rect 31297 10795 31355 10801
rect 31297 10792 31309 10795
rect 30616 10764 31309 10792
rect 30616 10752 30622 10764
rect 31297 10761 31309 10764
rect 31343 10761 31355 10795
rect 31297 10755 31355 10761
rect 24673 10727 24731 10733
rect 24320 10696 24532 10724
rect 21453 10659 21511 10665
rect 21453 10625 21465 10659
rect 21499 10625 21511 10659
rect 21453 10619 21511 10625
rect 21818 10616 21824 10668
rect 21876 10616 21882 10668
rect 22002 10616 22008 10668
rect 22060 10616 22066 10668
rect 22094 10616 22100 10668
rect 22152 10656 22158 10668
rect 22373 10659 22431 10665
rect 22373 10656 22385 10659
rect 22152 10628 22385 10656
rect 22152 10616 22158 10628
rect 22373 10625 22385 10628
rect 22419 10625 22431 10659
rect 22373 10619 22431 10625
rect 22646 10616 22652 10668
rect 22704 10616 22710 10668
rect 22922 10616 22928 10668
rect 22980 10616 22986 10668
rect 23477 10659 23535 10665
rect 23477 10625 23489 10659
rect 23523 10656 23535 10659
rect 23584 10656 23612 10684
rect 23523 10628 23980 10656
rect 23523 10625 23535 10628
rect 23477 10619 23535 10625
rect 22186 10588 22192 10600
rect 21008 10560 22192 10588
rect 22186 10548 22192 10560
rect 22244 10548 22250 10600
rect 22278 10548 22284 10600
rect 22336 10588 22342 10600
rect 22465 10591 22523 10597
rect 22465 10588 22477 10591
rect 22336 10560 22477 10588
rect 22336 10548 22342 10560
rect 22465 10557 22477 10560
rect 22511 10557 22523 10591
rect 23017 10591 23075 10597
rect 23017 10588 23029 10591
rect 22465 10551 22523 10557
rect 22572 10560 23029 10588
rect 22572 10532 22600 10560
rect 23017 10557 23029 10560
rect 23063 10557 23075 10591
rect 23017 10551 23075 10557
rect 23566 10548 23572 10600
rect 23624 10548 23630 10600
rect 20714 10520 20720 10532
rect 18472 10492 19840 10520
rect 20272 10492 20720 10520
rect 18472 10480 18478 10492
rect 15948 10424 16252 10452
rect 15841 10415 15899 10421
rect 16298 10412 16304 10464
rect 16356 10412 16362 10464
rect 16758 10412 16764 10464
rect 16816 10412 16822 10464
rect 17405 10455 17463 10461
rect 17405 10421 17417 10455
rect 17451 10452 17463 10455
rect 17494 10452 17500 10464
rect 17451 10424 17500 10452
rect 17451 10421 17463 10424
rect 17405 10415 17463 10421
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 17770 10412 17776 10464
rect 17828 10412 17834 10464
rect 19242 10412 19248 10464
rect 19300 10412 19306 10464
rect 19334 10412 19340 10464
rect 19392 10452 19398 10464
rect 19521 10455 19579 10461
rect 19521 10452 19533 10455
rect 19392 10424 19533 10452
rect 19392 10412 19398 10424
rect 19521 10421 19533 10424
rect 19567 10421 19579 10455
rect 19521 10415 19579 10421
rect 19886 10412 19892 10464
rect 19944 10412 19950 10464
rect 20272 10461 20300 10492
rect 20714 10480 20720 10492
rect 20772 10480 20778 10532
rect 21542 10520 21548 10532
rect 21100 10492 21548 10520
rect 20257 10455 20315 10461
rect 20257 10421 20269 10455
rect 20303 10421 20315 10455
rect 20257 10415 20315 10421
rect 20346 10412 20352 10464
rect 20404 10412 20410 10464
rect 20622 10412 20628 10464
rect 20680 10452 20686 10464
rect 20898 10452 20904 10464
rect 20680 10424 20904 10452
rect 20680 10412 20686 10424
rect 20898 10412 20904 10424
rect 20956 10412 20962 10464
rect 21100 10461 21128 10492
rect 21542 10480 21548 10492
rect 21600 10480 21606 10532
rect 21637 10523 21695 10529
rect 21637 10489 21649 10523
rect 21683 10520 21695 10523
rect 22554 10520 22560 10532
rect 21683 10492 22560 10520
rect 21683 10489 21695 10492
rect 21637 10483 21695 10489
rect 22554 10480 22560 10492
rect 22612 10480 22618 10532
rect 23293 10523 23351 10529
rect 23293 10520 23305 10523
rect 22664 10492 23305 10520
rect 21085 10455 21143 10461
rect 21085 10421 21097 10455
rect 21131 10421 21143 10455
rect 21085 10415 21143 10421
rect 21174 10412 21180 10464
rect 21232 10452 21238 10464
rect 21269 10455 21327 10461
rect 21269 10452 21281 10455
rect 21232 10424 21281 10452
rect 21232 10412 21238 10424
rect 21269 10421 21281 10424
rect 21315 10452 21327 10455
rect 21818 10452 21824 10464
rect 21315 10424 21824 10452
rect 21315 10421 21327 10424
rect 21269 10415 21327 10421
rect 21818 10412 21824 10424
rect 21876 10412 21882 10464
rect 22664 10461 22692 10492
rect 23293 10489 23305 10492
rect 23339 10489 23351 10523
rect 23293 10483 23351 10489
rect 23382 10480 23388 10532
rect 23440 10520 23446 10532
rect 23845 10523 23903 10529
rect 23845 10520 23857 10523
rect 23440 10492 23857 10520
rect 23440 10480 23446 10492
rect 23845 10489 23857 10492
rect 23891 10489 23903 10523
rect 23845 10483 23903 10489
rect 22649 10455 22707 10461
rect 22649 10421 22661 10455
rect 22695 10421 22707 10455
rect 22649 10415 22707 10421
rect 22922 10412 22928 10464
rect 22980 10412 22986 10464
rect 23014 10412 23020 10464
rect 23072 10452 23078 10464
rect 23400 10452 23428 10480
rect 23072 10424 23428 10452
rect 23072 10412 23078 10424
rect 23474 10412 23480 10464
rect 23532 10412 23538 10464
rect 23952 10461 23980 10628
rect 24118 10616 24124 10668
rect 24176 10616 24182 10668
rect 24213 10659 24271 10665
rect 24213 10625 24225 10659
rect 24259 10656 24271 10659
rect 24302 10656 24308 10668
rect 24259 10628 24308 10656
rect 24259 10625 24271 10628
rect 24213 10619 24271 10625
rect 24302 10616 24308 10628
rect 24360 10616 24366 10668
rect 24504 10588 24532 10696
rect 24673 10693 24685 10727
rect 24719 10693 24731 10727
rect 25501 10727 25559 10733
rect 24673 10687 24731 10693
rect 24780 10696 25084 10724
rect 24578 10616 24584 10668
rect 24636 10656 24642 10668
rect 24780 10656 24808 10696
rect 24636 10628 24808 10656
rect 24636 10616 24642 10628
rect 24946 10616 24952 10668
rect 25004 10616 25010 10668
rect 25056 10656 25084 10696
rect 25501 10693 25513 10727
rect 25547 10693 25559 10727
rect 25501 10687 25559 10693
rect 25608 10696 26096 10724
rect 25608 10656 25636 10696
rect 26068 10665 26096 10696
rect 26142 10684 26148 10736
rect 26200 10724 26206 10736
rect 30190 10724 30196 10736
rect 26200 10696 30196 10724
rect 26200 10684 26206 10696
rect 30190 10684 30196 10696
rect 30248 10684 30254 10736
rect 31386 10724 31392 10736
rect 30944 10696 31392 10724
rect 25056 10628 25636 10656
rect 25777 10659 25835 10665
rect 25777 10625 25789 10659
rect 25823 10625 25835 10659
rect 25777 10619 25835 10625
rect 26053 10659 26111 10665
rect 26053 10625 26065 10659
rect 26099 10625 26111 10659
rect 26053 10619 26111 10625
rect 24504 10560 24716 10588
rect 24688 10520 24716 10560
rect 24762 10548 24768 10600
rect 24820 10548 24826 10600
rect 24854 10548 24860 10600
rect 24912 10588 24918 10600
rect 25593 10591 25651 10597
rect 25593 10588 25605 10591
rect 24912 10560 25605 10588
rect 24912 10548 24918 10560
rect 25593 10557 25605 10560
rect 25639 10588 25651 10591
rect 25682 10588 25688 10600
rect 25639 10560 25688 10588
rect 25639 10557 25651 10560
rect 25593 10551 25651 10557
rect 25682 10548 25688 10560
rect 25740 10548 25746 10600
rect 25792 10520 25820 10619
rect 26786 10616 26792 10668
rect 26844 10656 26850 10668
rect 27065 10659 27123 10665
rect 27065 10656 27077 10659
rect 26844 10628 27077 10656
rect 26844 10616 26850 10628
rect 27065 10625 27077 10628
rect 27111 10656 27123 10659
rect 27111 10628 27292 10656
rect 27111 10625 27123 10628
rect 27065 10619 27123 10625
rect 25866 10548 25872 10600
rect 25924 10588 25930 10600
rect 26145 10591 26203 10597
rect 26145 10588 26157 10591
rect 25924 10560 26157 10588
rect 25924 10548 25930 10560
rect 26145 10557 26157 10560
rect 26191 10557 26203 10591
rect 26145 10551 26203 10557
rect 26970 10548 26976 10600
rect 27028 10588 27034 10600
rect 27157 10591 27215 10597
rect 27157 10588 27169 10591
rect 27028 10560 27169 10588
rect 27028 10548 27034 10560
rect 27157 10557 27169 10560
rect 27203 10557 27215 10591
rect 27264 10588 27292 10628
rect 27338 10616 27344 10668
rect 27396 10616 27402 10668
rect 27617 10659 27675 10665
rect 27617 10625 27629 10659
rect 27663 10625 27675 10659
rect 27617 10619 27675 10625
rect 27801 10659 27859 10665
rect 27801 10625 27813 10659
rect 27847 10625 27859 10659
rect 28077 10659 28135 10665
rect 28077 10656 28089 10659
rect 27801 10619 27859 10625
rect 27908 10628 28089 10656
rect 27632 10588 27660 10619
rect 27264 10560 27660 10588
rect 27157 10551 27215 10557
rect 25958 10520 25964 10532
rect 24688 10492 25728 10520
rect 25792 10492 25964 10520
rect 23937 10455 23995 10461
rect 23937 10421 23949 10455
rect 23983 10421 23995 10455
rect 23937 10415 23995 10421
rect 24949 10455 25007 10461
rect 24949 10421 24961 10455
rect 24995 10452 25007 10455
rect 25314 10452 25320 10464
rect 24995 10424 25320 10452
rect 24995 10421 25007 10424
rect 24949 10415 25007 10421
rect 25314 10412 25320 10424
rect 25372 10412 25378 10464
rect 25590 10412 25596 10464
rect 25648 10412 25654 10464
rect 25700 10452 25728 10492
rect 25958 10480 25964 10492
rect 26016 10520 26022 10532
rect 26421 10523 26479 10529
rect 26421 10520 26433 10523
rect 26016 10492 26433 10520
rect 26016 10480 26022 10492
rect 26421 10489 26433 10492
rect 26467 10489 26479 10523
rect 27172 10520 27200 10551
rect 27816 10520 27844 10619
rect 27172 10492 27844 10520
rect 26421 10483 26479 10489
rect 26142 10452 26148 10464
rect 25700 10424 26148 10452
rect 26142 10412 26148 10424
rect 26200 10412 26206 10464
rect 26234 10412 26240 10464
rect 26292 10412 26298 10464
rect 26602 10412 26608 10464
rect 26660 10452 26666 10464
rect 27065 10455 27123 10461
rect 27065 10452 27077 10455
rect 26660 10424 27077 10452
rect 26660 10412 26666 10424
rect 27065 10421 27077 10424
rect 27111 10452 27123 10455
rect 27908 10452 27936 10628
rect 28077 10625 28089 10628
rect 28123 10625 28135 10659
rect 28077 10619 28135 10625
rect 28258 10616 28264 10668
rect 28316 10616 28322 10668
rect 30377 10659 30435 10665
rect 30377 10625 30389 10659
rect 30423 10625 30435 10659
rect 30377 10619 30435 10625
rect 29546 10548 29552 10600
rect 29604 10588 29610 10600
rect 29730 10588 29736 10600
rect 29604 10560 29736 10588
rect 29604 10548 29610 10560
rect 29730 10548 29736 10560
rect 29788 10548 29794 10600
rect 30392 10588 30420 10619
rect 30466 10616 30472 10668
rect 30524 10656 30530 10668
rect 30944 10665 30972 10696
rect 31386 10684 31392 10696
rect 31444 10684 31450 10736
rect 30929 10659 30987 10665
rect 30524 10628 30696 10656
rect 30524 10616 30530 10628
rect 30392 10560 30604 10588
rect 30576 10464 30604 10560
rect 30668 10520 30696 10628
rect 30929 10625 30941 10659
rect 30975 10625 30987 10659
rect 30929 10619 30987 10625
rect 31018 10616 31024 10668
rect 31076 10616 31082 10668
rect 31478 10616 31484 10668
rect 31536 10656 31542 10668
rect 32217 10659 32275 10665
rect 32217 10656 32229 10659
rect 31536 10628 32229 10656
rect 31536 10616 31542 10628
rect 32217 10625 32229 10628
rect 32263 10625 32275 10659
rect 32217 10619 32275 10625
rect 31941 10591 31999 10597
rect 31941 10557 31953 10591
rect 31987 10588 31999 10591
rect 32122 10588 32128 10600
rect 31987 10560 32128 10588
rect 31987 10557 31999 10560
rect 31941 10551 31999 10557
rect 32122 10548 32128 10560
rect 32180 10548 32186 10600
rect 30745 10523 30803 10529
rect 30745 10520 30757 10523
rect 30668 10492 30757 10520
rect 30745 10489 30757 10492
rect 30791 10489 30803 10523
rect 30745 10483 30803 10489
rect 27111 10424 27936 10452
rect 27111 10421 27123 10424
rect 27065 10415 27123 10421
rect 29730 10412 29736 10464
rect 29788 10452 29794 10464
rect 30193 10455 30251 10461
rect 30193 10452 30205 10455
rect 29788 10424 30205 10452
rect 29788 10412 29794 10424
rect 30193 10421 30205 10424
rect 30239 10421 30251 10455
rect 30193 10415 30251 10421
rect 30558 10412 30564 10464
rect 30616 10452 30622 10464
rect 30653 10455 30711 10461
rect 30653 10452 30665 10455
rect 30616 10424 30665 10452
rect 30616 10412 30622 10424
rect 30653 10421 30665 10424
rect 30699 10421 30711 10455
rect 30653 10415 30711 10421
rect 31205 10455 31263 10461
rect 31205 10421 31217 10455
rect 31251 10452 31263 10455
rect 31570 10452 31576 10464
rect 31251 10424 31576 10452
rect 31251 10421 31263 10424
rect 31205 10415 31263 10421
rect 31570 10412 31576 10424
rect 31628 10412 31634 10464
rect 32398 10412 32404 10464
rect 32456 10412 32462 10464
rect 1104 10362 32844 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 32844 10362
rect 1104 10288 32844 10310
rect 4062 10248 4068 10260
rect 3436 10220 4068 10248
rect 3436 10053 3464 10220
rect 3605 10183 3663 10189
rect 3605 10149 3617 10183
rect 3651 10149 3663 10183
rect 3605 10143 3663 10149
rect 3620 10056 3648 10143
rect 3896 10112 3924 10220
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 4264 10220 5479 10248
rect 3970 10140 3976 10192
rect 4028 10180 4034 10192
rect 4264 10180 4292 10220
rect 4028 10152 4292 10180
rect 4341 10183 4399 10189
rect 4028 10140 4034 10152
rect 4341 10149 4353 10183
rect 4387 10180 4399 10183
rect 5350 10180 5356 10192
rect 4387 10152 5356 10180
rect 4387 10149 4399 10152
rect 4341 10143 4399 10149
rect 5350 10140 5356 10152
rect 5408 10140 5414 10192
rect 5451 10180 5479 10220
rect 5718 10208 5724 10260
rect 5776 10248 5782 10260
rect 5997 10251 6055 10257
rect 5997 10248 6009 10251
rect 5776 10220 6009 10248
rect 5776 10208 5782 10220
rect 5997 10217 6009 10220
rect 6043 10217 6055 10251
rect 5997 10211 6055 10217
rect 6086 10208 6092 10260
rect 6144 10248 6150 10260
rect 6730 10248 6736 10260
rect 6144 10220 6736 10248
rect 6144 10208 6150 10220
rect 6730 10208 6736 10220
rect 6788 10208 6794 10260
rect 8110 10248 8116 10260
rect 6932 10220 8116 10248
rect 6932 10192 6960 10220
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 9125 10251 9183 10257
rect 9125 10217 9137 10251
rect 9171 10248 9183 10251
rect 9214 10248 9220 10260
rect 9171 10220 9220 10248
rect 9171 10217 9183 10220
rect 9125 10211 9183 10217
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 9582 10208 9588 10260
rect 9640 10208 9646 10260
rect 9677 10251 9735 10257
rect 9677 10217 9689 10251
rect 9723 10248 9735 10251
rect 10134 10248 10140 10260
rect 9723 10220 10140 10248
rect 9723 10217 9735 10220
rect 9677 10211 9735 10217
rect 10134 10208 10140 10220
rect 10192 10208 10198 10260
rect 10410 10208 10416 10260
rect 10468 10248 10474 10260
rect 10781 10251 10839 10257
rect 10781 10248 10793 10251
rect 10468 10220 10793 10248
rect 10468 10208 10474 10220
rect 10781 10217 10793 10220
rect 10827 10217 10839 10251
rect 10781 10211 10839 10217
rect 12894 10208 12900 10260
rect 12952 10248 12958 10260
rect 15470 10248 15476 10260
rect 12952 10220 15476 10248
rect 12952 10208 12958 10220
rect 15470 10208 15476 10220
rect 15528 10208 15534 10260
rect 15565 10251 15623 10257
rect 15565 10217 15577 10251
rect 15611 10248 15623 10251
rect 15930 10248 15936 10260
rect 15611 10220 15936 10248
rect 15611 10217 15623 10220
rect 15565 10211 15623 10217
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 16022 10208 16028 10260
rect 16080 10208 16086 10260
rect 16942 10208 16948 10260
rect 17000 10208 17006 10260
rect 17402 10208 17408 10260
rect 17460 10208 17466 10260
rect 17494 10208 17500 10260
rect 17552 10248 17558 10260
rect 19794 10248 19800 10260
rect 17552 10220 19800 10248
rect 17552 10208 17558 10220
rect 19794 10208 19800 10220
rect 19852 10208 19858 10260
rect 19981 10251 20039 10257
rect 19981 10217 19993 10251
rect 20027 10248 20039 10251
rect 20714 10248 20720 10260
rect 20027 10220 20720 10248
rect 20027 10217 20039 10220
rect 19981 10211 20039 10217
rect 20714 10208 20720 10220
rect 20772 10208 20778 10260
rect 22278 10208 22284 10260
rect 22336 10248 22342 10260
rect 22465 10251 22523 10257
rect 22465 10248 22477 10251
rect 22336 10220 22477 10248
rect 22336 10208 22342 10220
rect 22465 10217 22477 10220
rect 22511 10248 22523 10251
rect 22511 10220 23060 10248
rect 22511 10217 22523 10220
rect 22465 10211 22523 10217
rect 6457 10183 6515 10189
rect 5451 10152 6040 10180
rect 4890 10112 4896 10124
rect 3896 10084 4896 10112
rect 4890 10072 4896 10084
rect 4948 10072 4954 10124
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10013 3479 10047
rect 3421 10007 3479 10013
rect 3602 10004 3608 10056
rect 3660 10044 3666 10056
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 3660 10016 3801 10044
rect 3660 10004 3666 10016
rect 3789 10013 3801 10016
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 3878 10004 3884 10056
rect 3936 10044 3942 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 3936 10016 4077 10044
rect 3936 10004 3942 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 4154 10004 4160 10056
rect 4212 10004 4218 10056
rect 4246 10004 4252 10056
rect 4304 10044 4310 10056
rect 5258 10044 5264 10056
rect 4304 10016 5264 10044
rect 4304 10004 4310 10016
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 5353 10047 5411 10053
rect 5353 10013 5365 10047
rect 5399 10013 5411 10047
rect 5353 10007 5411 10013
rect 3970 9936 3976 9988
rect 4028 9936 4034 9988
rect 5074 9976 5080 9988
rect 4080 9948 5080 9976
rect 3326 9868 3332 9920
rect 3384 9908 3390 9920
rect 4080 9908 4108 9948
rect 5074 9936 5080 9948
rect 5132 9936 5138 9988
rect 5368 9976 5396 10007
rect 5810 10004 5816 10056
rect 5868 10044 5874 10056
rect 5905 10047 5963 10053
rect 5905 10044 5917 10047
rect 5868 10016 5917 10044
rect 5868 10004 5874 10016
rect 5905 10013 5917 10016
rect 5951 10013 5963 10047
rect 6012 10044 6040 10152
rect 6457 10149 6469 10183
rect 6503 10180 6515 10183
rect 6638 10180 6644 10192
rect 6503 10152 6644 10180
rect 6503 10149 6515 10152
rect 6457 10143 6515 10149
rect 6638 10140 6644 10152
rect 6696 10140 6702 10192
rect 6914 10140 6920 10192
rect 6972 10140 6978 10192
rect 7101 10183 7159 10189
rect 7101 10149 7113 10183
rect 7147 10180 7159 10183
rect 7742 10180 7748 10192
rect 7147 10152 7748 10180
rect 7147 10149 7159 10152
rect 7101 10143 7159 10149
rect 7742 10140 7748 10152
rect 7800 10180 7806 10192
rect 12986 10180 12992 10192
rect 7800 10152 12992 10180
rect 7800 10140 7806 10152
rect 8478 10112 8484 10124
rect 7208 10084 8484 10112
rect 6181 10047 6239 10053
rect 6181 10044 6193 10047
rect 6012 10016 6193 10044
rect 5905 10007 5963 10013
rect 6181 10013 6193 10016
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 6270 10004 6276 10056
rect 6328 10044 6334 10056
rect 6328 10016 6868 10044
rect 6328 10004 6334 10016
rect 6840 9976 6868 10016
rect 6914 10004 6920 10056
rect 6972 10004 6978 10056
rect 7098 9976 7104 9988
rect 5368 9948 6132 9976
rect 6840 9948 7104 9976
rect 3384 9880 4108 9908
rect 3384 9868 3390 9880
rect 4890 9868 4896 9920
rect 4948 9908 4954 9920
rect 5442 9908 5448 9920
rect 4948 9880 5448 9908
rect 4948 9868 4954 9880
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 5537 9911 5595 9917
rect 5537 9877 5549 9911
rect 5583 9908 5595 9911
rect 5626 9908 5632 9920
rect 5583 9880 5632 9908
rect 5583 9877 5595 9880
rect 5537 9871 5595 9877
rect 5626 9868 5632 9880
rect 5684 9868 5690 9920
rect 5721 9911 5779 9917
rect 5721 9877 5733 9911
rect 5767 9908 5779 9911
rect 5810 9908 5816 9920
rect 5767 9880 5816 9908
rect 5767 9877 5779 9880
rect 5721 9871 5779 9877
rect 5810 9868 5816 9880
rect 5868 9868 5874 9920
rect 6104 9908 6132 9948
rect 7098 9936 7104 9948
rect 7156 9936 7162 9988
rect 7208 9908 7236 10084
rect 8478 10072 8484 10084
rect 8536 10072 8542 10124
rect 9324 10053 9352 10152
rect 12986 10140 12992 10152
rect 13044 10140 13050 10192
rect 15749 10183 15807 10189
rect 15749 10149 15761 10183
rect 15795 10180 15807 10183
rect 15795 10152 19840 10180
rect 15795 10149 15807 10152
rect 15749 10143 15807 10149
rect 9490 10072 9496 10124
rect 9548 10112 9554 10124
rect 9548 10084 9996 10112
rect 9548 10072 9554 10084
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10044 9459 10047
rect 9674 10044 9680 10056
rect 9447 10016 9680 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 6104 9880 7236 9908
rect 7558 9868 7564 9920
rect 7616 9868 7622 9920
rect 7760 9908 7788 10007
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 9858 10004 9864 10056
rect 9916 10004 9922 10056
rect 9968 10044 9996 10084
rect 10594 10072 10600 10124
rect 10652 10112 10658 10124
rect 10873 10115 10931 10121
rect 10873 10112 10885 10115
rect 10652 10084 10885 10112
rect 10652 10072 10658 10084
rect 10873 10081 10885 10084
rect 10919 10081 10931 10115
rect 10873 10075 10931 10081
rect 10962 10072 10968 10124
rect 11020 10112 11026 10124
rect 14550 10112 14556 10124
rect 11020 10084 14556 10112
rect 11020 10072 11026 10084
rect 14550 10072 14556 10084
rect 14608 10112 14614 10124
rect 15381 10115 15439 10121
rect 15381 10112 15393 10115
rect 14608 10084 15393 10112
rect 14608 10072 14614 10084
rect 15381 10081 15393 10084
rect 15427 10081 15439 10115
rect 17129 10115 17187 10121
rect 15381 10075 15439 10081
rect 15488 10084 16988 10112
rect 10781 10047 10839 10053
rect 10781 10044 10793 10047
rect 9968 10016 10793 10044
rect 10781 10013 10793 10016
rect 10827 10013 10839 10047
rect 10781 10007 10839 10013
rect 11057 10047 11115 10053
rect 11057 10013 11069 10047
rect 11103 10013 11115 10047
rect 11057 10007 11115 10013
rect 9030 9936 9036 9988
rect 9088 9976 9094 9988
rect 9585 9979 9643 9985
rect 9585 9976 9597 9979
rect 9088 9948 9597 9976
rect 9088 9936 9094 9948
rect 9585 9945 9597 9948
rect 9631 9945 9643 9979
rect 9585 9939 9643 9945
rect 10042 9936 10048 9988
rect 10100 9976 10106 9988
rect 10318 9976 10324 9988
rect 10100 9948 10324 9976
rect 10100 9936 10106 9948
rect 10318 9936 10324 9948
rect 10376 9976 10382 9988
rect 11072 9976 11100 10007
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 12710 10044 12716 10056
rect 12492 10016 12716 10044
rect 12492 10004 12498 10016
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 12894 10004 12900 10056
rect 12952 10044 12958 10056
rect 13262 10044 13268 10056
rect 12952 10016 13268 10044
rect 12952 10004 12958 10016
rect 13262 10004 13268 10016
rect 13320 10004 13326 10056
rect 15488 10044 15516 10084
rect 13372 10016 15516 10044
rect 15565 10047 15623 10053
rect 13372 9976 13400 10016
rect 15565 10013 15577 10047
rect 15611 10013 15623 10047
rect 15565 10007 15623 10013
rect 10376 9948 13400 9976
rect 10376 9936 10382 9948
rect 13814 9936 13820 9988
rect 13872 9976 13878 9988
rect 15289 9979 15347 9985
rect 15289 9976 15301 9979
rect 13872 9948 15301 9976
rect 13872 9936 13878 9948
rect 15289 9945 15301 9948
rect 15335 9945 15347 9979
rect 15580 9976 15608 10007
rect 15838 10004 15844 10056
rect 15896 10004 15902 10056
rect 16390 10004 16396 10056
rect 16448 10004 16454 10056
rect 16574 10004 16580 10056
rect 16632 10044 16638 10056
rect 16853 10047 16911 10053
rect 16853 10044 16865 10047
rect 16632 10016 16865 10044
rect 16632 10004 16638 10016
rect 16853 10013 16865 10016
rect 16899 10013 16911 10047
rect 16960 10044 16988 10084
rect 17129 10081 17141 10115
rect 17175 10112 17187 10115
rect 18046 10112 18052 10124
rect 17175 10084 18052 10112
rect 17175 10081 17187 10084
rect 17129 10075 17187 10081
rect 18046 10072 18052 10084
rect 18104 10072 18110 10124
rect 19610 10072 19616 10124
rect 19668 10072 19674 10124
rect 19812 10112 19840 10152
rect 20070 10140 20076 10192
rect 20128 10180 20134 10192
rect 20346 10180 20352 10192
rect 20128 10152 20352 10180
rect 20128 10140 20134 10152
rect 20346 10140 20352 10152
rect 20404 10140 20410 10192
rect 22097 10183 22155 10189
rect 22097 10149 22109 10183
rect 22143 10180 22155 10183
rect 22186 10180 22192 10192
rect 22143 10152 22192 10180
rect 22143 10149 22155 10152
rect 22097 10143 22155 10149
rect 22186 10140 22192 10152
rect 22244 10140 22250 10192
rect 23032 10180 23060 10220
rect 23382 10208 23388 10260
rect 23440 10248 23446 10260
rect 24673 10251 24731 10257
rect 24673 10248 24685 10251
rect 23440 10220 24685 10248
rect 23440 10208 23446 10220
rect 24673 10217 24685 10220
rect 24719 10248 24731 10251
rect 24719 10220 25360 10248
rect 24719 10217 24731 10220
rect 24673 10211 24731 10217
rect 25332 10180 25360 10220
rect 27706 10208 27712 10260
rect 27764 10208 27770 10260
rect 29638 10208 29644 10260
rect 29696 10208 29702 10260
rect 23032 10152 24716 10180
rect 25332 10152 28488 10180
rect 22646 10112 22652 10124
rect 19812 10084 21772 10112
rect 17221 10047 17279 10053
rect 17221 10044 17233 10047
rect 16960 10016 17233 10044
rect 16853 10007 16911 10013
rect 17221 10013 17233 10016
rect 17267 10013 17279 10047
rect 18509 10047 18567 10053
rect 18509 10044 18521 10047
rect 17221 10007 17279 10013
rect 17328 10016 18521 10044
rect 16022 9976 16028 9988
rect 15580 9948 16028 9976
rect 15289 9939 15347 9945
rect 16022 9936 16028 9948
rect 16080 9936 16086 9988
rect 16482 9936 16488 9988
rect 16540 9976 16546 9988
rect 16945 9979 17003 9985
rect 16945 9976 16957 9979
rect 16540 9948 16957 9976
rect 16540 9936 16546 9948
rect 16945 9945 16957 9948
rect 16991 9945 17003 9979
rect 16945 9939 17003 9945
rect 17126 9936 17132 9988
rect 17184 9976 17190 9988
rect 17328 9976 17356 10016
rect 18509 10013 18521 10016
rect 18555 10013 18567 10047
rect 18509 10007 18567 10013
rect 19150 10004 19156 10056
rect 19208 10044 19214 10056
rect 19245 10047 19303 10053
rect 19981 10047 20039 10053
rect 19245 10044 19257 10047
rect 19208 10016 19257 10044
rect 19208 10004 19214 10016
rect 19245 10013 19257 10016
rect 19291 10013 19303 10047
rect 19245 10007 19303 10013
rect 19802 10041 19860 10047
rect 19802 10007 19814 10041
rect 19848 10038 19860 10041
rect 19848 10010 19932 10038
rect 19848 10007 19860 10010
rect 19802 10001 19860 10007
rect 19334 9976 19340 9988
rect 17184 9948 17356 9976
rect 17926 9948 19340 9976
rect 17184 9936 17190 9948
rect 8846 9908 8852 9920
rect 7760 9880 8852 9908
rect 8846 9868 8852 9880
rect 8904 9908 8910 9920
rect 10870 9908 10876 9920
rect 8904 9880 10876 9908
rect 8904 9868 8910 9880
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 11238 9868 11244 9920
rect 11296 9868 11302 9920
rect 16574 9868 16580 9920
rect 16632 9868 16638 9920
rect 16666 9868 16672 9920
rect 16724 9908 16730 9920
rect 17926 9908 17954 9948
rect 19334 9936 19340 9948
rect 19392 9936 19398 9988
rect 19426 9936 19432 9988
rect 19484 9936 19490 9988
rect 19904 9976 19932 10010
rect 19981 10013 19993 10047
rect 20027 10044 20039 10047
rect 20346 10044 20352 10056
rect 20027 10016 20352 10044
rect 20027 10013 20039 10016
rect 19981 10007 20039 10013
rect 20346 10004 20352 10016
rect 20404 10004 20410 10056
rect 20070 9976 20076 9988
rect 19904 9948 20076 9976
rect 20070 9936 20076 9948
rect 20128 9936 20134 9988
rect 21744 9976 21772 10084
rect 22296 10084 22652 10112
rect 22296 10053 22324 10084
rect 22646 10072 22652 10084
rect 22704 10072 22710 10124
rect 22922 10072 22928 10124
rect 22980 10112 22986 10124
rect 22980 10084 24440 10112
rect 22980 10072 22986 10084
rect 22281 10047 22339 10053
rect 22281 10013 22293 10047
rect 22327 10013 22339 10047
rect 22281 10007 22339 10013
rect 22373 10047 22431 10053
rect 22373 10013 22385 10047
rect 22419 10013 22431 10047
rect 22373 10007 22431 10013
rect 22388 9976 22416 10007
rect 22554 10004 22560 10056
rect 22612 10004 22618 10056
rect 22830 10004 22836 10056
rect 22888 10044 22894 10056
rect 24210 10044 24216 10056
rect 22888 10016 24216 10044
rect 22888 10004 22894 10016
rect 24210 10004 24216 10016
rect 24268 10004 24274 10056
rect 24412 10053 24440 10084
rect 24486 10072 24492 10124
rect 24544 10072 24550 10124
rect 24688 10053 24716 10152
rect 27709 10115 27767 10121
rect 27709 10081 27721 10115
rect 27755 10112 27767 10115
rect 28350 10112 28356 10124
rect 27755 10084 28356 10112
rect 27755 10081 27767 10084
rect 27709 10075 27767 10081
rect 28350 10072 28356 10084
rect 28408 10072 28414 10124
rect 28460 10112 28488 10152
rect 28626 10140 28632 10192
rect 28684 10180 28690 10192
rect 28684 10152 30236 10180
rect 28684 10140 28690 10152
rect 29641 10115 29699 10121
rect 29641 10112 29653 10115
rect 28460 10084 29653 10112
rect 29641 10081 29653 10084
rect 29687 10081 29699 10115
rect 29641 10075 29699 10081
rect 24397 10047 24455 10053
rect 24397 10013 24409 10047
rect 24443 10013 24455 10047
rect 24397 10007 24455 10013
rect 24673 10047 24731 10053
rect 24673 10013 24685 10047
rect 24719 10013 24731 10047
rect 24673 10007 24731 10013
rect 26510 10004 26516 10056
rect 26568 10044 26574 10056
rect 27522 10044 27528 10056
rect 26568 10016 27528 10044
rect 26568 10004 26574 10016
rect 27522 10004 27528 10016
rect 27580 10004 27586 10056
rect 27982 10004 27988 10056
rect 28040 10044 28046 10056
rect 29549 10047 29607 10053
rect 29549 10044 29561 10047
rect 28040 10016 29561 10044
rect 28040 10004 28046 10016
rect 29549 10013 29561 10016
rect 29595 10013 29607 10047
rect 29549 10007 29607 10013
rect 29825 10047 29883 10053
rect 29825 10013 29837 10047
rect 29871 10044 29883 10047
rect 30098 10044 30104 10056
rect 29871 10016 30104 10044
rect 29871 10013 29883 10016
rect 29825 10007 29883 10013
rect 30098 10004 30104 10016
rect 30156 10004 30162 10056
rect 30208 10053 30236 10152
rect 31849 10115 31907 10121
rect 31849 10112 31861 10115
rect 30576 10084 31861 10112
rect 30576 10053 30604 10084
rect 31849 10081 31861 10084
rect 31895 10081 31907 10115
rect 31849 10075 31907 10081
rect 30193 10047 30251 10053
rect 30193 10013 30205 10047
rect 30239 10013 30251 10047
rect 30193 10007 30251 10013
rect 30561 10047 30619 10053
rect 30561 10013 30573 10047
rect 30607 10013 30619 10047
rect 30561 10007 30619 10013
rect 31478 10004 31484 10056
rect 31536 10004 31542 10056
rect 31570 10004 31576 10056
rect 31628 10004 31634 10056
rect 32490 10004 32496 10056
rect 32548 10004 32554 10056
rect 24762 9976 24768 9988
rect 21744 9948 24768 9976
rect 24762 9936 24768 9948
rect 24820 9936 24826 9988
rect 27154 9936 27160 9988
rect 27212 9976 27218 9988
rect 27801 9979 27859 9985
rect 27801 9976 27813 9979
rect 27212 9948 27813 9976
rect 27212 9936 27218 9948
rect 27801 9945 27813 9948
rect 27847 9945 27859 9979
rect 27801 9939 27859 9945
rect 29730 9936 29736 9988
rect 29788 9976 29794 9988
rect 30377 9979 30435 9985
rect 30377 9976 30389 9979
rect 29788 9948 30389 9976
rect 29788 9936 29794 9948
rect 30377 9945 30389 9948
rect 30423 9945 30435 9979
rect 30377 9939 30435 9945
rect 30466 9936 30472 9988
rect 30524 9936 30530 9988
rect 30650 9936 30656 9988
rect 30708 9976 30714 9988
rect 30837 9979 30895 9985
rect 30837 9976 30849 9979
rect 30708 9948 30849 9976
rect 30708 9936 30714 9948
rect 30837 9945 30849 9948
rect 30883 9945 30895 9979
rect 30837 9939 30895 9945
rect 16724 9880 17954 9908
rect 16724 9868 16730 9880
rect 18230 9868 18236 9920
rect 18288 9908 18294 9920
rect 18325 9911 18383 9917
rect 18325 9908 18337 9911
rect 18288 9880 18337 9908
rect 18288 9868 18294 9880
rect 18325 9877 18337 9880
rect 18371 9877 18383 9911
rect 18325 9871 18383 9877
rect 20165 9911 20223 9917
rect 20165 9877 20177 9911
rect 20211 9908 20223 9911
rect 20438 9908 20444 9920
rect 20211 9880 20444 9908
rect 20211 9877 20223 9880
rect 20165 9871 20223 9877
rect 20438 9868 20444 9880
rect 20496 9908 20502 9920
rect 24670 9908 24676 9920
rect 20496 9880 24676 9908
rect 20496 9868 20502 9880
rect 24670 9868 24676 9880
rect 24728 9868 24734 9920
rect 24857 9911 24915 9917
rect 24857 9877 24869 9911
rect 24903 9908 24915 9911
rect 25958 9908 25964 9920
rect 24903 9880 25964 9908
rect 24903 9877 24915 9880
rect 24857 9871 24915 9877
rect 25958 9868 25964 9880
rect 26016 9868 26022 9920
rect 27338 9868 27344 9920
rect 27396 9868 27402 9920
rect 29914 9868 29920 9920
rect 29972 9908 29978 9920
rect 30009 9911 30067 9917
rect 30009 9908 30021 9911
rect 29972 9880 30021 9908
rect 29972 9868 29978 9880
rect 30009 9877 30021 9880
rect 30055 9877 30067 9911
rect 30009 9871 30067 9877
rect 30742 9868 30748 9920
rect 30800 9868 30806 9920
rect 31757 9911 31815 9917
rect 31757 9877 31769 9911
rect 31803 9908 31815 9911
rect 31846 9908 31852 9920
rect 31803 9880 31852 9908
rect 31803 9877 31815 9880
rect 31757 9871 31815 9877
rect 31846 9868 31852 9880
rect 31904 9868 31910 9920
rect 1104 9818 32844 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 32844 9818
rect 1104 9744 32844 9766
rect 3878 9704 3884 9716
rect 3344 9676 3884 9704
rect 2774 9528 2780 9580
rect 2832 9568 2838 9580
rect 3344 9577 3372 9676
rect 3878 9664 3884 9676
rect 3936 9664 3942 9716
rect 4525 9707 4583 9713
rect 4525 9673 4537 9707
rect 4571 9704 4583 9707
rect 4706 9704 4712 9716
rect 4571 9676 4712 9704
rect 4571 9673 4583 9676
rect 4525 9667 4583 9673
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 5350 9704 5356 9716
rect 5276 9676 5356 9704
rect 3602 9596 3608 9648
rect 3660 9636 3666 9648
rect 4249 9639 4307 9645
rect 4249 9636 4261 9639
rect 3660 9608 4261 9636
rect 3660 9596 3666 9608
rect 4249 9605 4261 9608
rect 4295 9636 4307 9639
rect 4295 9608 4936 9636
rect 4295 9605 4307 9608
rect 4249 9599 4307 9605
rect 3053 9571 3111 9577
rect 3053 9568 3065 9571
rect 2832 9540 3065 9568
rect 2832 9528 2838 9540
rect 3053 9537 3065 9540
rect 3099 9537 3111 9571
rect 3053 9531 3111 9537
rect 3329 9571 3387 9577
rect 3329 9537 3341 9571
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 3510 9528 3516 9580
rect 3568 9528 3574 9580
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9537 3755 9571
rect 3697 9531 3755 9537
rect 3418 9460 3424 9512
rect 3476 9500 3482 9512
rect 3712 9500 3740 9531
rect 3878 9528 3884 9580
rect 3936 9568 3942 9580
rect 3973 9571 4031 9577
rect 3973 9568 3985 9571
rect 3936 9540 3985 9568
rect 3936 9528 3942 9540
rect 3973 9537 3985 9540
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9537 4215 9571
rect 4157 9531 4215 9537
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9568 4399 9571
rect 4798 9568 4804 9580
rect 4387 9540 4804 9568
rect 4387 9537 4399 9540
rect 4341 9531 4399 9537
rect 3476 9472 3740 9500
rect 3476 9460 3482 9472
rect 4062 9460 4068 9512
rect 4120 9500 4126 9512
rect 4172 9500 4200 9531
rect 4246 9500 4252 9512
rect 4120 9472 4252 9500
rect 4120 9460 4126 9472
rect 4246 9460 4252 9472
rect 4304 9460 4310 9512
rect 3237 9435 3295 9441
rect 3237 9401 3249 9435
rect 3283 9432 3295 9435
rect 4356 9432 4384 9531
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 4908 9500 4936 9608
rect 5276 9577 5304 9676
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 5718 9704 5724 9716
rect 5552 9676 5724 9704
rect 5552 9645 5580 9676
rect 5718 9664 5724 9676
rect 5776 9704 5782 9716
rect 5776 9676 5948 9704
rect 5776 9664 5782 9676
rect 5537 9639 5595 9645
rect 5537 9605 5549 9639
rect 5583 9605 5595 9639
rect 5537 9599 5595 9605
rect 5629 9639 5687 9645
rect 5629 9605 5641 9639
rect 5675 9636 5687 9639
rect 5810 9636 5816 9648
rect 5675 9608 5816 9636
rect 5675 9605 5687 9608
rect 5629 9599 5687 9605
rect 5810 9596 5816 9608
rect 5868 9596 5874 9648
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9537 5319 9571
rect 5261 9531 5319 9537
rect 5353 9571 5411 9577
rect 5353 9537 5365 9571
rect 5399 9537 5411 9571
rect 5721 9571 5779 9577
rect 5721 9568 5733 9571
rect 5353 9531 5411 9537
rect 5451 9540 5733 9568
rect 5368 9500 5396 9531
rect 4908 9472 5396 9500
rect 3283 9404 4384 9432
rect 3283 9401 3295 9404
rect 3237 9395 3295 9401
rect 3804 9376 3832 9404
rect 4706 9392 4712 9444
rect 4764 9432 4770 9444
rect 5077 9435 5135 9441
rect 5077 9432 5089 9435
rect 4764 9404 5089 9432
rect 4764 9392 4770 9404
rect 5077 9401 5089 9404
rect 5123 9401 5135 9435
rect 5077 9395 5135 9401
rect 5258 9392 5264 9444
rect 5316 9432 5322 9444
rect 5451 9432 5479 9540
rect 5721 9537 5733 9540
rect 5767 9568 5779 9571
rect 5920 9572 5948 9676
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 6730 9704 6736 9716
rect 6052 9676 6736 9704
rect 6052 9664 6058 9676
rect 6730 9664 6736 9676
rect 6788 9664 6794 9716
rect 6825 9707 6883 9713
rect 6825 9673 6837 9707
rect 6871 9673 6883 9707
rect 6825 9667 6883 9673
rect 8757 9707 8815 9713
rect 8757 9673 8769 9707
rect 8803 9704 8815 9707
rect 9214 9704 9220 9716
rect 8803 9676 9220 9704
rect 8803 9673 8815 9676
rect 8757 9667 8815 9673
rect 6270 9596 6276 9648
rect 6328 9636 6334 9648
rect 6840 9636 6868 9667
rect 9214 9664 9220 9676
rect 9272 9664 9278 9716
rect 9306 9664 9312 9716
rect 9364 9704 9370 9716
rect 10042 9704 10048 9716
rect 9364 9676 10048 9704
rect 9364 9664 9370 9676
rect 10042 9664 10048 9676
rect 10100 9664 10106 9716
rect 10689 9707 10747 9713
rect 10689 9673 10701 9707
rect 10735 9704 10747 9707
rect 10962 9704 10968 9716
rect 10735 9676 10968 9704
rect 10735 9673 10747 9676
rect 10689 9667 10747 9673
rect 10962 9664 10968 9676
rect 11020 9664 11026 9716
rect 11057 9707 11115 9713
rect 11057 9673 11069 9707
rect 11103 9673 11115 9707
rect 11057 9667 11115 9673
rect 12437 9707 12495 9713
rect 12437 9673 12449 9707
rect 12483 9704 12495 9707
rect 12526 9704 12532 9716
rect 12483 9676 12532 9704
rect 12483 9673 12495 9676
rect 12437 9667 12495 9673
rect 7193 9639 7251 9645
rect 7193 9636 7205 9639
rect 6328 9608 6800 9636
rect 6840 9608 7205 9636
rect 6328 9596 6334 9608
rect 5989 9575 6047 9581
rect 5989 9572 6001 9575
rect 5767 9540 5856 9568
rect 5920 9544 6001 9572
rect 5767 9537 5779 9540
rect 5721 9531 5779 9537
rect 5828 9500 5856 9540
rect 5989 9541 6001 9544
rect 6035 9541 6047 9575
rect 5989 9535 6047 9541
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9537 6423 9571
rect 6365 9531 6423 9537
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9537 6699 9571
rect 6772 9568 6800 9608
rect 7193 9605 7205 9608
rect 7239 9636 7251 9639
rect 8481 9639 8539 9645
rect 8481 9636 8493 9639
rect 7239 9608 8493 9636
rect 7239 9605 7251 9608
rect 7193 9599 7251 9605
rect 6917 9571 6975 9577
rect 6917 9568 6929 9571
rect 6772 9540 6929 9568
rect 6641 9531 6699 9537
rect 6917 9537 6929 9540
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 6380 9500 6408 9531
rect 5828 9472 6408 9500
rect 6656 9432 6684 9531
rect 6932 9500 6960 9531
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 7064 9540 7113 9568
rect 7064 9528 7070 9540
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 7282 9528 7288 9580
rect 7340 9528 7346 9580
rect 7576 9577 7604 9608
rect 8481 9605 8493 9608
rect 8527 9605 8539 9639
rect 8481 9599 8539 9605
rect 8938 9596 8944 9648
rect 8996 9636 9002 9648
rect 11072 9636 11100 9667
rect 12526 9664 12532 9676
rect 12584 9704 12590 9716
rect 15838 9704 15844 9716
rect 12584 9676 15844 9704
rect 12584 9664 12590 9676
rect 15838 9664 15844 9676
rect 15896 9664 15902 9716
rect 16482 9664 16488 9716
rect 16540 9664 16546 9716
rect 16666 9704 16672 9716
rect 16592 9676 16672 9704
rect 12894 9636 12900 9648
rect 8996 9608 10180 9636
rect 8996 9596 9002 9608
rect 7561 9571 7619 9577
rect 7561 9537 7573 9571
rect 7607 9537 7619 9571
rect 7561 9531 7619 9537
rect 7650 9528 7656 9580
rect 7708 9568 7714 9580
rect 7745 9571 7803 9577
rect 7745 9568 7757 9571
rect 7708 9540 7757 9568
rect 7708 9528 7714 9540
rect 7745 9537 7757 9540
rect 7791 9537 7803 9571
rect 7745 9531 7803 9537
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9537 7895 9571
rect 7837 9531 7895 9537
rect 7852 9500 7880 9531
rect 7926 9528 7932 9580
rect 7984 9528 7990 9580
rect 8205 9571 8263 9577
rect 8205 9537 8217 9571
rect 8251 9537 8263 9571
rect 8205 9531 8263 9537
rect 8389 9571 8447 9577
rect 8389 9537 8401 9571
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 8573 9571 8631 9577
rect 8573 9537 8585 9571
rect 8619 9568 8631 9571
rect 9858 9568 9864 9580
rect 8619 9540 9864 9568
rect 8619 9537 8631 9540
rect 8573 9531 8631 9537
rect 8220 9500 8248 9531
rect 6932 9472 8248 9500
rect 5316 9404 5479 9432
rect 5828 9404 6684 9432
rect 5316 9392 5322 9404
rect 3786 9324 3792 9376
rect 3844 9324 3850 9376
rect 3881 9367 3939 9373
rect 3881 9333 3893 9367
rect 3927 9364 3939 9367
rect 5166 9364 5172 9376
rect 3927 9336 5172 9364
rect 3927 9333 3939 9336
rect 3881 9327 3939 9333
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 5828 9364 5856 9404
rect 7282 9392 7288 9444
rect 7340 9432 7346 9444
rect 7742 9432 7748 9444
rect 7340 9404 7748 9432
rect 7340 9392 7346 9404
rect 7742 9392 7748 9404
rect 7800 9432 7806 9444
rect 7926 9432 7932 9444
rect 7800 9404 7932 9432
rect 7800 9392 7806 9404
rect 7926 9392 7932 9404
rect 7984 9392 7990 9444
rect 8113 9435 8171 9441
rect 8113 9401 8125 9435
rect 8159 9432 8171 9435
rect 8294 9432 8300 9444
rect 8159 9404 8300 9432
rect 8159 9401 8171 9404
rect 8113 9395 8171 9401
rect 8294 9392 8300 9404
rect 8352 9392 8358 9444
rect 5500 9336 5856 9364
rect 5905 9367 5963 9373
rect 5500 9324 5506 9336
rect 5905 9333 5917 9367
rect 5951 9364 5963 9367
rect 6086 9364 6092 9376
rect 5951 9336 6092 9364
rect 5951 9333 5963 9336
rect 5905 9327 5963 9333
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 6181 9367 6239 9373
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 6454 9364 6460 9376
rect 6227 9336 6460 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 6549 9367 6607 9373
rect 6549 9333 6561 9367
rect 6595 9364 6607 9367
rect 6638 9364 6644 9376
rect 6595 9336 6644 9364
rect 6595 9333 6607 9336
rect 6549 9327 6607 9333
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 7466 9324 7472 9376
rect 7524 9324 7530 9376
rect 7558 9324 7564 9376
rect 7616 9364 7622 9376
rect 8404 9364 8432 9531
rect 9858 9528 9864 9540
rect 9916 9528 9922 9580
rect 10042 9528 10048 9580
rect 10100 9528 10106 9580
rect 10152 9577 10180 9608
rect 10336 9608 11100 9636
rect 11992 9608 12900 9636
rect 10336 9580 10364 9608
rect 10137 9571 10195 9577
rect 10137 9537 10149 9571
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 10318 9528 10324 9580
rect 10376 9528 10382 9580
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 8938 9460 8944 9512
rect 8996 9460 9002 9512
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9500 9275 9503
rect 9490 9500 9496 9512
rect 9263 9472 9496 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 9582 9460 9588 9512
rect 9640 9500 9646 9512
rect 10428 9500 10456 9531
rect 10502 9528 10508 9580
rect 10560 9528 10566 9580
rect 10962 9528 10968 9580
rect 11020 9528 11026 9580
rect 11992 9577 12020 9608
rect 12894 9596 12900 9608
rect 12952 9596 12958 9648
rect 12986 9596 12992 9648
rect 13044 9636 13050 9648
rect 14366 9636 14372 9648
rect 13044 9608 14372 9636
rect 13044 9596 13050 9608
rect 14366 9596 14372 9608
rect 14424 9596 14430 9648
rect 16592 9636 16620 9676
rect 16666 9664 16672 9676
rect 16724 9664 16730 9716
rect 18601 9707 18659 9713
rect 18601 9673 18613 9707
rect 18647 9704 18659 9707
rect 19150 9704 19156 9716
rect 18647 9676 19156 9704
rect 18647 9673 18659 9676
rect 18601 9667 18659 9673
rect 19150 9664 19156 9676
rect 19208 9664 19214 9716
rect 20073 9707 20131 9713
rect 20073 9704 20085 9707
rect 20031 9676 20085 9704
rect 20073 9673 20085 9676
rect 20119 9704 20131 9707
rect 20530 9704 20536 9716
rect 20119 9676 20536 9704
rect 20119 9673 20131 9676
rect 20073 9667 20131 9673
rect 20088 9636 20116 9667
rect 20530 9664 20536 9676
rect 20588 9664 20594 9716
rect 30466 9704 30472 9716
rect 29840 9676 30472 9704
rect 15948 9608 16620 9636
rect 17604 9608 18368 9636
rect 11241 9571 11299 9577
rect 11241 9537 11253 9571
rect 11287 9537 11299 9571
rect 11241 9531 11299 9537
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9537 12035 9571
rect 12253 9571 12311 9577
rect 12253 9568 12265 9571
rect 11977 9531 12035 9537
rect 12084 9540 12265 9568
rect 9640 9472 10456 9500
rect 9640 9460 9646 9472
rect 10870 9460 10876 9512
rect 10928 9500 10934 9512
rect 11256 9500 11284 9531
rect 10928 9472 11284 9500
rect 10928 9460 10934 9472
rect 9122 9392 9128 9444
rect 9180 9432 9186 9444
rect 9180 9404 9904 9432
rect 9180 9392 9186 9404
rect 9674 9364 9680 9376
rect 7616 9336 9680 9364
rect 7616 9324 7622 9336
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 9876 9373 9904 9404
rect 10502 9392 10508 9444
rect 10560 9432 10566 9444
rect 10781 9435 10839 9441
rect 10781 9432 10793 9435
rect 10560 9404 10793 9432
rect 10560 9392 10566 9404
rect 10781 9401 10793 9404
rect 10827 9401 10839 9435
rect 10781 9395 10839 9401
rect 11146 9392 11152 9444
rect 11204 9432 11210 9444
rect 12084 9432 12112 9540
rect 12253 9537 12265 9540
rect 12299 9537 12311 9571
rect 12253 9531 12311 9537
rect 12802 9528 12808 9580
rect 12860 9528 12866 9580
rect 13078 9528 13084 9580
rect 13136 9528 13142 9580
rect 13354 9528 13360 9580
rect 13412 9528 13418 9580
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 13817 9571 13875 9577
rect 13817 9568 13829 9571
rect 13587 9540 13829 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 13817 9537 13829 9540
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9568 14059 9571
rect 15562 9568 15568 9580
rect 14047 9540 15568 9568
rect 14047 9537 14059 9540
rect 14001 9531 14059 9537
rect 12989 9503 13047 9509
rect 12989 9469 13001 9503
rect 13035 9500 13047 9503
rect 13170 9500 13176 9512
rect 13035 9472 13176 9500
rect 13035 9469 13047 9472
rect 12989 9463 13047 9469
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 13556 9500 13584 9531
rect 13280 9472 13584 9500
rect 11204 9404 12112 9432
rect 12161 9435 12219 9441
rect 11204 9392 11210 9404
rect 12161 9401 12173 9435
rect 12207 9432 12219 9435
rect 12434 9432 12440 9444
rect 12207 9404 12440 9432
rect 12207 9401 12219 9404
rect 12161 9395 12219 9401
rect 12434 9392 12440 9404
rect 12492 9392 12498 9444
rect 13280 9441 13308 9472
rect 13722 9460 13728 9512
rect 13780 9500 13786 9512
rect 14016 9500 14044 9531
rect 15562 9528 15568 9540
rect 15620 9528 15626 9580
rect 13780 9472 14044 9500
rect 15948 9500 15976 9608
rect 16022 9528 16028 9580
rect 16080 9528 16086 9580
rect 16301 9571 16359 9577
rect 16301 9537 16313 9571
rect 16347 9568 16359 9571
rect 16574 9568 16580 9580
rect 16347 9540 16580 9568
rect 16347 9537 16359 9540
rect 16301 9531 16359 9537
rect 16574 9528 16580 9540
rect 16632 9568 16638 9580
rect 17604 9568 17632 9608
rect 18340 9580 18368 9608
rect 19444 9608 20116 9636
rect 16632 9540 17632 9568
rect 17773 9571 17831 9577
rect 16632 9528 16638 9540
rect 17773 9537 17785 9571
rect 17819 9568 17831 9571
rect 17862 9568 17868 9580
rect 17819 9540 17868 9568
rect 17819 9537 17831 9540
rect 17773 9531 17831 9537
rect 17862 9528 17868 9540
rect 17920 9528 17926 9580
rect 17957 9571 18015 9577
rect 17957 9537 17969 9571
rect 18003 9568 18015 9571
rect 18138 9568 18144 9580
rect 18003 9540 18144 9568
rect 18003 9537 18015 9540
rect 17957 9531 18015 9537
rect 18138 9528 18144 9540
rect 18196 9528 18202 9580
rect 18230 9528 18236 9580
rect 18288 9528 18294 9580
rect 18322 9528 18328 9580
rect 18380 9568 18386 9580
rect 19444 9577 19472 9608
rect 20254 9596 20260 9648
rect 20312 9636 20318 9648
rect 25225 9639 25283 9645
rect 20312 9608 20944 9636
rect 20312 9596 20318 9608
rect 20916 9580 20944 9608
rect 21008 9608 25176 9636
rect 18417 9571 18475 9577
rect 18417 9568 18429 9571
rect 18380 9540 18429 9568
rect 18380 9528 18386 9540
rect 18417 9537 18429 9540
rect 18463 9537 18475 9571
rect 18417 9531 18475 9537
rect 19429 9571 19487 9577
rect 19429 9537 19441 9571
rect 19475 9537 19487 9571
rect 19429 9531 19487 9537
rect 19794 9528 19800 9580
rect 19852 9568 19858 9580
rect 19889 9571 19947 9577
rect 19889 9568 19901 9571
rect 19852 9540 19901 9568
rect 19852 9528 19858 9540
rect 19889 9537 19901 9540
rect 19935 9537 19947 9571
rect 19889 9531 19947 9537
rect 19978 9528 19984 9580
rect 20036 9568 20042 9580
rect 20438 9568 20444 9580
rect 20036 9540 20444 9568
rect 20036 9528 20042 9540
rect 20438 9528 20444 9540
rect 20496 9528 20502 9580
rect 20898 9528 20904 9580
rect 20956 9528 20962 9580
rect 16117 9503 16175 9509
rect 16117 9500 16129 9503
rect 15948 9472 16129 9500
rect 13780 9460 13786 9472
rect 16117 9469 16129 9472
rect 16163 9469 16175 9503
rect 16117 9463 16175 9469
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 16724 9472 17908 9500
rect 16724 9460 16730 9472
rect 13265 9435 13323 9441
rect 12912 9404 13216 9432
rect 9861 9367 9919 9373
rect 9861 9333 9873 9367
rect 9907 9364 9919 9367
rect 12912 9364 12940 9404
rect 9907 9336 12940 9364
rect 9907 9333 9919 9336
rect 9861 9327 9919 9333
rect 12986 9324 12992 9376
rect 13044 9324 13050 9376
rect 13188 9364 13216 9404
rect 13265 9401 13277 9435
rect 13311 9401 13323 9435
rect 17770 9432 17776 9444
rect 13265 9395 13323 9401
rect 13464 9404 17776 9432
rect 13464 9364 13492 9404
rect 17770 9392 17776 9404
rect 17828 9392 17834 9444
rect 17880 9432 17908 9472
rect 18966 9460 18972 9512
rect 19024 9500 19030 9512
rect 19521 9503 19579 9509
rect 19521 9500 19533 9503
rect 19024 9472 19533 9500
rect 19024 9460 19030 9472
rect 19521 9469 19533 9472
rect 19567 9469 19579 9503
rect 21008 9500 21036 9608
rect 21085 9571 21143 9577
rect 21085 9537 21097 9571
rect 21131 9568 21143 9571
rect 21174 9568 21180 9580
rect 21131 9540 21180 9568
rect 21131 9537 21143 9540
rect 21085 9531 21143 9537
rect 21174 9528 21180 9540
rect 21232 9528 21238 9580
rect 21450 9528 21456 9580
rect 21508 9528 21514 9580
rect 21910 9528 21916 9580
rect 21968 9528 21974 9580
rect 22186 9528 22192 9580
rect 22244 9528 22250 9580
rect 23014 9528 23020 9580
rect 23072 9528 23078 9580
rect 24949 9571 25007 9577
rect 24949 9568 24961 9571
rect 24412 9540 24961 9568
rect 19521 9463 19579 9469
rect 19628 9472 21036 9500
rect 21269 9503 21327 9509
rect 19628 9432 19656 9472
rect 21269 9469 21281 9503
rect 21315 9500 21327 9503
rect 21542 9500 21548 9512
rect 21315 9472 21548 9500
rect 21315 9469 21327 9472
rect 21269 9463 21327 9469
rect 21542 9460 21548 9472
rect 21600 9460 21606 9512
rect 22097 9503 22155 9509
rect 22097 9469 22109 9503
rect 22143 9500 22155 9503
rect 22738 9500 22744 9512
rect 22143 9472 22744 9500
rect 22143 9469 22155 9472
rect 22097 9463 22155 9469
rect 22738 9460 22744 9472
rect 22796 9460 22802 9512
rect 22925 9503 22983 9509
rect 22925 9469 22937 9503
rect 22971 9500 22983 9503
rect 24302 9500 24308 9512
rect 22971 9472 24308 9500
rect 22971 9469 22983 9472
rect 22925 9463 22983 9469
rect 24302 9460 24308 9472
rect 24360 9460 24366 9512
rect 17880 9404 19656 9432
rect 19797 9435 19855 9441
rect 19797 9401 19809 9435
rect 19843 9432 19855 9435
rect 19843 9404 19932 9432
rect 19843 9401 19855 9404
rect 19797 9395 19855 9401
rect 13188 9336 13492 9364
rect 13541 9367 13599 9373
rect 13541 9333 13553 9367
rect 13587 9364 13599 9367
rect 14090 9364 14096 9376
rect 13587 9336 14096 9364
rect 13587 9333 13599 9336
rect 13541 9327 13599 9333
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 14185 9367 14243 9373
rect 14185 9333 14197 9367
rect 14231 9364 14243 9367
rect 14826 9364 14832 9376
rect 14231 9336 14832 9364
rect 14231 9333 14243 9336
rect 14185 9327 14243 9333
rect 14826 9324 14832 9336
rect 14884 9324 14890 9376
rect 16114 9324 16120 9376
rect 16172 9364 16178 9376
rect 16301 9367 16359 9373
rect 16301 9364 16313 9367
rect 16172 9336 16313 9364
rect 16172 9324 16178 9336
rect 16301 9333 16313 9336
rect 16347 9364 16359 9367
rect 16574 9364 16580 9376
rect 16347 9336 16580 9364
rect 16347 9333 16359 9336
rect 16301 9327 16359 9333
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 18138 9324 18144 9376
rect 18196 9324 18202 9376
rect 19334 9324 19340 9376
rect 19392 9364 19398 9376
rect 19429 9367 19487 9373
rect 19429 9364 19441 9367
rect 19392 9336 19441 9364
rect 19392 9324 19398 9336
rect 19429 9333 19441 9336
rect 19475 9333 19487 9367
rect 19904 9364 19932 9404
rect 19978 9392 19984 9444
rect 20036 9432 20042 9444
rect 21726 9432 21732 9444
rect 20036 9404 21732 9432
rect 20036 9392 20042 9404
rect 21726 9392 21732 9404
rect 21784 9392 21790 9444
rect 22649 9435 22707 9441
rect 22649 9432 22661 9435
rect 22204 9404 22661 9432
rect 20990 9364 20996 9376
rect 19904 9336 20996 9364
rect 19429 9327 19487 9333
rect 20990 9324 20996 9336
rect 21048 9324 21054 9376
rect 21637 9367 21695 9373
rect 21637 9333 21649 9367
rect 21683 9364 21695 9367
rect 22002 9364 22008 9376
rect 21683 9336 22008 9364
rect 21683 9333 21695 9336
rect 21637 9327 21695 9333
rect 22002 9324 22008 9336
rect 22060 9324 22066 9376
rect 22204 9373 22232 9404
rect 22649 9401 22661 9404
rect 22695 9401 22707 9435
rect 22649 9395 22707 9401
rect 22189 9367 22247 9373
rect 22189 9333 22201 9367
rect 22235 9333 22247 9367
rect 22189 9327 22247 9333
rect 22278 9324 22284 9376
rect 22336 9364 22342 9376
rect 22373 9367 22431 9373
rect 22373 9364 22385 9367
rect 22336 9336 22385 9364
rect 22336 9324 22342 9336
rect 22373 9333 22385 9336
rect 22419 9333 22431 9367
rect 22373 9327 22431 9333
rect 22554 9324 22560 9376
rect 22612 9364 22618 9376
rect 22833 9367 22891 9373
rect 22833 9364 22845 9367
rect 22612 9336 22845 9364
rect 22612 9324 22618 9336
rect 22833 9333 22845 9336
rect 22879 9364 22891 9367
rect 24412 9364 24440 9540
rect 24949 9537 24961 9540
rect 24995 9537 25007 9571
rect 24949 9531 25007 9537
rect 24670 9460 24676 9512
rect 24728 9500 24734 9512
rect 25041 9503 25099 9509
rect 25041 9500 25053 9503
rect 24728 9472 25053 9500
rect 24728 9460 24734 9472
rect 25041 9469 25053 9472
rect 25087 9469 25099 9503
rect 25148 9500 25176 9608
rect 25225 9605 25237 9639
rect 25271 9636 25283 9639
rect 27338 9636 27344 9648
rect 25271 9608 27344 9636
rect 25271 9605 25283 9608
rect 25225 9599 25283 9605
rect 27338 9596 27344 9608
rect 27396 9596 27402 9648
rect 28994 9596 29000 9648
rect 29052 9636 29058 9648
rect 29730 9636 29736 9648
rect 29052 9608 29736 9636
rect 29052 9596 29058 9608
rect 29730 9596 29736 9608
rect 29788 9596 29794 9648
rect 29840 9645 29868 9676
rect 30466 9664 30472 9676
rect 30524 9704 30530 9716
rect 30524 9676 31248 9704
rect 30524 9664 30530 9676
rect 29825 9639 29883 9645
rect 29825 9605 29837 9639
rect 29871 9605 29883 9639
rect 30650 9636 30656 9648
rect 29825 9599 29883 9605
rect 29932 9608 30656 9636
rect 26234 9528 26240 9580
rect 26292 9568 26298 9580
rect 26329 9571 26387 9577
rect 26329 9568 26341 9571
rect 26292 9540 26341 9568
rect 26292 9528 26298 9540
rect 26329 9537 26341 9540
rect 26375 9537 26387 9571
rect 26329 9531 26387 9537
rect 29270 9528 29276 9580
rect 29328 9568 29334 9580
rect 29932 9577 29960 9608
rect 30650 9596 30656 9608
rect 30708 9596 30714 9648
rect 29549 9571 29607 9577
rect 29549 9568 29561 9571
rect 29328 9540 29561 9568
rect 29328 9528 29334 9540
rect 29549 9537 29561 9540
rect 29595 9537 29607 9571
rect 29549 9531 29607 9537
rect 29917 9571 29975 9577
rect 29917 9537 29929 9571
rect 29963 9537 29975 9571
rect 30449 9571 30507 9577
rect 30449 9568 30461 9571
rect 29917 9531 29975 9537
rect 30116 9540 30461 9568
rect 27430 9500 27436 9512
rect 25148 9472 27436 9500
rect 25041 9463 25099 9469
rect 27430 9460 27436 9472
rect 27488 9460 27494 9512
rect 24486 9392 24492 9444
rect 24544 9432 24550 9444
rect 24765 9435 24823 9441
rect 24765 9432 24777 9435
rect 24544 9404 24777 9432
rect 24544 9392 24550 9404
rect 24765 9401 24777 9404
rect 24811 9401 24823 9435
rect 24765 9395 24823 9401
rect 25130 9392 25136 9444
rect 25188 9432 25194 9444
rect 25682 9432 25688 9444
rect 25188 9404 25688 9432
rect 25188 9392 25194 9404
rect 25682 9392 25688 9404
rect 25740 9392 25746 9444
rect 27246 9432 27252 9444
rect 26528 9404 27252 9432
rect 26528 9376 26556 9404
rect 27246 9392 27252 9404
rect 27304 9392 27310 9444
rect 27338 9392 27344 9444
rect 27396 9432 27402 9444
rect 27706 9432 27712 9444
rect 27396 9404 27712 9432
rect 27396 9392 27402 9404
rect 27706 9392 27712 9404
rect 27764 9392 27770 9444
rect 30116 9441 30144 9540
rect 30449 9537 30461 9540
rect 30495 9537 30507 9571
rect 30449 9531 30507 9537
rect 30193 9503 30251 9509
rect 30193 9469 30205 9503
rect 30239 9469 30251 9503
rect 30193 9463 30251 9469
rect 30101 9435 30159 9441
rect 30101 9401 30113 9435
rect 30147 9401 30159 9435
rect 30101 9395 30159 9401
rect 24581 9367 24639 9373
rect 24581 9364 24593 9367
rect 22879 9336 24593 9364
rect 22879 9333 22891 9336
rect 22833 9327 22891 9333
rect 24581 9333 24593 9336
rect 24627 9333 24639 9367
rect 24581 9327 24639 9333
rect 25225 9367 25283 9373
rect 25225 9333 25237 9367
rect 25271 9364 25283 9367
rect 26326 9364 26332 9376
rect 25271 9336 26332 9364
rect 25271 9333 25283 9336
rect 25225 9327 25283 9333
rect 26326 9324 26332 9336
rect 26384 9324 26390 9376
rect 26510 9324 26516 9376
rect 26568 9324 26574 9376
rect 27062 9324 27068 9376
rect 27120 9364 27126 9376
rect 28350 9364 28356 9376
rect 27120 9336 28356 9364
rect 27120 9324 27126 9336
rect 28350 9324 28356 9336
rect 28408 9324 28414 9376
rect 30208 9364 30236 9463
rect 30834 9364 30840 9376
rect 30208 9336 30840 9364
rect 30834 9324 30840 9336
rect 30892 9364 30898 9376
rect 31110 9364 31116 9376
rect 30892 9336 31116 9364
rect 30892 9324 30898 9336
rect 31110 9324 31116 9336
rect 31168 9324 31174 9376
rect 31220 9364 31248 9676
rect 31478 9664 31484 9716
rect 31536 9704 31542 9716
rect 31573 9707 31631 9713
rect 31573 9704 31585 9707
rect 31536 9676 31585 9704
rect 31536 9664 31542 9676
rect 31573 9673 31585 9676
rect 31619 9673 31631 9707
rect 31573 9667 31631 9673
rect 31846 9528 31852 9580
rect 31904 9568 31910 9580
rect 31941 9571 31999 9577
rect 31941 9568 31953 9571
rect 31904 9540 31953 9568
rect 31904 9528 31910 9540
rect 31941 9537 31953 9540
rect 31987 9537 31999 9571
rect 31941 9531 31999 9537
rect 32490 9528 32496 9580
rect 32548 9528 32554 9580
rect 32306 9392 32312 9444
rect 32364 9392 32370 9444
rect 31757 9367 31815 9373
rect 31757 9364 31769 9367
rect 31220 9336 31769 9364
rect 31757 9333 31769 9336
rect 31803 9333 31815 9367
rect 31757 9327 31815 9333
rect 1104 9274 32844 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 32844 9274
rect 1104 9200 32844 9222
rect 3605 9163 3663 9169
rect 3605 9129 3617 9163
rect 3651 9160 3663 9163
rect 4062 9160 4068 9172
rect 3651 9132 4068 9160
rect 3651 9129 3663 9132
rect 3605 9123 3663 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 5074 9120 5080 9172
rect 5132 9160 5138 9172
rect 5537 9163 5595 9169
rect 5537 9160 5549 9163
rect 5132 9132 5549 9160
rect 5132 9120 5138 9132
rect 5537 9129 5549 9132
rect 5583 9129 5595 9163
rect 5537 9123 5595 9129
rect 5810 9120 5816 9172
rect 5868 9160 5874 9172
rect 6454 9160 6460 9172
rect 5868 9132 6460 9160
rect 5868 9120 5874 9132
rect 6454 9120 6460 9132
rect 6512 9120 6518 9172
rect 6730 9120 6736 9172
rect 6788 9160 6794 9172
rect 6825 9163 6883 9169
rect 6825 9160 6837 9163
rect 6788 9132 6837 9160
rect 6788 9120 6794 9132
rect 6825 9129 6837 9132
rect 6871 9129 6883 9163
rect 6825 9123 6883 9129
rect 8941 9163 8999 9169
rect 8941 9129 8953 9163
rect 8987 9160 8999 9163
rect 9030 9160 9036 9172
rect 8987 9132 9036 9160
rect 8987 9129 8999 9132
rect 8941 9123 8999 9129
rect 9030 9120 9036 9132
rect 9088 9120 9094 9172
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9129 9183 9163
rect 9125 9123 9183 9129
rect 4893 9095 4951 9101
rect 4893 9061 4905 9095
rect 4939 9092 4951 9095
rect 5442 9092 5448 9104
rect 4939 9064 5448 9092
rect 4939 9061 4951 9064
rect 4893 9055 4951 9061
rect 5442 9052 5448 9064
rect 5500 9052 5506 9104
rect 5994 9052 6000 9104
rect 6052 9052 6058 9104
rect 6181 9095 6239 9101
rect 6181 9061 6193 9095
rect 6227 9092 6239 9095
rect 7190 9092 7196 9104
rect 6227 9064 7196 9092
rect 6227 9061 6239 9064
rect 6181 9055 6239 9061
rect 7190 9052 7196 9064
rect 7248 9052 7254 9104
rect 9140 9092 9168 9123
rect 9214 9120 9220 9172
rect 9272 9160 9278 9172
rect 11790 9160 11796 9172
rect 9272 9132 11796 9160
rect 9272 9120 9278 9132
rect 11790 9120 11796 9132
rect 11848 9120 11854 9172
rect 12529 9163 12587 9169
rect 12529 9129 12541 9163
rect 12575 9129 12587 9163
rect 12529 9123 12587 9129
rect 12713 9163 12771 9169
rect 12713 9129 12725 9163
rect 12759 9160 12771 9163
rect 13722 9160 13728 9172
rect 12759 9132 13728 9160
rect 12759 9129 12771 9132
rect 12713 9123 12771 9129
rect 10134 9092 10140 9104
rect 9140 9064 10140 9092
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 12158 9052 12164 9104
rect 12216 9092 12222 9104
rect 12216 9064 12388 9092
rect 12216 9052 12222 9064
rect 5258 9024 5264 9036
rect 4448 8996 5264 9024
rect 4448 8968 4476 8996
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 6012 9024 6040 9052
rect 5368 8996 5764 9024
rect 6012 8996 6592 9024
rect 2958 8916 2964 8968
rect 3016 8956 3022 8968
rect 3421 8959 3479 8965
rect 3421 8956 3433 8959
rect 3016 8928 3433 8956
rect 3016 8916 3022 8928
rect 3421 8925 3433 8928
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 3936 8928 3985 8956
rect 3936 8916 3942 8928
rect 3973 8925 3985 8928
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8956 4123 8959
rect 4154 8956 4160 8968
rect 4111 8928 4160 8956
rect 4111 8925 4123 8928
rect 4065 8919 4123 8925
rect 4154 8916 4160 8928
rect 4212 8916 4218 8968
rect 4430 8916 4436 8968
rect 4488 8916 4494 8968
rect 4522 8916 4528 8968
rect 4580 8956 4586 8968
rect 4706 8956 4712 8968
rect 4580 8928 4712 8956
rect 4580 8916 4586 8928
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 4798 8916 4804 8968
rect 4856 8956 4862 8968
rect 5368 8965 5396 8996
rect 5736 8968 5764 8996
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 4856 8928 4997 8956
rect 4856 8916 4862 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 5353 8959 5411 8965
rect 5353 8925 5365 8959
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 5626 8916 5632 8968
rect 5684 8916 5690 8968
rect 5718 8916 5724 8968
rect 5776 8956 5782 8968
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5776 8928 6009 8956
rect 5776 8916 5782 8928
rect 5997 8925 6009 8928
rect 6043 8956 6055 8959
rect 6086 8956 6092 8968
rect 6043 8928 6092 8956
rect 6043 8925 6055 8928
rect 5997 8919 6055 8925
rect 6086 8916 6092 8928
rect 6144 8916 6150 8968
rect 6273 8959 6331 8965
rect 6273 8925 6285 8959
rect 6319 8925 6331 8959
rect 6273 8919 6331 8925
rect 3510 8848 3516 8900
rect 3568 8888 3574 8900
rect 4249 8891 4307 8897
rect 4249 8888 4261 8891
rect 3568 8860 4261 8888
rect 3568 8848 3574 8860
rect 4249 8857 4261 8860
rect 4295 8857 4307 8891
rect 4249 8851 4307 8857
rect 4338 8848 4344 8900
rect 4396 8848 4402 8900
rect 5169 8891 5227 8897
rect 5169 8857 5181 8891
rect 5215 8857 5227 8891
rect 5169 8851 5227 8857
rect 5261 8891 5319 8897
rect 5261 8857 5273 8891
rect 5307 8888 5319 8891
rect 5644 8888 5672 8916
rect 5307 8860 5672 8888
rect 5307 8857 5319 8860
rect 5261 8851 5319 8857
rect 3789 8823 3847 8829
rect 3789 8789 3801 8823
rect 3835 8820 3847 8823
rect 4356 8820 4384 8848
rect 3835 8792 4384 8820
rect 4617 8823 4675 8829
rect 3835 8789 3847 8792
rect 3789 8783 3847 8789
rect 4617 8789 4629 8823
rect 4663 8820 4675 8823
rect 4890 8820 4896 8832
rect 4663 8792 4896 8820
rect 4663 8789 4675 8792
rect 4617 8783 4675 8789
rect 4890 8780 4896 8792
rect 4948 8780 4954 8832
rect 5184 8820 5212 8851
rect 5810 8848 5816 8900
rect 5868 8848 5874 8900
rect 5902 8848 5908 8900
rect 5960 8848 5966 8900
rect 6288 8888 6316 8919
rect 6454 8916 6460 8968
rect 6512 8916 6518 8968
rect 6564 8965 6592 8996
rect 6914 8984 6920 9036
rect 6972 9024 6978 9036
rect 9766 9024 9772 9036
rect 6972 8996 7604 9024
rect 6972 8984 6978 8996
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 6638 8916 6644 8968
rect 6696 8916 6702 8968
rect 7576 8965 7604 8996
rect 8036 8996 9772 9024
rect 8036 8965 8064 8996
rect 9766 8984 9772 8996
rect 9824 9024 9830 9036
rect 10962 9024 10968 9036
rect 9824 8996 10968 9024
rect 9824 8984 9830 8996
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 11256 8996 11468 9024
rect 7285 8959 7343 8965
rect 7285 8956 7297 8959
rect 6886 8928 7297 8956
rect 6104 8860 6316 8888
rect 5442 8820 5448 8832
rect 5184 8792 5448 8820
rect 5442 8780 5448 8792
rect 5500 8820 5506 8832
rect 5828 8820 5856 8848
rect 6104 8832 6132 8860
rect 5500 8792 5856 8820
rect 5500 8780 5506 8792
rect 6086 8780 6092 8832
rect 6144 8780 6150 8832
rect 6638 8780 6644 8832
rect 6696 8820 6702 8832
rect 6886 8820 6914 8928
rect 7285 8925 7297 8928
rect 7331 8925 7343 8959
rect 7285 8919 7343 8925
rect 7561 8959 7619 8965
rect 7561 8925 7573 8959
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 8021 8959 8079 8965
rect 8021 8925 8033 8959
rect 8067 8925 8079 8959
rect 8021 8919 8079 8925
rect 9122 8916 9128 8968
rect 9180 8916 9186 8968
rect 9214 8916 9220 8968
rect 9272 8916 9278 8968
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 9950 8956 9956 8968
rect 9548 8928 9956 8956
rect 9548 8916 9554 8928
rect 9950 8916 9956 8928
rect 10008 8956 10014 8968
rect 11256 8956 11284 8996
rect 10008 8928 11284 8956
rect 10008 8916 10014 8928
rect 11330 8916 11336 8968
rect 11388 8916 11394 8968
rect 11440 8956 11468 8996
rect 11606 8984 11612 9036
rect 11664 9024 11670 9036
rect 12250 9024 12256 9036
rect 11664 8996 12256 9024
rect 11664 8984 11670 8996
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 12360 9033 12388 9064
rect 12434 9052 12440 9104
rect 12492 9092 12498 9104
rect 12544 9092 12572 9123
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 14550 9120 14556 9172
rect 14608 9120 14614 9172
rect 15930 9160 15936 9172
rect 14660 9132 15936 9160
rect 14660 9092 14688 9132
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 16390 9120 16396 9172
rect 16448 9160 16454 9172
rect 16850 9160 16856 9172
rect 16448 9132 16856 9160
rect 16448 9120 16454 9132
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 17034 9120 17040 9172
rect 17092 9160 17098 9172
rect 17405 9163 17463 9169
rect 17405 9160 17417 9163
rect 17092 9132 17417 9160
rect 17092 9120 17098 9132
rect 17405 9129 17417 9132
rect 17451 9129 17463 9163
rect 18414 9160 18420 9172
rect 17405 9123 17463 9129
rect 17926 9132 18420 9160
rect 12492 9064 14688 9092
rect 14737 9095 14795 9101
rect 12492 9052 12498 9064
rect 14737 9061 14749 9095
rect 14783 9061 14795 9095
rect 14737 9055 14795 9061
rect 12345 9027 12403 9033
rect 12345 8993 12357 9027
rect 12391 8993 12403 9027
rect 14752 9024 14780 9055
rect 15102 9052 15108 9104
rect 15160 9092 15166 9104
rect 17926 9092 17954 9132
rect 18414 9120 18420 9132
rect 18472 9120 18478 9172
rect 18598 9120 18604 9172
rect 18656 9120 18662 9172
rect 18690 9120 18696 9172
rect 18748 9160 18754 9172
rect 18748 9132 21864 9160
rect 18748 9120 18754 9132
rect 15160 9064 17954 9092
rect 15160 9052 15166 9064
rect 18138 9052 18144 9104
rect 18196 9092 18202 9104
rect 21836 9092 21864 9132
rect 21910 9120 21916 9172
rect 21968 9120 21974 9172
rect 22002 9120 22008 9172
rect 22060 9160 22066 9172
rect 22097 9163 22155 9169
rect 22097 9160 22109 9163
rect 22060 9132 22109 9160
rect 22060 9120 22066 9132
rect 22097 9129 22109 9132
rect 22143 9160 22155 9163
rect 22370 9160 22376 9172
rect 22143 9132 22376 9160
rect 22143 9129 22155 9132
rect 22097 9123 22155 9129
rect 22370 9120 22376 9132
rect 22428 9120 22434 9172
rect 25593 9163 25651 9169
rect 25593 9129 25605 9163
rect 25639 9129 25651 9163
rect 25593 9123 25651 9129
rect 18196 9064 20484 9092
rect 21836 9064 25452 9092
rect 18196 9052 18202 9064
rect 12345 8987 12403 8993
rect 12452 8996 14688 9024
rect 14752 8996 18460 9024
rect 12452 8956 12480 8996
rect 11440 8928 12480 8956
rect 12526 8916 12532 8968
rect 12584 8916 12590 8968
rect 12894 8916 12900 8968
rect 12952 8956 12958 8968
rect 13354 8956 13360 8968
rect 12952 8928 13360 8956
rect 12952 8916 12958 8928
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 14090 8916 14096 8968
rect 14148 8916 14154 8968
rect 14366 8916 14372 8968
rect 14424 8916 14430 8968
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8925 14611 8959
rect 14660 8956 14688 8996
rect 16666 8956 16672 8968
rect 14660 8928 16672 8956
rect 14553 8919 14611 8925
rect 8202 8848 8208 8900
rect 8260 8888 8266 8900
rect 9030 8888 9036 8900
rect 8260 8860 9036 8888
rect 8260 8848 8266 8860
rect 9030 8848 9036 8860
rect 9088 8848 9094 8900
rect 9398 8848 9404 8900
rect 9456 8848 9462 8900
rect 9674 8848 9680 8900
rect 9732 8888 9738 8900
rect 10962 8888 10968 8900
rect 9732 8860 10968 8888
rect 9732 8848 9738 8860
rect 10962 8848 10968 8860
rect 11020 8848 11026 8900
rect 11422 8848 11428 8900
rect 11480 8888 11486 8900
rect 12253 8891 12311 8897
rect 12253 8888 12265 8891
rect 11480 8860 12265 8888
rect 11480 8848 11486 8860
rect 12253 8857 12265 8860
rect 12299 8857 12311 8891
rect 12253 8851 12311 8857
rect 6696 8792 6914 8820
rect 6696 8780 6702 8792
rect 7006 8780 7012 8832
rect 7064 8820 7070 8832
rect 7469 8823 7527 8829
rect 7469 8820 7481 8823
rect 7064 8792 7481 8820
rect 7064 8780 7070 8792
rect 7469 8789 7481 8792
rect 7515 8820 7527 8823
rect 7650 8820 7656 8832
rect 7515 8792 7656 8820
rect 7515 8789 7527 8792
rect 7469 8783 7527 8789
rect 7650 8780 7656 8792
rect 7708 8780 7714 8832
rect 7742 8780 7748 8832
rect 7800 8780 7806 8832
rect 7834 8780 7840 8832
rect 7892 8820 7898 8832
rect 9858 8820 9864 8832
rect 7892 8792 9864 8820
rect 7892 8780 7898 8792
rect 9858 8780 9864 8792
rect 9916 8820 9922 8832
rect 11146 8820 11152 8832
rect 9916 8792 11152 8820
rect 9916 8780 9922 8792
rect 11146 8780 11152 8792
rect 11204 8780 11210 8832
rect 12268 8820 12296 8851
rect 12342 8848 12348 8900
rect 12400 8888 12406 8900
rect 14568 8888 14596 8919
rect 16666 8916 16672 8928
rect 16724 8916 16730 8968
rect 16850 8916 16856 8968
rect 16908 8956 16914 8968
rect 18432 8965 18460 8996
rect 18506 8984 18512 9036
rect 18564 8984 18570 9036
rect 20456 9024 20484 9064
rect 23382 9024 23388 9036
rect 18616 8996 19334 9024
rect 20456 8996 23388 9024
rect 17129 8959 17187 8965
rect 17129 8956 17141 8959
rect 16908 8928 17141 8956
rect 16908 8916 16914 8928
rect 17129 8925 17141 8928
rect 17175 8925 17187 8959
rect 17129 8919 17187 8925
rect 17589 8959 17647 8965
rect 17589 8925 17601 8959
rect 17635 8956 17647 8959
rect 18417 8959 18475 8965
rect 17635 8928 18368 8956
rect 17635 8925 17647 8928
rect 17589 8919 17647 8925
rect 17218 8888 17224 8900
rect 12400 8860 14596 8888
rect 14660 8860 17224 8888
rect 12400 8848 12406 8860
rect 12894 8820 12900 8832
rect 12268 8792 12900 8820
rect 12894 8780 12900 8792
rect 12952 8780 12958 8832
rect 13170 8780 13176 8832
rect 13228 8820 13234 8832
rect 14660 8820 14688 8860
rect 17218 8848 17224 8860
rect 17276 8848 17282 8900
rect 13228 8792 14688 8820
rect 13228 8780 13234 8792
rect 14826 8780 14832 8832
rect 14884 8820 14890 8832
rect 16390 8820 16396 8832
rect 14884 8792 16396 8820
rect 14884 8780 14890 8792
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 16850 8780 16856 8832
rect 16908 8820 16914 8832
rect 16945 8823 17003 8829
rect 16945 8820 16957 8823
rect 16908 8792 16957 8820
rect 16908 8780 16914 8792
rect 16945 8789 16957 8792
rect 16991 8789 17003 8823
rect 16945 8783 17003 8789
rect 17313 8823 17371 8829
rect 17313 8789 17325 8823
rect 17359 8820 17371 8823
rect 17604 8820 17632 8919
rect 17770 8848 17776 8900
rect 17828 8848 17834 8900
rect 18340 8888 18368 8928
rect 18417 8925 18429 8959
rect 18463 8925 18475 8959
rect 18417 8919 18475 8925
rect 18616 8888 18644 8996
rect 18693 8959 18751 8965
rect 18693 8925 18705 8959
rect 18739 8925 18751 8959
rect 19306 8956 19334 8996
rect 23382 8984 23388 8996
rect 23440 8984 23446 9036
rect 25424 9024 25452 9064
rect 25608 9024 25636 9123
rect 25682 9120 25688 9172
rect 25740 9160 25746 9172
rect 25961 9163 26019 9169
rect 25961 9160 25973 9163
rect 25740 9132 25973 9160
rect 25740 9120 25746 9132
rect 25961 9129 25973 9132
rect 26007 9160 26019 9163
rect 26050 9160 26056 9172
rect 26007 9132 26056 9160
rect 26007 9129 26019 9132
rect 25961 9123 26019 9129
rect 26050 9120 26056 9132
rect 26108 9120 26114 9172
rect 26145 9163 26203 9169
rect 26145 9129 26157 9163
rect 26191 9129 26203 9163
rect 26145 9123 26203 9129
rect 25866 9052 25872 9104
rect 25924 9092 25930 9104
rect 26160 9092 26188 9123
rect 26602 9120 26608 9172
rect 26660 9120 26666 9172
rect 26973 9163 27031 9169
rect 26973 9129 26985 9163
rect 27019 9160 27031 9163
rect 27614 9160 27620 9172
rect 27019 9132 27620 9160
rect 27019 9129 27031 9132
rect 26973 9123 27031 9129
rect 26510 9092 26516 9104
rect 25924 9064 26188 9092
rect 26344 9064 26516 9092
rect 25924 9052 25930 9064
rect 26142 9024 26148 9036
rect 25424 8996 26148 9024
rect 26142 8984 26148 8996
rect 26200 8984 26206 9036
rect 26344 9033 26372 9064
rect 26510 9052 26516 9064
rect 26568 9052 26574 9104
rect 26988 9092 27016 9123
rect 27614 9120 27620 9132
rect 27672 9120 27678 9172
rect 27709 9163 27767 9169
rect 27709 9129 27721 9163
rect 27755 9129 27767 9163
rect 27709 9123 27767 9129
rect 28077 9163 28135 9169
rect 28077 9129 28089 9163
rect 28123 9160 28135 9163
rect 28166 9160 28172 9172
rect 28123 9132 28172 9160
rect 28123 9129 28135 9132
rect 28077 9123 28135 9129
rect 26620 9064 27016 9092
rect 26329 9027 26387 9033
rect 26329 8993 26341 9027
rect 26375 8993 26387 9027
rect 26620 9024 26648 9064
rect 27246 9052 27252 9104
rect 27304 9092 27310 9104
rect 27724 9092 27752 9123
rect 28166 9120 28172 9132
rect 28224 9120 28230 9172
rect 29270 9120 29276 9172
rect 29328 9120 29334 9172
rect 32490 9120 32496 9172
rect 32548 9120 32554 9172
rect 27304 9064 27752 9092
rect 27304 9052 27310 9064
rect 26329 8987 26387 8993
rect 26429 8996 26648 9024
rect 19306 8928 21956 8956
rect 18693 8919 18751 8925
rect 18340 8860 18644 8888
rect 18708 8888 18736 8919
rect 21928 8888 21956 8928
rect 22002 8916 22008 8968
rect 22060 8956 22066 8968
rect 22097 8959 22155 8965
rect 22097 8956 22109 8959
rect 22060 8928 22109 8956
rect 22060 8916 22066 8928
rect 22097 8925 22109 8928
rect 22143 8925 22155 8959
rect 22097 8919 22155 8925
rect 22189 8959 22247 8965
rect 22189 8925 22201 8959
rect 22235 8956 22247 8959
rect 22278 8956 22284 8968
rect 22235 8928 22284 8956
rect 22235 8925 22247 8928
rect 22189 8919 22247 8925
rect 22278 8916 22284 8928
rect 22336 8916 22342 8968
rect 22384 8959 22442 8965
rect 22384 8925 22396 8959
rect 22430 8956 22442 8959
rect 22554 8956 22560 8968
rect 22430 8928 22560 8956
rect 22430 8925 22442 8928
rect 22384 8919 22442 8925
rect 22554 8916 22560 8928
rect 22612 8916 22618 8968
rect 25501 8959 25559 8965
rect 25501 8956 25513 8959
rect 24136 8928 25513 8956
rect 24136 8888 24164 8928
rect 25501 8925 25513 8928
rect 25547 8956 25559 8959
rect 25590 8956 25596 8968
rect 25547 8928 25596 8956
rect 25547 8925 25559 8928
rect 25501 8919 25559 8925
rect 25590 8916 25596 8928
rect 25648 8916 25654 8968
rect 25682 8916 25688 8968
rect 25740 8916 25746 8968
rect 25774 8916 25780 8968
rect 25832 8916 25838 8968
rect 26429 8965 26457 8996
rect 26786 8984 26792 9036
rect 26844 9024 26850 9036
rect 26844 8996 27016 9024
rect 26844 8984 26850 8996
rect 26414 8959 26472 8965
rect 26414 8925 26426 8959
rect 26460 8925 26472 8959
rect 26414 8919 26472 8925
rect 26602 8916 26608 8968
rect 26660 8956 26666 8968
rect 26988 8965 27016 8996
rect 27522 8984 27528 9036
rect 27580 9024 27586 9036
rect 27709 9027 27767 9033
rect 27709 9024 27721 9027
rect 27580 8996 27721 9024
rect 27580 8984 27586 8996
rect 27709 8993 27721 8996
rect 27755 8993 27767 9027
rect 27709 8987 27767 8993
rect 27798 8984 27804 9036
rect 27856 9024 27862 9036
rect 28810 9024 28816 9036
rect 27856 8996 28816 9024
rect 27856 8984 27862 8996
rect 27908 8965 27936 8996
rect 28810 8984 28816 8996
rect 28868 8984 28874 9036
rect 26881 8959 26939 8965
rect 26881 8956 26893 8959
rect 26660 8928 26893 8956
rect 26660 8916 26666 8928
rect 26881 8925 26893 8928
rect 26927 8925 26939 8959
rect 26881 8919 26939 8925
rect 26973 8959 27031 8965
rect 26973 8925 26985 8959
rect 27019 8925 27031 8959
rect 27893 8959 27951 8965
rect 26973 8919 27031 8925
rect 27080 8928 27752 8956
rect 18708 8860 20300 8888
rect 21928 8860 24164 8888
rect 17359 8792 17632 8820
rect 17359 8789 17371 8792
rect 17313 8783 17371 8789
rect 18230 8780 18236 8832
rect 18288 8820 18294 8832
rect 18877 8823 18935 8829
rect 18877 8820 18889 8823
rect 18288 8792 18889 8820
rect 18288 8780 18294 8792
rect 18877 8789 18889 8792
rect 18923 8789 18935 8823
rect 20272 8820 20300 8860
rect 24578 8848 24584 8900
rect 24636 8888 24642 8900
rect 24636 8860 26096 8888
rect 24636 8848 24642 8860
rect 24946 8820 24952 8832
rect 20272 8792 24952 8820
rect 18877 8783 18935 8789
rect 24946 8780 24952 8792
rect 25004 8820 25010 8832
rect 25317 8823 25375 8829
rect 25317 8820 25329 8823
rect 25004 8792 25329 8820
rect 25004 8780 25010 8792
rect 25317 8789 25329 8792
rect 25363 8789 25375 8823
rect 26068 8820 26096 8860
rect 26142 8848 26148 8900
rect 26200 8888 26206 8900
rect 26697 8891 26755 8897
rect 26697 8888 26709 8891
rect 26200 8860 26709 8888
rect 26200 8848 26206 8860
rect 26697 8857 26709 8860
rect 26743 8857 26755 8891
rect 26697 8851 26755 8857
rect 27080 8820 27108 8928
rect 27338 8848 27344 8900
rect 27396 8888 27402 8900
rect 27617 8891 27675 8897
rect 27617 8888 27629 8891
rect 27396 8860 27629 8888
rect 27396 8848 27402 8860
rect 27617 8857 27629 8860
rect 27663 8857 27675 8891
rect 27724 8888 27752 8928
rect 27893 8925 27905 8959
rect 27939 8925 27951 8959
rect 27893 8919 27951 8925
rect 28350 8916 28356 8968
rect 28408 8916 28414 8968
rect 29086 8916 29092 8968
rect 29144 8916 29150 8968
rect 31110 8916 31116 8968
rect 31168 8916 31174 8968
rect 28905 8891 28963 8897
rect 28905 8888 28917 8891
rect 27724 8860 28917 8888
rect 27617 8851 27675 8857
rect 28905 8857 28917 8860
rect 28951 8857 28963 8891
rect 28905 8851 28963 8857
rect 30742 8848 30748 8900
rect 30800 8888 30806 8900
rect 31358 8891 31416 8897
rect 31358 8888 31370 8891
rect 30800 8860 31370 8888
rect 30800 8848 30806 8860
rect 31358 8857 31370 8860
rect 31404 8857 31416 8891
rect 31358 8851 31416 8857
rect 26068 8792 27108 8820
rect 25317 8783 25375 8789
rect 27154 8780 27160 8832
rect 27212 8780 27218 8832
rect 27522 8780 27528 8832
rect 27580 8820 27586 8832
rect 28169 8823 28227 8829
rect 28169 8820 28181 8823
rect 27580 8792 28181 8820
rect 27580 8780 27586 8792
rect 28169 8789 28181 8792
rect 28215 8789 28227 8823
rect 28169 8783 28227 8789
rect 1104 8730 32844 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 32844 8730
rect 1104 8656 32844 8678
rect 4065 8619 4123 8625
rect 4065 8585 4077 8619
rect 4111 8585 4123 8619
rect 4065 8579 4123 8585
rect 4080 8548 4108 8579
rect 4430 8576 4436 8628
rect 4488 8616 4494 8628
rect 4617 8619 4675 8625
rect 4617 8616 4629 8619
rect 4488 8588 4629 8616
rect 4488 8576 4494 8588
rect 4617 8585 4629 8588
rect 4663 8585 4675 8619
rect 4617 8579 4675 8585
rect 4798 8576 4804 8628
rect 4856 8616 4862 8628
rect 5902 8616 5908 8628
rect 4856 8588 5908 8616
rect 4856 8576 4862 8588
rect 5902 8576 5908 8588
rect 5960 8616 5966 8628
rect 6270 8616 6276 8628
rect 5960 8588 6276 8616
rect 5960 8576 5966 8588
rect 6270 8576 6276 8588
rect 6328 8616 6334 8628
rect 6822 8616 6828 8628
rect 6328 8588 6828 8616
rect 6328 8576 6334 8588
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 7466 8576 7472 8628
rect 7524 8616 7530 8628
rect 7524 8588 8064 8616
rect 7524 8576 7530 8588
rect 4154 8548 4160 8560
rect 4080 8520 4160 8548
rect 4154 8508 4160 8520
rect 4212 8548 4218 8560
rect 4212 8520 5396 8548
rect 4212 8508 4218 8520
rect 3142 8440 3148 8492
rect 3200 8480 3206 8492
rect 4249 8483 4307 8489
rect 4249 8480 4261 8483
rect 3200 8452 4261 8480
rect 3200 8440 3206 8452
rect 4249 8449 4261 8452
rect 4295 8449 4307 8483
rect 4249 8443 4307 8449
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 4614 8480 4620 8492
rect 4479 8452 4620 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 4264 8412 4292 8443
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 5258 8440 5264 8492
rect 5316 8440 5322 8492
rect 4982 8412 4988 8424
rect 4264 8384 4988 8412
rect 4982 8372 4988 8384
rect 5040 8372 5046 8424
rect 5368 8412 5396 8520
rect 5442 8508 5448 8560
rect 5500 8508 5506 8560
rect 7374 8508 7380 8560
rect 7432 8508 7438 8560
rect 8036 8548 8064 8588
rect 8754 8576 8760 8628
rect 8812 8576 8818 8628
rect 9214 8576 9220 8628
rect 9272 8616 9278 8628
rect 9401 8619 9459 8625
rect 9401 8616 9413 8619
rect 9272 8588 9413 8616
rect 9272 8576 9278 8588
rect 9401 8585 9413 8588
rect 9447 8616 9459 8619
rect 9447 8588 10640 8616
rect 9447 8585 9459 8588
rect 9401 8579 9459 8585
rect 8772 8548 8800 8576
rect 8036 8520 8708 8548
rect 8772 8520 9260 8548
rect 5534 8440 5540 8492
rect 5592 8440 5598 8492
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8480 5687 8483
rect 5718 8480 5724 8492
rect 5675 8452 5724 8480
rect 5675 8449 5687 8452
rect 5629 8443 5687 8449
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 5994 8480 6000 8492
rect 5951 8452 6000 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 7193 8483 7251 8489
rect 7193 8449 7205 8483
rect 7239 8449 7251 8483
rect 7193 8443 7251 8449
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8449 7527 8483
rect 7469 8443 7527 8449
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8480 7619 8483
rect 7834 8480 7840 8492
rect 7607 8452 7840 8480
rect 7607 8449 7619 8452
rect 7561 8443 7619 8449
rect 7208 8412 7236 8443
rect 5368 8384 7236 8412
rect 4338 8304 4344 8356
rect 4396 8344 4402 8356
rect 4706 8344 4712 8356
rect 4396 8316 4712 8344
rect 4396 8304 4402 8316
rect 4706 8304 4712 8316
rect 4764 8344 4770 8356
rect 7484 8344 7512 8443
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 8036 8489 8064 8520
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 8202 8440 8208 8492
rect 8260 8480 8266 8492
rect 8297 8483 8355 8489
rect 8573 8484 8631 8489
rect 8297 8480 8309 8483
rect 8260 8452 8309 8480
rect 8260 8440 8266 8452
rect 8297 8449 8309 8452
rect 8343 8449 8355 8483
rect 8496 8483 8631 8484
rect 8496 8480 8585 8483
rect 8297 8443 8355 8449
rect 8404 8456 8585 8480
rect 8404 8452 8524 8456
rect 7650 8372 7656 8424
rect 7708 8412 7714 8424
rect 8220 8412 8248 8440
rect 8404 8424 8432 8452
rect 8573 8449 8585 8456
rect 8619 8449 8631 8483
rect 8680 8484 8708 8520
rect 8757 8484 8815 8489
rect 8680 8483 8815 8484
rect 8680 8456 8769 8483
rect 8573 8443 8631 8449
rect 8757 8449 8769 8456
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 8846 8440 8852 8492
rect 8904 8440 8910 8492
rect 8941 8484 8999 8489
rect 9030 8484 9036 8492
rect 8941 8483 9036 8484
rect 8941 8449 8953 8483
rect 8987 8456 9036 8483
rect 8987 8449 8999 8456
rect 8941 8443 8999 8449
rect 9030 8440 9036 8456
rect 9088 8440 9094 8492
rect 9232 8489 9260 8520
rect 9306 8508 9312 8560
rect 9364 8548 9370 8560
rect 9364 8520 9628 8548
rect 9364 8508 9370 8520
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 9600 8480 9628 8520
rect 9674 8508 9680 8560
rect 9732 8508 9738 8560
rect 10244 8548 10272 8588
rect 10413 8551 10471 8557
rect 10413 8548 10425 8551
rect 10244 8520 10425 8548
rect 10413 8517 10425 8520
rect 10459 8517 10471 8551
rect 10612 8548 10640 8588
rect 11330 8576 11336 8628
rect 11388 8576 11394 8628
rect 11698 8576 11704 8628
rect 11756 8576 11762 8628
rect 11882 8576 11888 8628
rect 11940 8576 11946 8628
rect 12529 8619 12587 8625
rect 12529 8585 12541 8619
rect 12575 8616 12587 8619
rect 13722 8616 13728 8628
rect 12575 8588 13728 8616
rect 12575 8585 12587 8588
rect 12529 8579 12587 8585
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 14001 8619 14059 8625
rect 14001 8585 14013 8619
rect 14047 8616 14059 8619
rect 14366 8616 14372 8628
rect 14047 8588 14372 8616
rect 14047 8585 14059 8588
rect 14001 8579 14059 8585
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 15473 8619 15531 8625
rect 15473 8616 15485 8619
rect 14936 8588 15485 8616
rect 10612 8520 10824 8548
rect 10413 8511 10471 8517
rect 9769 8483 9827 8489
rect 9769 8480 9781 8483
rect 9600 8452 9781 8480
rect 9769 8449 9781 8452
rect 9815 8449 9827 8483
rect 9769 8443 9827 8449
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 10183 8486 10241 8489
rect 10060 8483 10272 8486
rect 10060 8480 10195 8483
rect 9968 8458 10195 8480
rect 9968 8452 10088 8458
rect 9968 8424 9996 8452
rect 10183 8449 10195 8458
rect 10229 8452 10272 8483
rect 10229 8449 10241 8452
rect 10183 8443 10241 8449
rect 10318 8440 10324 8492
rect 10376 8440 10382 8492
rect 10796 8489 10824 8520
rect 10962 8508 10968 8560
rect 11020 8508 11026 8560
rect 11054 8508 11060 8560
rect 11112 8508 11118 8560
rect 11716 8548 11744 8576
rect 14936 8557 14964 8588
rect 15473 8585 15485 8588
rect 15519 8585 15531 8619
rect 15473 8579 15531 8585
rect 16853 8619 16911 8625
rect 16853 8585 16865 8619
rect 16899 8616 16911 8619
rect 16942 8616 16948 8628
rect 16899 8588 16948 8616
rect 16899 8585 16911 8588
rect 16853 8579 16911 8585
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 17313 8619 17371 8625
rect 17313 8585 17325 8619
rect 17359 8585 17371 8619
rect 17313 8579 17371 8585
rect 11532 8520 11744 8548
rect 12069 8551 12127 8557
rect 10505 8483 10563 8489
rect 10505 8464 10517 8483
rect 10428 8449 10517 8464
rect 10551 8449 10563 8483
rect 10428 8443 10563 8449
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 10428 8436 10548 8443
rect 11146 8440 11152 8492
rect 11204 8440 11210 8492
rect 11532 8489 11560 8520
rect 12069 8517 12081 8551
rect 12115 8548 12127 8551
rect 14921 8551 14979 8557
rect 12115 8520 13676 8548
rect 12115 8517 12127 8520
rect 12069 8511 12127 8517
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 11698 8440 11704 8492
rect 11756 8440 11762 8492
rect 12250 8440 12256 8492
rect 12308 8440 12314 8492
rect 12345 8483 12403 8489
rect 12345 8449 12357 8483
rect 12391 8480 12403 8483
rect 12526 8480 12532 8492
rect 12391 8452 12532 8480
rect 12391 8449 12403 8452
rect 12345 8443 12403 8449
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 12713 8483 12771 8489
rect 12713 8449 12725 8483
rect 12759 8480 12771 8483
rect 12805 8483 12863 8489
rect 12805 8480 12817 8483
rect 12759 8452 12817 8480
rect 12759 8449 12771 8452
rect 12713 8443 12771 8449
rect 12805 8449 12817 8452
rect 12851 8480 12863 8483
rect 12894 8480 12900 8492
rect 12851 8452 12900 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 12986 8440 12992 8492
rect 13044 8480 13050 8492
rect 13170 8480 13176 8492
rect 13044 8452 13176 8480
rect 13044 8440 13050 8452
rect 13170 8440 13176 8452
rect 13228 8440 13234 8492
rect 13538 8440 13544 8492
rect 13596 8440 13602 8492
rect 7708 8384 8248 8412
rect 7708 8372 7714 8384
rect 8386 8372 8392 8424
rect 8444 8372 8450 8424
rect 9582 8412 9588 8424
rect 9048 8384 9588 8412
rect 4764 8316 7512 8344
rect 7745 8347 7803 8353
rect 4764 8304 4770 8316
rect 7745 8313 7757 8347
rect 7791 8344 7803 8347
rect 8018 8344 8024 8356
rect 7791 8316 8024 8344
rect 7791 8313 7803 8316
rect 7745 8307 7803 8313
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 8846 8304 8852 8356
rect 8904 8344 8910 8356
rect 9048 8344 9076 8384
rect 9582 8372 9588 8384
rect 9640 8412 9646 8424
rect 9950 8412 9956 8424
rect 9640 8384 9956 8412
rect 9640 8372 9646 8384
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 8904 8316 9076 8344
rect 9125 8347 9183 8353
rect 8904 8304 8910 8316
rect 9125 8313 9137 8347
rect 9171 8344 9183 8347
rect 9398 8344 9404 8356
rect 9171 8316 9404 8344
rect 9171 8313 9183 8316
rect 9125 8307 9183 8313
rect 9398 8304 9404 8316
rect 9456 8304 9462 8356
rect 10428 8344 10456 8436
rect 10870 8372 10876 8424
rect 10928 8412 10934 8424
rect 13262 8412 13268 8424
rect 10928 8384 13268 8412
rect 10928 8372 10934 8384
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 10502 8344 10508 8356
rect 10428 8316 10508 8344
rect 10502 8304 10508 8316
rect 10560 8304 10566 8356
rect 10689 8347 10747 8353
rect 10689 8313 10701 8347
rect 10735 8344 10747 8347
rect 11422 8344 11428 8356
rect 10735 8316 11428 8344
rect 10735 8313 10747 8316
rect 10689 8307 10747 8313
rect 11422 8304 11428 8316
rect 11480 8304 11486 8356
rect 12342 8304 12348 8356
rect 12400 8344 12406 8356
rect 12618 8344 12624 8356
rect 12400 8316 12624 8344
rect 12400 8304 12406 8316
rect 12618 8304 12624 8316
rect 12676 8304 12682 8356
rect 12989 8347 13047 8353
rect 12728 8316 12940 8344
rect 5810 8236 5816 8288
rect 5868 8236 5874 8288
rect 5902 8236 5908 8288
rect 5960 8276 5966 8288
rect 6089 8279 6147 8285
rect 6089 8276 6101 8279
rect 5960 8248 6101 8276
rect 5960 8236 5966 8248
rect 6089 8245 6101 8248
rect 6135 8245 6147 8279
rect 6089 8239 6147 8245
rect 8110 8236 8116 8288
rect 8168 8276 8174 8288
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 8168 8248 8217 8276
rect 8168 8236 8174 8248
rect 8205 8245 8217 8248
rect 8251 8245 8263 8279
rect 8205 8239 8263 8245
rect 8478 8236 8484 8288
rect 8536 8236 8542 8288
rect 10045 8279 10103 8285
rect 10045 8245 10057 8279
rect 10091 8276 10103 8279
rect 10870 8276 10876 8288
rect 10091 8248 10876 8276
rect 10091 8245 10103 8248
rect 10045 8239 10103 8245
rect 10870 8236 10876 8248
rect 10928 8236 10934 8288
rect 11514 8236 11520 8288
rect 11572 8236 11578 8288
rect 12158 8236 12164 8288
rect 12216 8236 12222 8288
rect 12250 8236 12256 8288
rect 12308 8276 12314 8288
rect 12728 8276 12756 8316
rect 12308 8248 12756 8276
rect 12912 8276 12940 8316
rect 12989 8313 13001 8347
rect 13035 8344 13047 8347
rect 13648 8344 13676 8520
rect 14921 8517 14933 8551
rect 14967 8517 14979 8551
rect 17328 8548 17356 8579
rect 17402 8576 17408 8628
rect 17460 8616 17466 8628
rect 19794 8616 19800 8628
rect 17460 8588 19800 8616
rect 17460 8576 17466 8588
rect 19794 8576 19800 8588
rect 19852 8576 19858 8628
rect 19886 8576 19892 8628
rect 19944 8616 19950 8628
rect 20073 8619 20131 8625
rect 20073 8616 20085 8619
rect 19944 8588 20085 8616
rect 19944 8576 19950 8588
rect 20073 8585 20085 8588
rect 20119 8585 20131 8619
rect 20073 8579 20131 8585
rect 20717 8619 20775 8625
rect 20717 8585 20729 8619
rect 20763 8616 20775 8619
rect 20763 8588 24256 8616
rect 20763 8585 20775 8588
rect 20717 8579 20775 8585
rect 19426 8548 19432 8560
rect 14921 8511 14979 8517
rect 15028 8520 16988 8548
rect 17328 8520 19432 8548
rect 13817 8483 13875 8489
rect 13817 8449 13829 8483
rect 13863 8480 13875 8483
rect 13906 8480 13912 8492
rect 13863 8452 13912 8480
rect 13863 8449 13875 8452
rect 13817 8443 13875 8449
rect 13906 8440 13912 8452
rect 13964 8440 13970 8492
rect 14090 8440 14096 8492
rect 14148 8480 14154 8492
rect 15028 8480 15056 8520
rect 14148 8452 15056 8480
rect 14148 8440 14154 8452
rect 15102 8440 15108 8492
rect 15160 8440 15166 8492
rect 15194 8440 15200 8492
rect 15252 8440 15258 8492
rect 15562 8440 15568 8492
rect 15620 8480 15626 8492
rect 15657 8483 15715 8489
rect 15657 8480 15669 8483
rect 15620 8452 15669 8480
rect 15620 8440 15626 8452
rect 15657 8449 15669 8452
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 15746 8440 15752 8492
rect 15804 8440 15810 8492
rect 15838 8440 15844 8492
rect 15896 8480 15902 8492
rect 15933 8483 15991 8489
rect 15933 8480 15945 8483
rect 15896 8452 15945 8480
rect 15896 8440 15902 8452
rect 15933 8449 15945 8452
rect 15979 8449 15991 8483
rect 15933 8443 15991 8449
rect 16666 8440 16672 8492
rect 16724 8440 16730 8492
rect 16960 8489 16988 8520
rect 19426 8508 19432 8520
rect 19484 8508 19490 8560
rect 20898 8548 20904 8560
rect 20456 8520 20904 8548
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 17126 8440 17132 8492
rect 17184 8480 17190 8492
rect 17497 8483 17555 8489
rect 17497 8480 17509 8483
rect 17184 8452 17509 8480
rect 17184 8440 17190 8452
rect 17497 8449 17509 8452
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 17678 8440 17684 8492
rect 17736 8440 17742 8492
rect 19794 8480 19800 8492
rect 19306 8452 19800 8480
rect 13722 8372 13728 8424
rect 13780 8372 13786 8424
rect 14752 8384 15516 8412
rect 14752 8344 14780 8384
rect 13035 8316 14780 8344
rect 13035 8313 13047 8316
rect 12989 8307 13047 8313
rect 15378 8304 15384 8356
rect 15436 8304 15442 8356
rect 15488 8344 15516 8384
rect 16574 8372 16580 8424
rect 16632 8412 16638 8424
rect 17037 8415 17095 8421
rect 17037 8412 17049 8415
rect 16632 8384 17049 8412
rect 16632 8372 16638 8384
rect 17037 8381 17049 8384
rect 17083 8381 17095 8415
rect 19306 8412 19334 8452
rect 19794 8440 19800 8452
rect 19852 8440 19858 8492
rect 20282 8483 20340 8489
rect 20282 8449 20294 8483
rect 20328 8480 20340 8483
rect 20456 8480 20484 8520
rect 20898 8508 20904 8520
rect 20956 8508 20962 8560
rect 23474 8508 23480 8560
rect 23532 8508 23538 8560
rect 23566 8508 23572 8560
rect 23624 8548 23630 8560
rect 24228 8557 24256 8588
rect 24670 8576 24676 8628
rect 24728 8576 24734 8628
rect 24762 8576 24768 8628
rect 24820 8616 24826 8628
rect 29546 8616 29552 8628
rect 24820 8588 29552 8616
rect 24820 8576 24826 8588
rect 29546 8576 29552 8588
rect 29604 8576 29610 8628
rect 24213 8551 24271 8557
rect 23624 8520 23980 8548
rect 23624 8508 23630 8520
rect 20328 8452 20484 8480
rect 20533 8483 20591 8489
rect 20328 8449 20340 8452
rect 20282 8443 20340 8449
rect 20533 8449 20545 8483
rect 20579 8480 20591 8483
rect 20990 8480 20996 8492
rect 20579 8452 20996 8480
rect 20579 8449 20591 8452
rect 20533 8443 20591 8449
rect 20990 8440 20996 8452
rect 21048 8440 21054 8492
rect 23492 8480 23520 8508
rect 23952 8492 23980 8520
rect 24213 8517 24225 8551
rect 24259 8517 24271 8551
rect 24213 8511 24271 8517
rect 27614 8508 27620 8560
rect 27672 8548 27678 8560
rect 27672 8520 30144 8548
rect 27672 8508 27678 8520
rect 23661 8483 23719 8489
rect 23661 8480 23673 8483
rect 23492 8452 23673 8480
rect 23661 8449 23673 8452
rect 23707 8449 23719 8483
rect 23661 8443 23719 8449
rect 23934 8440 23940 8492
rect 23992 8440 23998 8492
rect 24489 8483 24547 8489
rect 24044 8452 24440 8480
rect 17037 8375 17095 8381
rect 17144 8384 19334 8412
rect 17144 8344 17172 8384
rect 20162 8372 20168 8424
rect 20220 8412 20226 8424
rect 20441 8415 20499 8421
rect 20441 8412 20453 8415
rect 20220 8384 20453 8412
rect 20220 8372 20226 8384
rect 20441 8381 20453 8384
rect 20487 8381 20499 8415
rect 20441 8375 20499 8381
rect 20898 8372 20904 8424
rect 20956 8412 20962 8424
rect 23753 8415 23811 8421
rect 23753 8412 23765 8415
rect 20956 8384 23765 8412
rect 20956 8372 20962 8384
rect 23753 8381 23765 8384
rect 23799 8381 23811 8415
rect 23753 8375 23811 8381
rect 15488 8316 17172 8344
rect 17865 8347 17923 8353
rect 17865 8313 17877 8347
rect 17911 8344 17923 8347
rect 24044 8344 24072 8452
rect 24305 8415 24363 8421
rect 24305 8381 24317 8415
rect 24351 8381 24363 8415
rect 24412 8412 24440 8452
rect 24489 8449 24501 8483
rect 24535 8480 24547 8483
rect 24762 8480 24768 8492
rect 24535 8452 24768 8480
rect 24535 8449 24547 8452
rect 24489 8443 24547 8449
rect 24762 8440 24768 8452
rect 24820 8440 24826 8492
rect 29733 8483 29791 8489
rect 29733 8449 29745 8483
rect 29779 8480 29791 8483
rect 30006 8480 30012 8492
rect 29779 8452 30012 8480
rect 29779 8449 29791 8452
rect 29733 8443 29791 8449
rect 30006 8440 30012 8452
rect 30064 8440 30070 8492
rect 30116 8480 30144 8520
rect 30558 8508 30564 8560
rect 30616 8548 30622 8560
rect 30837 8551 30895 8557
rect 30837 8548 30849 8551
rect 30616 8520 30849 8548
rect 30616 8508 30622 8520
rect 30837 8517 30849 8520
rect 30883 8517 30895 8551
rect 30837 8511 30895 8517
rect 30929 8551 30987 8557
rect 30929 8517 30941 8551
rect 30975 8548 30987 8551
rect 31846 8548 31852 8560
rect 30975 8520 31852 8548
rect 30975 8517 30987 8520
rect 30929 8511 30987 8517
rect 31846 8508 31852 8520
rect 31904 8508 31910 8560
rect 30653 8483 30711 8489
rect 30653 8480 30665 8483
rect 30116 8452 30665 8480
rect 30653 8449 30665 8452
rect 30699 8449 30711 8483
rect 30653 8443 30711 8449
rect 31021 8483 31079 8489
rect 31021 8449 31033 8483
rect 31067 8480 31079 8483
rect 31297 8483 31355 8489
rect 31297 8480 31309 8483
rect 31067 8452 31309 8480
rect 31067 8449 31079 8452
rect 31021 8443 31079 8449
rect 31297 8449 31309 8452
rect 31343 8449 31355 8483
rect 31297 8443 31355 8449
rect 31941 8483 31999 8489
rect 31941 8449 31953 8483
rect 31987 8480 31999 8483
rect 32214 8480 32220 8492
rect 31987 8452 32220 8480
rect 31987 8449 31999 8452
rect 31941 8443 31999 8449
rect 32214 8440 32220 8452
rect 32272 8440 32278 8492
rect 29825 8415 29883 8421
rect 29825 8412 29837 8415
rect 24412 8384 29837 8412
rect 24305 8375 24363 8381
rect 29825 8381 29837 8384
rect 29871 8381 29883 8415
rect 29825 8375 29883 8381
rect 17911 8316 24072 8344
rect 24121 8347 24179 8353
rect 17911 8313 17923 8316
rect 17865 8307 17923 8313
rect 24121 8313 24133 8347
rect 24167 8344 24179 8347
rect 24320 8344 24348 8375
rect 24167 8316 24348 8344
rect 24167 8313 24179 8316
rect 24121 8307 24179 8313
rect 30098 8304 30104 8356
rect 30156 8304 30162 8356
rect 32398 8304 32404 8356
rect 32456 8304 32462 8356
rect 13541 8279 13599 8285
rect 13541 8276 13553 8279
rect 12912 8248 13553 8276
rect 12308 8236 12314 8248
rect 13541 8245 13553 8248
rect 13587 8245 13599 8279
rect 13541 8239 13599 8245
rect 14918 8236 14924 8288
rect 14976 8236 14982 8288
rect 15102 8236 15108 8288
rect 15160 8276 15166 8288
rect 15286 8276 15292 8288
rect 15160 8248 15292 8276
rect 15160 8236 15166 8248
rect 15286 8236 15292 8248
rect 15344 8276 15350 8288
rect 15562 8276 15568 8288
rect 15344 8248 15568 8276
rect 15344 8236 15350 8248
rect 15562 8236 15568 8248
rect 15620 8236 15626 8288
rect 15930 8236 15936 8288
rect 15988 8236 15994 8288
rect 16022 8236 16028 8288
rect 16080 8276 16086 8288
rect 16945 8279 17003 8285
rect 16945 8276 16957 8279
rect 16080 8248 16957 8276
rect 16080 8236 16086 8248
rect 16945 8245 16957 8248
rect 16991 8245 17003 8279
rect 16945 8239 17003 8245
rect 17494 8236 17500 8288
rect 17552 8236 17558 8288
rect 19886 8236 19892 8288
rect 19944 8276 19950 8288
rect 20257 8279 20315 8285
rect 20257 8276 20269 8279
rect 19944 8248 20269 8276
rect 19944 8236 19950 8248
rect 20257 8245 20269 8248
rect 20303 8245 20315 8279
rect 20257 8239 20315 8245
rect 21818 8236 21824 8288
rect 21876 8276 21882 8288
rect 22646 8276 22652 8288
rect 21876 8248 22652 8276
rect 21876 8236 21882 8248
rect 22646 8236 22652 8248
rect 22704 8236 22710 8288
rect 23750 8236 23756 8288
rect 23808 8236 23814 8288
rect 24026 8236 24032 8288
rect 24084 8276 24090 8288
rect 24213 8279 24271 8285
rect 24213 8276 24225 8279
rect 24084 8248 24225 8276
rect 24084 8236 24090 8248
rect 24213 8245 24225 8248
rect 24259 8245 24271 8279
rect 24213 8239 24271 8245
rect 24302 8236 24308 8288
rect 24360 8276 24366 8288
rect 27338 8276 27344 8288
rect 24360 8248 27344 8276
rect 24360 8236 24366 8248
rect 27338 8236 27344 8248
rect 27396 8236 27402 8288
rect 29914 8236 29920 8288
rect 29972 8236 29978 8288
rect 31202 8236 31208 8288
rect 31260 8236 31266 8288
rect 31294 8236 31300 8288
rect 31352 8276 31358 8288
rect 31754 8276 31760 8288
rect 31352 8248 31760 8276
rect 31352 8236 31358 8248
rect 31754 8236 31760 8248
rect 31812 8236 31818 8288
rect 1104 8186 32844 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 32844 8186
rect 1104 8112 32844 8134
rect 4798 8032 4804 8084
rect 4856 8072 4862 8084
rect 7926 8072 7932 8084
rect 4856 8044 7932 8072
rect 4856 8032 4862 8044
rect 7926 8032 7932 8044
rect 7984 8032 7990 8084
rect 8573 8075 8631 8081
rect 8573 8041 8585 8075
rect 8619 8072 8631 8075
rect 8846 8072 8852 8084
rect 8619 8044 8852 8072
rect 8619 8041 8631 8044
rect 8573 8035 8631 8041
rect 8846 8032 8852 8044
rect 8904 8032 8910 8084
rect 8938 8032 8944 8084
rect 8996 8032 9002 8084
rect 9030 8032 9036 8084
rect 9088 8072 9094 8084
rect 10870 8072 10876 8084
rect 9088 8044 10876 8072
rect 9088 8032 9094 8044
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 11241 8075 11299 8081
rect 11241 8041 11253 8075
rect 11287 8072 11299 8075
rect 11514 8072 11520 8084
rect 11287 8044 11520 8072
rect 11287 8041 11299 8044
rect 11241 8035 11299 8041
rect 11514 8032 11520 8044
rect 11572 8032 11578 8084
rect 11698 8032 11704 8084
rect 11756 8072 11762 8084
rect 11756 8044 12434 8072
rect 11756 8032 11762 8044
rect 5258 7964 5264 8016
rect 5316 8004 5322 8016
rect 5902 8004 5908 8016
rect 5316 7976 5908 8004
rect 5316 7964 5322 7976
rect 5902 7964 5908 7976
rect 5960 7964 5966 8016
rect 5994 7964 6000 8016
rect 6052 8004 6058 8016
rect 7834 8004 7840 8016
rect 6052 7976 7840 8004
rect 6052 7964 6058 7976
rect 7834 7964 7840 7976
rect 7892 8004 7898 8016
rect 9306 8004 9312 8016
rect 7892 7976 9312 8004
rect 7892 7964 7898 7976
rect 9306 7964 9312 7976
rect 9364 7964 9370 8016
rect 10778 7964 10784 8016
rect 10836 8004 10842 8016
rect 12250 8004 12256 8016
rect 10836 7976 12256 8004
rect 10836 7964 10842 7976
rect 12250 7964 12256 7976
rect 12308 7964 12314 8016
rect 12406 8004 12434 8044
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 13173 8075 13231 8081
rect 13173 8072 13185 8075
rect 12676 8044 13185 8072
rect 12676 8032 12682 8044
rect 13173 8041 13185 8044
rect 13219 8072 13231 8075
rect 13630 8072 13636 8084
rect 13219 8044 13636 8072
rect 13219 8041 13231 8044
rect 13173 8035 13231 8041
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 14645 8075 14703 8081
rect 14645 8041 14657 8075
rect 14691 8072 14703 8075
rect 14829 8075 14887 8081
rect 14691 8044 14780 8072
rect 14691 8041 14703 8044
rect 14645 8035 14703 8041
rect 14458 8004 14464 8016
rect 12406 7976 14464 8004
rect 14458 7964 14464 7976
rect 14516 7964 14522 8016
rect 14752 8004 14780 8044
rect 14829 8041 14841 8075
rect 14875 8072 14887 8075
rect 15838 8072 15844 8084
rect 14875 8044 15844 8072
rect 14875 8041 14887 8044
rect 14829 8035 14887 8041
rect 15838 8032 15844 8044
rect 15896 8032 15902 8084
rect 16666 8032 16672 8084
rect 16724 8032 16730 8084
rect 16776 8044 17080 8072
rect 16776 8004 16804 8044
rect 16942 8004 16948 8016
rect 14752 7976 16804 8004
rect 16868 7976 16948 8004
rect 5626 7896 5632 7948
rect 5684 7936 5690 7948
rect 5684 7908 6500 7936
rect 5684 7896 5690 7908
rect 6181 7871 6239 7877
rect 6181 7837 6193 7871
rect 6227 7868 6239 7871
rect 6270 7868 6276 7880
rect 6227 7840 6276 7868
rect 6227 7837 6239 7840
rect 6181 7831 6239 7837
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 6472 7877 6500 7908
rect 8110 7896 8116 7948
rect 8168 7936 8174 7948
rect 11606 7936 11612 7948
rect 8168 7908 9352 7936
rect 8168 7896 8174 7908
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 6730 7868 6736 7880
rect 6595 7840 6736 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 8389 7871 8447 7877
rect 8389 7868 8401 7871
rect 7156 7840 8401 7868
rect 7156 7828 7162 7840
rect 8389 7837 8401 7840
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 8938 7868 8944 7880
rect 8536 7840 8944 7868
rect 8536 7828 8542 7840
rect 8938 7828 8944 7840
rect 8996 7868 9002 7880
rect 9125 7871 9183 7877
rect 9125 7868 9137 7871
rect 8996 7840 9137 7868
rect 8996 7828 9002 7840
rect 9125 7837 9137 7840
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 9214 7828 9220 7880
rect 9272 7828 9278 7880
rect 9324 7877 9352 7908
rect 11440 7908 11612 7936
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7837 9367 7871
rect 9309 7831 9367 7837
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7868 9551 7871
rect 9582 7868 9588 7880
rect 9539 7840 9588 7868
rect 9539 7837 9551 7840
rect 9493 7831 9551 7837
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 10410 7868 10416 7880
rect 9692 7840 10416 7868
rect 6362 7760 6368 7812
rect 6420 7760 6426 7812
rect 6914 7760 6920 7812
rect 6972 7800 6978 7812
rect 9692 7800 9720 7840
rect 10410 7828 10416 7840
rect 10468 7828 10474 7880
rect 11440 7877 11468 7908
rect 11606 7896 11612 7908
rect 11664 7896 11670 7948
rect 13354 7896 13360 7948
rect 13412 7936 13418 7948
rect 13630 7936 13636 7948
rect 13412 7908 13636 7936
rect 13412 7896 13418 7908
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 14550 7896 14556 7948
rect 14608 7896 14614 7948
rect 15746 7896 15752 7948
rect 15804 7936 15810 7948
rect 16868 7945 16896 7976
rect 16942 7964 16948 7976
rect 17000 7964 17006 8016
rect 17052 8004 17080 8044
rect 17126 8032 17132 8084
rect 17184 8032 17190 8084
rect 17862 8072 17868 8084
rect 17512 8044 17868 8072
rect 17512 8004 17540 8044
rect 17862 8032 17868 8044
rect 17920 8032 17926 8084
rect 19521 8075 19579 8081
rect 19521 8041 19533 8075
rect 19567 8072 19579 8075
rect 19978 8072 19984 8084
rect 19567 8044 19984 8072
rect 19567 8041 19579 8044
rect 19521 8035 19579 8041
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 20073 8075 20131 8081
rect 20073 8041 20085 8075
rect 20119 8072 20131 8075
rect 20162 8072 20168 8084
rect 20119 8044 20168 8072
rect 20119 8041 20131 8044
rect 20073 8035 20131 8041
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 20990 8032 20996 8084
rect 21048 8072 21054 8084
rect 21726 8072 21732 8084
rect 21048 8044 21732 8072
rect 21048 8032 21054 8044
rect 21726 8032 21732 8044
rect 21784 8032 21790 8084
rect 22189 8075 22247 8081
rect 22189 8072 22201 8075
rect 21836 8044 22201 8072
rect 17052 7976 17540 8004
rect 17589 8007 17647 8013
rect 17589 7973 17601 8007
rect 17635 8004 17647 8007
rect 21836 8004 21864 8044
rect 22189 8041 22201 8044
rect 22235 8041 22247 8075
rect 22189 8035 22247 8041
rect 22830 8032 22836 8084
rect 22888 8032 22894 8084
rect 25774 8032 25780 8084
rect 25832 8032 25838 8084
rect 31294 8072 31300 8084
rect 25884 8044 31300 8072
rect 17635 7976 19932 8004
rect 17635 7973 17647 7976
rect 17589 7967 17647 7973
rect 16853 7939 16911 7945
rect 15804 7908 16804 7936
rect 15804 7896 15810 7908
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7868 11575 7871
rect 11790 7868 11796 7880
rect 11563 7840 11796 7868
rect 11563 7837 11575 7840
rect 11517 7831 11575 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 12618 7828 12624 7880
rect 12676 7868 12682 7880
rect 12713 7871 12771 7877
rect 12713 7868 12725 7871
rect 12676 7840 12725 7868
rect 12676 7828 12682 7840
rect 12713 7837 12725 7840
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 12986 7828 12992 7880
rect 13044 7828 13050 7880
rect 14366 7828 14372 7880
rect 14424 7864 14430 7880
rect 14461 7871 14519 7877
rect 14461 7864 14473 7871
rect 14424 7837 14473 7864
rect 14507 7837 14519 7871
rect 14424 7836 14519 7837
rect 14424 7828 14430 7836
rect 14461 7831 14519 7836
rect 16206 7828 16212 7880
rect 16264 7828 16270 7880
rect 6972 7772 9720 7800
rect 6972 7760 6978 7772
rect 9950 7760 9956 7812
rect 10008 7800 10014 7812
rect 10008 7772 13952 7800
rect 10008 7760 10014 7772
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 6638 7732 6644 7744
rect 5592 7704 6644 7732
rect 5592 7692 5598 7704
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 6733 7735 6791 7741
rect 6733 7701 6745 7735
rect 6779 7732 6791 7735
rect 10962 7732 10968 7744
rect 6779 7704 10968 7732
rect 6779 7701 6791 7704
rect 6733 7695 6791 7701
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 12897 7735 12955 7741
rect 12897 7701 12909 7735
rect 12943 7732 12955 7735
rect 13814 7732 13820 7744
rect 12943 7704 13820 7732
rect 12943 7701 12955 7704
rect 12897 7695 12955 7701
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 13924 7732 13952 7772
rect 14090 7760 14096 7812
rect 14148 7800 14154 7812
rect 14550 7800 14556 7812
rect 14148 7772 14556 7800
rect 14148 7760 14154 7772
rect 14550 7760 14556 7772
rect 14608 7800 14614 7812
rect 16025 7803 16083 7809
rect 16025 7800 16037 7803
rect 14608 7772 16037 7800
rect 14608 7760 14614 7772
rect 16025 7769 16037 7772
rect 16071 7769 16083 7803
rect 16025 7763 16083 7769
rect 16298 7760 16304 7812
rect 16356 7800 16362 7812
rect 16669 7803 16727 7809
rect 16669 7800 16681 7803
rect 16356 7772 16681 7800
rect 16356 7760 16362 7772
rect 16669 7769 16681 7772
rect 16715 7769 16727 7803
rect 16669 7763 16727 7769
rect 15838 7732 15844 7744
rect 13924 7704 15844 7732
rect 15838 7692 15844 7704
rect 15896 7692 15902 7744
rect 16390 7692 16396 7744
rect 16448 7692 16454 7744
rect 16776 7732 16804 7908
rect 16853 7905 16865 7939
rect 16899 7905 16911 7939
rect 16853 7899 16911 7905
rect 17126 7896 17132 7948
rect 17184 7936 17190 7948
rect 17604 7936 17632 7967
rect 17184 7908 17632 7936
rect 17184 7896 17190 7908
rect 17954 7896 17960 7948
rect 18012 7936 18018 7948
rect 19904 7945 19932 7976
rect 21744 7976 21864 8004
rect 22097 8007 22155 8013
rect 19337 7939 19395 7945
rect 19337 7936 19349 7939
rect 18012 7908 19349 7936
rect 18012 7896 18018 7908
rect 19337 7905 19349 7908
rect 19383 7905 19395 7939
rect 19337 7899 19395 7905
rect 19889 7939 19947 7945
rect 19889 7905 19901 7939
rect 19935 7905 19947 7939
rect 19889 7899 19947 7905
rect 19978 7896 19984 7948
rect 20036 7936 20042 7948
rect 21634 7936 21640 7948
rect 20036 7908 21640 7936
rect 20036 7896 20042 7908
rect 21634 7896 21640 7908
rect 21692 7896 21698 7948
rect 16945 7871 17003 7877
rect 16945 7837 16957 7871
rect 16991 7868 17003 7871
rect 17034 7868 17040 7880
rect 16991 7840 17040 7868
rect 16991 7837 17003 7840
rect 16945 7831 17003 7837
rect 17034 7828 17040 7840
rect 17092 7828 17098 7880
rect 17218 7828 17224 7880
rect 17276 7828 17282 7880
rect 19521 7871 19579 7877
rect 19521 7868 19533 7871
rect 19352 7840 19533 7868
rect 19352 7812 19380 7840
rect 19521 7837 19533 7840
rect 19567 7837 19579 7871
rect 20073 7871 20131 7877
rect 19521 7831 19579 7837
rect 19628 7840 20024 7868
rect 17405 7803 17463 7809
rect 17405 7769 17417 7803
rect 17451 7800 17463 7803
rect 17586 7800 17592 7812
rect 17451 7772 17592 7800
rect 17451 7769 17463 7772
rect 17405 7763 17463 7769
rect 17586 7760 17592 7772
rect 17644 7760 17650 7812
rect 18506 7760 18512 7812
rect 18564 7800 18570 7812
rect 19245 7803 19303 7809
rect 19245 7800 19257 7803
rect 18564 7772 19257 7800
rect 18564 7760 18570 7772
rect 19245 7769 19257 7772
rect 19291 7769 19303 7803
rect 19245 7763 19303 7769
rect 19334 7760 19340 7812
rect 19392 7760 19398 7812
rect 19628 7732 19656 7840
rect 19797 7803 19855 7809
rect 19797 7769 19809 7803
rect 19843 7769 19855 7803
rect 19996 7800 20024 7840
rect 20073 7837 20085 7871
rect 20119 7868 20131 7871
rect 20162 7868 20168 7880
rect 20119 7840 20168 7868
rect 20119 7837 20131 7840
rect 20073 7831 20131 7837
rect 20162 7828 20168 7840
rect 20220 7868 20226 7880
rect 20622 7868 20628 7880
rect 20220 7840 20628 7868
rect 20220 7828 20226 7840
rect 20622 7828 20628 7840
rect 20680 7828 20686 7880
rect 21744 7877 21772 7976
rect 22097 7973 22109 8007
rect 22143 8004 22155 8007
rect 22554 8004 22560 8016
rect 22143 7976 22560 8004
rect 22143 7973 22155 7976
rect 22097 7967 22155 7973
rect 22554 7964 22560 7976
rect 22612 7964 22618 8016
rect 22848 8004 22876 8032
rect 25884 8004 25912 8044
rect 31294 8032 31300 8044
rect 31352 8032 31358 8084
rect 32214 8032 32220 8084
rect 32272 8072 32278 8084
rect 32493 8075 32551 8081
rect 32493 8072 32505 8075
rect 32272 8044 32505 8072
rect 32272 8032 32278 8044
rect 32493 8041 32505 8044
rect 32539 8041 32551 8075
rect 32493 8035 32551 8041
rect 22848 7976 25912 8004
rect 29365 8007 29423 8013
rect 29365 7973 29377 8007
rect 29411 7973 29423 8007
rect 29365 7967 29423 7973
rect 21818 7896 21824 7948
rect 21876 7896 21882 7948
rect 22204 7908 25452 7936
rect 22204 7877 22232 7908
rect 21729 7871 21787 7877
rect 21729 7837 21741 7871
rect 21775 7837 21787 7871
rect 21729 7831 21787 7837
rect 22189 7871 22247 7877
rect 22189 7837 22201 7871
rect 22235 7837 22247 7871
rect 22189 7831 22247 7837
rect 22281 7871 22339 7877
rect 22281 7837 22293 7871
rect 22327 7837 22339 7871
rect 22649 7871 22707 7877
rect 22649 7868 22661 7871
rect 22281 7831 22339 7837
rect 22572 7840 22661 7868
rect 21744 7800 21772 7831
rect 19996 7772 21772 7800
rect 19797 7763 19855 7769
rect 16776 7704 19656 7732
rect 19705 7735 19763 7741
rect 19705 7701 19717 7735
rect 19751 7732 19763 7735
rect 19812 7732 19840 7763
rect 21818 7760 21824 7812
rect 21876 7800 21882 7812
rect 22296 7800 22324 7831
rect 21876 7772 22324 7800
rect 21876 7760 21882 7772
rect 19751 7704 19840 7732
rect 20257 7735 20315 7741
rect 19751 7701 19763 7704
rect 19705 7695 19763 7701
rect 20257 7701 20269 7735
rect 20303 7732 20315 7735
rect 21910 7732 21916 7744
rect 20303 7704 21916 7732
rect 20303 7701 20315 7704
rect 20257 7695 20315 7701
rect 21910 7692 21916 7704
rect 21968 7692 21974 7744
rect 22572 7741 22600 7840
rect 22649 7837 22661 7840
rect 22695 7837 22707 7871
rect 22649 7831 22707 7837
rect 22738 7828 22744 7880
rect 22796 7828 22802 7880
rect 25424 7868 25452 7908
rect 25498 7896 25504 7948
rect 25556 7936 25562 7948
rect 25869 7939 25927 7945
rect 25869 7936 25881 7939
rect 25556 7908 25881 7936
rect 25556 7896 25562 7908
rect 25869 7905 25881 7908
rect 25915 7905 25927 7939
rect 27154 7936 27160 7948
rect 25869 7899 25927 7905
rect 25976 7908 27160 7936
rect 25976 7868 26004 7908
rect 27154 7896 27160 7908
rect 27212 7896 27218 7948
rect 25424 7840 26004 7868
rect 26053 7871 26111 7877
rect 26053 7837 26065 7871
rect 26099 7868 26111 7871
rect 26878 7868 26884 7880
rect 26099 7840 26884 7868
rect 26099 7837 26111 7840
rect 26053 7831 26111 7837
rect 26878 7828 26884 7840
rect 26936 7828 26942 7880
rect 28810 7828 28816 7880
rect 28868 7828 28874 7880
rect 29178 7828 29184 7880
rect 29236 7828 29242 7880
rect 22922 7760 22928 7812
rect 22980 7800 22986 7812
rect 25777 7803 25835 7809
rect 25777 7800 25789 7803
rect 22980 7772 25789 7800
rect 22980 7760 22986 7772
rect 25777 7769 25789 7772
rect 25823 7769 25835 7803
rect 25777 7763 25835 7769
rect 28994 7760 29000 7812
rect 29052 7760 29058 7812
rect 29089 7803 29147 7809
rect 29089 7769 29101 7803
rect 29135 7769 29147 7803
rect 29380 7800 29408 7967
rect 29546 7828 29552 7880
rect 29604 7868 29610 7880
rect 31110 7868 31116 7880
rect 29604 7840 31116 7868
rect 29604 7828 29610 7840
rect 31110 7828 31116 7840
rect 31168 7828 31174 7880
rect 31202 7828 31208 7880
rect 31260 7868 31266 7880
rect 31369 7871 31427 7877
rect 31369 7868 31381 7871
rect 31260 7840 31381 7868
rect 31260 7828 31266 7840
rect 31369 7837 31381 7840
rect 31415 7837 31427 7871
rect 31369 7831 31427 7837
rect 29794 7803 29852 7809
rect 29794 7800 29806 7803
rect 29380 7772 29806 7800
rect 29089 7763 29147 7769
rect 29794 7769 29806 7772
rect 29840 7769 29852 7803
rect 29794 7763 29852 7769
rect 22557 7735 22615 7741
rect 22557 7701 22569 7735
rect 22603 7701 22615 7735
rect 22557 7695 22615 7701
rect 23017 7735 23075 7741
rect 23017 7701 23029 7735
rect 23063 7732 23075 7735
rect 23106 7732 23112 7744
rect 23063 7704 23112 7732
rect 23063 7701 23075 7704
rect 23017 7695 23075 7701
rect 23106 7692 23112 7704
rect 23164 7692 23170 7744
rect 26050 7692 26056 7744
rect 26108 7732 26114 7744
rect 26237 7735 26295 7741
rect 26237 7732 26249 7735
rect 26108 7704 26249 7732
rect 26108 7692 26114 7704
rect 26237 7701 26249 7704
rect 26283 7701 26295 7735
rect 29104 7732 29132 7763
rect 30466 7732 30472 7744
rect 29104 7704 30472 7732
rect 26237 7695 26295 7701
rect 30466 7692 30472 7704
rect 30524 7732 30530 7744
rect 30742 7732 30748 7744
rect 30524 7704 30748 7732
rect 30524 7692 30530 7704
rect 30742 7692 30748 7704
rect 30800 7692 30806 7744
rect 30926 7692 30932 7744
rect 30984 7692 30990 7744
rect 1104 7642 32844 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 32844 7642
rect 1104 7568 32844 7590
rect 6362 7488 6368 7540
rect 6420 7488 6426 7540
rect 6914 7488 6920 7540
rect 6972 7488 6978 7540
rect 7193 7531 7251 7537
rect 7193 7497 7205 7531
rect 7239 7528 7251 7531
rect 7837 7531 7895 7537
rect 7239 7500 7512 7528
rect 7239 7497 7251 7500
rect 7193 7491 7251 7497
rect 3970 7420 3976 7472
rect 4028 7460 4034 7472
rect 4065 7463 4123 7469
rect 4065 7460 4077 7463
rect 4028 7432 4077 7460
rect 4028 7420 4034 7432
rect 4065 7429 4077 7432
rect 4111 7429 4123 7463
rect 4065 7423 4123 7429
rect 4154 7420 4160 7472
rect 4212 7460 4218 7472
rect 5813 7463 5871 7469
rect 5813 7460 5825 7463
rect 4212 7432 4568 7460
rect 4212 7420 4218 7432
rect 3881 7395 3939 7401
rect 3881 7361 3893 7395
rect 3927 7361 3939 7395
rect 3881 7355 3939 7361
rect 3896 7324 3924 7355
rect 4246 7352 4252 7404
rect 4304 7352 4310 7404
rect 4540 7401 4568 7432
rect 4724 7432 5825 7460
rect 4724 7404 4752 7432
rect 5813 7429 5825 7432
rect 5859 7460 5871 7463
rect 6380 7460 6408 7488
rect 7484 7472 7512 7500
rect 7837 7497 7849 7531
rect 7883 7497 7895 7531
rect 7837 7491 7895 7497
rect 8481 7531 8539 7537
rect 8481 7497 8493 7531
rect 8527 7528 8539 7531
rect 12986 7528 12992 7540
rect 8527 7500 12992 7528
rect 8527 7497 8539 7500
rect 8481 7491 8539 7497
rect 6549 7463 6607 7469
rect 6549 7460 6561 7463
rect 5859 7432 6561 7460
rect 5859 7429 5871 7432
rect 5813 7423 5871 7429
rect 6549 7429 6561 7432
rect 6595 7429 6607 7463
rect 6549 7423 6607 7429
rect 6638 7420 6644 7472
rect 6696 7460 6702 7472
rect 6696 7432 7328 7460
rect 6696 7420 6702 7432
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 4706 7352 4712 7404
rect 4764 7352 4770 7404
rect 4798 7352 4804 7404
rect 4856 7352 4862 7404
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7361 4951 7395
rect 4893 7355 4951 7361
rect 4816 7324 4844 7352
rect 3896 7296 4844 7324
rect 4908 7324 4936 7355
rect 4982 7352 4988 7404
rect 5040 7392 5046 7404
rect 5353 7395 5411 7401
rect 5353 7392 5365 7395
rect 5040 7364 5365 7392
rect 5040 7352 5046 7364
rect 5353 7361 5365 7364
rect 5399 7361 5411 7395
rect 5353 7355 5411 7361
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 5592 7364 5641 7392
rect 5592 7352 5598 7364
rect 5629 7361 5641 7364
rect 5675 7361 5687 7395
rect 5629 7355 5687 7361
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 6012 7324 6040 7355
rect 6362 7352 6368 7404
rect 6420 7352 6426 7404
rect 6730 7352 6736 7404
rect 6788 7352 6794 7404
rect 7006 7352 7012 7404
rect 7064 7352 7070 7404
rect 7300 7401 7328 7432
rect 7466 7420 7472 7472
rect 7524 7420 7530 7472
rect 7852 7460 7880 7491
rect 12986 7488 12992 7500
rect 13044 7488 13050 7540
rect 13262 7488 13268 7540
rect 13320 7528 13326 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 13320 7500 13461 7528
rect 13320 7488 13326 7500
rect 13449 7497 13461 7500
rect 13495 7528 13507 7531
rect 14366 7528 14372 7540
rect 13495 7500 14372 7528
rect 13495 7497 13507 7500
rect 13449 7491 13507 7497
rect 14366 7488 14372 7500
rect 14424 7488 14430 7540
rect 16206 7488 16212 7540
rect 16264 7528 16270 7540
rect 16301 7531 16359 7537
rect 16301 7528 16313 7531
rect 16264 7500 16313 7528
rect 16264 7488 16270 7500
rect 16301 7497 16313 7500
rect 16347 7497 16359 7531
rect 16301 7491 16359 7497
rect 18782 7488 18788 7540
rect 18840 7528 18846 7540
rect 21913 7531 21971 7537
rect 21913 7528 21925 7531
rect 18840 7500 21925 7528
rect 18840 7488 18846 7500
rect 21913 7497 21925 7500
rect 21959 7528 21971 7531
rect 21959 7500 22140 7528
rect 21959 7497 21971 7500
rect 21913 7491 21971 7497
rect 7852 7432 9904 7460
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7361 7619 7395
rect 7561 7355 7619 7361
rect 6748 7324 6776 7352
rect 4908 7296 6776 7324
rect 4433 7259 4491 7265
rect 4433 7225 4445 7259
rect 4479 7225 4491 7259
rect 4433 7219 4491 7225
rect 4448 7188 4476 7219
rect 5074 7216 5080 7268
rect 5132 7216 5138 7268
rect 5184 7265 5212 7296
rect 5169 7259 5227 7265
rect 5169 7225 5181 7259
rect 5215 7225 5227 7259
rect 5169 7219 5227 7225
rect 5902 7216 5908 7268
rect 5960 7256 5966 7268
rect 6362 7256 6368 7268
rect 5960 7228 6368 7256
rect 5960 7216 5966 7228
rect 6362 7216 6368 7228
rect 6420 7256 6426 7268
rect 7576 7256 7604 7355
rect 7650 7352 7656 7404
rect 7708 7352 7714 7404
rect 7834 7352 7840 7404
rect 7892 7392 7898 7404
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 7892 7364 7941 7392
rect 7892 7352 7898 7364
rect 7929 7361 7941 7364
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 8110 7352 8116 7404
rect 8168 7352 8174 7404
rect 8202 7352 8208 7404
rect 8260 7352 8266 7404
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7392 8355 7395
rect 8478 7392 8484 7404
rect 8343 7364 8484 7392
rect 8343 7361 8355 7364
rect 8297 7355 8355 7361
rect 8478 7352 8484 7364
rect 8536 7352 8542 7404
rect 8570 7352 8576 7404
rect 8628 7352 8634 7404
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 8128 7324 8156 7352
rect 8772 7324 8800 7355
rect 8846 7352 8852 7404
rect 8904 7352 8910 7404
rect 8938 7352 8944 7404
rect 8996 7352 9002 7404
rect 9030 7352 9036 7404
rect 9088 7392 9094 7404
rect 9217 7395 9275 7401
rect 9217 7392 9229 7395
rect 9088 7364 9229 7392
rect 9088 7352 9094 7364
rect 9217 7361 9229 7364
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7361 9459 7395
rect 9401 7355 9459 7361
rect 9416 7324 9444 7355
rect 9490 7352 9496 7404
rect 9548 7352 9554 7404
rect 9876 7401 9904 7432
rect 10502 7420 10508 7472
rect 10560 7460 10566 7472
rect 10560 7432 13216 7460
rect 10560 7420 10566 7432
rect 9585 7395 9643 7401
rect 9585 7361 9597 7395
rect 9631 7361 9643 7395
rect 9585 7355 9643 7361
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 9600 7324 9628 7355
rect 10410 7352 10416 7404
rect 10468 7352 10474 7404
rect 12526 7352 12532 7404
rect 12584 7352 12590 7404
rect 12805 7395 12863 7401
rect 12805 7361 12817 7395
rect 12851 7392 12863 7395
rect 13078 7392 13084 7404
rect 12851 7364 13084 7392
rect 12851 7361 12863 7364
rect 12805 7355 12863 7361
rect 13078 7352 13084 7364
rect 13136 7352 13142 7404
rect 13188 7401 13216 7432
rect 13354 7420 13360 7472
rect 13412 7420 13418 7472
rect 14458 7420 14464 7472
rect 14516 7460 14522 7472
rect 15470 7460 15476 7472
rect 14516 7432 15476 7460
rect 14516 7420 14522 7432
rect 15470 7420 15476 7432
rect 15528 7460 15534 7472
rect 17586 7460 17592 7472
rect 15528 7432 17592 7460
rect 15528 7420 15534 7432
rect 17586 7420 17592 7432
rect 17644 7420 17650 7472
rect 19334 7420 19340 7472
rect 19392 7420 19398 7472
rect 22112 7469 22140 7500
rect 23382 7488 23388 7540
rect 23440 7528 23446 7540
rect 24305 7531 24363 7537
rect 23440 7500 24256 7528
rect 23440 7488 23446 7500
rect 22097 7463 22155 7469
rect 22097 7429 22109 7463
rect 22143 7429 22155 7463
rect 23845 7463 23903 7469
rect 23845 7460 23857 7463
rect 22097 7423 22155 7429
rect 22296 7432 23857 7460
rect 13173 7395 13231 7401
rect 13173 7361 13185 7395
rect 13219 7392 13231 7395
rect 13538 7392 13544 7404
rect 13219 7364 13544 7392
rect 13219 7361 13231 7364
rect 13173 7355 13231 7361
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 13633 7395 13691 7401
rect 13633 7361 13645 7395
rect 13679 7392 13691 7395
rect 13814 7392 13820 7404
rect 13679 7364 13820 7392
rect 13679 7361 13691 7364
rect 13633 7355 13691 7361
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 16485 7395 16543 7401
rect 16485 7392 16497 7395
rect 13924 7364 16497 7392
rect 9950 7324 9956 7336
rect 8128 7296 9444 7324
rect 9508 7296 9628 7324
rect 9784 7296 9956 7324
rect 6420 7228 7604 7256
rect 6420 7216 6426 7228
rect 8938 7216 8944 7268
rect 8996 7256 9002 7268
rect 9508 7256 9536 7296
rect 9784 7265 9812 7296
rect 9950 7284 9956 7296
rect 10008 7284 10014 7336
rect 12345 7327 12403 7333
rect 12345 7293 12357 7327
rect 12391 7324 12403 7327
rect 12618 7324 12624 7336
rect 12391 7296 12624 7324
rect 12391 7293 12403 7296
rect 12345 7287 12403 7293
rect 12618 7284 12624 7296
rect 12676 7284 12682 7336
rect 12728 7296 13308 7324
rect 8996 7228 9536 7256
rect 9769 7259 9827 7265
rect 8996 7216 9002 7228
rect 9769 7225 9781 7259
rect 9815 7225 9827 7259
rect 9769 7219 9827 7225
rect 9858 7216 9864 7268
rect 9916 7256 9922 7268
rect 10045 7259 10103 7265
rect 10045 7256 10057 7259
rect 9916 7228 10057 7256
rect 9916 7216 9922 7228
rect 10045 7225 10057 7228
rect 10091 7256 10103 7259
rect 12728 7256 12756 7296
rect 13170 7256 13176 7268
rect 10091 7228 12756 7256
rect 12820 7228 13176 7256
rect 10091 7225 10103 7228
rect 10045 7219 10103 7225
rect 5534 7188 5540 7200
rect 4448 7160 5540 7188
rect 5534 7148 5540 7160
rect 5592 7188 5598 7200
rect 6086 7188 6092 7200
rect 5592 7160 6092 7188
rect 5592 7148 5598 7160
rect 6086 7148 6092 7160
rect 6144 7148 6150 7200
rect 6181 7191 6239 7197
rect 6181 7157 6193 7191
rect 6227 7188 6239 7191
rect 6822 7188 6828 7200
rect 6227 7160 6828 7188
rect 6227 7157 6239 7160
rect 6181 7151 6239 7157
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 7006 7148 7012 7200
rect 7064 7188 7070 7200
rect 9030 7188 9036 7200
rect 7064 7160 9036 7188
rect 7064 7148 7070 7160
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 9125 7191 9183 7197
rect 9125 7157 9137 7191
rect 9171 7188 9183 7191
rect 10502 7188 10508 7200
rect 9171 7160 10508 7188
rect 9171 7157 9183 7160
rect 9125 7151 9183 7157
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 10597 7191 10655 7197
rect 10597 7157 10609 7191
rect 10643 7188 10655 7191
rect 10686 7188 10692 7200
rect 10643 7160 10692 7188
rect 10643 7157 10655 7160
rect 10597 7151 10655 7157
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 10870 7148 10876 7200
rect 10928 7188 10934 7200
rect 12618 7188 12624 7200
rect 10928 7160 12624 7188
rect 10928 7148 10934 7160
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 12820 7197 12848 7228
rect 13170 7216 13176 7228
rect 13228 7216 13234 7268
rect 12805 7191 12863 7197
rect 12805 7157 12817 7191
rect 12851 7157 12863 7191
rect 12805 7151 12863 7157
rect 12986 7148 12992 7200
rect 13044 7148 13050 7200
rect 13280 7188 13308 7296
rect 13446 7284 13452 7336
rect 13504 7324 13510 7336
rect 13924 7324 13952 7364
rect 16485 7361 16497 7364
rect 16531 7361 16543 7395
rect 16485 7355 16543 7361
rect 16574 7352 16580 7404
rect 16632 7392 16638 7404
rect 22296 7392 22324 7432
rect 23845 7429 23857 7432
rect 23891 7429 23903 7463
rect 23845 7423 23903 7429
rect 16632 7364 22324 7392
rect 22373 7395 22431 7401
rect 16632 7352 16638 7364
rect 22373 7361 22385 7395
rect 22419 7392 22431 7395
rect 23658 7392 23664 7404
rect 22419 7364 23664 7392
rect 22419 7361 22431 7364
rect 22373 7355 22431 7361
rect 23658 7352 23664 7364
rect 23716 7352 23722 7404
rect 24121 7395 24179 7401
rect 24121 7392 24133 7395
rect 23860 7364 24133 7392
rect 23860 7336 23888 7364
rect 24121 7361 24133 7364
rect 24167 7361 24179 7395
rect 24228 7392 24256 7500
rect 24305 7497 24317 7531
rect 24351 7497 24363 7531
rect 24305 7491 24363 7497
rect 26237 7531 26295 7537
rect 26237 7497 26249 7531
rect 26283 7528 26295 7531
rect 27614 7528 27620 7540
rect 26283 7500 27620 7528
rect 26283 7497 26295 7500
rect 26237 7491 26295 7497
rect 24320 7460 24348 7491
rect 27614 7488 27620 7500
rect 27672 7488 27678 7540
rect 29178 7488 29184 7540
rect 29236 7528 29242 7540
rect 30101 7531 30159 7537
rect 30101 7528 30113 7531
rect 29236 7500 30113 7528
rect 29236 7488 29242 7500
rect 30101 7497 30113 7500
rect 30147 7497 30159 7531
rect 30101 7491 30159 7497
rect 24320 7432 25912 7460
rect 25884 7401 25912 7432
rect 27890 7420 27896 7472
rect 27948 7420 27954 7472
rect 28077 7463 28135 7469
rect 28077 7429 28089 7463
rect 28123 7460 28135 7463
rect 28166 7460 28172 7472
rect 28123 7432 28172 7460
rect 28123 7429 28135 7432
rect 28077 7423 28135 7429
rect 28166 7420 28172 7432
rect 28224 7420 28230 7472
rect 25869 7395 25927 7401
rect 24228 7364 24348 7392
rect 24121 7355 24179 7361
rect 13504 7296 13952 7324
rect 13504 7284 13510 7296
rect 16390 7284 16396 7336
rect 16448 7324 16454 7336
rect 20162 7324 20168 7336
rect 16448 7296 20168 7324
rect 16448 7284 16454 7296
rect 20162 7284 20168 7296
rect 20220 7284 20226 7336
rect 22281 7327 22339 7333
rect 22281 7293 22293 7327
rect 22327 7293 22339 7327
rect 22281 7287 22339 7293
rect 13906 7216 13912 7268
rect 13964 7256 13970 7268
rect 14274 7256 14280 7268
rect 13964 7228 14280 7256
rect 13964 7216 13970 7228
rect 14274 7216 14280 7228
rect 14332 7256 14338 7268
rect 22296 7256 22324 7287
rect 23842 7284 23848 7336
rect 23900 7284 23906 7336
rect 24029 7327 24087 7333
rect 24029 7293 24041 7327
rect 24075 7324 24087 7327
rect 24210 7324 24216 7336
rect 24075 7296 24216 7324
rect 24075 7293 24087 7296
rect 24029 7287 24087 7293
rect 24210 7284 24216 7296
rect 24268 7284 24274 7336
rect 24320 7324 24348 7364
rect 25869 7361 25881 7395
rect 25915 7361 25927 7395
rect 25869 7355 25927 7361
rect 25958 7352 25964 7404
rect 26016 7352 26022 7404
rect 27801 7395 27859 7401
rect 27801 7361 27813 7395
rect 27847 7392 27859 7395
rect 27908 7392 27936 7420
rect 27847 7364 27936 7392
rect 31941 7395 31999 7401
rect 27847 7361 27859 7364
rect 27801 7355 27859 7361
rect 31941 7361 31953 7395
rect 31987 7392 31999 7395
rect 32125 7395 32183 7401
rect 32125 7392 32137 7395
rect 31987 7364 32137 7392
rect 31987 7361 31999 7364
rect 31941 7355 31999 7361
rect 32125 7361 32137 7364
rect 32171 7392 32183 7395
rect 32490 7392 32496 7404
rect 32171 7364 32496 7392
rect 32171 7361 32183 7364
rect 32125 7355 32183 7361
rect 32490 7352 32496 7364
rect 32548 7352 32554 7404
rect 27893 7327 27951 7333
rect 27893 7324 27905 7327
rect 24320 7296 27905 7324
rect 27893 7293 27905 7296
rect 27939 7293 27951 7327
rect 27893 7287 27951 7293
rect 30745 7327 30803 7333
rect 30745 7293 30757 7327
rect 30791 7324 30803 7327
rect 30926 7324 30932 7336
rect 30791 7296 30932 7324
rect 30791 7293 30803 7296
rect 30745 7287 30803 7293
rect 30926 7284 30932 7296
rect 30984 7324 30990 7336
rect 32214 7324 32220 7336
rect 30984 7296 32220 7324
rect 30984 7284 30990 7296
rect 32214 7284 32220 7296
rect 32272 7284 32278 7336
rect 27617 7259 27675 7265
rect 27617 7256 27629 7259
rect 14332 7228 22140 7256
rect 22296 7228 27629 7256
rect 14332 7216 14338 7228
rect 19242 7188 19248 7200
rect 13280 7160 19248 7188
rect 19242 7148 19248 7160
rect 19300 7148 19306 7200
rect 22112 7197 22140 7228
rect 27617 7225 27629 7228
rect 27663 7225 27675 7259
rect 27617 7219 27675 7225
rect 22097 7191 22155 7197
rect 22097 7157 22109 7191
rect 22143 7157 22155 7191
rect 22097 7151 22155 7157
rect 22370 7148 22376 7200
rect 22428 7188 22434 7200
rect 22557 7191 22615 7197
rect 22557 7188 22569 7191
rect 22428 7160 22569 7188
rect 22428 7148 22434 7160
rect 22557 7157 22569 7160
rect 22603 7157 22615 7191
rect 22557 7151 22615 7157
rect 24118 7148 24124 7200
rect 24176 7148 24182 7200
rect 26050 7148 26056 7200
rect 26108 7148 26114 7200
rect 27798 7148 27804 7200
rect 27856 7148 27862 7200
rect 30834 7148 30840 7200
rect 30892 7188 30898 7200
rect 31297 7191 31355 7197
rect 31297 7188 31309 7191
rect 30892 7160 31309 7188
rect 30892 7148 30898 7160
rect 31297 7157 31309 7160
rect 31343 7157 31355 7191
rect 31297 7151 31355 7157
rect 32306 7148 32312 7200
rect 32364 7148 32370 7200
rect 1104 7098 32844 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 32844 7098
rect 1104 7024 32844 7046
rect 4706 6944 4712 6996
rect 4764 6944 4770 6996
rect 5074 6944 5080 6996
rect 5132 6984 5138 6996
rect 5132 6956 7144 6984
rect 5132 6944 5138 6956
rect 3970 6876 3976 6928
rect 4028 6916 4034 6928
rect 4028 6888 4660 6916
rect 4028 6876 4034 6888
rect 4632 6780 4660 6888
rect 5442 6876 5448 6928
rect 5500 6916 5506 6928
rect 7006 6916 7012 6928
rect 5500 6888 7012 6916
rect 5500 6876 5506 6888
rect 7006 6876 7012 6888
rect 7064 6876 7070 6928
rect 7116 6916 7144 6956
rect 7650 6944 7656 6996
rect 7708 6984 7714 6996
rect 7837 6987 7895 6993
rect 7837 6984 7849 6987
rect 7708 6956 7849 6984
rect 7708 6944 7714 6956
rect 7837 6953 7849 6956
rect 7883 6953 7895 6987
rect 7837 6947 7895 6953
rect 7926 6944 7932 6996
rect 7984 6984 7990 6996
rect 9490 6984 9496 6996
rect 7984 6956 9496 6984
rect 7984 6944 7990 6956
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 9585 6987 9643 6993
rect 9585 6953 9597 6987
rect 9631 6984 9643 6987
rect 9858 6984 9864 6996
rect 9631 6956 9864 6984
rect 9631 6953 9643 6956
rect 9585 6947 9643 6953
rect 9858 6944 9864 6956
rect 9916 6944 9922 6996
rect 10505 6987 10563 6993
rect 10505 6953 10517 6987
rect 10551 6984 10563 6987
rect 10686 6984 10692 6996
rect 10551 6956 10692 6984
rect 10551 6953 10563 6956
rect 10505 6947 10563 6953
rect 10686 6944 10692 6956
rect 10744 6944 10750 6996
rect 11238 6944 11244 6996
rect 11296 6984 11302 6996
rect 11422 6984 11428 6996
rect 11296 6956 11428 6984
rect 11296 6944 11302 6956
rect 11422 6944 11428 6956
rect 11480 6944 11486 6996
rect 12989 6987 13047 6993
rect 12989 6953 13001 6987
rect 13035 6984 13047 6987
rect 13078 6984 13084 6996
rect 13035 6956 13084 6984
rect 13035 6953 13047 6956
rect 12989 6947 13047 6953
rect 13078 6944 13084 6956
rect 13136 6944 13142 6996
rect 13630 6944 13636 6996
rect 13688 6944 13694 6996
rect 14826 6984 14832 6996
rect 13740 6956 14832 6984
rect 11514 6916 11520 6928
rect 7116 6888 11520 6916
rect 11514 6876 11520 6888
rect 11572 6876 11578 6928
rect 13446 6916 13452 6928
rect 12406 6888 13452 6916
rect 9582 6808 9588 6860
rect 9640 6848 9646 6860
rect 10321 6851 10379 6857
rect 10321 6848 10333 6851
rect 9640 6820 10333 6848
rect 9640 6808 9646 6820
rect 10321 6817 10333 6820
rect 10367 6817 10379 6851
rect 10321 6811 10379 6817
rect 10428 6820 11652 6848
rect 4893 6783 4951 6789
rect 4893 6780 4905 6783
rect 4632 6752 4905 6780
rect 4893 6749 4905 6752
rect 4939 6749 4951 6783
rect 4893 6743 4951 6749
rect 7653 6783 7711 6789
rect 7653 6749 7665 6783
rect 7699 6780 7711 6783
rect 7742 6780 7748 6792
rect 7699 6752 7748 6780
rect 7699 6749 7711 6752
rect 7653 6743 7711 6749
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 9306 6740 9312 6792
rect 9364 6740 9370 6792
rect 9398 6740 9404 6792
rect 9456 6740 9462 6792
rect 10428 6780 10456 6820
rect 9600 6752 10456 6780
rect 10505 6783 10563 6789
rect 9600 6721 9628 6752
rect 10505 6749 10517 6783
rect 10551 6780 10563 6783
rect 10594 6780 10600 6792
rect 10551 6752 10600 6780
rect 10551 6749 10563 6752
rect 10505 6743 10563 6749
rect 10594 6740 10600 6752
rect 10652 6740 10658 6792
rect 10778 6740 10784 6792
rect 10836 6780 10842 6792
rect 10873 6783 10931 6789
rect 10873 6780 10885 6783
rect 10836 6752 10885 6780
rect 10836 6740 10842 6752
rect 10873 6749 10885 6752
rect 10919 6749 10931 6783
rect 10873 6743 10931 6749
rect 11149 6783 11207 6789
rect 11149 6749 11161 6783
rect 11195 6749 11207 6783
rect 11149 6743 11207 6749
rect 9585 6715 9643 6721
rect 9585 6681 9597 6715
rect 9631 6681 9643 6715
rect 9585 6675 9643 6681
rect 10229 6715 10287 6721
rect 10229 6681 10241 6715
rect 10275 6712 10287 6715
rect 10962 6712 10968 6724
rect 10275 6684 10968 6712
rect 10275 6681 10287 6684
rect 10229 6675 10287 6681
rect 10962 6672 10968 6684
rect 11020 6712 11026 6724
rect 11164 6712 11192 6743
rect 11238 6740 11244 6792
rect 11296 6780 11302 6792
rect 11425 6783 11483 6789
rect 11425 6780 11437 6783
rect 11296 6752 11437 6780
rect 11296 6740 11302 6752
rect 11425 6749 11437 6752
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 11514 6740 11520 6792
rect 11572 6740 11578 6792
rect 11624 6780 11652 6820
rect 11698 6808 11704 6860
rect 11756 6848 11762 6860
rect 12406 6848 12434 6888
rect 13446 6876 13452 6888
rect 13504 6916 13510 6928
rect 13740 6916 13768 6956
rect 14826 6944 14832 6956
rect 14884 6944 14890 6996
rect 15120 6956 15332 6984
rect 13504 6888 13768 6916
rect 13817 6919 13875 6925
rect 13504 6876 13510 6888
rect 13817 6885 13829 6919
rect 13863 6916 13875 6919
rect 13863 6888 13952 6916
rect 13863 6885 13875 6888
rect 13817 6879 13875 6885
rect 13354 6848 13360 6860
rect 11756 6820 12434 6848
rect 12820 6820 13360 6848
rect 11756 6808 11762 6820
rect 12820 6789 12848 6820
rect 13354 6808 13360 6820
rect 13412 6808 13418 6860
rect 13541 6851 13599 6857
rect 13541 6817 13553 6851
rect 13587 6848 13599 6851
rect 13924 6848 13952 6888
rect 15120 6848 15148 6956
rect 13587 6820 13768 6848
rect 13924 6820 15148 6848
rect 15304 6848 15332 6956
rect 15470 6944 15476 6996
rect 15528 6984 15534 6996
rect 17957 6987 18015 6993
rect 15528 6956 16068 6984
rect 15528 6944 15534 6956
rect 16040 6916 16068 6956
rect 17957 6953 17969 6987
rect 18003 6984 18015 6987
rect 18506 6984 18512 6996
rect 18003 6956 18512 6984
rect 18003 6953 18015 6956
rect 17957 6947 18015 6953
rect 18506 6944 18512 6956
rect 18564 6944 18570 6996
rect 20349 6987 20407 6993
rect 20349 6953 20361 6987
rect 20395 6984 20407 6987
rect 20622 6984 20628 6996
rect 20395 6956 20628 6984
rect 20395 6953 20407 6956
rect 20349 6947 20407 6953
rect 20622 6944 20628 6956
rect 20680 6944 20686 6996
rect 22189 6987 22247 6993
rect 22189 6953 22201 6987
rect 22235 6984 22247 6987
rect 22557 6987 22615 6993
rect 22557 6984 22569 6987
rect 22235 6956 22569 6984
rect 22235 6953 22247 6956
rect 22189 6947 22247 6953
rect 22557 6953 22569 6956
rect 22603 6984 22615 6987
rect 23198 6984 23204 6996
rect 22603 6956 23204 6984
rect 22603 6953 22615 6956
rect 22557 6947 22615 6953
rect 23198 6944 23204 6956
rect 23256 6944 23262 6996
rect 26421 6987 26479 6993
rect 26421 6953 26433 6987
rect 26467 6953 26479 6987
rect 26421 6947 26479 6953
rect 15764 6888 15976 6916
rect 16040 6888 18460 6916
rect 15764 6848 15792 6888
rect 15304 6820 15792 6848
rect 15948 6848 15976 6888
rect 16574 6848 16580 6860
rect 15948 6820 16580 6848
rect 13587 6817 13599 6820
rect 13541 6811 13599 6817
rect 12805 6783 12863 6789
rect 11624 6752 11836 6780
rect 11532 6712 11560 6740
rect 11020 6684 11100 6712
rect 11164 6684 11560 6712
rect 11020 6672 11026 6684
rect 9125 6647 9183 6653
rect 9125 6613 9137 6647
rect 9171 6644 9183 6647
rect 9490 6644 9496 6656
rect 9171 6616 9496 6644
rect 9171 6613 9183 6616
rect 9125 6607 9183 6613
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 10689 6647 10747 6653
rect 10689 6613 10701 6647
rect 10735 6644 10747 6647
rect 10870 6644 10876 6656
rect 10735 6616 10876 6644
rect 10735 6613 10747 6616
rect 10689 6607 10747 6613
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 11072 6653 11100 6684
rect 11057 6647 11115 6653
rect 11057 6613 11069 6647
rect 11103 6613 11115 6647
rect 11057 6607 11115 6613
rect 11333 6647 11391 6653
rect 11333 6613 11345 6647
rect 11379 6644 11391 6647
rect 11514 6644 11520 6656
rect 11379 6616 11520 6644
rect 11379 6613 11391 6616
rect 11333 6607 11391 6613
rect 11514 6604 11520 6616
rect 11572 6604 11578 6656
rect 11808 6644 11836 6752
rect 12805 6749 12817 6783
rect 12851 6749 12863 6783
rect 12805 6743 12863 6749
rect 12986 6740 12992 6792
rect 13044 6780 13050 6792
rect 13449 6783 13507 6789
rect 13449 6780 13461 6783
rect 13044 6752 13461 6780
rect 13044 6740 13050 6752
rect 13449 6749 13461 6752
rect 13495 6749 13507 6783
rect 13449 6743 13507 6749
rect 11882 6672 11888 6724
rect 11940 6712 11946 6724
rect 13556 6712 13584 6811
rect 11940 6684 13584 6712
rect 13740 6712 13768 6820
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 18432 6857 18460 6888
rect 18874 6876 18880 6928
rect 18932 6916 18938 6928
rect 18932 6888 19196 6916
rect 18932 6876 18938 6888
rect 18417 6851 18475 6857
rect 18417 6817 18429 6851
rect 18463 6848 18475 6851
rect 19168 6848 19196 6888
rect 19242 6876 19248 6928
rect 19300 6916 19306 6928
rect 26436 6916 26464 6947
rect 32490 6944 32496 6996
rect 32548 6944 32554 6996
rect 19300 6888 26464 6916
rect 19300 6876 19306 6888
rect 18463 6820 18920 6848
rect 19168 6820 20208 6848
rect 18463 6817 18475 6820
rect 18417 6811 18475 6817
rect 15841 6799 15899 6805
rect 13906 6740 13912 6792
rect 13964 6780 13970 6792
rect 15102 6780 15108 6792
rect 13964 6752 15108 6780
rect 13964 6740 13970 6752
rect 15102 6740 15108 6752
rect 15160 6740 15166 6792
rect 15194 6740 15200 6792
rect 15252 6740 15258 6792
rect 15841 6765 15853 6799
rect 15887 6765 15899 6799
rect 15841 6759 15899 6765
rect 15856 6724 15884 6759
rect 16206 6740 16212 6792
rect 16264 6740 16270 6792
rect 17770 6740 17776 6792
rect 17828 6740 17834 6792
rect 17954 6740 17960 6792
rect 18012 6780 18018 6792
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 18012 6752 18245 6780
rect 18012 6740 18018 6752
rect 18233 6749 18245 6752
rect 18279 6749 18291 6783
rect 18233 6743 18291 6749
rect 18785 6783 18843 6789
rect 18785 6749 18797 6783
rect 18831 6749 18843 6783
rect 18892 6780 18920 6820
rect 19978 6780 19984 6792
rect 18892 6752 19984 6780
rect 18785 6743 18843 6749
rect 14458 6712 14464 6724
rect 13740 6684 14464 6712
rect 11940 6672 11946 6684
rect 14458 6672 14464 6684
rect 14516 6672 14522 6724
rect 15381 6715 15439 6721
rect 15381 6681 15393 6715
rect 15427 6681 15439 6715
rect 15381 6675 15439 6681
rect 12342 6644 12348 6656
rect 11808 6616 12348 6644
rect 12342 6604 12348 6616
rect 12400 6644 12406 6656
rect 15396 6644 15424 6675
rect 15470 6672 15476 6724
rect 15528 6712 15534 6724
rect 15565 6715 15623 6721
rect 15565 6712 15577 6715
rect 15528 6684 15577 6712
rect 15528 6672 15534 6684
rect 15565 6681 15577 6684
rect 15611 6681 15623 6715
rect 15565 6675 15623 6681
rect 15838 6672 15844 6724
rect 15896 6672 15902 6724
rect 16022 6672 16028 6724
rect 16080 6672 16086 6724
rect 17586 6672 17592 6724
rect 17644 6672 17650 6724
rect 18509 6715 18567 6721
rect 18509 6681 18521 6715
rect 18555 6712 18567 6715
rect 18690 6712 18696 6724
rect 18555 6684 18696 6712
rect 18555 6681 18567 6684
rect 18509 6675 18567 6681
rect 18690 6672 18696 6684
rect 18748 6672 18754 6724
rect 12400 6616 15424 6644
rect 12400 6604 12406 6616
rect 15654 6604 15660 6656
rect 15712 6604 15718 6656
rect 16393 6647 16451 6653
rect 16393 6613 16405 6647
rect 16439 6644 16451 6647
rect 17678 6644 17684 6656
rect 16439 6616 17684 6644
rect 16439 6613 16451 6616
rect 16393 6607 16451 6613
rect 17678 6604 17684 6616
rect 17736 6604 17742 6656
rect 18046 6604 18052 6656
rect 18104 6604 18110 6656
rect 18414 6604 18420 6656
rect 18472 6644 18478 6656
rect 18601 6647 18659 6653
rect 18601 6644 18613 6647
rect 18472 6616 18613 6644
rect 18472 6604 18478 6616
rect 18601 6613 18613 6616
rect 18647 6644 18659 6647
rect 18800 6644 18828 6743
rect 19978 6740 19984 6752
rect 20036 6740 20042 6792
rect 20070 6740 20076 6792
rect 20128 6740 20134 6792
rect 20180 6780 20208 6820
rect 20254 6808 20260 6860
rect 20312 6808 20318 6860
rect 21634 6808 21640 6860
rect 21692 6848 21698 6860
rect 22094 6848 22100 6860
rect 21692 6820 22100 6848
rect 21692 6808 21698 6820
rect 22094 6808 22100 6820
rect 22152 6848 22158 6860
rect 22152 6820 24440 6848
rect 22152 6808 22158 6820
rect 20349 6783 20407 6789
rect 20349 6780 20361 6783
rect 20180 6752 20361 6780
rect 20349 6749 20361 6752
rect 20395 6749 20407 6783
rect 20349 6743 20407 6749
rect 22370 6740 22376 6792
rect 22428 6740 22434 6792
rect 22462 6740 22468 6792
rect 22520 6740 22526 6792
rect 22554 6740 22560 6792
rect 22612 6740 22618 6792
rect 24412 6789 24440 6820
rect 24762 6808 24768 6860
rect 24820 6808 24826 6860
rect 26142 6808 26148 6860
rect 26200 6848 26206 6860
rect 29546 6848 29552 6860
rect 26200 6820 29552 6848
rect 26200 6808 26206 6820
rect 29546 6808 29552 6820
rect 29604 6848 29610 6860
rect 31113 6851 31171 6857
rect 31113 6848 31125 6851
rect 29604 6820 31125 6848
rect 29604 6808 29610 6820
rect 31113 6817 31125 6820
rect 31159 6817 31171 6851
rect 31113 6811 31171 6817
rect 24397 6783 24455 6789
rect 24397 6749 24409 6783
rect 24443 6749 24455 6783
rect 24397 6743 24455 6749
rect 25314 6740 25320 6792
rect 25372 6780 25378 6792
rect 26421 6783 26479 6789
rect 26421 6780 26433 6783
rect 25372 6752 26433 6780
rect 25372 6740 25378 6752
rect 26421 6749 26433 6752
rect 26467 6749 26479 6783
rect 26421 6743 26479 6749
rect 26510 6740 26516 6792
rect 26568 6740 26574 6792
rect 30098 6740 30104 6792
rect 30156 6780 30162 6792
rect 30469 6783 30527 6789
rect 30469 6780 30481 6783
rect 30156 6752 30481 6780
rect 30156 6740 30162 6752
rect 30469 6749 30481 6752
rect 30515 6749 30527 6783
rect 30469 6743 30527 6749
rect 30742 6740 30748 6792
rect 30800 6740 30806 6792
rect 30834 6740 30840 6792
rect 30892 6740 30898 6792
rect 18874 6672 18880 6724
rect 18932 6712 18938 6724
rect 20088 6712 20116 6740
rect 18932 6684 20116 6712
rect 22281 6715 22339 6721
rect 18932 6672 18938 6684
rect 22281 6681 22293 6715
rect 22327 6712 22339 6715
rect 22388 6712 22416 6740
rect 22327 6684 22416 6712
rect 22327 6681 22339 6684
rect 22281 6675 22339 6681
rect 24578 6672 24584 6724
rect 24636 6672 24642 6724
rect 28994 6672 29000 6724
rect 29052 6712 29058 6724
rect 30653 6715 30711 6721
rect 30653 6712 30665 6715
rect 29052 6684 30665 6712
rect 29052 6672 29058 6684
rect 30653 6681 30665 6684
rect 30699 6681 30711 6715
rect 31358 6715 31416 6721
rect 31358 6712 31370 6715
rect 30653 6675 30711 6681
rect 31036 6684 31370 6712
rect 18647 6616 18828 6644
rect 18647 6613 18659 6616
rect 18601 6607 18659 6613
rect 18966 6604 18972 6656
rect 19024 6604 19030 6656
rect 20530 6604 20536 6656
rect 20588 6604 20594 6656
rect 20622 6604 20628 6656
rect 20680 6644 20686 6656
rect 22646 6644 22652 6656
rect 20680 6616 22652 6644
rect 20680 6604 20686 6616
rect 22646 6604 22652 6616
rect 22704 6604 22710 6656
rect 22741 6647 22799 6653
rect 22741 6613 22753 6647
rect 22787 6644 22799 6647
rect 23566 6644 23572 6656
rect 22787 6616 23572 6644
rect 22787 6613 22799 6616
rect 22741 6607 22799 6613
rect 23566 6604 23572 6616
rect 23624 6604 23630 6656
rect 26789 6647 26847 6653
rect 26789 6613 26801 6647
rect 26835 6644 26847 6647
rect 27890 6644 27896 6656
rect 26835 6616 27896 6644
rect 26835 6613 26847 6616
rect 26789 6607 26847 6613
rect 27890 6604 27896 6616
rect 27948 6604 27954 6656
rect 31036 6653 31064 6684
rect 31358 6681 31370 6684
rect 31404 6681 31416 6715
rect 31358 6675 31416 6681
rect 31021 6647 31079 6653
rect 31021 6613 31033 6647
rect 31067 6613 31079 6647
rect 31021 6607 31079 6613
rect 1104 6554 32844 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 32844 6554
rect 1104 6480 32844 6502
rect 10134 6400 10140 6452
rect 10192 6440 10198 6452
rect 14090 6440 14096 6452
rect 10192 6412 14096 6440
rect 10192 6400 10198 6412
rect 14090 6400 14096 6412
rect 14148 6400 14154 6452
rect 14182 6400 14188 6452
rect 14240 6400 14246 6452
rect 14553 6443 14611 6449
rect 14553 6409 14565 6443
rect 14599 6440 14611 6443
rect 14918 6440 14924 6452
rect 14599 6412 14924 6440
rect 14599 6409 14611 6412
rect 14553 6403 14611 6409
rect 14918 6400 14924 6412
rect 14976 6400 14982 6452
rect 15746 6400 15752 6452
rect 15804 6400 15810 6452
rect 18598 6400 18604 6452
rect 18656 6400 18662 6452
rect 22281 6443 22339 6449
rect 19306 6412 22232 6440
rect 2746 6344 11836 6372
rect 2590 6196 2596 6248
rect 2648 6236 2654 6248
rect 2746 6236 2774 6344
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6304 10655 6307
rect 10686 6304 10692 6316
rect 10643 6276 10692 6304
rect 10643 6273 10655 6276
rect 10597 6267 10655 6273
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 10796 6236 10824 6267
rect 11514 6264 11520 6316
rect 11572 6264 11578 6316
rect 11808 6304 11836 6344
rect 14200 6335 14228 6400
rect 19306 6372 19334 6412
rect 15672 6344 19334 6372
rect 14185 6329 14243 6335
rect 13906 6304 13912 6316
rect 11808 6276 13912 6304
rect 13906 6264 13912 6276
rect 13964 6264 13970 6316
rect 14185 6295 14197 6329
rect 14231 6295 14243 6329
rect 15672 6316 15700 6344
rect 14185 6289 14243 6295
rect 15102 6264 15108 6316
rect 15160 6304 15166 6316
rect 15381 6307 15439 6313
rect 15381 6304 15393 6307
rect 15160 6276 15393 6304
rect 15160 6264 15166 6276
rect 15381 6273 15393 6276
rect 15427 6273 15439 6307
rect 15381 6267 15439 6273
rect 15565 6307 15623 6313
rect 15565 6273 15577 6307
rect 15611 6304 15623 6307
rect 15654 6304 15660 6316
rect 15611 6276 15660 6304
rect 15611 6273 15623 6276
rect 15565 6267 15623 6273
rect 15654 6264 15660 6276
rect 15712 6264 15718 6316
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17126 6304 17132 6316
rect 17083 6276 17132 6304
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 17126 6264 17132 6276
rect 17184 6264 17190 6316
rect 17310 6264 17316 6316
rect 17368 6264 17374 6316
rect 17589 6307 17647 6313
rect 17589 6273 17601 6307
rect 17635 6273 17647 6307
rect 17589 6267 17647 6273
rect 2648 6208 2774 6236
rect 10612 6208 10824 6236
rect 2648 6196 2654 6208
rect 10612 6180 10640 6208
rect 11422 6196 11428 6248
rect 11480 6236 11486 6248
rect 11609 6239 11667 6245
rect 11609 6236 11621 6239
rect 11480 6208 11621 6236
rect 11480 6196 11486 6208
rect 11609 6205 11621 6208
rect 11655 6205 11667 6239
rect 11609 6199 11667 6205
rect 14277 6239 14335 6245
rect 14277 6205 14289 6239
rect 14323 6236 14335 6239
rect 15470 6236 15476 6248
rect 14323 6208 15476 6236
rect 14323 6205 14335 6208
rect 14277 6199 14335 6205
rect 15470 6196 15476 6208
rect 15528 6196 15534 6248
rect 17218 6196 17224 6248
rect 17276 6196 17282 6248
rect 10594 6128 10600 6180
rect 10652 6128 10658 6180
rect 11238 6128 11244 6180
rect 11296 6168 11302 6180
rect 17604 6168 17632 6267
rect 17770 6264 17776 6316
rect 17828 6304 17834 6316
rect 18892 6313 18920 6344
rect 19702 6332 19708 6384
rect 19760 6372 19766 6384
rect 19889 6375 19947 6381
rect 19889 6372 19901 6375
rect 19760 6344 19901 6372
rect 19760 6332 19766 6344
rect 19889 6341 19901 6344
rect 19935 6341 19947 6375
rect 19889 6335 19947 6341
rect 19978 6332 19984 6384
rect 20036 6372 20042 6384
rect 20036 6344 20208 6372
rect 20036 6332 20042 6344
rect 17865 6307 17923 6313
rect 17865 6304 17877 6307
rect 17828 6276 17877 6304
rect 17828 6264 17834 6276
rect 17865 6273 17877 6276
rect 17911 6273 17923 6307
rect 17865 6267 17923 6273
rect 18877 6307 18935 6313
rect 18877 6273 18889 6307
rect 18923 6273 18935 6307
rect 18877 6267 18935 6273
rect 18969 6307 19027 6313
rect 18969 6273 18981 6307
rect 19015 6304 19027 6307
rect 19015 6276 19104 6304
rect 19015 6273 19027 6276
rect 18969 6267 19027 6273
rect 17678 6196 17684 6248
rect 17736 6236 17742 6248
rect 18782 6236 18788 6248
rect 17736 6208 18788 6236
rect 17736 6196 17742 6208
rect 18782 6196 18788 6208
rect 18840 6196 18846 6248
rect 19076 6177 19104 6276
rect 19242 6264 19248 6316
rect 19300 6264 19306 6316
rect 19610 6264 19616 6316
rect 19668 6304 19674 6316
rect 20180 6313 20208 6344
rect 20714 6332 20720 6384
rect 20772 6372 20778 6384
rect 20901 6375 20959 6381
rect 20901 6372 20913 6375
rect 20772 6344 20913 6372
rect 20772 6332 20778 6344
rect 20901 6341 20913 6344
rect 20947 6341 20959 6375
rect 20901 6335 20959 6341
rect 21174 6332 21180 6384
rect 21232 6372 21238 6384
rect 22204 6372 22232 6412
rect 22281 6409 22293 6443
rect 22327 6440 22339 6443
rect 22554 6440 22560 6452
rect 22327 6412 22560 6440
rect 22327 6409 22339 6412
rect 22281 6403 22339 6409
rect 22554 6400 22560 6412
rect 22612 6400 22618 6452
rect 22741 6443 22799 6449
rect 22741 6409 22753 6443
rect 22787 6440 22799 6443
rect 23014 6440 23020 6452
rect 22787 6412 23020 6440
rect 22787 6409 22799 6412
rect 22741 6403 22799 6409
rect 23014 6400 23020 6412
rect 23072 6400 23078 6452
rect 23385 6443 23443 6449
rect 23385 6409 23397 6443
rect 23431 6440 23443 6443
rect 26418 6440 26424 6452
rect 23431 6412 26424 6440
rect 23431 6409 23443 6412
rect 23385 6403 23443 6409
rect 21232 6344 22140 6372
rect 22204 6344 22600 6372
rect 21232 6332 21238 6344
rect 20165 6307 20223 6313
rect 19668 6276 20116 6304
rect 19668 6264 19674 6276
rect 19518 6196 19524 6248
rect 19576 6236 19582 6248
rect 19981 6239 20039 6245
rect 19981 6236 19993 6239
rect 19576 6208 19993 6236
rect 19576 6196 19582 6208
rect 19981 6205 19993 6208
rect 20027 6205 20039 6239
rect 20088 6236 20116 6276
rect 20165 6273 20177 6307
rect 20211 6273 20223 6307
rect 20165 6267 20223 6273
rect 20530 6264 20536 6316
rect 20588 6304 20594 6316
rect 22112 6313 22140 6344
rect 21085 6307 21143 6313
rect 21085 6304 21097 6307
rect 20588 6276 21097 6304
rect 20588 6264 20594 6276
rect 21085 6273 21097 6276
rect 21131 6273 21143 6307
rect 21821 6307 21879 6313
rect 21821 6304 21833 6307
rect 21085 6267 21143 6273
rect 21192 6276 21833 6304
rect 21192 6236 21220 6276
rect 21821 6273 21833 6276
rect 21867 6273 21879 6307
rect 21821 6267 21879 6273
rect 22097 6307 22155 6313
rect 22097 6273 22109 6307
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 22370 6264 22376 6316
rect 22428 6264 22434 6316
rect 22572 6304 22600 6344
rect 22646 6332 22652 6384
rect 22704 6372 22710 6384
rect 22704 6344 23428 6372
rect 22704 6332 22710 6344
rect 22572 6276 23152 6304
rect 20088 6208 21220 6236
rect 21269 6239 21327 6245
rect 19981 6199 20039 6205
rect 21269 6205 21281 6239
rect 21315 6236 21327 6239
rect 21913 6239 21971 6245
rect 21913 6236 21925 6239
rect 21315 6208 21925 6236
rect 21315 6205 21327 6208
rect 21269 6199 21327 6205
rect 21913 6205 21925 6208
rect 21959 6236 21971 6239
rect 22465 6239 22523 6245
rect 21959 6208 22416 6236
rect 21959 6205 21971 6208
rect 21913 6199 21971 6205
rect 11296 6140 17632 6168
rect 19061 6171 19119 6177
rect 11296 6128 11302 6140
rect 19061 6137 19073 6171
rect 19107 6168 19119 6171
rect 20622 6168 20628 6180
rect 19107 6140 20628 6168
rect 19107 6137 19119 6140
rect 19061 6131 19119 6137
rect 20622 6128 20628 6140
rect 20680 6128 20686 6180
rect 10965 6103 11023 6109
rect 10965 6069 10977 6103
rect 11011 6100 11023 6103
rect 11330 6100 11336 6112
rect 11011 6072 11336 6100
rect 11011 6069 11023 6072
rect 10965 6063 11023 6069
rect 11330 6060 11336 6072
rect 11388 6060 11394 6112
rect 11698 6060 11704 6112
rect 11756 6060 11762 6112
rect 11885 6103 11943 6109
rect 11885 6069 11897 6103
rect 11931 6100 11943 6103
rect 11974 6100 11980 6112
rect 11931 6072 11980 6100
rect 11931 6069 11943 6072
rect 11885 6063 11943 6069
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 13998 6060 14004 6112
rect 14056 6100 14062 6112
rect 14185 6103 14243 6109
rect 14185 6100 14197 6103
rect 14056 6072 14197 6100
rect 14056 6060 14062 6072
rect 14185 6069 14197 6072
rect 14231 6069 14243 6103
rect 14185 6063 14243 6069
rect 15470 6060 15476 6112
rect 15528 6100 15534 6112
rect 17037 6103 17095 6109
rect 17037 6100 17049 6103
rect 15528 6072 17049 6100
rect 15528 6060 15534 6072
rect 17037 6069 17049 6072
rect 17083 6069 17095 6103
rect 17037 6063 17095 6069
rect 17494 6060 17500 6112
rect 17552 6060 17558 6112
rect 17770 6060 17776 6112
rect 17828 6060 17834 6112
rect 17862 6060 17868 6112
rect 17920 6100 17926 6112
rect 18049 6103 18107 6109
rect 18049 6100 18061 6103
rect 17920 6072 18061 6100
rect 17920 6060 17926 6072
rect 18049 6069 18061 6072
rect 18095 6069 18107 6103
rect 18049 6063 18107 6069
rect 18966 6060 18972 6112
rect 19024 6060 19030 6112
rect 20070 6060 20076 6112
rect 20128 6060 20134 6112
rect 20346 6060 20352 6112
rect 20404 6060 20410 6112
rect 22094 6060 22100 6112
rect 22152 6060 22158 6112
rect 22388 6109 22416 6208
rect 22465 6205 22477 6239
rect 22511 6236 22523 6239
rect 23014 6236 23020 6248
rect 22511 6208 23020 6236
rect 22511 6205 22523 6208
rect 22465 6199 22523 6205
rect 23014 6196 23020 6208
rect 23072 6196 23078 6248
rect 23124 6168 23152 6276
rect 23198 6264 23204 6316
rect 23256 6264 23262 6316
rect 23400 6236 23428 6344
rect 23492 6313 23520 6412
rect 26418 6400 26424 6412
rect 26476 6400 26482 6452
rect 26605 6443 26663 6449
rect 26605 6409 26617 6443
rect 26651 6440 26663 6443
rect 26970 6440 26976 6452
rect 26651 6412 26976 6440
rect 26651 6409 26663 6412
rect 26605 6403 26663 6409
rect 26970 6400 26976 6412
rect 27028 6400 27034 6452
rect 31662 6400 31668 6452
rect 31720 6440 31726 6452
rect 32401 6443 32459 6449
rect 32401 6440 32413 6443
rect 31720 6412 32413 6440
rect 31720 6400 31726 6412
rect 32401 6409 32413 6412
rect 32447 6409 32459 6443
rect 32401 6403 32459 6409
rect 24857 6375 24915 6381
rect 24857 6372 24869 6375
rect 24412 6344 24869 6372
rect 23477 6307 23535 6313
rect 23477 6273 23489 6307
rect 23523 6273 23535 6307
rect 23477 6267 23535 6273
rect 24412 6236 24440 6344
rect 24857 6341 24869 6344
rect 24903 6372 24915 6375
rect 24903 6344 26372 6372
rect 24903 6341 24915 6344
rect 24857 6335 24915 6341
rect 25038 6264 25044 6316
rect 25096 6264 25102 6316
rect 25222 6264 25228 6316
rect 25280 6304 25286 6316
rect 25317 6307 25375 6313
rect 25317 6304 25329 6307
rect 25280 6276 25329 6304
rect 25280 6264 25286 6276
rect 25317 6273 25329 6276
rect 25363 6273 25375 6307
rect 25317 6267 25375 6273
rect 25409 6307 25467 6313
rect 25409 6273 25421 6307
rect 25455 6304 25467 6307
rect 25774 6304 25780 6316
rect 25455 6276 25780 6304
rect 25455 6273 25467 6276
rect 25409 6267 25467 6273
rect 25774 6264 25780 6276
rect 25832 6264 25838 6316
rect 25958 6264 25964 6316
rect 26016 6264 26022 6316
rect 26344 6313 26372 6344
rect 26145 6307 26203 6313
rect 26145 6273 26157 6307
rect 26191 6273 26203 6307
rect 26145 6267 26203 6273
rect 26329 6307 26387 6313
rect 26329 6273 26341 6307
rect 26375 6273 26387 6307
rect 26329 6267 26387 6273
rect 26421 6307 26479 6313
rect 26421 6273 26433 6307
rect 26467 6304 26479 6307
rect 26510 6304 26516 6316
rect 26467 6276 26516 6304
rect 26467 6273 26479 6276
rect 26421 6267 26479 6273
rect 23400 6208 24440 6236
rect 25498 6196 25504 6248
rect 25556 6236 25562 6248
rect 26160 6236 26188 6267
rect 25556 6208 26188 6236
rect 25556 6196 25562 6208
rect 26436 6168 26464 6267
rect 26510 6264 26516 6276
rect 26568 6264 26574 6316
rect 32214 6264 32220 6316
rect 32272 6264 32278 6316
rect 23124 6140 26464 6168
rect 22373 6103 22431 6109
rect 22373 6069 22385 6103
rect 22419 6069 22431 6103
rect 22373 6063 22431 6069
rect 23382 6060 23388 6112
rect 23440 6100 23446 6112
rect 23661 6103 23719 6109
rect 23661 6100 23673 6103
rect 23440 6072 23673 6100
rect 23440 6060 23446 6072
rect 23661 6069 23673 6072
rect 23707 6100 23719 6103
rect 24302 6100 24308 6112
rect 23707 6072 24308 6100
rect 23707 6069 23719 6072
rect 23661 6063 23719 6069
rect 24302 6060 24308 6072
rect 24360 6060 24366 6112
rect 25222 6060 25228 6112
rect 25280 6060 25286 6112
rect 25314 6060 25320 6112
rect 25372 6060 25378 6112
rect 25682 6060 25688 6112
rect 25740 6060 25746 6112
rect 25958 6060 25964 6112
rect 26016 6100 26022 6112
rect 26145 6103 26203 6109
rect 26145 6100 26157 6103
rect 26016 6072 26157 6100
rect 26016 6060 26022 6072
rect 26145 6069 26157 6072
rect 26191 6069 26203 6103
rect 26145 6063 26203 6069
rect 1104 6010 32844 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 32844 6010
rect 1104 5936 32844 5958
rect 6825 5899 6883 5905
rect 6825 5865 6837 5899
rect 6871 5896 6883 5899
rect 8202 5896 8208 5908
rect 6871 5868 8208 5896
rect 6871 5865 6883 5868
rect 6825 5859 6883 5865
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 9398 5856 9404 5908
rect 9456 5896 9462 5908
rect 13541 5899 13599 5905
rect 9456 5868 13492 5896
rect 9456 5856 9462 5868
rect 8478 5788 8484 5840
rect 8536 5828 8542 5840
rect 9217 5831 9275 5837
rect 9217 5828 9229 5831
rect 8536 5800 9229 5828
rect 8536 5788 8542 5800
rect 9217 5797 9229 5800
rect 9263 5828 9275 5831
rect 11054 5828 11060 5840
rect 9263 5800 11060 5828
rect 9263 5797 9275 5800
rect 9217 5791 9275 5797
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 11514 5788 11520 5840
rect 11572 5828 11578 5840
rect 13262 5828 13268 5840
rect 11572 5800 13268 5828
rect 11572 5788 11578 5800
rect 13262 5788 13268 5800
rect 13320 5788 13326 5840
rect 13464 5828 13492 5868
rect 13541 5865 13553 5899
rect 13587 5896 13599 5899
rect 14182 5896 14188 5908
rect 13587 5868 14188 5896
rect 13587 5865 13599 5868
rect 13541 5859 13599 5865
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 14458 5856 14464 5908
rect 14516 5896 14522 5908
rect 14516 5868 15240 5896
rect 14516 5856 14522 5868
rect 15102 5828 15108 5840
rect 13464 5800 15108 5828
rect 15102 5788 15108 5800
rect 15160 5788 15166 5840
rect 15212 5828 15240 5868
rect 16666 5856 16672 5908
rect 16724 5896 16730 5908
rect 18046 5896 18052 5908
rect 16724 5868 18052 5896
rect 16724 5856 16730 5868
rect 18046 5856 18052 5868
rect 18104 5896 18110 5908
rect 18233 5899 18291 5905
rect 18233 5896 18245 5899
rect 18104 5868 18245 5896
rect 18104 5856 18110 5868
rect 18233 5865 18245 5868
rect 18279 5865 18291 5899
rect 18233 5859 18291 5865
rect 18693 5899 18751 5905
rect 18693 5865 18705 5899
rect 18739 5896 18751 5899
rect 19058 5896 19064 5908
rect 18739 5868 19064 5896
rect 18739 5865 18751 5868
rect 18693 5859 18751 5865
rect 19058 5856 19064 5868
rect 19116 5856 19122 5908
rect 20898 5896 20904 5908
rect 19306 5868 20904 5896
rect 19306 5828 19334 5868
rect 20898 5856 20904 5868
rect 20956 5856 20962 5908
rect 20990 5856 20996 5908
rect 21048 5896 21054 5908
rect 22370 5896 22376 5908
rect 21048 5868 22376 5896
rect 21048 5856 21054 5868
rect 22370 5856 22376 5868
rect 22428 5856 22434 5908
rect 23014 5856 23020 5908
rect 23072 5896 23078 5908
rect 23477 5899 23535 5905
rect 23477 5896 23489 5899
rect 23072 5868 23489 5896
rect 23072 5856 23078 5868
rect 23477 5865 23489 5868
rect 23523 5865 23535 5899
rect 23477 5859 23535 5865
rect 23937 5899 23995 5905
rect 23937 5865 23949 5899
rect 23983 5896 23995 5899
rect 24394 5896 24400 5908
rect 23983 5868 24400 5896
rect 23983 5865 23995 5868
rect 23937 5859 23995 5865
rect 24394 5856 24400 5868
rect 24452 5856 24458 5908
rect 15212 5800 19334 5828
rect 20346 5788 20352 5840
rect 20404 5828 20410 5840
rect 23290 5828 23296 5840
rect 20404 5800 23296 5828
rect 20404 5788 20410 5800
rect 23290 5788 23296 5800
rect 23348 5788 23354 5840
rect 25038 5828 25044 5840
rect 23584 5800 25044 5828
rect 5350 5720 5356 5772
rect 5408 5760 5414 5772
rect 5408 5732 9076 5760
rect 5408 5720 5414 5732
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 5592 5664 7236 5692
rect 5592 5652 5598 5664
rect 6917 5627 6975 5633
rect 6917 5593 6929 5627
rect 6963 5593 6975 5627
rect 6917 5587 6975 5593
rect 6932 5556 6960 5587
rect 7098 5584 7104 5636
rect 7156 5584 7162 5636
rect 7208 5624 7236 5664
rect 7374 5652 7380 5704
rect 7432 5652 7438 5704
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5692 8631 5695
rect 8662 5692 8668 5704
rect 8619 5664 8668 5692
rect 8619 5661 8631 5664
rect 8573 5655 8631 5661
rect 8128 5624 8156 5655
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 9048 5701 9076 5732
rect 9306 5720 9312 5772
rect 9364 5760 9370 5772
rect 11606 5760 11612 5772
rect 9364 5732 11612 5760
rect 9364 5720 9370 5732
rect 11606 5720 11612 5732
rect 11664 5720 11670 5772
rect 12526 5720 12532 5772
rect 12584 5760 12590 5772
rect 17126 5760 17132 5772
rect 12584 5732 17132 5760
rect 12584 5720 12590 5732
rect 17126 5720 17132 5732
rect 17184 5720 17190 5772
rect 17218 5720 17224 5772
rect 17276 5760 17282 5772
rect 17313 5763 17371 5769
rect 17313 5760 17325 5763
rect 17276 5732 17325 5760
rect 17276 5720 17282 5732
rect 17313 5729 17325 5732
rect 17359 5760 17371 5763
rect 18325 5763 18383 5769
rect 18325 5760 18337 5763
rect 17359 5732 18337 5760
rect 17359 5729 17371 5732
rect 17313 5723 17371 5729
rect 18325 5729 18337 5732
rect 18371 5729 18383 5763
rect 18325 5723 18383 5729
rect 18966 5720 18972 5772
rect 19024 5760 19030 5772
rect 23584 5760 23612 5800
rect 25038 5788 25044 5800
rect 25096 5788 25102 5840
rect 19024 5732 23612 5760
rect 23661 5763 23719 5769
rect 19024 5720 19030 5732
rect 23661 5729 23673 5763
rect 23707 5760 23719 5763
rect 25222 5760 25228 5772
rect 23707 5732 25228 5760
rect 23707 5729 23719 5732
rect 23661 5723 23719 5729
rect 25222 5720 25228 5732
rect 25280 5720 25286 5772
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5661 9091 5695
rect 9033 5655 9091 5661
rect 9122 5652 9128 5704
rect 9180 5692 9186 5704
rect 11238 5692 11244 5704
rect 9180 5664 11244 5692
rect 9180 5652 9186 5664
rect 11238 5652 11244 5664
rect 11296 5652 11302 5704
rect 12066 5652 12072 5704
rect 12124 5692 12130 5704
rect 15286 5692 15292 5704
rect 12124 5664 15292 5692
rect 12124 5652 12130 5664
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 18506 5652 18512 5704
rect 18564 5652 18570 5704
rect 18782 5652 18788 5704
rect 18840 5692 18846 5704
rect 20438 5692 20444 5704
rect 18840 5664 20444 5692
rect 18840 5652 18846 5664
rect 20438 5652 20444 5664
rect 20496 5692 20502 5704
rect 20990 5692 20996 5704
rect 20496 5664 20996 5692
rect 20496 5652 20502 5664
rect 20990 5652 20996 5664
rect 21048 5652 21054 5704
rect 23382 5652 23388 5704
rect 23440 5652 23446 5704
rect 23753 5695 23811 5701
rect 23753 5661 23765 5695
rect 23799 5692 23811 5695
rect 31754 5692 31760 5704
rect 23799 5664 31760 5692
rect 23799 5661 23811 5664
rect 23753 5655 23811 5661
rect 31754 5652 31760 5664
rect 31812 5652 31818 5704
rect 11422 5624 11428 5636
rect 7208 5596 8156 5624
rect 8220 5596 11428 5624
rect 7193 5559 7251 5565
rect 7193 5556 7205 5559
rect 6932 5528 7205 5556
rect 7193 5525 7205 5528
rect 7239 5556 7251 5559
rect 8220 5556 8248 5596
rect 11422 5584 11428 5596
rect 11480 5584 11486 5636
rect 11606 5584 11612 5636
rect 11664 5624 11670 5636
rect 13173 5627 13231 5633
rect 13173 5624 13185 5627
rect 11664 5596 13185 5624
rect 11664 5584 11670 5596
rect 13173 5593 13185 5596
rect 13219 5593 13231 5627
rect 13173 5587 13231 5593
rect 13357 5627 13415 5633
rect 13357 5593 13369 5627
rect 13403 5624 13415 5627
rect 13446 5624 13452 5636
rect 13403 5596 13452 5624
rect 13403 5593 13415 5596
rect 13357 5587 13415 5593
rect 13446 5584 13452 5596
rect 13504 5584 13510 5636
rect 16945 5627 17003 5633
rect 16945 5624 16957 5627
rect 13556 5596 16957 5624
rect 7239 5528 8248 5556
rect 7239 5525 7251 5528
rect 7193 5519 7251 5525
rect 8294 5516 8300 5568
rect 8352 5516 8358 5568
rect 8386 5516 8392 5568
rect 8444 5556 8450 5568
rect 11882 5556 11888 5568
rect 8444 5528 11888 5556
rect 8444 5516 8450 5528
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 13262 5516 13268 5568
rect 13320 5556 13326 5568
rect 13556 5556 13584 5596
rect 16945 5593 16957 5596
rect 16991 5624 17003 5627
rect 17034 5624 17040 5636
rect 16991 5596 17040 5624
rect 16991 5593 17003 5596
rect 16945 5587 17003 5593
rect 17034 5584 17040 5596
rect 17092 5584 17098 5636
rect 17129 5627 17187 5633
rect 17129 5593 17141 5627
rect 17175 5624 17187 5627
rect 17862 5624 17868 5636
rect 17175 5596 17868 5624
rect 17175 5593 17187 5596
rect 17129 5587 17187 5593
rect 13320 5528 13584 5556
rect 13320 5516 13326 5528
rect 14090 5516 14096 5568
rect 14148 5556 14154 5568
rect 14458 5556 14464 5568
rect 14148 5528 14464 5556
rect 14148 5516 14154 5528
rect 14458 5516 14464 5528
rect 14516 5556 14522 5568
rect 16666 5556 16672 5568
rect 14516 5528 16672 5556
rect 14516 5516 14522 5528
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 16758 5516 16764 5568
rect 16816 5556 16822 5568
rect 17144 5556 17172 5587
rect 17862 5584 17868 5596
rect 17920 5584 17926 5636
rect 18233 5627 18291 5633
rect 18233 5593 18245 5627
rect 18279 5624 18291 5627
rect 19610 5624 19616 5636
rect 18279 5596 19616 5624
rect 18279 5593 18291 5596
rect 18233 5587 18291 5593
rect 19610 5584 19616 5596
rect 19668 5584 19674 5636
rect 23198 5584 23204 5636
rect 23256 5584 23262 5636
rect 23474 5584 23480 5636
rect 23532 5584 23538 5636
rect 16816 5528 17172 5556
rect 16816 5516 16822 5528
rect 17218 5516 17224 5568
rect 17276 5556 17282 5568
rect 24578 5556 24584 5568
rect 17276 5528 24584 5556
rect 17276 5516 17282 5528
rect 24578 5516 24584 5528
rect 24636 5516 24642 5568
rect 1104 5466 32844 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 32844 5466
rect 1104 5392 32844 5414
rect 1302 5312 1308 5364
rect 1360 5352 1366 5364
rect 8665 5355 8723 5361
rect 8665 5352 8677 5355
rect 1360 5324 8677 5352
rect 1360 5312 1366 5324
rect 8665 5321 8677 5324
rect 8711 5321 8723 5355
rect 8665 5315 8723 5321
rect 12066 5312 12072 5364
rect 12124 5312 12130 5364
rect 21082 5352 21088 5364
rect 14200 5324 21088 5352
rect 8202 5244 8208 5296
rect 8260 5244 8266 5296
rect 8312 5256 8616 5284
rect 3234 5176 3240 5228
rect 3292 5216 3298 5228
rect 8312 5216 8340 5256
rect 3292 5188 8340 5216
rect 3292 5176 3298 5188
rect 8478 5176 8484 5228
rect 8536 5176 8542 5228
rect 8588 5216 8616 5256
rect 10962 5244 10968 5296
rect 11020 5284 11026 5296
rect 11609 5287 11667 5293
rect 11609 5284 11621 5287
rect 11020 5256 11621 5284
rect 11020 5244 11026 5256
rect 11609 5253 11621 5256
rect 11655 5253 11667 5287
rect 14200 5284 14228 5324
rect 21082 5312 21088 5324
rect 21140 5312 21146 5364
rect 23109 5355 23167 5361
rect 23109 5321 23121 5355
rect 23155 5352 23167 5355
rect 23198 5352 23204 5364
rect 23155 5324 23204 5352
rect 23155 5321 23167 5324
rect 23109 5315 23167 5321
rect 23198 5312 23204 5324
rect 23256 5312 23262 5364
rect 31570 5352 31576 5364
rect 24596 5324 31576 5352
rect 11609 5247 11667 5253
rect 11808 5256 14228 5284
rect 11808 5216 11836 5256
rect 14366 5244 14372 5296
rect 14424 5284 14430 5296
rect 16114 5284 16120 5296
rect 14424 5256 16120 5284
rect 14424 5244 14430 5256
rect 8588 5188 11836 5216
rect 11882 5176 11888 5228
rect 11940 5176 11946 5228
rect 14274 5216 14280 5228
rect 14200 5188 14280 5216
rect 8294 5108 8300 5160
rect 8352 5148 8358 5160
rect 8389 5151 8447 5157
rect 8389 5148 8401 5151
rect 8352 5120 8401 5148
rect 8352 5108 8358 5120
rect 8389 5117 8401 5120
rect 8435 5148 8447 5151
rect 9582 5148 9588 5160
rect 8435 5120 9588 5148
rect 8435 5117 8447 5120
rect 8389 5111 8447 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 11330 5108 11336 5160
rect 11388 5148 11394 5160
rect 11701 5151 11759 5157
rect 11701 5148 11713 5151
rect 11388 5120 11713 5148
rect 11388 5108 11394 5120
rect 11701 5117 11713 5120
rect 11747 5117 11759 5151
rect 11701 5111 11759 5117
rect 8018 5040 8024 5092
rect 8076 5080 8082 5092
rect 8076 5052 8524 5080
rect 8076 5040 8082 5052
rect 8386 4972 8392 5024
rect 8444 4972 8450 5024
rect 8496 5012 8524 5052
rect 10042 5040 10048 5092
rect 10100 5080 10106 5092
rect 14200 5089 14228 5188
rect 14274 5176 14280 5188
rect 14332 5176 14338 5228
rect 14458 5176 14464 5228
rect 14516 5176 14522 5228
rect 14568 5225 14596 5256
rect 16114 5244 16120 5256
rect 16172 5284 16178 5296
rect 18049 5287 18107 5293
rect 18049 5284 18061 5287
rect 16172 5256 18061 5284
rect 16172 5244 16178 5256
rect 18049 5253 18061 5256
rect 18095 5253 18107 5287
rect 18049 5247 18107 5253
rect 23845 5287 23903 5293
rect 23845 5253 23857 5287
rect 23891 5284 23903 5287
rect 23891 5256 24155 5284
rect 23891 5253 23903 5256
rect 23845 5247 23903 5253
rect 14553 5219 14611 5225
rect 14553 5185 14565 5219
rect 14599 5185 14611 5219
rect 14553 5179 14611 5185
rect 14829 5219 14887 5225
rect 14829 5185 14841 5219
rect 14875 5216 14887 5219
rect 15010 5216 15016 5228
rect 14875 5188 15016 5216
rect 14875 5185 14887 5188
rect 14829 5179 14887 5185
rect 15010 5176 15016 5188
rect 15068 5176 15074 5228
rect 18325 5219 18383 5225
rect 18325 5185 18337 5219
rect 18371 5216 18383 5219
rect 18506 5216 18512 5228
rect 18371 5188 18512 5216
rect 18371 5185 18383 5188
rect 18325 5179 18383 5185
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 23566 5176 23572 5228
rect 23624 5176 23630 5228
rect 23750 5176 23756 5228
rect 23808 5176 23814 5228
rect 23934 5176 23940 5228
rect 23992 5176 23998 5228
rect 24127 5216 24155 5256
rect 24210 5216 24216 5228
rect 24127 5188 24216 5216
rect 24210 5176 24216 5188
rect 24268 5176 24274 5228
rect 24397 5219 24455 5225
rect 24397 5216 24409 5219
rect 24320 5188 24409 5216
rect 15746 5108 15752 5160
rect 15804 5148 15810 5160
rect 16022 5148 16028 5160
rect 15804 5120 16028 5148
rect 15804 5108 15810 5120
rect 16022 5108 16028 5120
rect 16080 5108 16086 5160
rect 18138 5108 18144 5160
rect 18196 5108 18202 5160
rect 24320 5148 24348 5188
rect 24397 5185 24409 5188
rect 24443 5185 24455 5219
rect 24397 5179 24455 5185
rect 24486 5176 24492 5228
rect 24544 5176 24550 5228
rect 24596 5216 24624 5324
rect 31570 5312 31576 5324
rect 31628 5312 31634 5364
rect 24673 5287 24731 5293
rect 24673 5253 24685 5287
rect 24719 5284 24731 5287
rect 30374 5284 30380 5296
rect 24719 5256 30380 5284
rect 24719 5253 24731 5256
rect 24673 5247 24731 5253
rect 30374 5244 30380 5256
rect 30432 5244 30438 5296
rect 24765 5219 24823 5225
rect 24765 5216 24777 5219
rect 24596 5188 24777 5216
rect 24765 5185 24777 5188
rect 24811 5185 24823 5219
rect 24765 5179 24823 5185
rect 24857 5219 24915 5225
rect 24857 5185 24869 5219
rect 24903 5216 24915 5219
rect 25133 5219 25191 5225
rect 25133 5216 25145 5219
rect 24903 5188 25145 5216
rect 24903 5185 24915 5188
rect 24857 5179 24915 5185
rect 25133 5185 25145 5188
rect 25179 5185 25191 5219
rect 29822 5216 29828 5228
rect 25133 5179 25191 5185
rect 25608 5188 29828 5216
rect 25608 5148 25636 5188
rect 29822 5176 29828 5188
rect 29880 5176 29886 5228
rect 24320 5120 25636 5148
rect 25682 5108 25688 5160
rect 25740 5108 25746 5160
rect 14185 5083 14243 5089
rect 10100 5052 11744 5080
rect 10100 5040 10106 5052
rect 11609 5015 11667 5021
rect 11609 5012 11621 5015
rect 8496 4984 11621 5012
rect 11609 4981 11621 4984
rect 11655 4981 11667 5015
rect 11716 5012 11744 5052
rect 14185 5049 14197 5083
rect 14231 5049 14243 5083
rect 14185 5043 14243 5049
rect 14642 5040 14648 5092
rect 14700 5040 14706 5092
rect 18509 5083 18567 5089
rect 18509 5049 18521 5083
rect 18555 5080 18567 5083
rect 18555 5052 24348 5080
rect 18555 5049 18567 5052
rect 18509 5043 18567 5049
rect 14366 5012 14372 5024
rect 11716 4984 14372 5012
rect 11609 4975 11667 4981
rect 14366 4972 14372 4984
rect 14424 4972 14430 5024
rect 14553 5015 14611 5021
rect 14553 4981 14565 5015
rect 14599 5012 14611 5015
rect 16206 5012 16212 5024
rect 14599 4984 16212 5012
rect 14599 4981 14611 4984
rect 14553 4975 14611 4981
rect 16206 4972 16212 4984
rect 16264 4972 16270 5024
rect 18046 4972 18052 5024
rect 18104 4972 18110 5024
rect 24118 4972 24124 5024
rect 24176 4972 24182 5024
rect 24210 4972 24216 5024
rect 24268 4972 24274 5024
rect 24320 5012 24348 5052
rect 24762 5012 24768 5024
rect 24320 4984 24768 5012
rect 24762 4972 24768 4984
rect 24820 4972 24826 5024
rect 24946 4972 24952 5024
rect 25004 5012 25010 5024
rect 25041 5015 25099 5021
rect 25041 5012 25053 5015
rect 25004 4984 25053 5012
rect 25004 4972 25010 4984
rect 25041 4981 25053 4984
rect 25087 4981 25099 5015
rect 25041 4975 25099 4981
rect 1104 4922 32844 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 32844 4922
rect 1104 4848 32844 4870
rect 12345 4811 12403 4817
rect 12345 4777 12357 4811
rect 12391 4777 12403 4811
rect 14458 4808 14464 4820
rect 12345 4771 12403 4777
rect 12452 4780 14464 4808
rect 9582 4632 9588 4684
rect 9640 4672 9646 4684
rect 12253 4675 12311 4681
rect 12253 4672 12265 4675
rect 9640 4644 12265 4672
rect 9640 4632 9646 4644
rect 9950 4564 9956 4616
rect 10008 4564 10014 4616
rect 10152 4613 10180 4644
rect 12253 4641 12265 4644
rect 12299 4641 12311 4675
rect 12253 4635 12311 4641
rect 10137 4607 10195 4613
rect 10137 4573 10149 4607
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4604 10379 4607
rect 10962 4604 10968 4616
rect 10367 4576 10968 4604
rect 10367 4573 10379 4576
rect 10321 4567 10379 4573
rect 10962 4564 10968 4576
rect 11020 4604 11026 4616
rect 12161 4607 12219 4613
rect 12161 4604 12173 4607
rect 11020 4576 12173 4604
rect 11020 4564 11026 4576
rect 12161 4573 12173 4576
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 12360 4536 12388 4771
rect 12452 4613 12480 4780
rect 14458 4768 14464 4780
rect 14516 4768 14522 4820
rect 14553 4811 14611 4817
rect 14553 4777 14565 4811
rect 14599 4808 14611 4811
rect 14642 4808 14648 4820
rect 14599 4780 14648 4808
rect 14599 4777 14611 4780
rect 14553 4771 14611 4777
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 14734 4768 14740 4820
rect 14792 4768 14798 4820
rect 15856 4780 16068 4808
rect 12618 4700 12624 4752
rect 12676 4700 12682 4752
rect 12989 4743 13047 4749
rect 12989 4709 13001 4743
rect 13035 4709 13047 4743
rect 12989 4703 13047 4709
rect 13004 4672 13032 4703
rect 14366 4700 14372 4752
rect 14424 4740 14430 4752
rect 15856 4740 15884 4780
rect 14424 4712 15884 4740
rect 16040 4740 16068 4780
rect 16114 4768 16120 4820
rect 16172 4768 16178 4820
rect 16298 4768 16304 4820
rect 16356 4768 16362 4820
rect 26234 4808 26240 4820
rect 22066 4780 26240 4808
rect 22066 4740 22094 4780
rect 26234 4768 26240 4780
rect 26292 4768 26298 4820
rect 16040 4712 22094 4740
rect 14424 4700 14430 4712
rect 22462 4700 22468 4752
rect 22520 4740 22526 4752
rect 22833 4743 22891 4749
rect 22833 4740 22845 4743
rect 22520 4712 22845 4740
rect 22520 4700 22526 4712
rect 22833 4709 22845 4712
rect 22879 4709 22891 4743
rect 22833 4703 22891 4709
rect 23753 4743 23811 4749
rect 23753 4709 23765 4743
rect 23799 4709 23811 4743
rect 24397 4743 24455 4749
rect 24397 4740 24409 4743
rect 23753 4703 23811 4709
rect 23952 4712 24409 4740
rect 15746 4672 15752 4684
rect 13004 4644 15752 4672
rect 12437 4607 12495 4613
rect 12437 4573 12449 4607
rect 12483 4573 12495 4607
rect 12437 4567 12495 4573
rect 12802 4564 12808 4616
rect 12860 4564 12866 4616
rect 13004 4536 13032 4644
rect 14384 4613 14412 4644
rect 15746 4632 15752 4644
rect 15804 4672 15810 4684
rect 15933 4675 15991 4681
rect 15804 4644 15884 4672
rect 15804 4632 15810 4644
rect 14369 4607 14427 4613
rect 14369 4573 14381 4607
rect 14415 4573 14427 4607
rect 14369 4567 14427 4573
rect 14550 4564 14556 4616
rect 14608 4564 14614 4616
rect 14642 4564 14648 4616
rect 14700 4604 14706 4616
rect 15856 4613 15884 4644
rect 15933 4641 15945 4675
rect 15979 4641 15991 4675
rect 23768 4672 23796 4703
rect 15933 4635 15991 4641
rect 21008 4644 23796 4672
rect 15841 4607 15899 4613
rect 14700 4576 15792 4604
rect 14700 4564 14706 4576
rect 12360 4508 13032 4536
rect 15764 4536 15792 4576
rect 15841 4573 15853 4607
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 15948 4536 15976 4635
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4604 16175 4607
rect 16206 4604 16212 4616
rect 16163 4576 16212 4604
rect 16163 4573 16175 4576
rect 16117 4567 16175 4573
rect 16206 4564 16212 4576
rect 16264 4604 16270 4616
rect 18138 4604 18144 4616
rect 16264 4576 18144 4604
rect 16264 4564 16270 4576
rect 18138 4564 18144 4576
rect 18196 4564 18202 4616
rect 19702 4564 19708 4616
rect 19760 4604 19766 4616
rect 19797 4607 19855 4613
rect 19797 4604 19809 4607
rect 19760 4576 19809 4604
rect 19760 4564 19766 4576
rect 19797 4573 19809 4576
rect 19843 4573 19855 4607
rect 19797 4567 19855 4573
rect 20806 4564 20812 4616
rect 20864 4564 20870 4616
rect 21008 4548 21036 4644
rect 21174 4564 21180 4616
rect 21232 4564 21238 4616
rect 22186 4564 22192 4616
rect 22244 4604 22250 4616
rect 22480 4613 22508 4644
rect 22281 4607 22339 4613
rect 22281 4604 22293 4607
rect 22244 4576 22293 4604
rect 22244 4564 22250 4576
rect 22281 4573 22293 4576
rect 22327 4573 22339 4607
rect 22281 4567 22339 4573
rect 22465 4607 22523 4613
rect 22465 4573 22477 4607
rect 22511 4573 22523 4607
rect 22465 4567 22523 4573
rect 22649 4607 22707 4613
rect 22649 4573 22661 4607
rect 22695 4604 22707 4607
rect 23017 4607 23075 4613
rect 23017 4604 23029 4607
rect 22695 4576 23029 4604
rect 22695 4573 22707 4576
rect 22649 4567 22707 4573
rect 23017 4573 23029 4576
rect 23063 4573 23075 4607
rect 23017 4567 23075 4573
rect 23566 4564 23572 4616
rect 23624 4564 23630 4616
rect 23750 4564 23756 4616
rect 23808 4604 23814 4616
rect 23952 4613 23980 4712
rect 24397 4709 24409 4712
rect 24443 4709 24455 4743
rect 24397 4703 24455 4709
rect 23937 4607 23995 4613
rect 23937 4604 23949 4607
rect 23808 4576 23949 4604
rect 23808 4564 23814 4576
rect 23937 4573 23949 4576
rect 23983 4573 23995 4607
rect 23937 4567 23995 4573
rect 24210 4564 24216 4616
rect 24268 4564 24274 4616
rect 24578 4564 24584 4616
rect 24636 4564 24642 4616
rect 24854 4564 24860 4616
rect 24912 4564 24918 4616
rect 24946 4564 24952 4616
rect 25004 4604 25010 4616
rect 25113 4607 25171 4613
rect 25113 4604 25125 4607
rect 25004 4576 25125 4604
rect 25004 4564 25010 4576
rect 25113 4573 25125 4576
rect 25159 4573 25171 4607
rect 25113 4567 25171 4573
rect 15764 4508 15976 4536
rect 20990 4496 20996 4548
rect 21048 4496 21054 4548
rect 21082 4496 21088 4548
rect 21140 4536 21146 4548
rect 22557 4539 22615 4545
rect 21140 4508 22094 4536
rect 21140 4496 21146 4508
rect 18506 4428 18512 4480
rect 18564 4468 18570 4480
rect 19245 4471 19303 4477
rect 19245 4468 19257 4471
rect 18564 4440 19257 4468
rect 18564 4428 18570 4440
rect 19245 4437 19257 4440
rect 19291 4437 19303 4471
rect 19245 4431 19303 4437
rect 21358 4428 21364 4480
rect 21416 4428 21422 4480
rect 22066 4468 22094 4508
rect 22557 4505 22569 4539
rect 22603 4536 22615 4539
rect 24872 4536 24900 4564
rect 26142 4536 26148 4548
rect 22603 4508 24072 4536
rect 24872 4508 26148 4536
rect 22603 4505 22615 4508
rect 22557 4499 22615 4505
rect 22572 4468 22600 4499
rect 24044 4477 24072 4508
rect 26142 4496 26148 4508
rect 26200 4496 26206 4548
rect 22066 4440 22600 4468
rect 24029 4471 24087 4477
rect 24029 4437 24041 4471
rect 24075 4437 24087 4471
rect 24029 4431 24087 4437
rect 25682 4428 25688 4480
rect 25740 4468 25746 4480
rect 26237 4471 26295 4477
rect 26237 4468 26249 4471
rect 25740 4440 26249 4468
rect 25740 4428 25746 4440
rect 26237 4437 26249 4440
rect 26283 4437 26295 4471
rect 26237 4431 26295 4437
rect 1104 4378 32844 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 32844 4378
rect 1104 4304 32844 4326
rect 1118 4224 1124 4276
rect 1176 4264 1182 4276
rect 12802 4264 12808 4276
rect 1176 4236 12808 4264
rect 1176 4224 1182 4236
rect 12802 4224 12808 4236
rect 12860 4224 12866 4276
rect 18877 4267 18935 4273
rect 18877 4233 18889 4267
rect 18923 4264 18935 4267
rect 19702 4264 19708 4276
rect 18923 4236 19708 4264
rect 18923 4233 18935 4236
rect 18877 4227 18935 4233
rect 19702 4224 19708 4236
rect 19760 4224 19766 4276
rect 21174 4224 21180 4276
rect 21232 4264 21238 4276
rect 21545 4267 21603 4273
rect 21545 4264 21557 4267
rect 21232 4236 21557 4264
rect 21232 4224 21238 4236
rect 21545 4233 21557 4236
rect 21591 4233 21603 4267
rect 21545 4227 21603 4233
rect 23934 4224 23940 4276
rect 23992 4264 23998 4276
rect 25317 4267 25375 4273
rect 25317 4264 25329 4267
rect 23992 4236 25329 4264
rect 23992 4224 23998 4236
rect 25317 4233 25329 4236
rect 25363 4233 25375 4267
rect 25317 4227 25375 4233
rect 22296 4168 22600 4196
rect 2406 4088 2412 4140
rect 2464 4128 2470 4140
rect 16574 4128 16580 4140
rect 2464 4100 16580 4128
rect 2464 4088 2470 4100
rect 16574 4088 16580 4100
rect 16632 4088 16638 4140
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 16925 4131 16983 4137
rect 16925 4128 16937 4131
rect 16816 4100 16937 4128
rect 16816 4088 16822 4100
rect 16925 4097 16937 4100
rect 16971 4097 16983 4131
rect 16925 4091 16983 4097
rect 18782 4088 18788 4140
rect 18840 4128 18846 4140
rect 19990 4131 20048 4137
rect 19990 4128 20002 4131
rect 18840 4100 20002 4128
rect 18840 4088 18846 4100
rect 19990 4097 20002 4100
rect 20036 4097 20048 4131
rect 19990 4091 20048 4097
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4128 20315 4131
rect 21910 4128 21916 4140
rect 20303 4100 21916 4128
rect 20303 4097 20315 4100
rect 20257 4091 20315 4097
rect 21910 4088 21916 4100
rect 21968 4128 21974 4140
rect 22189 4131 22247 4137
rect 22189 4128 22201 4131
rect 21968 4100 22201 4128
rect 21968 4088 21974 4100
rect 22189 4097 22201 4100
rect 22235 4128 22247 4131
rect 22296 4128 22324 4168
rect 22462 4137 22468 4140
rect 22456 4128 22468 4137
rect 22235 4100 22324 4128
rect 22423 4100 22468 4128
rect 22235 4097 22247 4100
rect 22189 4091 22247 4097
rect 22456 4091 22468 4100
rect 22462 4088 22468 4091
rect 22520 4088 22526 4140
rect 22572 4128 22600 4168
rect 23952 4168 24256 4196
rect 23845 4131 23903 4137
rect 23845 4128 23857 4131
rect 22572 4100 23857 4128
rect 23845 4097 23857 4100
rect 23891 4128 23903 4131
rect 23952 4128 23980 4168
rect 24118 4137 24124 4140
rect 24112 4128 24124 4137
rect 23891 4100 23980 4128
rect 24079 4100 24124 4128
rect 23891 4097 23903 4100
rect 23845 4091 23903 4097
rect 24112 4091 24124 4100
rect 24118 4088 24124 4091
rect 24176 4088 24182 4140
rect 24228 4128 24256 4168
rect 24854 4128 24860 4140
rect 24228 4100 24860 4128
rect 24854 4088 24860 4100
rect 24912 4088 24918 4140
rect 16669 4063 16727 4069
rect 16669 4029 16681 4063
rect 16715 4029 16727 4063
rect 16669 4023 16727 4029
rect 16684 3924 16712 4023
rect 20898 4020 20904 4072
rect 20956 4020 20962 4072
rect 25222 4020 25228 4072
rect 25280 4060 25286 4072
rect 25866 4060 25872 4072
rect 25280 4032 25872 4060
rect 25280 4020 25286 4032
rect 25866 4020 25872 4032
rect 25924 4020 25930 4072
rect 18233 3995 18291 4001
rect 18233 3992 18245 3995
rect 17604 3964 18245 3992
rect 17604 3924 17632 3964
rect 18233 3961 18245 3964
rect 18279 3992 18291 3995
rect 31018 3992 31024 4004
rect 18279 3964 19012 3992
rect 18279 3961 18291 3964
rect 18233 3955 18291 3961
rect 16684 3896 17632 3924
rect 17678 3884 17684 3936
rect 17736 3924 17742 3936
rect 18049 3927 18107 3933
rect 18049 3924 18061 3927
rect 17736 3896 18061 3924
rect 17736 3884 17742 3896
rect 18049 3893 18061 3896
rect 18095 3893 18107 3927
rect 18984 3924 19012 3964
rect 20272 3964 22094 3992
rect 20272 3924 20300 3964
rect 18984 3896 20300 3924
rect 22066 3924 22094 3964
rect 23124 3964 23888 3992
rect 23124 3924 23152 3964
rect 22066 3896 23152 3924
rect 18049 3887 18107 3893
rect 23566 3884 23572 3936
rect 23624 3884 23630 3936
rect 23860 3924 23888 3964
rect 24780 3964 31024 3992
rect 24780 3924 24808 3964
rect 31018 3952 31024 3964
rect 31076 3952 31082 4004
rect 23860 3896 24808 3924
rect 25222 3884 25228 3936
rect 25280 3884 25286 3936
rect 1104 3834 32844 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 32844 3834
rect 1104 3760 32844 3782
rect 10226 3680 10232 3732
rect 10284 3720 10290 3732
rect 31386 3720 31392 3732
rect 10284 3692 31392 3720
rect 10284 3680 10290 3692
rect 31386 3680 31392 3692
rect 31444 3680 31450 3732
rect 16758 3612 16764 3664
rect 16816 3612 16822 3664
rect 18782 3612 18788 3664
rect 18840 3612 18846 3664
rect 16482 3584 16488 3596
rect 16408 3556 16488 3584
rect 16408 3525 16436 3556
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 17497 3587 17555 3593
rect 17497 3553 17509 3587
rect 17543 3584 17555 3587
rect 17678 3584 17684 3596
rect 17543 3556 17684 3584
rect 17543 3553 17555 3556
rect 17497 3547 17555 3553
rect 17678 3544 17684 3556
rect 17736 3544 17742 3596
rect 18340 3556 18644 3584
rect 16209 3519 16267 3525
rect 16209 3485 16221 3519
rect 16255 3485 16267 3519
rect 16209 3479 16267 3485
rect 16393 3519 16451 3525
rect 16393 3485 16405 3519
rect 16439 3485 16451 3519
rect 16393 3479 16451 3485
rect 16577 3519 16635 3525
rect 16577 3485 16589 3519
rect 16623 3516 16635 3519
rect 16853 3519 16911 3525
rect 16853 3516 16865 3519
rect 16623 3488 16865 3516
rect 16623 3485 16635 3488
rect 16577 3479 16635 3485
rect 16853 3485 16865 3488
rect 16899 3485 16911 3519
rect 16853 3479 16911 3485
rect 16224 3380 16252 3479
rect 18230 3476 18236 3528
rect 18288 3476 18294 3528
rect 16485 3451 16543 3457
rect 16485 3417 16497 3451
rect 16531 3448 16543 3451
rect 18340 3448 18368 3556
rect 18506 3476 18512 3528
rect 18564 3476 18570 3528
rect 18616 3525 18644 3556
rect 21910 3544 21916 3596
rect 21968 3544 21974 3596
rect 18601 3519 18659 3525
rect 18601 3485 18613 3519
rect 18647 3516 18659 3519
rect 21082 3516 21088 3528
rect 18647 3488 21088 3516
rect 18647 3485 18659 3488
rect 18601 3479 18659 3485
rect 21082 3476 21088 3488
rect 21140 3476 21146 3528
rect 21358 3476 21364 3528
rect 21416 3516 21422 3528
rect 21646 3519 21704 3525
rect 21646 3516 21658 3519
rect 21416 3488 21658 3516
rect 21416 3476 21422 3488
rect 21646 3485 21658 3488
rect 21692 3485 21704 3519
rect 21646 3479 21704 3485
rect 16531 3420 18368 3448
rect 18417 3451 18475 3457
rect 16531 3417 16543 3420
rect 16485 3411 16543 3417
rect 18417 3417 18429 3451
rect 18463 3448 18475 3451
rect 20990 3448 20996 3460
rect 18463 3420 20996 3448
rect 18463 3417 18475 3420
rect 18417 3411 18475 3417
rect 18432 3380 18460 3411
rect 20990 3408 20996 3420
rect 21048 3408 21054 3460
rect 16224 3352 18460 3380
rect 20533 3383 20591 3389
rect 20533 3349 20545 3383
rect 20579 3380 20591 3383
rect 20898 3380 20904 3392
rect 20579 3352 20904 3380
rect 20579 3349 20591 3352
rect 20533 3343 20591 3349
rect 20898 3340 20904 3352
rect 20956 3380 20962 3392
rect 21358 3380 21364 3392
rect 20956 3352 21364 3380
rect 20956 3340 20962 3352
rect 21358 3340 21364 3352
rect 21416 3340 21422 3392
rect 1104 3290 32844 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 32844 3290
rect 1104 3216 32844 3238
rect 16574 3136 16580 3188
rect 16632 3176 16638 3188
rect 28442 3176 28448 3188
rect 16632 3148 28448 3176
rect 16632 3136 16638 3148
rect 28442 3136 28448 3148
rect 28500 3136 28506 3188
rect 5810 3068 5816 3120
rect 5868 3108 5874 3120
rect 28074 3108 28080 3120
rect 5868 3080 28080 3108
rect 5868 3068 5874 3080
rect 28074 3068 28080 3080
rect 28132 3068 28138 3120
rect 1104 2746 32844 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 32844 2746
rect 1104 2672 32844 2694
rect 17678 2388 17684 2440
rect 17736 2428 17742 2440
rect 17773 2431 17831 2437
rect 17773 2428 17785 2431
rect 17736 2400 17785 2428
rect 17736 2388 17742 2400
rect 17773 2397 17785 2400
rect 17819 2397 17831 2431
rect 17773 2391 17831 2397
rect 19702 2388 19708 2440
rect 19760 2388 19766 2440
rect 21358 2388 21364 2440
rect 21416 2388 21422 2440
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2428 22983 2431
rect 23566 2428 23572 2440
rect 22971 2400 23572 2428
rect 22971 2397 22983 2400
rect 22925 2391 22983 2397
rect 23566 2388 23572 2400
rect 23624 2388 23630 2440
rect 24857 2431 24915 2437
rect 24857 2397 24869 2431
rect 24903 2428 24915 2431
rect 25682 2428 25688 2440
rect 24903 2400 25688 2428
rect 24903 2397 24915 2400
rect 24857 2391 24915 2397
rect 25682 2388 25688 2400
rect 25740 2388 25746 2440
rect 25866 2388 25872 2440
rect 25924 2388 25930 2440
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29696 2400 29745 2428
rect 29696 2388 29702 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17589 2295 17647 2301
rect 17589 2292 17601 2295
rect 17460 2264 17601 2292
rect 17460 2252 17466 2264
rect 17589 2261 17601 2264
rect 17635 2261 17647 2295
rect 17589 2255 17647 2261
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 19521 2295 19579 2301
rect 19521 2292 19533 2295
rect 19392 2264 19533 2292
rect 19392 2252 19398 2264
rect 19521 2261 19533 2264
rect 19567 2261 19579 2295
rect 19521 2255 19579 2261
rect 21266 2252 21272 2304
rect 21324 2292 21330 2304
rect 21545 2295 21603 2301
rect 21545 2292 21557 2295
rect 21324 2264 21557 2292
rect 21324 2252 21330 2264
rect 21545 2261 21557 2264
rect 21591 2261 21603 2295
rect 21545 2255 21603 2261
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22741 2295 22799 2301
rect 22741 2292 22753 2295
rect 22612 2264 22753 2292
rect 22612 2252 22618 2264
rect 22741 2261 22753 2264
rect 22787 2261 22799 2295
rect 22741 2255 22799 2261
rect 24486 2252 24492 2304
rect 24544 2292 24550 2304
rect 24673 2295 24731 2301
rect 24673 2292 24685 2295
rect 24544 2264 24685 2292
rect 24544 2252 24550 2264
rect 24673 2261 24685 2264
rect 24719 2261 24731 2295
rect 24673 2255 24731 2261
rect 25774 2252 25780 2304
rect 25832 2292 25838 2304
rect 26053 2295 26111 2301
rect 26053 2292 26065 2295
rect 25832 2264 26065 2292
rect 25832 2252 25838 2264
rect 26053 2261 26065 2264
rect 26099 2261 26111 2295
rect 26053 2255 26111 2261
rect 1104 2202 32844 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 32844 2202
rect 1104 2128 32844 2150
<< via1 >>
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 18696 31424 18748 31476
rect 21272 31424 21324 31476
rect 25136 31424 25188 31476
rect 16764 31356 16816 31408
rect 23204 31356 23256 31408
rect 17132 31288 17184 31340
rect 19340 31331 19392 31340
rect 19340 31297 19349 31331
rect 19349 31297 19383 31331
rect 19383 31297 19392 31331
rect 19340 31288 19392 31297
rect 21916 31331 21968 31340
rect 21916 31297 21925 31331
rect 21925 31297 21959 31331
rect 21959 31297 21968 31331
rect 21916 31288 21968 31297
rect 23664 31331 23716 31340
rect 23664 31297 23673 31331
rect 23673 31297 23707 31331
rect 23707 31297 23716 31331
rect 23664 31288 23716 31297
rect 25320 31331 25372 31340
rect 25320 31297 25329 31331
rect 25329 31297 25363 31331
rect 25363 31297 25372 31331
rect 25320 31288 25372 31297
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 13452 30744 13504 30796
rect 26976 30744 27028 30796
rect 1308 30540 1360 30592
rect 18512 30676 18564 30728
rect 14832 30608 14884 30660
rect 32312 30608 32364 30660
rect 14096 30540 14148 30592
rect 28264 30540 28316 30592
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 6092 30336 6144 30388
rect 14096 30336 14148 30388
rect 21916 30336 21968 30388
rect 17316 30200 17368 30252
rect 18696 30200 18748 30252
rect 19340 30200 19392 30252
rect 20536 30243 20588 30252
rect 20536 30209 20570 30243
rect 20570 30209 20588 30243
rect 20536 30200 20588 30209
rect 26148 30200 26200 30252
rect 940 29996 992 30048
rect 10692 29996 10744 30048
rect 18880 30039 18932 30048
rect 18880 30005 18889 30039
rect 18889 30005 18923 30039
rect 18923 30005 18932 30039
rect 18880 29996 18932 30005
rect 20628 29996 20680 30048
rect 20904 29996 20956 30048
rect 22192 29996 22244 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 1216 29792 1268 29844
rect 8852 29792 8904 29844
rect 9864 29792 9916 29844
rect 17132 29792 17184 29844
rect 1032 29724 1084 29776
rect 7196 29724 7248 29776
rect 9404 29724 9456 29776
rect 11704 29724 11756 29776
rect 5632 29656 5684 29708
rect 3240 29631 3292 29640
rect 3240 29597 3249 29631
rect 3249 29597 3283 29631
rect 3283 29597 3292 29631
rect 3240 29588 3292 29597
rect 7012 29588 7064 29640
rect 17316 29699 17368 29708
rect 17316 29665 17325 29699
rect 17325 29665 17359 29699
rect 17359 29665 17368 29699
rect 17316 29656 17368 29665
rect 18696 29835 18748 29844
rect 18696 29801 18705 29835
rect 18705 29801 18739 29835
rect 18739 29801 18748 29835
rect 18696 29792 18748 29801
rect 20536 29792 20588 29844
rect 23664 29792 23716 29844
rect 20628 29656 20680 29708
rect 9128 29520 9180 29572
rect 3332 29452 3384 29504
rect 3424 29495 3476 29504
rect 3424 29461 3433 29495
rect 3433 29461 3467 29495
rect 3467 29461 3476 29495
rect 3424 29452 3476 29461
rect 5264 29452 5316 29504
rect 10232 29520 10284 29572
rect 10692 29588 10744 29640
rect 16580 29588 16632 29640
rect 17500 29588 17552 29640
rect 18880 29588 18932 29640
rect 20904 29631 20956 29640
rect 20904 29597 20913 29631
rect 20913 29597 20947 29631
rect 20947 29597 20956 29631
rect 20904 29588 20956 29597
rect 17224 29520 17276 29572
rect 10508 29452 10560 29504
rect 16856 29452 16908 29504
rect 17408 29495 17460 29504
rect 17408 29461 17417 29495
rect 17417 29461 17451 29495
rect 17451 29461 17460 29495
rect 17408 29452 17460 29461
rect 18420 29563 18472 29572
rect 18420 29529 18429 29563
rect 18429 29529 18463 29563
rect 18463 29529 18472 29563
rect 18420 29520 18472 29529
rect 21272 29631 21324 29640
rect 21272 29597 21281 29631
rect 21281 29597 21315 29631
rect 21315 29597 21324 29631
rect 21272 29588 21324 29597
rect 22468 29520 22520 29572
rect 24492 29520 24544 29572
rect 25780 29631 25832 29640
rect 25780 29597 25789 29631
rect 25789 29597 25823 29631
rect 25823 29597 25832 29631
rect 25780 29588 25832 29597
rect 29000 29520 29052 29572
rect 22100 29452 22152 29504
rect 22192 29452 22244 29504
rect 22376 29452 22428 29504
rect 25320 29452 25372 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 1400 29155 1452 29164
rect 1400 29121 1409 29155
rect 1409 29121 1443 29155
rect 1443 29121 1452 29155
rect 1400 29112 1452 29121
rect 3516 29248 3568 29300
rect 2780 29180 2832 29232
rect 3056 29112 3108 29164
rect 3424 29180 3476 29232
rect 2228 29044 2280 29096
rect 4344 29112 4396 29164
rect 4712 29155 4764 29164
rect 4712 29121 4721 29155
rect 4721 29121 4755 29155
rect 4755 29121 4764 29155
rect 4712 29112 4764 29121
rect 4620 29044 4672 29096
rect 2872 28976 2924 29028
rect 7196 29155 7248 29164
rect 7196 29121 7205 29155
rect 7205 29121 7239 29155
rect 7239 29121 7248 29155
rect 7196 29112 7248 29121
rect 7472 29155 7524 29164
rect 7472 29121 7481 29155
rect 7481 29121 7515 29155
rect 7515 29121 7524 29155
rect 7472 29112 7524 29121
rect 7564 29112 7616 29164
rect 1676 28908 1728 28960
rect 2964 28908 3016 28960
rect 3148 28908 3200 28960
rect 3792 28951 3844 28960
rect 3792 28917 3801 28951
rect 3801 28917 3835 28951
rect 3835 28917 3844 28951
rect 3792 28908 3844 28917
rect 3884 28908 3936 28960
rect 4252 28908 4304 28960
rect 4896 28951 4948 28960
rect 4896 28917 4905 28951
rect 4905 28917 4939 28951
rect 4939 28917 4948 28951
rect 4896 28908 4948 28917
rect 4988 28951 5040 28960
rect 4988 28917 4997 28951
rect 4997 28917 5031 28951
rect 5031 28917 5040 28951
rect 4988 28908 5040 28917
rect 5448 28951 5500 28960
rect 5448 28917 5457 28951
rect 5457 28917 5491 28951
rect 5491 28917 5500 28951
rect 5448 28908 5500 28917
rect 6736 28976 6788 29028
rect 8024 29155 8076 29164
rect 8024 29121 8033 29155
rect 8033 29121 8067 29155
rect 8067 29121 8076 29155
rect 8024 29112 8076 29121
rect 8852 29155 8904 29164
rect 8852 29121 8861 29155
rect 8861 29121 8895 29155
rect 8895 29121 8904 29155
rect 8852 29112 8904 29121
rect 9128 29291 9180 29300
rect 9128 29257 9137 29291
rect 9137 29257 9171 29291
rect 9171 29257 9180 29291
rect 9128 29248 9180 29257
rect 9680 29291 9732 29300
rect 9680 29257 9689 29291
rect 9689 29257 9723 29291
rect 9723 29257 9732 29291
rect 9680 29248 9732 29257
rect 9772 29248 9824 29300
rect 9036 29180 9088 29232
rect 9404 29155 9456 29164
rect 9404 29121 9413 29155
rect 9413 29121 9447 29155
rect 9447 29121 9456 29155
rect 9404 29112 9456 29121
rect 8668 29044 8720 29096
rect 9772 29112 9824 29164
rect 9864 29155 9916 29164
rect 9864 29121 9873 29155
rect 9873 29121 9907 29155
rect 9907 29121 9916 29155
rect 9864 29112 9916 29121
rect 10048 29180 10100 29232
rect 10600 29112 10652 29164
rect 9680 29044 9732 29096
rect 10968 29112 11020 29164
rect 15936 29291 15988 29300
rect 15936 29257 15945 29291
rect 15945 29257 15979 29291
rect 15979 29257 15988 29291
rect 15936 29248 15988 29257
rect 16396 29248 16448 29300
rect 8392 28976 8444 29028
rect 12716 29155 12768 29164
rect 12716 29121 12725 29155
rect 12725 29121 12759 29155
rect 12759 29121 12768 29155
rect 12716 29112 12768 29121
rect 13268 29112 13320 29164
rect 16856 29223 16908 29232
rect 16856 29189 16865 29223
rect 16865 29189 16899 29223
rect 16899 29189 16908 29223
rect 16856 29180 16908 29189
rect 18420 29180 18472 29232
rect 22468 29291 22520 29300
rect 22468 29257 22477 29291
rect 22477 29257 22511 29291
rect 22511 29257 22520 29291
rect 22468 29248 22520 29257
rect 24492 29291 24544 29300
rect 24492 29257 24501 29291
rect 24501 29257 24535 29291
rect 24535 29257 24544 29291
rect 24492 29248 24544 29257
rect 16304 29112 16356 29164
rect 17408 29112 17460 29164
rect 11152 29044 11204 29096
rect 22100 29223 22152 29232
rect 22100 29189 22109 29223
rect 22109 29189 22143 29223
rect 22143 29189 22152 29223
rect 22100 29180 22152 29189
rect 20168 29155 20220 29164
rect 20168 29121 20177 29155
rect 20177 29121 20211 29155
rect 20211 29121 20220 29155
rect 20168 29112 20220 29121
rect 21916 29155 21968 29164
rect 21916 29121 21925 29155
rect 21925 29121 21959 29155
rect 21959 29121 21968 29155
rect 21916 29112 21968 29121
rect 22192 29155 22244 29164
rect 22192 29121 22201 29155
rect 22201 29121 22235 29155
rect 22235 29121 22244 29155
rect 22192 29112 22244 29121
rect 22376 29112 22428 29164
rect 11244 29019 11296 29028
rect 11244 28985 11253 29019
rect 11253 28985 11287 29019
rect 11287 28985 11296 29019
rect 11244 28976 11296 28985
rect 12072 28976 12124 29028
rect 12900 28976 12952 29028
rect 17224 29019 17276 29028
rect 17224 28985 17233 29019
rect 17233 28985 17267 29019
rect 17267 28985 17276 29019
rect 17224 28976 17276 28985
rect 18144 29019 18196 29028
rect 18144 28985 18153 29019
rect 18153 28985 18187 29019
rect 18187 28985 18196 29019
rect 18144 28976 18196 28985
rect 23756 29044 23808 29096
rect 29920 29180 29972 29232
rect 25320 29112 25372 29164
rect 24400 29044 24452 29096
rect 5908 28908 5960 28960
rect 7104 28908 7156 28960
rect 8208 28908 8260 28960
rect 9220 28951 9272 28960
rect 9220 28917 9229 28951
rect 9229 28917 9263 28951
rect 9263 28917 9272 28951
rect 9220 28908 9272 28917
rect 9864 28908 9916 28960
rect 10692 28908 10744 28960
rect 10784 28908 10836 28960
rect 11520 28951 11572 28960
rect 11520 28917 11529 28951
rect 11529 28917 11563 28951
rect 11563 28917 11572 28951
rect 11520 28908 11572 28917
rect 11980 28951 12032 28960
rect 11980 28917 11989 28951
rect 11989 28917 12023 28951
rect 12023 28917 12032 28951
rect 11980 28908 12032 28917
rect 12808 28908 12860 28960
rect 15844 28908 15896 28960
rect 18420 28951 18472 28960
rect 18420 28917 18429 28951
rect 18429 28917 18463 28951
rect 18463 28917 18472 28951
rect 18420 28908 18472 28917
rect 30380 28976 30432 29028
rect 19616 28908 19668 28960
rect 19892 28908 19944 28960
rect 23756 28908 23808 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 2872 28704 2924 28756
rect 4068 28704 4120 28756
rect 4344 28704 4396 28756
rect 4896 28704 4948 28756
rect 5816 28704 5868 28756
rect 8024 28704 8076 28756
rect 4620 28636 4672 28688
rect 5356 28679 5408 28688
rect 5356 28645 5365 28679
rect 5365 28645 5399 28679
rect 5399 28645 5408 28679
rect 5356 28636 5408 28645
rect 3148 28611 3200 28620
rect 3148 28577 3157 28611
rect 3157 28577 3191 28611
rect 3191 28577 3200 28611
rect 3148 28568 3200 28577
rect 4804 28568 4856 28620
rect 4988 28568 5040 28620
rect 1400 28543 1452 28552
rect 1400 28509 1409 28543
rect 1409 28509 1443 28543
rect 1443 28509 1452 28543
rect 1400 28500 1452 28509
rect 1676 28543 1728 28552
rect 1676 28509 1710 28543
rect 1710 28509 1728 28543
rect 1676 28500 1728 28509
rect 2504 28500 2556 28552
rect 3332 28543 3384 28552
rect 3332 28509 3341 28543
rect 3341 28509 3375 28543
rect 3375 28509 3384 28543
rect 3332 28500 3384 28509
rect 2964 28432 3016 28484
rect 2320 28364 2372 28416
rect 2688 28364 2740 28416
rect 3700 28432 3752 28484
rect 4252 28543 4304 28552
rect 4252 28509 4261 28543
rect 4261 28509 4295 28543
rect 4295 28509 4304 28543
rect 4252 28500 4304 28509
rect 4344 28543 4396 28552
rect 4344 28509 4353 28543
rect 4353 28509 4387 28543
rect 4387 28509 4396 28543
rect 4344 28500 4396 28509
rect 3332 28364 3384 28416
rect 4068 28407 4120 28416
rect 4068 28373 4077 28407
rect 4077 28373 4111 28407
rect 4111 28373 4120 28407
rect 5816 28611 5868 28620
rect 5816 28577 5825 28611
rect 5825 28577 5859 28611
rect 5859 28577 5868 28611
rect 5816 28568 5868 28577
rect 5908 28611 5960 28620
rect 5908 28577 5917 28611
rect 5917 28577 5951 28611
rect 5951 28577 5960 28611
rect 5908 28568 5960 28577
rect 6644 28568 6696 28620
rect 10416 28704 10468 28756
rect 10784 28704 10836 28756
rect 12440 28704 12492 28756
rect 12532 28747 12584 28756
rect 12532 28713 12541 28747
rect 12541 28713 12575 28747
rect 12575 28713 12584 28747
rect 12532 28704 12584 28713
rect 12716 28704 12768 28756
rect 8576 28636 8628 28688
rect 4068 28364 4120 28373
rect 4528 28407 4580 28416
rect 4528 28373 4537 28407
rect 4537 28373 4571 28407
rect 4571 28373 4580 28407
rect 4528 28364 4580 28373
rect 4620 28407 4672 28416
rect 4620 28373 4629 28407
rect 4629 28373 4663 28407
rect 4663 28373 4672 28407
rect 4620 28364 4672 28373
rect 6000 28500 6052 28552
rect 6736 28500 6788 28552
rect 7104 28500 7156 28552
rect 7196 28543 7248 28552
rect 7196 28509 7205 28543
rect 7205 28509 7239 28543
rect 7239 28509 7248 28543
rect 7196 28500 7248 28509
rect 5724 28432 5776 28484
rect 8208 28500 8260 28552
rect 8300 28543 8352 28552
rect 8300 28509 8309 28543
rect 8309 28509 8343 28543
rect 8343 28509 8352 28543
rect 8300 28500 8352 28509
rect 9220 28568 9272 28620
rect 8760 28500 8812 28552
rect 11152 28636 11204 28688
rect 11888 28679 11940 28688
rect 11888 28645 11897 28679
rect 11897 28645 11931 28679
rect 11931 28645 11940 28679
rect 11888 28636 11940 28645
rect 12072 28636 12124 28688
rect 9772 28543 9824 28552
rect 9772 28509 9781 28543
rect 9781 28509 9815 28543
rect 9815 28509 9824 28543
rect 9772 28500 9824 28509
rect 10508 28543 10560 28552
rect 10508 28509 10517 28543
rect 10517 28509 10551 28543
rect 10551 28509 10560 28543
rect 10508 28500 10560 28509
rect 10784 28543 10836 28552
rect 10784 28509 10793 28543
rect 10793 28509 10827 28543
rect 10827 28509 10836 28543
rect 10784 28500 10836 28509
rect 10876 28543 10928 28552
rect 10876 28509 10885 28543
rect 10885 28509 10919 28543
rect 10919 28509 10928 28543
rect 10876 28500 10928 28509
rect 11428 28500 11480 28552
rect 11520 28543 11572 28552
rect 11520 28509 11529 28543
rect 11529 28509 11563 28543
rect 11563 28509 11572 28543
rect 11520 28500 11572 28509
rect 11980 28543 12032 28552
rect 11980 28509 11989 28543
rect 11989 28509 12023 28543
rect 12023 28509 12032 28543
rect 11980 28500 12032 28509
rect 12348 28543 12400 28552
rect 12348 28509 12357 28543
rect 12357 28509 12391 28543
rect 12391 28509 12400 28543
rect 12348 28500 12400 28509
rect 12716 28568 12768 28620
rect 13176 28636 13228 28688
rect 12900 28543 12952 28552
rect 12900 28509 12909 28543
rect 12909 28509 12943 28543
rect 12943 28509 12952 28543
rect 12900 28500 12952 28509
rect 12992 28543 13044 28552
rect 12992 28509 13001 28543
rect 13001 28509 13035 28543
rect 13035 28509 13044 28543
rect 12992 28500 13044 28509
rect 16028 28704 16080 28756
rect 17316 28704 17368 28756
rect 19432 28704 19484 28756
rect 19892 28747 19944 28756
rect 19892 28713 19901 28747
rect 19901 28713 19935 28747
rect 19935 28713 19944 28747
rect 19892 28704 19944 28713
rect 19984 28704 20036 28756
rect 13912 28636 13964 28688
rect 17960 28636 18012 28688
rect 13544 28568 13596 28620
rect 18236 28568 18288 28620
rect 14280 28543 14332 28552
rect 6644 28407 6696 28416
rect 6644 28373 6653 28407
rect 6653 28373 6687 28407
rect 6687 28373 6696 28407
rect 6644 28364 6696 28373
rect 7196 28364 7248 28416
rect 7472 28364 7524 28416
rect 7748 28364 7800 28416
rect 8300 28364 8352 28416
rect 9036 28364 9088 28416
rect 9588 28432 9640 28484
rect 10140 28432 10192 28484
rect 9404 28364 9456 28416
rect 9956 28407 10008 28416
rect 9956 28373 9965 28407
rect 9965 28373 9999 28407
rect 9999 28373 10008 28407
rect 9956 28364 10008 28373
rect 11060 28407 11112 28416
rect 11060 28373 11069 28407
rect 11069 28373 11103 28407
rect 11103 28373 11112 28407
rect 11060 28364 11112 28373
rect 11612 28475 11664 28484
rect 11612 28441 11621 28475
rect 11621 28441 11655 28475
rect 11655 28441 11664 28475
rect 11612 28432 11664 28441
rect 11980 28364 12032 28416
rect 12532 28432 12584 28484
rect 14280 28509 14289 28543
rect 14289 28509 14323 28543
rect 14323 28509 14332 28543
rect 14280 28500 14332 28509
rect 14556 28543 14608 28552
rect 14556 28509 14565 28543
rect 14565 28509 14599 28543
rect 14599 28509 14608 28543
rect 14556 28500 14608 28509
rect 15292 28500 15344 28552
rect 12440 28364 12492 28416
rect 14096 28407 14148 28416
rect 14096 28373 14105 28407
rect 14105 28373 14139 28407
rect 14139 28373 14148 28407
rect 15844 28475 15896 28484
rect 15844 28441 15853 28475
rect 15853 28441 15887 28475
rect 15887 28441 15896 28475
rect 15844 28432 15896 28441
rect 16028 28475 16080 28484
rect 16028 28441 16037 28475
rect 16037 28441 16071 28475
rect 16071 28441 16080 28475
rect 16028 28432 16080 28441
rect 16396 28500 16448 28552
rect 17316 28475 17368 28484
rect 17316 28441 17325 28475
rect 17325 28441 17359 28475
rect 17359 28441 17368 28475
rect 17316 28432 17368 28441
rect 18052 28500 18104 28552
rect 18420 28636 18472 28688
rect 19340 28636 19392 28688
rect 18420 28500 18472 28552
rect 20168 28568 20220 28620
rect 20352 28636 20404 28688
rect 21732 28568 21784 28620
rect 20536 28543 20588 28552
rect 20536 28509 20545 28543
rect 20545 28509 20579 28543
rect 20579 28509 20588 28543
rect 20536 28500 20588 28509
rect 23204 28543 23256 28552
rect 23204 28509 23213 28543
rect 23213 28509 23247 28543
rect 23247 28509 23256 28543
rect 23204 28500 23256 28509
rect 23388 28543 23440 28552
rect 23388 28509 23397 28543
rect 23397 28509 23431 28543
rect 23431 28509 23440 28543
rect 23388 28500 23440 28509
rect 23756 28543 23808 28552
rect 23756 28509 23765 28543
rect 23765 28509 23799 28543
rect 23799 28509 23808 28543
rect 23756 28500 23808 28509
rect 24492 28500 24544 28552
rect 14096 28364 14148 28373
rect 14464 28364 14516 28416
rect 15016 28364 15068 28416
rect 16212 28407 16264 28416
rect 16212 28373 16221 28407
rect 16221 28373 16255 28407
rect 16255 28373 16264 28407
rect 16212 28364 16264 28373
rect 17684 28407 17736 28416
rect 17684 28373 17693 28407
rect 17693 28373 17727 28407
rect 17727 28373 17736 28407
rect 17684 28364 17736 28373
rect 18236 28432 18288 28484
rect 23480 28432 23532 28484
rect 29092 28432 29144 28484
rect 18972 28364 19024 28416
rect 19432 28364 19484 28416
rect 19984 28364 20036 28416
rect 20168 28407 20220 28416
rect 20168 28373 20177 28407
rect 20177 28373 20211 28407
rect 20211 28373 20220 28407
rect 20168 28364 20220 28373
rect 23572 28407 23624 28416
rect 23572 28373 23581 28407
rect 23581 28373 23615 28407
rect 23615 28373 23624 28407
rect 23572 28364 23624 28373
rect 23940 28364 23992 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 3240 28160 3292 28212
rect 5356 28203 5408 28212
rect 5356 28169 5365 28203
rect 5365 28169 5399 28203
rect 5399 28169 5408 28203
rect 5356 28160 5408 28169
rect 3332 28135 3384 28144
rect 3332 28101 3341 28135
rect 3341 28101 3375 28135
rect 3375 28101 3384 28135
rect 3332 28092 3384 28101
rect 3792 28092 3844 28144
rect 4344 28092 4396 28144
rect 4804 28092 4856 28144
rect 1676 28067 1728 28076
rect 1676 28033 1710 28067
rect 1710 28033 1728 28067
rect 1676 28024 1728 28033
rect 3148 28024 3200 28076
rect 4252 28024 4304 28076
rect 5448 28067 5500 28076
rect 5448 28033 5457 28067
rect 5457 28033 5491 28067
rect 5491 28033 5500 28067
rect 5448 28024 5500 28033
rect 6644 28160 6696 28212
rect 6184 28067 6236 28076
rect 6184 28033 6193 28067
rect 6193 28033 6227 28067
rect 6227 28033 6236 28067
rect 6184 28024 6236 28033
rect 6460 28024 6512 28076
rect 6644 28067 6696 28076
rect 6644 28033 6653 28067
rect 6653 28033 6687 28067
rect 6687 28033 6696 28067
rect 6644 28024 6696 28033
rect 7196 28160 7248 28212
rect 8392 28160 8444 28212
rect 9772 28160 9824 28212
rect 9864 28160 9916 28212
rect 11060 28160 11112 28212
rect 1400 27999 1452 28008
rect 1400 27965 1409 27999
rect 1409 27965 1443 27999
rect 1443 27965 1452 27999
rect 1400 27956 1452 27965
rect 2964 27956 3016 28008
rect 3240 27956 3292 28008
rect 7564 28092 7616 28144
rect 4068 27888 4120 27940
rect 4620 27888 4672 27940
rect 4988 27888 5040 27940
rect 6000 27888 6052 27940
rect 7196 28067 7248 28076
rect 7196 28033 7205 28067
rect 7205 28033 7239 28067
rect 7239 28033 7248 28067
rect 7196 28024 7248 28033
rect 7472 28067 7524 28076
rect 7472 28033 7481 28067
rect 7481 28033 7515 28067
rect 7515 28033 7524 28067
rect 7472 28024 7524 28033
rect 7748 28067 7800 28076
rect 7748 28033 7757 28067
rect 7757 28033 7791 28067
rect 7791 28033 7800 28067
rect 7748 28024 7800 28033
rect 8024 28067 8076 28076
rect 8024 28033 8033 28067
rect 8033 28033 8067 28067
rect 8067 28033 8076 28067
rect 8024 28024 8076 28033
rect 8668 28092 8720 28144
rect 8760 28135 8812 28144
rect 8760 28101 8769 28135
rect 8769 28101 8803 28135
rect 8803 28101 8812 28135
rect 8760 28092 8812 28101
rect 9404 28092 9456 28144
rect 9588 28092 9640 28144
rect 8576 28067 8628 28076
rect 8576 28033 8585 28067
rect 8585 28033 8619 28067
rect 8619 28033 8628 28067
rect 8576 28024 8628 28033
rect 9036 28024 9088 28076
rect 9496 28067 9548 28076
rect 9496 28033 9505 28067
rect 9505 28033 9539 28067
rect 9539 28033 9548 28067
rect 9496 28024 9548 28033
rect 9864 28024 9916 28076
rect 10048 28067 10100 28076
rect 10048 28033 10057 28067
rect 10057 28033 10091 28067
rect 10091 28033 10100 28067
rect 10048 28024 10100 28033
rect 11244 28092 11296 28144
rect 7104 27956 7156 28008
rect 7564 27956 7616 28008
rect 10232 27956 10284 28008
rect 8668 27888 8720 27940
rect 9128 27931 9180 27940
rect 9128 27897 9137 27931
rect 9137 27897 9171 27931
rect 9171 27897 9180 27931
rect 9128 27888 9180 27897
rect 3608 27820 3660 27872
rect 5816 27820 5868 27872
rect 6920 27863 6972 27872
rect 6920 27829 6929 27863
rect 6929 27829 6963 27863
rect 6963 27829 6972 27863
rect 6920 27820 6972 27829
rect 7840 27820 7892 27872
rect 8760 27820 8812 27872
rect 9680 27888 9732 27940
rect 10140 27888 10192 27940
rect 10784 28067 10836 28076
rect 10784 28033 10793 28067
rect 10793 28033 10827 28067
rect 10827 28033 10836 28067
rect 10784 28024 10836 28033
rect 11152 28067 11204 28076
rect 11152 28033 11161 28067
rect 11161 28033 11195 28067
rect 11195 28033 11204 28067
rect 11152 28024 11204 28033
rect 11428 28160 11480 28212
rect 12532 28160 12584 28212
rect 12992 28160 13044 28212
rect 13360 28160 13412 28212
rect 14556 28160 14608 28212
rect 22376 28160 22428 28212
rect 11520 28024 11572 28076
rect 9312 27863 9364 27872
rect 9312 27829 9321 27863
rect 9321 27829 9355 27863
rect 9355 27829 9364 27863
rect 9312 27820 9364 27829
rect 9588 27863 9640 27872
rect 9588 27829 9597 27863
rect 9597 27829 9631 27863
rect 9631 27829 9640 27863
rect 9588 27820 9640 27829
rect 10416 27820 10468 27872
rect 11244 27956 11296 28008
rect 14280 28092 14332 28144
rect 12532 28067 12584 28076
rect 12532 28033 12541 28067
rect 12541 28033 12575 28067
rect 12575 28033 12584 28067
rect 12532 28024 12584 28033
rect 12716 28024 12768 28076
rect 14096 28024 14148 28076
rect 12808 27956 12860 28008
rect 13728 27956 13780 28008
rect 14832 28067 14884 28076
rect 14832 28033 14841 28067
rect 14841 28033 14875 28067
rect 14875 28033 14884 28067
rect 14832 28024 14884 28033
rect 15016 28067 15068 28076
rect 15016 28033 15025 28067
rect 15025 28033 15059 28067
rect 15059 28033 15068 28067
rect 15016 28024 15068 28033
rect 15108 28024 15160 28076
rect 16580 28024 16632 28076
rect 18328 28092 18380 28144
rect 19156 28024 19208 28076
rect 19616 28024 19668 28076
rect 20260 28092 20312 28144
rect 20536 28024 20588 28076
rect 22284 28067 22336 28076
rect 22284 28033 22293 28067
rect 22293 28033 22327 28067
rect 22327 28033 22336 28067
rect 22284 28024 22336 28033
rect 22560 28067 22612 28076
rect 22560 28033 22569 28067
rect 22569 28033 22603 28067
rect 22603 28033 22612 28067
rect 22560 28024 22612 28033
rect 23296 28135 23348 28144
rect 23296 28101 23305 28135
rect 23305 28101 23339 28135
rect 23339 28101 23348 28135
rect 23296 28092 23348 28101
rect 25596 28135 25648 28144
rect 25596 28101 25605 28135
rect 25605 28101 25639 28135
rect 25639 28101 25648 28135
rect 25596 28092 25648 28101
rect 23756 28024 23808 28076
rect 24860 28067 24912 28076
rect 24860 28033 24869 28067
rect 24869 28033 24903 28067
rect 24903 28033 24912 28067
rect 24860 28024 24912 28033
rect 25504 28024 25556 28076
rect 15292 27956 15344 28008
rect 16672 27956 16724 28008
rect 11428 27888 11480 27940
rect 10876 27820 10928 27872
rect 12164 27863 12216 27872
rect 12164 27829 12173 27863
rect 12173 27829 12207 27863
rect 12207 27829 12216 27863
rect 12164 27820 12216 27829
rect 12256 27863 12308 27872
rect 12256 27829 12265 27863
rect 12265 27829 12299 27863
rect 12299 27829 12308 27863
rect 12256 27820 12308 27829
rect 12808 27863 12860 27872
rect 12808 27829 12817 27863
rect 12817 27829 12851 27863
rect 12851 27829 12860 27863
rect 12808 27820 12860 27829
rect 12992 27820 13044 27872
rect 13544 27820 13596 27872
rect 13912 27863 13964 27872
rect 13912 27829 13921 27863
rect 13921 27829 13955 27863
rect 13955 27829 13964 27863
rect 13912 27820 13964 27829
rect 14372 27820 14424 27872
rect 14464 27820 14516 27872
rect 14648 27820 14700 27872
rect 16856 27820 16908 27872
rect 18144 27956 18196 28008
rect 19248 27956 19300 28008
rect 20352 27956 20404 28008
rect 22100 27999 22152 28008
rect 22100 27965 22109 27999
rect 22109 27965 22143 27999
rect 22143 27965 22152 27999
rect 22100 27956 22152 27965
rect 24768 27956 24820 28008
rect 17776 27888 17828 27940
rect 21732 27888 21784 27940
rect 21824 27931 21876 27940
rect 21824 27897 21833 27931
rect 21833 27897 21867 27931
rect 21867 27897 21876 27931
rect 21824 27888 21876 27897
rect 17960 27820 18012 27872
rect 18604 27863 18656 27872
rect 18604 27829 18613 27863
rect 18613 27829 18647 27863
rect 18647 27829 18656 27863
rect 18604 27820 18656 27829
rect 19892 27820 19944 27872
rect 20444 27820 20496 27872
rect 23388 27863 23440 27872
rect 23388 27829 23397 27863
rect 23397 27829 23431 27863
rect 23431 27829 23440 27863
rect 23388 27820 23440 27829
rect 25596 27888 25648 27940
rect 24768 27820 24820 27872
rect 25136 27863 25188 27872
rect 25136 27829 25145 27863
rect 25145 27829 25179 27863
rect 25179 27829 25188 27863
rect 25136 27820 25188 27829
rect 25320 27863 25372 27872
rect 25320 27829 25329 27863
rect 25329 27829 25363 27863
rect 25363 27829 25372 27863
rect 25320 27820 25372 27829
rect 25504 27863 25556 27872
rect 25504 27829 25513 27863
rect 25513 27829 25547 27863
rect 25547 27829 25556 27863
rect 25504 27820 25556 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 1676 27616 1728 27668
rect 4804 27616 4856 27668
rect 5172 27616 5224 27668
rect 7288 27659 7340 27668
rect 7288 27625 7297 27659
rect 7297 27625 7331 27659
rect 7331 27625 7340 27659
rect 7288 27616 7340 27625
rect 7380 27659 7432 27668
rect 7380 27625 7389 27659
rect 7389 27625 7423 27659
rect 7423 27625 7432 27659
rect 7380 27616 7432 27625
rect 7840 27616 7892 27668
rect 2228 27591 2280 27600
rect 2228 27557 2237 27591
rect 2237 27557 2271 27591
rect 2271 27557 2280 27591
rect 2228 27548 2280 27557
rect 2504 27523 2556 27532
rect 2504 27489 2513 27523
rect 2513 27489 2547 27523
rect 2547 27489 2556 27523
rect 2504 27480 2556 27489
rect 2964 27548 3016 27600
rect 2872 27523 2924 27532
rect 2872 27489 2881 27523
rect 2881 27489 2915 27523
rect 2915 27489 2924 27523
rect 2872 27480 2924 27489
rect 3700 27548 3752 27600
rect 4068 27548 4120 27600
rect 3332 27523 3384 27532
rect 3332 27489 3366 27523
rect 3366 27489 3384 27523
rect 3332 27480 3384 27489
rect 1492 27412 1544 27464
rect 3056 27412 3108 27464
rect 4252 27412 4304 27464
rect 4988 27548 5040 27600
rect 5632 27591 5684 27600
rect 5632 27557 5641 27591
rect 5641 27557 5675 27591
rect 5675 27557 5684 27591
rect 5632 27548 5684 27557
rect 4620 27480 4672 27532
rect 6552 27548 6604 27600
rect 7472 27548 7524 27600
rect 3148 27387 3200 27396
rect 3148 27353 3157 27387
rect 3157 27353 3191 27387
rect 3191 27353 3200 27387
rect 3148 27344 3200 27353
rect 3884 27344 3936 27396
rect 3240 27276 3292 27328
rect 3424 27276 3476 27328
rect 4988 27344 5040 27396
rect 5540 27344 5592 27396
rect 6368 27412 6420 27464
rect 6920 27412 6972 27464
rect 7380 27412 7432 27464
rect 6460 27344 6512 27396
rect 8024 27548 8076 27600
rect 7932 27412 7984 27464
rect 9588 27548 9640 27600
rect 9312 27480 9364 27532
rect 8484 27412 8536 27464
rect 9956 27480 10008 27532
rect 9588 27412 9640 27464
rect 9680 27412 9732 27464
rect 10140 27455 10192 27464
rect 10140 27421 10149 27455
rect 10149 27421 10183 27455
rect 10183 27421 10192 27455
rect 10140 27412 10192 27421
rect 10232 27412 10284 27464
rect 5080 27276 5132 27328
rect 5632 27276 5684 27328
rect 6276 27319 6328 27328
rect 6276 27285 6285 27319
rect 6285 27285 6319 27319
rect 6319 27285 6328 27319
rect 6276 27276 6328 27285
rect 7196 27276 7248 27328
rect 7932 27319 7984 27328
rect 7932 27285 7941 27319
rect 7941 27285 7975 27319
rect 7975 27285 7984 27319
rect 7932 27276 7984 27285
rect 9128 27276 9180 27328
rect 9864 27344 9916 27396
rect 9404 27276 9456 27328
rect 10416 27344 10468 27396
rect 10600 27455 10652 27464
rect 10600 27421 10609 27455
rect 10609 27421 10643 27455
rect 10643 27421 10652 27455
rect 10600 27412 10652 27421
rect 11060 27616 11112 27668
rect 12532 27616 12584 27668
rect 14556 27659 14608 27668
rect 14556 27625 14565 27659
rect 14565 27625 14599 27659
rect 14599 27625 14608 27659
rect 14556 27616 14608 27625
rect 15016 27616 15068 27668
rect 15200 27659 15252 27668
rect 15200 27625 15209 27659
rect 15209 27625 15243 27659
rect 15243 27625 15252 27659
rect 15200 27616 15252 27625
rect 16028 27659 16080 27668
rect 16028 27625 16037 27659
rect 16037 27625 16071 27659
rect 16071 27625 16080 27659
rect 16028 27616 16080 27625
rect 16396 27616 16448 27668
rect 10968 27548 11020 27600
rect 11336 27548 11388 27600
rect 12256 27548 12308 27600
rect 12624 27548 12676 27600
rect 12992 27591 13044 27600
rect 12992 27557 13001 27591
rect 13001 27557 13035 27591
rect 13035 27557 13044 27591
rect 12992 27548 13044 27557
rect 11336 27412 11388 27464
rect 11520 27455 11572 27464
rect 11520 27421 11529 27455
rect 11529 27421 11563 27455
rect 11563 27421 11572 27455
rect 11520 27412 11572 27421
rect 10876 27387 10928 27396
rect 10876 27353 10885 27387
rect 10885 27353 10919 27387
rect 10919 27353 10928 27387
rect 10876 27344 10928 27353
rect 11060 27276 11112 27328
rect 11152 27319 11204 27328
rect 11152 27285 11161 27319
rect 11161 27285 11195 27319
rect 11195 27285 11204 27319
rect 11152 27276 11204 27285
rect 11428 27276 11480 27328
rect 11980 27455 12032 27464
rect 11980 27421 11989 27455
rect 11989 27421 12023 27455
rect 12023 27421 12032 27455
rect 11980 27412 12032 27421
rect 12348 27412 12400 27464
rect 12532 27412 12584 27464
rect 12808 27455 12860 27464
rect 12808 27421 12817 27455
rect 12817 27421 12851 27455
rect 12851 27421 12860 27455
rect 12808 27412 12860 27421
rect 11888 27344 11940 27396
rect 13360 27276 13412 27328
rect 14924 27480 14976 27532
rect 16304 27591 16356 27600
rect 16304 27557 16313 27591
rect 16313 27557 16347 27591
rect 16347 27557 16356 27591
rect 16304 27548 16356 27557
rect 17592 27616 17644 27668
rect 17960 27616 18012 27668
rect 18880 27659 18932 27668
rect 18880 27625 18889 27659
rect 18889 27625 18923 27659
rect 18923 27625 18932 27659
rect 18880 27616 18932 27625
rect 19340 27616 19392 27668
rect 20260 27616 20312 27668
rect 20444 27659 20496 27668
rect 20444 27625 20453 27659
rect 20453 27625 20487 27659
rect 20487 27625 20496 27659
rect 20444 27616 20496 27625
rect 22468 27659 22520 27668
rect 22468 27625 22477 27659
rect 22477 27625 22511 27659
rect 22511 27625 22520 27659
rect 22468 27616 22520 27625
rect 14556 27276 14608 27328
rect 14648 27276 14700 27328
rect 15200 27412 15252 27464
rect 15384 27455 15436 27464
rect 15384 27421 15393 27455
rect 15393 27421 15427 27455
rect 15427 27421 15436 27455
rect 15384 27412 15436 27421
rect 14924 27344 14976 27396
rect 16488 27455 16540 27464
rect 16488 27421 16497 27455
rect 16497 27421 16531 27455
rect 16531 27421 16540 27455
rect 16488 27412 16540 27421
rect 18420 27480 18472 27532
rect 19248 27523 19300 27532
rect 19248 27489 19257 27523
rect 19257 27489 19291 27523
rect 19291 27489 19300 27523
rect 19248 27480 19300 27489
rect 16304 27276 16356 27328
rect 16948 27344 17000 27396
rect 17224 27412 17276 27464
rect 17776 27455 17828 27464
rect 17776 27421 17785 27455
rect 17785 27421 17819 27455
rect 17819 27421 17828 27455
rect 17776 27412 17828 27421
rect 18696 27455 18748 27464
rect 18696 27421 18705 27455
rect 18705 27421 18739 27455
rect 18739 27421 18748 27455
rect 18696 27412 18748 27421
rect 19524 27523 19576 27532
rect 19524 27489 19533 27523
rect 19533 27489 19567 27523
rect 19567 27489 19576 27523
rect 19524 27480 19576 27489
rect 24216 27659 24268 27668
rect 24216 27625 24225 27659
rect 24225 27625 24259 27659
rect 24259 27625 24268 27659
rect 24216 27616 24268 27625
rect 25596 27659 25648 27668
rect 25596 27625 25605 27659
rect 25605 27625 25639 27659
rect 25639 27625 25648 27659
rect 25596 27616 25648 27625
rect 26148 27616 26200 27668
rect 29736 27616 29788 27668
rect 20260 27480 20312 27532
rect 19984 27412 20036 27464
rect 22376 27523 22428 27532
rect 22376 27489 22385 27523
rect 22385 27489 22419 27523
rect 22419 27489 22428 27523
rect 22376 27480 22428 27489
rect 25320 27548 25372 27600
rect 17316 27276 17368 27328
rect 17868 27344 17920 27396
rect 17592 27319 17644 27328
rect 17592 27285 17601 27319
rect 17601 27285 17635 27319
rect 17635 27285 17644 27319
rect 19432 27344 19484 27396
rect 23572 27412 23624 27464
rect 23940 27455 23992 27464
rect 23940 27421 23949 27455
rect 23949 27421 23983 27455
rect 23983 27421 23992 27455
rect 23940 27412 23992 27421
rect 26516 27480 26568 27532
rect 17592 27276 17644 27285
rect 19248 27276 19300 27328
rect 19616 27276 19668 27328
rect 19708 27276 19760 27328
rect 19984 27276 20036 27328
rect 22008 27276 22060 27328
rect 22284 27387 22336 27396
rect 22284 27353 22293 27387
rect 22293 27353 22327 27387
rect 22327 27353 22336 27387
rect 22284 27344 22336 27353
rect 23848 27344 23900 27396
rect 25964 27412 26016 27464
rect 24124 27344 24176 27396
rect 22928 27276 22980 27328
rect 23940 27276 23992 27328
rect 26792 27387 26844 27396
rect 26792 27353 26801 27387
rect 26801 27353 26835 27387
rect 26835 27353 26844 27387
rect 26792 27344 26844 27353
rect 26884 27276 26936 27328
rect 27344 27276 27396 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 3056 27072 3108 27124
rect 3516 27072 3568 27124
rect 2780 27004 2832 27056
rect 4712 27072 4764 27124
rect 5080 27072 5132 27124
rect 6460 27072 6512 27124
rect 6644 27072 6696 27124
rect 2320 26979 2372 26988
rect 2320 26945 2329 26979
rect 2329 26945 2363 26979
rect 2363 26945 2372 26979
rect 2320 26936 2372 26945
rect 2872 26979 2924 26988
rect 2872 26945 2881 26979
rect 2881 26945 2915 26979
rect 2915 26945 2924 26979
rect 2872 26936 2924 26945
rect 3240 26979 3292 26988
rect 3240 26945 3249 26979
rect 3249 26945 3283 26979
rect 3283 26945 3292 26979
rect 3240 26936 3292 26945
rect 3516 26979 3568 26988
rect 3516 26945 3525 26979
rect 3525 26945 3559 26979
rect 3559 26945 3568 26979
rect 3516 26936 3568 26945
rect 3792 26979 3844 26988
rect 3792 26945 3801 26979
rect 3801 26945 3835 26979
rect 3835 26945 3844 26979
rect 3792 26936 3844 26945
rect 3884 26936 3936 26988
rect 4712 26979 4764 26988
rect 4712 26945 4721 26979
rect 4721 26945 4755 26979
rect 4755 26945 4764 26979
rect 4712 26936 4764 26945
rect 4896 26936 4948 26988
rect 6184 27004 6236 27056
rect 2596 26911 2648 26920
rect 2596 26877 2605 26911
rect 2605 26877 2639 26911
rect 2639 26877 2648 26911
rect 2596 26868 2648 26877
rect 3056 26911 3108 26920
rect 3056 26877 3065 26911
rect 3065 26877 3099 26911
rect 3099 26877 3108 26911
rect 3056 26868 3108 26877
rect 2964 26800 3016 26852
rect 3976 26868 4028 26920
rect 4620 26868 4672 26920
rect 4068 26800 4120 26852
rect 5632 26936 5684 26988
rect 6552 26936 6604 26988
rect 7012 27072 7064 27124
rect 7288 27072 7340 27124
rect 7472 27072 7524 27124
rect 7104 27004 7156 27056
rect 9496 27072 9548 27124
rect 6828 26868 6880 26920
rect 7012 26979 7064 26988
rect 7012 26945 7021 26979
rect 7021 26945 7055 26979
rect 7055 26945 7064 26979
rect 7012 26936 7064 26945
rect 7196 26936 7248 26988
rect 7472 26979 7524 26988
rect 7472 26945 7481 26979
rect 7481 26945 7515 26979
rect 7515 26945 7524 26979
rect 7472 26936 7524 26945
rect 7656 26979 7708 26988
rect 7656 26945 7665 26979
rect 7665 26945 7699 26979
rect 7699 26945 7708 26979
rect 7656 26936 7708 26945
rect 7840 26936 7892 26988
rect 8760 27004 8812 27056
rect 7748 26868 7800 26920
rect 3148 26732 3200 26784
rect 3516 26732 3568 26784
rect 8116 26800 8168 26852
rect 8392 26936 8444 26988
rect 9036 26979 9088 26988
rect 9036 26945 9045 26979
rect 9045 26945 9079 26979
rect 9079 26945 9088 26979
rect 9036 26936 9088 26945
rect 9128 26936 9180 26988
rect 9312 26979 9364 26988
rect 9312 26945 9321 26979
rect 9321 26945 9355 26979
rect 9355 26945 9364 26979
rect 9312 26936 9364 26945
rect 9772 27004 9824 27056
rect 9956 26979 10008 26988
rect 9404 26868 9456 26920
rect 9956 26945 9965 26979
rect 9965 26945 9999 26979
rect 9999 26945 10008 26979
rect 9956 26936 10008 26945
rect 10232 27072 10284 27124
rect 10416 27072 10468 27124
rect 11244 27004 11296 27056
rect 9772 26868 9824 26920
rect 10968 26936 11020 26988
rect 11060 26979 11112 26988
rect 11060 26945 11069 26979
rect 11069 26945 11103 26979
rect 11103 26945 11112 26979
rect 11704 27072 11756 27124
rect 11796 27072 11848 27124
rect 12532 27072 12584 27124
rect 13728 27072 13780 27124
rect 11060 26936 11112 26945
rect 10416 26868 10468 26920
rect 13360 27004 13412 27056
rect 12440 26936 12492 26988
rect 13176 26936 13228 26988
rect 13636 27004 13688 27056
rect 14464 27047 14516 27056
rect 14464 27013 14473 27047
rect 14473 27013 14507 27047
rect 14507 27013 14516 27047
rect 14464 27004 14516 27013
rect 12992 26868 13044 26920
rect 13728 26936 13780 26988
rect 14004 26979 14056 26988
rect 14004 26945 14013 26979
rect 14013 26945 14047 26979
rect 14047 26945 14056 26979
rect 14004 26936 14056 26945
rect 14188 26979 14240 26988
rect 14188 26945 14197 26979
rect 14197 26945 14231 26979
rect 14231 26945 14240 26979
rect 14188 26936 14240 26945
rect 14924 27115 14976 27124
rect 14924 27081 14933 27115
rect 14933 27081 14967 27115
rect 14967 27081 14976 27115
rect 14924 27072 14976 27081
rect 15016 27072 15068 27124
rect 22284 27072 22336 27124
rect 22560 27072 22612 27124
rect 14832 27004 14884 27056
rect 13360 26868 13412 26920
rect 15936 26936 15988 26988
rect 16856 26979 16908 26988
rect 16856 26945 16865 26979
rect 16865 26945 16899 26979
rect 16899 26945 16908 26979
rect 16856 26936 16908 26945
rect 17316 27047 17368 27056
rect 17316 27013 17325 27047
rect 17325 27013 17359 27047
rect 17359 27013 17368 27047
rect 17316 27004 17368 27013
rect 18512 27047 18564 27056
rect 18512 27013 18521 27047
rect 18521 27013 18555 27047
rect 18555 27013 18564 27047
rect 18512 27004 18564 27013
rect 18604 27004 18656 27056
rect 18236 26936 18288 26988
rect 19524 27004 19576 27056
rect 20720 27004 20772 27056
rect 19248 26936 19300 26988
rect 19616 26979 19668 26994
rect 19616 26945 19625 26979
rect 19625 26945 19659 26979
rect 19659 26945 19668 26979
rect 19616 26942 19668 26945
rect 19984 26936 20036 26988
rect 20444 26936 20496 26988
rect 4252 26775 4304 26784
rect 4252 26741 4261 26775
rect 4261 26741 4295 26775
rect 4295 26741 4304 26775
rect 4252 26732 4304 26741
rect 4712 26732 4764 26784
rect 4804 26732 4856 26784
rect 5908 26732 5960 26784
rect 6000 26775 6052 26784
rect 6000 26741 6009 26775
rect 6009 26741 6043 26775
rect 6043 26741 6052 26775
rect 6000 26732 6052 26741
rect 6828 26732 6880 26784
rect 7656 26732 7708 26784
rect 13912 26800 13964 26852
rect 14004 26800 14056 26852
rect 15568 26868 15620 26920
rect 17132 26868 17184 26920
rect 19892 26868 19944 26920
rect 8484 26775 8536 26784
rect 8484 26741 8493 26775
rect 8493 26741 8527 26775
rect 8527 26741 8536 26775
rect 8484 26732 8536 26741
rect 8576 26732 8628 26784
rect 9864 26775 9916 26784
rect 9864 26741 9873 26775
rect 9873 26741 9907 26775
rect 9907 26741 9916 26775
rect 9864 26732 9916 26741
rect 10232 26732 10284 26784
rect 10784 26732 10836 26784
rect 12992 26775 13044 26784
rect 12992 26741 13001 26775
rect 13001 26741 13035 26775
rect 13035 26741 13044 26775
rect 12992 26732 13044 26741
rect 13544 26775 13596 26784
rect 13544 26741 13553 26775
rect 13553 26741 13587 26775
rect 13587 26741 13596 26775
rect 13544 26732 13596 26741
rect 13820 26732 13872 26784
rect 14740 26800 14792 26852
rect 16488 26800 16540 26852
rect 16028 26732 16080 26784
rect 17408 26775 17460 26784
rect 17408 26741 17417 26775
rect 17417 26741 17451 26775
rect 17451 26741 17460 26775
rect 17408 26732 17460 26741
rect 17776 26775 17828 26784
rect 17776 26741 17785 26775
rect 17785 26741 17819 26775
rect 17819 26741 17828 26775
rect 17776 26732 17828 26741
rect 18788 26800 18840 26852
rect 19248 26843 19300 26852
rect 19248 26809 19257 26843
rect 19257 26809 19291 26843
rect 19291 26809 19300 26843
rect 19248 26800 19300 26809
rect 20812 26868 20864 26920
rect 21456 26936 21508 26988
rect 22560 26936 22612 26988
rect 23296 26979 23348 26988
rect 23296 26945 23305 26979
rect 23305 26945 23339 26979
rect 23339 26945 23348 26979
rect 23296 26936 23348 26945
rect 23756 27004 23808 27056
rect 28264 27115 28316 27124
rect 28264 27081 28273 27115
rect 28273 27081 28307 27115
rect 28307 27081 28316 27115
rect 28264 27072 28316 27081
rect 22008 26800 22060 26852
rect 25412 26936 25464 26988
rect 25596 26979 25648 26988
rect 25596 26945 25605 26979
rect 25605 26945 25639 26979
rect 25639 26945 25648 26979
rect 25596 26936 25648 26945
rect 25964 26936 26016 26988
rect 26976 26979 27028 26988
rect 26976 26945 26985 26979
rect 26985 26945 27019 26979
rect 27019 26945 27028 26979
rect 26976 26936 27028 26945
rect 27252 26979 27304 26988
rect 27252 26945 27261 26979
rect 27261 26945 27295 26979
rect 27295 26945 27304 26979
rect 27252 26936 27304 26945
rect 29920 27004 29972 27056
rect 30932 26979 30984 26988
rect 30932 26945 30941 26979
rect 30941 26945 30975 26979
rect 30975 26945 30984 26979
rect 30932 26936 30984 26945
rect 30380 26868 30432 26920
rect 31300 26979 31352 26988
rect 31300 26945 31309 26979
rect 31309 26945 31343 26979
rect 31343 26945 31352 26979
rect 31300 26936 31352 26945
rect 32496 26979 32548 26988
rect 32496 26945 32505 26979
rect 32505 26945 32539 26979
rect 32539 26945 32548 26979
rect 32496 26936 32548 26945
rect 27068 26800 27120 26852
rect 29828 26800 29880 26852
rect 19156 26732 19208 26784
rect 19524 26775 19576 26784
rect 19524 26741 19533 26775
rect 19533 26741 19567 26775
rect 19567 26741 19576 26775
rect 19524 26732 19576 26741
rect 19616 26732 19668 26784
rect 19800 26732 19852 26784
rect 19892 26775 19944 26784
rect 19892 26741 19901 26775
rect 19901 26741 19935 26775
rect 19935 26741 19944 26775
rect 19892 26732 19944 26741
rect 20168 26732 20220 26784
rect 22468 26732 22520 26784
rect 22836 26775 22888 26784
rect 22836 26741 22845 26775
rect 22845 26741 22879 26775
rect 22879 26741 22888 26775
rect 22836 26732 22888 26741
rect 23204 26732 23256 26784
rect 23756 26775 23808 26784
rect 23756 26741 23765 26775
rect 23765 26741 23799 26775
rect 23799 26741 23808 26775
rect 23756 26732 23808 26741
rect 25228 26775 25280 26784
rect 25228 26741 25237 26775
rect 25237 26741 25271 26775
rect 25271 26741 25280 26775
rect 25228 26732 25280 26741
rect 25688 26775 25740 26784
rect 25688 26741 25697 26775
rect 25697 26741 25731 26775
rect 25731 26741 25740 26775
rect 25688 26732 25740 26741
rect 26056 26775 26108 26784
rect 26056 26741 26065 26775
rect 26065 26741 26099 26775
rect 26099 26741 26108 26775
rect 26056 26732 26108 26741
rect 27160 26775 27212 26784
rect 27160 26741 27169 26775
rect 27169 26741 27203 26775
rect 27203 26741 27212 26775
rect 27160 26732 27212 26741
rect 27436 26775 27488 26784
rect 27436 26741 27445 26775
rect 27445 26741 27479 26775
rect 27479 26741 27488 26775
rect 27436 26732 27488 26741
rect 28356 26732 28408 26784
rect 31392 26732 31444 26784
rect 31668 26732 31720 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 3792 26528 3844 26580
rect 4160 26528 4212 26580
rect 4896 26571 4948 26580
rect 4896 26537 4905 26571
rect 4905 26537 4939 26571
rect 4939 26537 4948 26571
rect 4896 26528 4948 26537
rect 5540 26528 5592 26580
rect 3700 26460 3752 26512
rect 3976 26460 4028 26512
rect 5080 26460 5132 26512
rect 6736 26528 6788 26580
rect 7012 26528 7064 26580
rect 7840 26571 7892 26580
rect 7840 26537 7849 26571
rect 7849 26537 7883 26571
rect 7883 26537 7892 26571
rect 7840 26528 7892 26537
rect 8116 26571 8168 26580
rect 8116 26537 8125 26571
rect 8125 26537 8159 26571
rect 8159 26537 8168 26571
rect 8116 26528 8168 26537
rect 8944 26528 8996 26580
rect 9404 26528 9456 26580
rect 9864 26528 9916 26580
rect 2872 26392 2924 26444
rect 1400 26367 1452 26376
rect 1400 26333 1409 26367
rect 1409 26333 1443 26367
rect 1443 26333 1452 26367
rect 1400 26324 1452 26333
rect 2964 26367 3016 26376
rect 2964 26333 2973 26367
rect 2973 26333 3007 26367
rect 3007 26333 3016 26367
rect 2964 26324 3016 26333
rect 4068 26392 4120 26444
rect 4528 26392 4580 26444
rect 1676 26299 1728 26308
rect 1676 26265 1710 26299
rect 1710 26265 1728 26299
rect 1676 26256 1728 26265
rect 2780 26256 2832 26308
rect 3700 26256 3752 26308
rect 4620 26324 4672 26376
rect 4712 26367 4764 26376
rect 4712 26333 4721 26367
rect 4721 26333 4755 26367
rect 4755 26333 4764 26367
rect 4712 26324 4764 26333
rect 5356 26392 5408 26444
rect 5264 26367 5316 26376
rect 5264 26333 5273 26367
rect 5273 26333 5307 26367
rect 5307 26333 5316 26367
rect 5264 26324 5316 26333
rect 5540 26367 5592 26376
rect 5540 26333 5549 26367
rect 5549 26333 5583 26367
rect 5583 26333 5592 26367
rect 5540 26324 5592 26333
rect 6184 26460 6236 26512
rect 6368 26460 6420 26512
rect 6184 26324 6236 26376
rect 6460 26324 6512 26376
rect 7288 26392 7340 26444
rect 9312 26392 9364 26444
rect 10140 26392 10192 26444
rect 11060 26460 11112 26512
rect 12256 26460 12308 26512
rect 13084 26460 13136 26512
rect 13636 26571 13688 26580
rect 13636 26537 13645 26571
rect 13645 26537 13679 26571
rect 13679 26537 13688 26571
rect 13636 26528 13688 26537
rect 14832 26528 14884 26580
rect 15016 26571 15068 26580
rect 15016 26537 15025 26571
rect 15025 26537 15059 26571
rect 15059 26537 15068 26571
rect 15016 26528 15068 26537
rect 15200 26571 15252 26580
rect 15200 26537 15209 26571
rect 15209 26537 15243 26571
rect 15243 26537 15252 26571
rect 15200 26528 15252 26537
rect 16028 26571 16080 26580
rect 16028 26537 16037 26571
rect 16037 26537 16071 26571
rect 16071 26537 16080 26571
rect 16028 26528 16080 26537
rect 14188 26460 14240 26512
rect 14464 26460 14516 26512
rect 17408 26460 17460 26512
rect 18420 26528 18472 26580
rect 19524 26528 19576 26580
rect 3148 26188 3200 26240
rect 3976 26188 4028 26240
rect 5632 26188 5684 26240
rect 5724 26188 5776 26240
rect 6184 26188 6236 26240
rect 6920 26256 6972 26308
rect 7748 26324 7800 26376
rect 8300 26324 8352 26376
rect 9220 26367 9272 26376
rect 9220 26333 9229 26367
rect 9229 26333 9263 26367
rect 9263 26333 9272 26367
rect 9220 26324 9272 26333
rect 6644 26188 6696 26240
rect 6736 26188 6788 26240
rect 7288 26299 7340 26308
rect 7288 26265 7297 26299
rect 7297 26265 7331 26299
rect 7331 26265 7340 26299
rect 7288 26256 7340 26265
rect 8116 26256 8168 26308
rect 10692 26324 10744 26376
rect 10784 26324 10836 26376
rect 11244 26324 11296 26376
rect 9496 26256 9548 26308
rect 7472 26188 7524 26240
rect 8300 26188 8352 26240
rect 8760 26188 8812 26240
rect 9220 26188 9272 26240
rect 10048 26231 10100 26240
rect 10048 26197 10057 26231
rect 10057 26197 10091 26231
rect 10091 26197 10100 26231
rect 10048 26188 10100 26197
rect 11704 26367 11756 26376
rect 11704 26333 11713 26367
rect 11713 26333 11747 26367
rect 11747 26333 11756 26367
rect 11704 26324 11756 26333
rect 14832 26435 14884 26444
rect 14832 26401 14841 26435
rect 14841 26401 14875 26435
rect 14875 26401 14884 26435
rect 14832 26392 14884 26401
rect 11888 26324 11940 26376
rect 12716 26324 12768 26376
rect 11428 26299 11480 26308
rect 11428 26265 11437 26299
rect 11437 26265 11471 26299
rect 11471 26265 11480 26299
rect 11428 26256 11480 26265
rect 11520 26299 11572 26308
rect 11520 26265 11529 26299
rect 11529 26265 11563 26299
rect 11563 26265 11572 26299
rect 11520 26256 11572 26265
rect 12808 26256 12860 26308
rect 13360 26324 13412 26376
rect 13728 26367 13780 26376
rect 13728 26333 13737 26367
rect 13737 26333 13771 26367
rect 13771 26333 13780 26367
rect 13728 26324 13780 26333
rect 15016 26367 15068 26376
rect 15016 26333 15025 26367
rect 15025 26333 15059 26367
rect 15059 26333 15068 26367
rect 15016 26324 15068 26333
rect 15292 26324 15344 26376
rect 11336 26188 11388 26240
rect 11888 26188 11940 26240
rect 13176 26188 13228 26240
rect 14832 26256 14884 26308
rect 16120 26256 16172 26308
rect 16304 26367 16356 26376
rect 16304 26333 16313 26367
rect 16313 26333 16347 26367
rect 16347 26333 16356 26367
rect 16304 26324 16356 26333
rect 18236 26324 18288 26376
rect 16488 26256 16540 26308
rect 17224 26256 17276 26308
rect 17592 26256 17644 26308
rect 18696 26460 18748 26512
rect 20168 26460 20220 26512
rect 22836 26528 22888 26580
rect 21364 26460 21416 26512
rect 21732 26460 21784 26512
rect 24860 26528 24912 26580
rect 25596 26528 25648 26580
rect 26976 26571 27028 26580
rect 26976 26537 26985 26571
rect 26985 26537 27019 26571
rect 27019 26537 27028 26571
rect 26976 26528 27028 26537
rect 27436 26528 27488 26580
rect 23480 26460 23532 26512
rect 25688 26460 25740 26512
rect 25964 26460 26016 26512
rect 27896 26571 27948 26580
rect 27896 26537 27905 26571
rect 27905 26537 27939 26571
rect 27939 26537 27948 26571
rect 27896 26528 27948 26537
rect 28356 26571 28408 26580
rect 28356 26537 28365 26571
rect 28365 26537 28399 26571
rect 28399 26537 28408 26571
rect 28356 26528 28408 26537
rect 31300 26528 31352 26580
rect 19892 26392 19944 26444
rect 19984 26392 20036 26444
rect 21916 26392 21968 26444
rect 22744 26392 22796 26444
rect 18696 26324 18748 26376
rect 18788 26367 18840 26376
rect 18788 26333 18797 26367
rect 18797 26333 18831 26367
rect 18831 26333 18840 26367
rect 18788 26324 18840 26333
rect 18880 26324 18932 26376
rect 20444 26324 20496 26376
rect 21180 26299 21232 26308
rect 21180 26265 21189 26299
rect 21189 26265 21223 26299
rect 21223 26265 21232 26299
rect 21180 26256 21232 26265
rect 21732 26324 21784 26376
rect 21824 26367 21876 26376
rect 21824 26333 21833 26367
rect 21833 26333 21867 26367
rect 21867 26333 21876 26367
rect 21824 26324 21876 26333
rect 23204 26435 23256 26444
rect 23204 26401 23213 26435
rect 23213 26401 23247 26435
rect 23247 26401 23256 26435
rect 23204 26392 23256 26401
rect 23756 26392 23808 26444
rect 26976 26392 27028 26444
rect 24308 26324 24360 26376
rect 27160 26324 27212 26376
rect 27896 26392 27948 26444
rect 28448 26460 28500 26512
rect 21548 26299 21600 26308
rect 21548 26265 21557 26299
rect 21557 26265 21591 26299
rect 21591 26265 21600 26299
rect 21548 26256 21600 26265
rect 23296 26256 23348 26308
rect 25320 26256 25372 26308
rect 27068 26299 27120 26308
rect 27068 26265 27077 26299
rect 27077 26265 27111 26299
rect 27111 26265 27120 26299
rect 27068 26256 27120 26265
rect 27712 26367 27764 26376
rect 27712 26333 27721 26367
rect 27721 26333 27755 26367
rect 27755 26333 27764 26367
rect 27712 26324 27764 26333
rect 18328 26231 18380 26240
rect 18328 26197 18337 26231
rect 18337 26197 18371 26231
rect 18371 26197 18380 26231
rect 18328 26188 18380 26197
rect 18512 26188 18564 26240
rect 22836 26188 22888 26240
rect 27252 26231 27304 26240
rect 27252 26197 27261 26231
rect 27261 26197 27295 26231
rect 27295 26197 27304 26231
rect 27252 26188 27304 26197
rect 29276 26324 29328 26376
rect 31760 26324 31812 26376
rect 32496 26367 32548 26376
rect 32496 26333 32505 26367
rect 32505 26333 32539 26367
rect 32539 26333 32548 26367
rect 32496 26324 32548 26333
rect 30932 26231 30984 26240
rect 30932 26197 30941 26231
rect 30941 26197 30975 26231
rect 30975 26197 30984 26231
rect 30932 26188 30984 26197
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 1676 25984 1728 26036
rect 2872 25984 2924 26036
rect 2964 25916 3016 25968
rect 5632 25984 5684 26036
rect 6552 25984 6604 26036
rect 6644 25984 6696 26036
rect 8392 25984 8444 26036
rect 9036 25984 9088 26036
rect 9496 25984 9548 26036
rect 5540 25916 5592 25968
rect 848 25848 900 25900
rect 2780 25848 2832 25900
rect 3148 25891 3200 25900
rect 3148 25857 3157 25891
rect 3157 25857 3191 25891
rect 3191 25857 3200 25891
rect 3148 25848 3200 25857
rect 3332 25848 3384 25900
rect 3700 25891 3752 25900
rect 3700 25857 3709 25891
rect 3709 25857 3743 25891
rect 3743 25857 3752 25891
rect 3700 25848 3752 25857
rect 4160 25848 4212 25900
rect 4528 25891 4580 25900
rect 4528 25857 4537 25891
rect 4537 25857 4571 25891
rect 4571 25857 4580 25891
rect 4528 25848 4580 25857
rect 4988 25848 5040 25900
rect 5080 25891 5132 25900
rect 5080 25857 5089 25891
rect 5089 25857 5123 25891
rect 5123 25857 5132 25891
rect 5080 25848 5132 25857
rect 5172 25848 5224 25900
rect 5908 25848 5960 25900
rect 6092 25848 6144 25900
rect 6368 25891 6420 25900
rect 6368 25857 6377 25891
rect 6377 25857 6411 25891
rect 6411 25857 6420 25891
rect 6368 25848 6420 25857
rect 6552 25891 6604 25900
rect 6552 25857 6561 25891
rect 6561 25857 6595 25891
rect 6595 25857 6604 25891
rect 6552 25848 6604 25857
rect 7656 25916 7708 25968
rect 8300 25916 8352 25968
rect 11428 25984 11480 26036
rect 11796 25984 11848 26036
rect 12532 25984 12584 26036
rect 13728 25984 13780 26036
rect 19800 25984 19852 26036
rect 11520 25916 11572 25968
rect 5816 25780 5868 25832
rect 6920 25848 6972 25900
rect 7196 25891 7248 25900
rect 7196 25857 7205 25891
rect 7205 25857 7239 25891
rect 7239 25857 7248 25891
rect 7196 25848 7248 25857
rect 5264 25712 5316 25764
rect 7104 25780 7156 25832
rect 8116 25848 8168 25900
rect 8392 25848 8444 25900
rect 8760 25891 8812 25900
rect 8760 25857 8769 25891
rect 8769 25857 8803 25891
rect 8803 25857 8812 25891
rect 8760 25848 8812 25857
rect 8300 25780 8352 25832
rect 8944 25780 8996 25832
rect 3700 25644 3752 25696
rect 4068 25644 4120 25696
rect 5172 25644 5224 25696
rect 6828 25712 6880 25764
rect 9404 25848 9456 25900
rect 9680 25891 9732 25900
rect 9680 25857 9689 25891
rect 9689 25857 9723 25891
rect 9723 25857 9732 25891
rect 9680 25848 9732 25857
rect 10324 25848 10376 25900
rect 10508 25848 10560 25900
rect 9496 25780 9548 25832
rect 11336 25848 11388 25900
rect 11428 25848 11480 25900
rect 11520 25780 11572 25832
rect 11704 25780 11756 25832
rect 12624 25780 12676 25832
rect 14280 25848 14332 25900
rect 16672 25916 16724 25968
rect 16764 25891 16816 25900
rect 16764 25857 16773 25891
rect 16773 25857 16807 25891
rect 16807 25857 16816 25891
rect 16764 25848 16816 25857
rect 16948 25891 17000 25900
rect 16948 25857 16957 25891
rect 16957 25857 16991 25891
rect 16991 25857 17000 25891
rect 16948 25848 17000 25857
rect 17408 25916 17460 25968
rect 20812 25984 20864 26036
rect 21916 25984 21968 26036
rect 22836 25984 22888 26036
rect 25412 25984 25464 26036
rect 30104 25984 30156 26036
rect 18420 25848 18472 25900
rect 19340 25848 19392 25900
rect 19616 25848 19668 25900
rect 19892 25891 19944 25900
rect 19892 25857 19901 25891
rect 19901 25857 19935 25891
rect 19935 25857 19944 25891
rect 19892 25848 19944 25857
rect 20260 25891 20312 25900
rect 20260 25857 20269 25891
rect 20269 25857 20303 25891
rect 20303 25857 20312 25891
rect 20260 25848 20312 25857
rect 20444 25891 20496 25900
rect 20444 25857 20453 25891
rect 20453 25857 20487 25891
rect 20487 25857 20496 25891
rect 20444 25848 20496 25857
rect 20996 25891 21048 25900
rect 20996 25857 21005 25891
rect 21005 25857 21039 25891
rect 21039 25857 21048 25891
rect 20996 25848 21048 25857
rect 21180 25848 21232 25900
rect 18696 25780 18748 25832
rect 7104 25644 7156 25696
rect 7196 25644 7248 25696
rect 8300 25644 8352 25696
rect 8576 25644 8628 25696
rect 9128 25712 9180 25764
rect 15752 25712 15804 25764
rect 17224 25712 17276 25764
rect 17500 25712 17552 25764
rect 10784 25644 10836 25696
rect 10968 25687 11020 25696
rect 10968 25653 10977 25687
rect 10977 25653 11011 25687
rect 11011 25653 11020 25687
rect 10968 25644 11020 25653
rect 12992 25687 13044 25696
rect 12992 25653 13001 25687
rect 13001 25653 13035 25687
rect 13035 25653 13044 25687
rect 12992 25644 13044 25653
rect 13084 25644 13136 25696
rect 13912 25644 13964 25696
rect 20720 25780 20772 25832
rect 20812 25780 20864 25832
rect 21916 25848 21968 25900
rect 22652 25848 22704 25900
rect 23112 25848 23164 25900
rect 23480 25848 23532 25900
rect 29920 25959 29972 25968
rect 29920 25925 29929 25959
rect 29929 25925 29963 25959
rect 29963 25925 29972 25959
rect 29920 25916 29972 25925
rect 24584 25848 24636 25900
rect 29644 25891 29696 25900
rect 29644 25857 29653 25891
rect 29653 25857 29687 25891
rect 29687 25857 29696 25891
rect 29644 25848 29696 25857
rect 30932 25848 30984 25900
rect 32128 25848 32180 25900
rect 19524 25712 19576 25764
rect 19340 25687 19392 25696
rect 19340 25653 19349 25687
rect 19349 25653 19383 25687
rect 19383 25653 19392 25687
rect 19340 25644 19392 25653
rect 19984 25687 20036 25696
rect 19984 25653 19993 25687
rect 19993 25653 20027 25687
rect 20027 25653 20036 25687
rect 25504 25780 25556 25832
rect 25780 25780 25832 25832
rect 19984 25644 20036 25653
rect 20260 25687 20312 25696
rect 20260 25653 20269 25687
rect 20269 25653 20303 25687
rect 20303 25653 20312 25687
rect 20260 25644 20312 25653
rect 20444 25644 20496 25696
rect 23848 25712 23900 25764
rect 29460 25712 29512 25764
rect 20996 25644 21048 25696
rect 21364 25644 21416 25696
rect 21456 25687 21508 25696
rect 21456 25653 21465 25687
rect 21465 25653 21499 25687
rect 21499 25653 21508 25687
rect 21456 25644 21508 25653
rect 21548 25644 21600 25696
rect 22928 25644 22980 25696
rect 23664 25687 23716 25696
rect 23664 25653 23673 25687
rect 23673 25653 23707 25687
rect 23707 25653 23716 25687
rect 23664 25644 23716 25653
rect 24216 25687 24268 25696
rect 24216 25653 24225 25687
rect 24225 25653 24259 25687
rect 24259 25653 24268 25687
rect 24216 25644 24268 25653
rect 24952 25644 25004 25696
rect 25964 25644 26016 25696
rect 31760 25780 31812 25832
rect 32220 25712 32272 25764
rect 30932 25644 30984 25696
rect 31760 25644 31812 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 3884 25440 3936 25492
rect 6184 25440 6236 25492
rect 6552 25440 6604 25492
rect 6736 25483 6788 25492
rect 6736 25449 6745 25483
rect 6745 25449 6779 25483
rect 6779 25449 6788 25483
rect 6736 25440 6788 25449
rect 6920 25440 6972 25492
rect 8484 25440 8536 25492
rect 8760 25440 8812 25492
rect 9312 25440 9364 25492
rect 4620 25372 4672 25424
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 3056 25279 3108 25288
rect 3056 25245 3065 25279
rect 3065 25245 3099 25279
rect 3099 25245 3108 25279
rect 3056 25236 3108 25245
rect 3148 25279 3200 25288
rect 3148 25245 3157 25279
rect 3157 25245 3191 25279
rect 3191 25245 3200 25279
rect 3148 25236 3200 25245
rect 3608 25279 3660 25288
rect 3608 25245 3617 25279
rect 3617 25245 3651 25279
rect 3651 25245 3660 25279
rect 3608 25236 3660 25245
rect 4344 25304 4396 25356
rect 6092 25372 6144 25424
rect 9680 25440 9732 25492
rect 11428 25440 11480 25492
rect 12808 25483 12860 25492
rect 12808 25449 12817 25483
rect 12817 25449 12851 25483
rect 12851 25449 12860 25483
rect 12808 25440 12860 25449
rect 13084 25440 13136 25492
rect 13728 25440 13780 25492
rect 17500 25440 17552 25492
rect 19708 25440 19760 25492
rect 20168 25440 20220 25492
rect 20444 25440 20496 25492
rect 20812 25440 20864 25492
rect 21364 25483 21416 25492
rect 21364 25449 21373 25483
rect 21373 25449 21407 25483
rect 21407 25449 21416 25483
rect 21364 25440 21416 25449
rect 22744 25483 22796 25492
rect 22744 25449 22753 25483
rect 22753 25449 22787 25483
rect 22787 25449 22796 25483
rect 22744 25440 22796 25449
rect 23664 25483 23716 25492
rect 23664 25449 23673 25483
rect 23673 25449 23707 25483
rect 23707 25449 23716 25483
rect 23664 25440 23716 25449
rect 24216 25483 24268 25492
rect 24216 25449 24225 25483
rect 24225 25449 24259 25483
rect 24259 25449 24268 25483
rect 24216 25440 24268 25449
rect 9588 25415 9640 25424
rect 9588 25381 9597 25415
rect 9597 25381 9631 25415
rect 9631 25381 9640 25415
rect 9588 25372 9640 25381
rect 4160 25279 4212 25288
rect 4160 25245 4169 25279
rect 4169 25245 4203 25279
rect 4203 25245 4212 25279
rect 4160 25236 4212 25245
rect 1676 25211 1728 25220
rect 1676 25177 1710 25211
rect 1710 25177 1728 25211
rect 1676 25168 1728 25177
rect 5264 25279 5316 25288
rect 5264 25245 5273 25279
rect 5273 25245 5307 25279
rect 5307 25245 5316 25279
rect 5264 25236 5316 25245
rect 6460 25304 6512 25356
rect 8576 25304 8628 25356
rect 5816 25279 5868 25288
rect 5816 25245 5825 25279
rect 5825 25245 5859 25279
rect 5859 25245 5868 25279
rect 5816 25236 5868 25245
rect 2872 25143 2924 25152
rect 2872 25109 2881 25143
rect 2881 25109 2915 25143
rect 2915 25109 2924 25143
rect 2872 25100 2924 25109
rect 3332 25143 3384 25152
rect 3332 25109 3341 25143
rect 3341 25109 3375 25143
rect 3375 25109 3384 25143
rect 3332 25100 3384 25109
rect 3424 25143 3476 25152
rect 3424 25109 3433 25143
rect 3433 25109 3467 25143
rect 3467 25109 3476 25143
rect 3424 25100 3476 25109
rect 4712 25168 4764 25220
rect 5632 25168 5684 25220
rect 6184 25279 6236 25288
rect 6184 25245 6193 25279
rect 6193 25245 6227 25279
rect 6227 25245 6236 25279
rect 6184 25236 6236 25245
rect 6552 25236 6604 25288
rect 6644 25279 6696 25288
rect 6644 25245 6653 25279
rect 6653 25245 6687 25279
rect 6687 25245 6696 25279
rect 6644 25236 6696 25245
rect 6828 25236 6880 25288
rect 8392 25236 8444 25288
rect 8944 25279 8996 25288
rect 8944 25245 8953 25279
rect 8953 25245 8987 25279
rect 8987 25245 8996 25279
rect 8944 25236 8996 25245
rect 9036 25236 9088 25288
rect 9496 25236 9548 25288
rect 11244 25372 11296 25424
rect 11704 25372 11756 25424
rect 9956 25304 10008 25356
rect 10140 25236 10192 25288
rect 10508 25279 10560 25288
rect 10508 25245 10517 25279
rect 10517 25245 10551 25279
rect 10551 25245 10560 25279
rect 10508 25236 10560 25245
rect 11152 25304 11204 25356
rect 4804 25100 4856 25152
rect 5816 25100 5868 25152
rect 6460 25100 6512 25152
rect 7932 25100 7984 25152
rect 9956 25211 10008 25220
rect 9956 25177 9965 25211
rect 9965 25177 9999 25211
rect 9999 25177 10008 25211
rect 9956 25168 10008 25177
rect 10140 25100 10192 25152
rect 10416 25100 10468 25152
rect 11244 25236 11296 25288
rect 11428 25279 11480 25288
rect 11428 25245 11437 25279
rect 11437 25245 11471 25279
rect 11471 25245 11480 25279
rect 11428 25236 11480 25245
rect 11520 25236 11572 25288
rect 11796 25279 11848 25288
rect 11796 25245 11805 25279
rect 11805 25245 11839 25279
rect 11839 25245 11848 25279
rect 11796 25236 11848 25245
rect 12348 25279 12400 25288
rect 12348 25245 12357 25279
rect 12357 25245 12391 25279
rect 12391 25245 12400 25279
rect 12348 25236 12400 25245
rect 12624 25415 12676 25424
rect 12624 25381 12633 25415
rect 12633 25381 12667 25415
rect 12667 25381 12676 25415
rect 12624 25372 12676 25381
rect 15292 25372 15344 25424
rect 16120 25372 16172 25424
rect 17224 25372 17276 25424
rect 13728 25304 13780 25356
rect 17040 25304 17092 25356
rect 12624 25236 12676 25288
rect 12992 25279 13044 25288
rect 12992 25245 13001 25279
rect 13001 25245 13035 25279
rect 13035 25245 13044 25279
rect 12992 25236 13044 25245
rect 13084 25279 13136 25288
rect 13084 25245 13093 25279
rect 13093 25245 13127 25279
rect 13127 25245 13136 25279
rect 13084 25236 13136 25245
rect 14372 25236 14424 25288
rect 14556 25236 14608 25288
rect 15200 25236 15252 25288
rect 16028 25236 16080 25288
rect 16396 25236 16448 25288
rect 16672 25279 16724 25288
rect 16672 25245 16681 25279
rect 16681 25245 16715 25279
rect 16715 25245 16724 25279
rect 16672 25236 16724 25245
rect 17224 25279 17276 25288
rect 17224 25245 17233 25279
rect 17233 25245 17267 25279
rect 17267 25245 17276 25279
rect 17224 25236 17276 25245
rect 12256 25211 12308 25220
rect 12256 25177 12265 25211
rect 12265 25177 12299 25211
rect 12299 25177 12308 25211
rect 12256 25168 12308 25177
rect 11796 25100 11848 25152
rect 12532 25100 12584 25152
rect 13360 25211 13412 25220
rect 13360 25177 13369 25211
rect 13369 25177 13403 25211
rect 13403 25177 13412 25211
rect 13360 25168 13412 25177
rect 16120 25211 16172 25220
rect 16120 25177 16129 25211
rect 16129 25177 16163 25211
rect 16163 25177 16172 25211
rect 16120 25168 16172 25177
rect 18420 25304 18472 25356
rect 19156 25304 19208 25356
rect 19892 25372 19944 25424
rect 20720 25415 20772 25424
rect 20720 25381 20729 25415
rect 20729 25381 20763 25415
rect 20763 25381 20772 25415
rect 20720 25372 20772 25381
rect 21088 25372 21140 25424
rect 21180 25372 21232 25424
rect 17408 25279 17460 25288
rect 17408 25245 17417 25279
rect 17417 25245 17451 25279
rect 17451 25245 17460 25279
rect 17408 25236 17460 25245
rect 17500 25236 17552 25288
rect 17776 25279 17828 25288
rect 17776 25245 17785 25279
rect 17785 25245 17819 25279
rect 17819 25245 17828 25279
rect 17776 25236 17828 25245
rect 18512 25236 18564 25288
rect 19432 25279 19484 25288
rect 19432 25245 19441 25279
rect 19441 25245 19475 25279
rect 19475 25245 19484 25279
rect 19432 25236 19484 25245
rect 19708 25236 19760 25288
rect 19984 25236 20036 25288
rect 20536 25279 20588 25288
rect 20536 25245 20545 25279
rect 20545 25245 20579 25279
rect 20579 25245 20588 25279
rect 20536 25236 20588 25245
rect 21180 25236 21232 25288
rect 21456 25304 21508 25356
rect 22652 25372 22704 25424
rect 23480 25372 23532 25424
rect 24860 25440 24912 25492
rect 25780 25440 25832 25492
rect 25964 25483 26016 25492
rect 25964 25449 25973 25483
rect 25973 25449 26007 25483
rect 26007 25449 26016 25483
rect 25964 25440 26016 25449
rect 29552 25483 29604 25492
rect 29552 25449 29561 25483
rect 29561 25449 29595 25483
rect 29595 25449 29604 25483
rect 29552 25440 29604 25449
rect 29644 25440 29696 25492
rect 32496 25483 32548 25492
rect 32496 25449 32505 25483
rect 32505 25449 32539 25483
rect 32539 25449 32548 25483
rect 32496 25440 32548 25449
rect 21548 25236 21600 25288
rect 21916 25279 21968 25288
rect 21916 25245 21925 25279
rect 21925 25245 21959 25279
rect 21959 25245 21968 25279
rect 21916 25236 21968 25245
rect 22652 25236 22704 25288
rect 22744 25236 22796 25288
rect 23112 25236 23164 25288
rect 24952 25304 25004 25356
rect 12992 25100 13044 25152
rect 14188 25100 14240 25152
rect 14372 25100 14424 25152
rect 16396 25143 16448 25152
rect 16396 25109 16405 25143
rect 16405 25109 16439 25143
rect 16439 25109 16448 25143
rect 16396 25100 16448 25109
rect 16580 25100 16632 25152
rect 16856 25100 16908 25152
rect 18052 25100 18104 25152
rect 18236 25143 18288 25152
rect 18236 25109 18245 25143
rect 18245 25109 18279 25143
rect 18279 25109 18288 25143
rect 18236 25100 18288 25109
rect 18420 25100 18472 25152
rect 24216 25211 24268 25220
rect 24216 25177 24225 25211
rect 24225 25177 24259 25211
rect 24259 25177 24268 25211
rect 24216 25168 24268 25177
rect 25044 25211 25096 25220
rect 25044 25177 25053 25211
rect 25053 25177 25087 25211
rect 25087 25177 25096 25211
rect 25044 25168 25096 25177
rect 25596 25304 25648 25356
rect 26516 25347 26568 25356
rect 26516 25313 26525 25347
rect 26525 25313 26559 25347
rect 26559 25313 26568 25347
rect 26516 25304 26568 25313
rect 27436 25304 27488 25356
rect 30932 25304 30984 25356
rect 25504 25236 25556 25288
rect 26608 25279 26660 25288
rect 26608 25245 26617 25279
rect 26617 25245 26651 25279
rect 26651 25245 26660 25279
rect 26608 25236 26660 25245
rect 29460 25236 29512 25288
rect 29644 25279 29696 25288
rect 29644 25245 29653 25279
rect 29653 25245 29687 25279
rect 29687 25245 29696 25279
rect 29644 25236 29696 25245
rect 31392 25279 31444 25288
rect 31392 25245 31426 25279
rect 31426 25245 31444 25279
rect 22100 25143 22152 25152
rect 22100 25109 22109 25143
rect 22109 25109 22143 25143
rect 22143 25109 22152 25143
rect 22100 25100 22152 25109
rect 23204 25100 23256 25152
rect 23388 25143 23440 25152
rect 23388 25109 23397 25143
rect 23397 25109 23431 25143
rect 23431 25109 23440 25143
rect 23388 25100 23440 25109
rect 24124 25100 24176 25152
rect 24768 25100 24820 25152
rect 26240 25168 26292 25220
rect 26516 25168 26568 25220
rect 31392 25236 31444 25245
rect 31852 25168 31904 25220
rect 26148 25143 26200 25152
rect 26148 25109 26157 25143
rect 26157 25109 26191 25143
rect 26191 25109 26200 25143
rect 26148 25100 26200 25109
rect 26792 25143 26844 25152
rect 26792 25109 26801 25143
rect 26801 25109 26835 25143
rect 26835 25109 26844 25143
rect 26792 25100 26844 25109
rect 30840 25143 30892 25152
rect 30840 25109 30849 25143
rect 30849 25109 30883 25143
rect 30883 25109 30892 25143
rect 30840 25100 30892 25109
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 3516 24939 3568 24948
rect 3516 24905 3525 24939
rect 3525 24905 3559 24939
rect 3559 24905 3568 24939
rect 3516 24896 3568 24905
rect 3976 24939 4028 24948
rect 3976 24905 3985 24939
rect 3985 24905 4019 24939
rect 4019 24905 4028 24939
rect 3976 24896 4028 24905
rect 5264 24896 5316 24948
rect 6000 24896 6052 24948
rect 6644 24896 6696 24948
rect 2688 24828 2740 24880
rect 2872 24828 2924 24880
rect 2044 24760 2096 24812
rect 2320 24760 2372 24812
rect 2412 24803 2464 24812
rect 2412 24769 2421 24803
rect 2421 24769 2455 24803
rect 2455 24769 2464 24803
rect 2412 24760 2464 24769
rect 3792 24803 3844 24812
rect 3792 24769 3801 24803
rect 3801 24769 3835 24803
rect 3835 24769 3844 24803
rect 3792 24760 3844 24769
rect 4068 24803 4120 24812
rect 4068 24769 4077 24803
rect 4077 24769 4111 24803
rect 4111 24769 4120 24803
rect 4068 24760 4120 24769
rect 5540 24871 5592 24880
rect 5540 24837 5549 24871
rect 5549 24837 5583 24871
rect 5583 24837 5592 24871
rect 5540 24828 5592 24837
rect 3148 24624 3200 24676
rect 2596 24599 2648 24608
rect 2596 24565 2605 24599
rect 2605 24565 2639 24599
rect 2639 24565 2648 24599
rect 4160 24692 4212 24744
rect 4344 24735 4396 24744
rect 4344 24701 4353 24735
rect 4353 24701 4387 24735
rect 4387 24701 4396 24735
rect 4344 24692 4396 24701
rect 5632 24803 5684 24812
rect 5632 24769 5641 24803
rect 5641 24769 5675 24803
rect 5675 24769 5684 24803
rect 5632 24760 5684 24769
rect 5816 24760 5868 24812
rect 6092 24760 6144 24812
rect 6184 24803 6236 24812
rect 6184 24769 6193 24803
rect 6193 24769 6227 24803
rect 6227 24769 6236 24803
rect 9036 24896 9088 24948
rect 7196 24871 7248 24880
rect 7196 24837 7205 24871
rect 7205 24837 7239 24871
rect 7239 24837 7248 24871
rect 7196 24828 7248 24837
rect 6184 24760 6236 24769
rect 3608 24624 3660 24676
rect 4068 24624 4120 24676
rect 5908 24667 5960 24676
rect 5908 24633 5917 24667
rect 5917 24633 5951 24667
rect 5951 24633 5960 24667
rect 5908 24624 5960 24633
rect 6000 24667 6052 24676
rect 6000 24633 6009 24667
rect 6009 24633 6043 24667
rect 6043 24633 6052 24667
rect 6000 24624 6052 24633
rect 6920 24624 6972 24676
rect 7840 24760 7892 24812
rect 8668 24828 8720 24880
rect 9956 24896 10008 24948
rect 11520 24896 11572 24948
rect 12256 24896 12308 24948
rect 10048 24828 10100 24880
rect 16396 24896 16448 24948
rect 16672 24939 16724 24948
rect 16672 24905 16681 24939
rect 16681 24905 16715 24939
rect 16715 24905 16724 24939
rect 16672 24896 16724 24905
rect 17868 24896 17920 24948
rect 19892 24896 19944 24948
rect 20168 24896 20220 24948
rect 8484 24803 8536 24812
rect 8484 24769 8493 24803
rect 8493 24769 8527 24803
rect 8527 24769 8536 24803
rect 8484 24760 8536 24769
rect 8576 24760 8628 24812
rect 9680 24760 9732 24812
rect 11520 24803 11572 24812
rect 11520 24769 11529 24803
rect 11529 24769 11563 24803
rect 11563 24769 11572 24803
rect 11520 24760 11572 24769
rect 11704 24803 11756 24812
rect 11704 24769 11713 24803
rect 11713 24769 11747 24803
rect 11747 24769 11756 24803
rect 11704 24760 11756 24769
rect 11796 24803 11848 24812
rect 11796 24769 11805 24803
rect 11805 24769 11839 24803
rect 11839 24769 11848 24803
rect 11796 24760 11848 24769
rect 12348 24760 12400 24812
rect 9772 24692 9824 24744
rect 12256 24692 12308 24744
rect 13912 24828 13964 24880
rect 14188 24828 14240 24880
rect 16120 24828 16172 24880
rect 2596 24556 2648 24565
rect 3700 24556 3752 24608
rect 6552 24556 6604 24608
rect 8484 24624 8536 24676
rect 7748 24556 7800 24608
rect 11520 24624 11572 24676
rect 13268 24803 13320 24812
rect 13268 24769 13277 24803
rect 13277 24769 13311 24803
rect 13311 24769 13320 24803
rect 13268 24760 13320 24769
rect 13452 24803 13504 24812
rect 13452 24769 13461 24803
rect 13461 24769 13495 24803
rect 13495 24769 13504 24803
rect 13452 24760 13504 24769
rect 13820 24760 13872 24812
rect 14648 24760 14700 24812
rect 14832 24803 14884 24812
rect 14832 24769 14841 24803
rect 14841 24769 14875 24803
rect 14875 24769 14884 24803
rect 14832 24760 14884 24769
rect 15108 24760 15160 24812
rect 16304 24760 16356 24812
rect 16672 24760 16724 24812
rect 16856 24803 16908 24812
rect 16856 24769 16865 24803
rect 16865 24769 16899 24803
rect 16899 24769 16908 24803
rect 16856 24760 16908 24769
rect 16948 24803 17000 24812
rect 16948 24769 16957 24803
rect 16957 24769 16991 24803
rect 16991 24769 17000 24803
rect 16948 24760 17000 24769
rect 13084 24667 13136 24676
rect 9496 24599 9548 24608
rect 9496 24565 9505 24599
rect 9505 24565 9539 24599
rect 9539 24565 9548 24599
rect 9496 24556 9548 24565
rect 9956 24556 10008 24608
rect 10692 24556 10744 24608
rect 11336 24556 11388 24608
rect 12256 24556 12308 24608
rect 12440 24556 12492 24608
rect 13084 24633 13093 24667
rect 13093 24633 13127 24667
rect 13127 24633 13136 24667
rect 13084 24624 13136 24633
rect 13912 24692 13964 24744
rect 14924 24692 14976 24744
rect 15936 24624 15988 24676
rect 18236 24828 18288 24880
rect 17592 24803 17644 24812
rect 17592 24769 17601 24803
rect 17601 24769 17635 24803
rect 17635 24769 17644 24803
rect 17592 24760 17644 24769
rect 18052 24760 18104 24812
rect 18144 24803 18196 24812
rect 18144 24769 18153 24803
rect 18153 24769 18187 24803
rect 18187 24769 18196 24803
rect 18144 24760 18196 24769
rect 20260 24828 20312 24880
rect 18420 24803 18472 24812
rect 18420 24769 18429 24803
rect 18429 24769 18463 24803
rect 18463 24769 18472 24803
rect 18420 24760 18472 24769
rect 18052 24624 18104 24676
rect 19156 24803 19208 24812
rect 19156 24769 19165 24803
rect 19165 24769 19199 24803
rect 19199 24769 19208 24803
rect 19156 24760 19208 24769
rect 19340 24760 19392 24812
rect 19616 24760 19668 24812
rect 19892 24803 19944 24812
rect 19892 24769 19901 24803
rect 19901 24769 19935 24803
rect 19935 24769 19944 24803
rect 19892 24760 19944 24769
rect 19984 24760 20036 24812
rect 22560 24896 22612 24948
rect 22744 24939 22796 24948
rect 22744 24905 22753 24939
rect 22753 24905 22787 24939
rect 22787 24905 22796 24939
rect 22744 24896 22796 24905
rect 21364 24760 21416 24812
rect 21456 24827 21508 24836
rect 21456 24793 21465 24827
rect 21465 24793 21499 24827
rect 21499 24793 21508 24827
rect 21456 24784 21508 24793
rect 22100 24828 22152 24880
rect 22928 24828 22980 24880
rect 23756 24939 23808 24948
rect 23756 24905 23765 24939
rect 23765 24905 23799 24939
rect 23799 24905 23808 24939
rect 23756 24896 23808 24905
rect 24860 24896 24912 24948
rect 22192 24803 22244 24812
rect 22192 24769 22201 24803
rect 22201 24769 22235 24803
rect 22235 24769 22244 24803
rect 22192 24760 22244 24769
rect 22468 24803 22520 24812
rect 22468 24769 22477 24803
rect 22477 24769 22511 24803
rect 22511 24769 22520 24803
rect 22468 24760 22520 24769
rect 22560 24803 22612 24812
rect 22560 24769 22569 24803
rect 22569 24769 22603 24803
rect 22603 24769 22612 24803
rect 22560 24760 22612 24769
rect 23112 24760 23164 24812
rect 21456 24692 21508 24744
rect 12992 24599 13044 24608
rect 12992 24565 13001 24599
rect 13001 24565 13035 24599
rect 13035 24565 13044 24599
rect 12992 24556 13044 24565
rect 14372 24599 14424 24608
rect 14372 24565 14381 24599
rect 14381 24565 14415 24599
rect 14415 24565 14424 24599
rect 14372 24556 14424 24565
rect 14556 24599 14608 24608
rect 14556 24565 14565 24599
rect 14565 24565 14599 24599
rect 14599 24565 14608 24599
rect 14556 24556 14608 24565
rect 14648 24599 14700 24608
rect 14648 24565 14657 24599
rect 14657 24565 14691 24599
rect 14691 24565 14700 24599
rect 14648 24556 14700 24565
rect 17408 24556 17460 24608
rect 18236 24599 18288 24608
rect 18236 24565 18245 24599
rect 18245 24565 18279 24599
rect 18279 24565 18288 24599
rect 18236 24556 18288 24565
rect 19248 24599 19300 24608
rect 19248 24565 19257 24599
rect 19257 24565 19291 24599
rect 19291 24565 19300 24599
rect 19248 24556 19300 24565
rect 19432 24599 19484 24608
rect 19432 24565 19441 24599
rect 19441 24565 19475 24599
rect 19475 24565 19484 24599
rect 19432 24556 19484 24565
rect 19892 24556 19944 24608
rect 20168 24599 20220 24608
rect 20168 24565 20177 24599
rect 20177 24565 20211 24599
rect 20211 24565 20220 24599
rect 20168 24556 20220 24565
rect 20536 24556 20588 24608
rect 20720 24599 20772 24608
rect 20720 24565 20729 24599
rect 20729 24565 20763 24599
rect 20763 24565 20772 24599
rect 20720 24556 20772 24565
rect 21272 24624 21324 24676
rect 21824 24667 21876 24676
rect 21824 24633 21833 24667
rect 21833 24633 21867 24667
rect 21867 24633 21876 24667
rect 21824 24624 21876 24633
rect 22100 24624 22152 24676
rect 22744 24624 22796 24676
rect 23204 24735 23256 24744
rect 23204 24701 23213 24735
rect 23213 24701 23247 24735
rect 23247 24701 23256 24735
rect 23204 24692 23256 24701
rect 23480 24803 23532 24812
rect 23480 24769 23489 24803
rect 23489 24769 23523 24803
rect 23523 24769 23532 24803
rect 23480 24760 23532 24769
rect 24216 24828 24268 24880
rect 26700 24828 26752 24880
rect 23940 24760 23992 24812
rect 26792 24760 26844 24812
rect 24308 24692 24360 24744
rect 23848 24624 23900 24676
rect 25964 24624 26016 24676
rect 28080 24760 28132 24812
rect 28172 24803 28224 24812
rect 28172 24769 28181 24803
rect 28181 24769 28215 24803
rect 28215 24769 28224 24803
rect 28172 24760 28224 24769
rect 28264 24760 28316 24812
rect 29368 24760 29420 24812
rect 31576 24760 31628 24812
rect 31852 24803 31904 24812
rect 31852 24769 31861 24803
rect 31861 24769 31895 24803
rect 31895 24769 31904 24803
rect 31852 24760 31904 24769
rect 32220 24803 32272 24812
rect 32220 24769 32229 24803
rect 32229 24769 32263 24803
rect 32263 24769 32272 24803
rect 32220 24760 32272 24769
rect 28540 24692 28592 24744
rect 30472 24735 30524 24744
rect 30472 24701 30481 24735
rect 30481 24701 30515 24735
rect 30515 24701 30524 24735
rect 30472 24692 30524 24701
rect 28264 24624 28316 24676
rect 29644 24624 29696 24676
rect 21640 24599 21692 24608
rect 21640 24565 21649 24599
rect 21649 24565 21683 24599
rect 21683 24565 21692 24599
rect 21640 24556 21692 24565
rect 22836 24556 22888 24608
rect 23296 24599 23348 24608
rect 23296 24565 23305 24599
rect 23305 24565 23339 24599
rect 23339 24565 23348 24599
rect 23296 24556 23348 24565
rect 23388 24599 23440 24608
rect 23388 24565 23397 24599
rect 23397 24565 23431 24599
rect 23431 24565 23440 24599
rect 23388 24556 23440 24565
rect 24308 24556 24360 24608
rect 24492 24556 24544 24608
rect 25136 24556 25188 24608
rect 29184 24556 29236 24608
rect 32496 24556 32548 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 1676 24352 1728 24404
rect 2136 24395 2188 24404
rect 2136 24361 2145 24395
rect 2145 24361 2179 24395
rect 2179 24361 2188 24395
rect 2136 24352 2188 24361
rect 2688 24284 2740 24336
rect 3424 24352 3476 24404
rect 3700 24352 3752 24404
rect 4344 24352 4396 24404
rect 4712 24352 4764 24404
rect 5356 24395 5408 24404
rect 5356 24361 5365 24395
rect 5365 24361 5399 24395
rect 5399 24361 5408 24395
rect 5356 24352 5408 24361
rect 4160 24284 4212 24336
rect 6184 24352 6236 24404
rect 5632 24284 5684 24336
rect 6920 24352 6972 24404
rect 8944 24352 8996 24404
rect 9312 24352 9364 24404
rect 3148 24216 3200 24268
rect 3332 24216 3384 24268
rect 3976 24216 4028 24268
rect 848 24148 900 24200
rect 1860 24191 1912 24200
rect 1860 24157 1869 24191
rect 1869 24157 1903 24191
rect 1903 24157 1912 24191
rect 1860 24148 1912 24157
rect 2596 24191 2648 24200
rect 2596 24157 2605 24191
rect 2605 24157 2639 24191
rect 2639 24157 2648 24191
rect 2596 24148 2648 24157
rect 2688 24148 2740 24200
rect 2780 24080 2832 24132
rect 5448 24191 5500 24200
rect 5448 24157 5457 24191
rect 5457 24157 5491 24191
rect 5491 24157 5500 24191
rect 5448 24148 5500 24157
rect 6736 24284 6788 24336
rect 7656 24284 7708 24336
rect 9680 24284 9732 24336
rect 6000 24191 6052 24200
rect 6000 24157 6009 24191
rect 6009 24157 6043 24191
rect 6043 24157 6052 24191
rect 6000 24148 6052 24157
rect 6092 24191 6144 24200
rect 6092 24157 6101 24191
rect 6101 24157 6135 24191
rect 6135 24157 6144 24191
rect 6092 24148 6144 24157
rect 6552 24191 6604 24200
rect 6552 24157 6561 24191
rect 6561 24157 6595 24191
rect 6595 24157 6604 24191
rect 6552 24148 6604 24157
rect 6920 24191 6972 24200
rect 6920 24157 6929 24191
rect 6929 24157 6963 24191
rect 6963 24157 6972 24191
rect 6920 24148 6972 24157
rect 7012 24148 7064 24200
rect 7380 24148 7432 24200
rect 8668 24148 8720 24200
rect 8944 24191 8996 24200
rect 8944 24157 8953 24191
rect 8953 24157 8987 24191
rect 8987 24157 8996 24191
rect 8944 24148 8996 24157
rect 4804 24080 4856 24132
rect 3332 24055 3384 24064
rect 3332 24021 3341 24055
rect 3341 24021 3375 24055
rect 3375 24021 3384 24055
rect 3332 24012 3384 24021
rect 3424 24012 3476 24064
rect 5540 24080 5592 24132
rect 6736 24080 6788 24132
rect 6184 24012 6236 24064
rect 8852 24080 8904 24132
rect 7472 24055 7524 24064
rect 7472 24021 7481 24055
rect 7481 24021 7515 24055
rect 7515 24021 7524 24055
rect 7472 24012 7524 24021
rect 8484 24012 8536 24064
rect 9128 24123 9180 24132
rect 9128 24089 9137 24123
rect 9137 24089 9171 24123
rect 9171 24089 9180 24123
rect 9128 24080 9180 24089
rect 9312 24191 9364 24200
rect 9312 24157 9321 24191
rect 9321 24157 9355 24191
rect 9355 24157 9364 24191
rect 9312 24148 9364 24157
rect 10140 24216 10192 24268
rect 11152 24352 11204 24404
rect 11428 24352 11480 24404
rect 12992 24352 13044 24404
rect 16304 24352 16356 24404
rect 16396 24352 16448 24404
rect 18144 24352 18196 24404
rect 19340 24352 19392 24404
rect 20536 24352 20588 24404
rect 20812 24352 20864 24404
rect 11520 24284 11572 24336
rect 14464 24284 14516 24336
rect 15108 24284 15160 24336
rect 19616 24284 19668 24336
rect 21548 24352 21600 24404
rect 22192 24352 22244 24404
rect 22652 24352 22704 24404
rect 24860 24352 24912 24404
rect 25228 24352 25280 24404
rect 27896 24352 27948 24404
rect 28080 24395 28132 24404
rect 28080 24361 28089 24395
rect 28089 24361 28123 24395
rect 28123 24361 28132 24395
rect 28080 24352 28132 24361
rect 21180 24284 21232 24336
rect 9956 24012 10008 24064
rect 10508 24191 10560 24200
rect 10508 24157 10517 24191
rect 10517 24157 10551 24191
rect 10551 24157 10560 24191
rect 10508 24148 10560 24157
rect 10600 24191 10652 24200
rect 10600 24157 10609 24191
rect 10609 24157 10643 24191
rect 10643 24157 10652 24191
rect 10600 24148 10652 24157
rect 10692 24148 10744 24200
rect 10784 24080 10836 24132
rect 11244 24148 11296 24200
rect 13176 24216 13228 24268
rect 20168 24216 20220 24268
rect 21640 24216 21692 24268
rect 24216 24216 24268 24268
rect 14096 24148 14148 24200
rect 14188 24148 14240 24200
rect 20812 24148 20864 24200
rect 21180 24148 21232 24200
rect 11888 24080 11940 24132
rect 11428 24012 11480 24064
rect 11796 24055 11848 24064
rect 11796 24021 11805 24055
rect 11805 24021 11839 24055
rect 11839 24021 11848 24055
rect 11796 24012 11848 24021
rect 12624 24080 12676 24132
rect 13084 24080 13136 24132
rect 14280 24080 14332 24132
rect 23020 24148 23072 24200
rect 23664 24148 23716 24200
rect 25412 24191 25464 24200
rect 25412 24157 25421 24191
rect 25421 24157 25455 24191
rect 25455 24157 25464 24191
rect 25412 24148 25464 24157
rect 29920 24284 29972 24336
rect 28264 24259 28316 24268
rect 28264 24225 28273 24259
rect 28273 24225 28307 24259
rect 28307 24225 28316 24259
rect 28264 24216 28316 24225
rect 12808 24012 12860 24064
rect 13728 24012 13780 24064
rect 18880 24012 18932 24064
rect 19524 24012 19576 24064
rect 20996 24012 21048 24064
rect 21272 24055 21324 24064
rect 21272 24021 21281 24055
rect 21281 24021 21315 24055
rect 21315 24021 21324 24055
rect 21272 24012 21324 24021
rect 23572 24123 23624 24132
rect 23572 24089 23581 24123
rect 23581 24089 23615 24123
rect 23615 24089 23624 24123
rect 23572 24080 23624 24089
rect 23756 24123 23808 24132
rect 23756 24089 23765 24123
rect 23765 24089 23799 24123
rect 23799 24089 23808 24123
rect 23756 24080 23808 24089
rect 24676 24080 24728 24132
rect 28816 24191 28868 24200
rect 28816 24157 28825 24191
rect 28825 24157 28859 24191
rect 28859 24157 28868 24191
rect 28816 24148 28868 24157
rect 29368 24216 29420 24268
rect 32128 24259 32180 24268
rect 32128 24225 32137 24259
rect 32137 24225 32171 24259
rect 32171 24225 32180 24259
rect 32128 24216 32180 24225
rect 29184 24191 29236 24200
rect 29184 24157 29193 24191
rect 29193 24157 29227 24191
rect 29227 24157 29236 24191
rect 29184 24148 29236 24157
rect 29644 24148 29696 24200
rect 30656 24148 30708 24200
rect 30932 24148 30984 24200
rect 21916 24055 21968 24064
rect 21916 24021 21925 24055
rect 21925 24021 21959 24055
rect 21959 24021 21968 24055
rect 21916 24012 21968 24021
rect 23112 24012 23164 24064
rect 25136 24012 25188 24064
rect 25688 24012 25740 24064
rect 27712 24012 27764 24064
rect 27804 24012 27856 24064
rect 28540 24055 28592 24064
rect 28540 24021 28549 24055
rect 28549 24021 28583 24055
rect 28583 24021 28592 24055
rect 28540 24012 28592 24021
rect 30472 24080 30524 24132
rect 29184 24012 29236 24064
rect 29368 24055 29420 24064
rect 29368 24021 29377 24055
rect 29377 24021 29411 24055
rect 29411 24021 29420 24055
rect 29368 24012 29420 24021
rect 30288 24012 30340 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 2412 23808 2464 23860
rect 2964 23851 3016 23860
rect 2964 23817 2973 23851
rect 2973 23817 3007 23851
rect 3007 23817 3016 23851
rect 2964 23808 3016 23817
rect 3056 23851 3108 23860
rect 3056 23817 3065 23851
rect 3065 23817 3099 23851
rect 3099 23817 3108 23851
rect 3056 23808 3108 23817
rect 1860 23740 1912 23792
rect 3332 23740 3384 23792
rect 3976 23808 4028 23860
rect 5448 23808 5500 23860
rect 5908 23808 5960 23860
rect 10692 23808 10744 23860
rect 4344 23740 4396 23792
rect 4620 23740 4672 23792
rect 4712 23740 4764 23792
rect 2228 23672 2280 23724
rect 940 23604 992 23656
rect 1308 23604 1360 23656
rect 2412 23604 2464 23656
rect 2872 23672 2924 23724
rect 4068 23672 4120 23724
rect 2320 23536 2372 23588
rect 2780 23536 2832 23588
rect 3424 23579 3476 23588
rect 3424 23545 3433 23579
rect 3433 23545 3467 23579
rect 3467 23545 3476 23579
rect 3424 23536 3476 23545
rect 4344 23647 4396 23656
rect 4344 23613 4353 23647
rect 4353 23613 4387 23647
rect 4387 23613 4396 23647
rect 4344 23604 4396 23613
rect 4160 23536 4212 23588
rect 4804 23604 4856 23656
rect 5172 23715 5224 23724
rect 5172 23681 5181 23715
rect 5181 23681 5215 23715
rect 5215 23681 5224 23715
rect 5172 23672 5224 23681
rect 5356 23672 5408 23724
rect 5908 23715 5960 23724
rect 5908 23681 5917 23715
rect 5917 23681 5951 23715
rect 5951 23681 5960 23715
rect 5908 23672 5960 23681
rect 10140 23740 10192 23792
rect 6368 23672 6420 23724
rect 6920 23672 6972 23724
rect 7564 23672 7616 23724
rect 8484 23672 8536 23724
rect 8852 23672 8904 23724
rect 9036 23715 9088 23724
rect 9036 23681 9045 23715
rect 9045 23681 9079 23715
rect 9079 23681 9088 23715
rect 9036 23672 9088 23681
rect 9404 23672 9456 23724
rect 10508 23672 10560 23724
rect 11704 23808 11756 23860
rect 11428 23740 11480 23792
rect 12072 23851 12124 23860
rect 12072 23817 12081 23851
rect 12081 23817 12115 23851
rect 12115 23817 12124 23851
rect 12072 23808 12124 23817
rect 12992 23851 13044 23860
rect 12992 23817 13001 23851
rect 13001 23817 13035 23851
rect 13035 23817 13044 23851
rect 12992 23808 13044 23817
rect 14832 23808 14884 23860
rect 12440 23740 12492 23792
rect 16488 23740 16540 23792
rect 5264 23604 5316 23656
rect 9772 23604 9824 23656
rect 9956 23604 10008 23656
rect 10324 23604 10376 23656
rect 10968 23672 11020 23724
rect 17684 23740 17736 23792
rect 18144 23808 18196 23860
rect 20720 23808 20772 23860
rect 21732 23740 21784 23792
rect 25228 23808 25280 23860
rect 11612 23672 11664 23724
rect 11704 23715 11756 23724
rect 11704 23681 11713 23715
rect 11713 23681 11747 23715
rect 11747 23681 11756 23715
rect 11704 23672 11756 23681
rect 11888 23715 11940 23724
rect 11888 23681 11897 23715
rect 11897 23681 11931 23715
rect 11931 23681 11940 23715
rect 11888 23672 11940 23681
rect 11980 23672 12032 23724
rect 12624 23672 12676 23724
rect 12992 23672 13044 23724
rect 13176 23715 13228 23724
rect 13176 23681 13185 23715
rect 13185 23681 13219 23715
rect 13219 23681 13228 23715
rect 13176 23672 13228 23681
rect 13728 23672 13780 23724
rect 14188 23672 14240 23724
rect 14280 23715 14332 23724
rect 14280 23681 14289 23715
rect 14289 23681 14323 23715
rect 14323 23681 14332 23715
rect 14280 23672 14332 23681
rect 15108 23672 15160 23724
rect 15660 23715 15712 23724
rect 15660 23681 15669 23715
rect 15669 23681 15703 23715
rect 15703 23681 15712 23715
rect 15660 23672 15712 23681
rect 16120 23672 16172 23724
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 18972 23672 19024 23724
rect 19064 23672 19116 23724
rect 6368 23579 6420 23588
rect 6368 23545 6377 23579
rect 6377 23545 6411 23579
rect 6411 23545 6420 23579
rect 6368 23536 6420 23545
rect 7472 23536 7524 23588
rect 4896 23511 4948 23520
rect 4896 23477 4905 23511
rect 4905 23477 4939 23511
rect 4939 23477 4948 23511
rect 4896 23468 4948 23477
rect 5080 23468 5132 23520
rect 5356 23511 5408 23520
rect 5356 23477 5365 23511
rect 5365 23477 5399 23511
rect 5399 23477 5408 23511
rect 5356 23468 5408 23477
rect 5448 23511 5500 23520
rect 5448 23477 5457 23511
rect 5457 23477 5491 23511
rect 5491 23477 5500 23511
rect 5448 23468 5500 23477
rect 5724 23511 5776 23520
rect 5724 23477 5733 23511
rect 5733 23477 5767 23511
rect 5767 23477 5776 23511
rect 5724 23468 5776 23477
rect 6736 23468 6788 23520
rect 7564 23468 7616 23520
rect 8300 23468 8352 23520
rect 8760 23468 8812 23520
rect 9036 23468 9088 23520
rect 9772 23468 9824 23520
rect 11704 23468 11756 23520
rect 18604 23604 18656 23656
rect 18696 23604 18748 23656
rect 22284 23672 22336 23724
rect 14464 23536 14516 23588
rect 15108 23536 15160 23588
rect 15568 23536 15620 23588
rect 18052 23536 18104 23588
rect 13728 23468 13780 23520
rect 14188 23468 14240 23520
rect 15292 23468 15344 23520
rect 15752 23468 15804 23520
rect 17500 23468 17552 23520
rect 18788 23536 18840 23588
rect 18880 23536 18932 23588
rect 23940 23672 23992 23724
rect 24860 23740 24912 23792
rect 27804 23808 27856 23860
rect 28080 23808 28132 23860
rect 28356 23808 28408 23860
rect 30472 23851 30524 23860
rect 30472 23817 30481 23851
rect 30481 23817 30515 23851
rect 30515 23817 30524 23851
rect 30472 23808 30524 23817
rect 31852 23808 31904 23860
rect 26240 23740 26292 23792
rect 28816 23740 28868 23792
rect 29368 23740 29420 23792
rect 23296 23604 23348 23656
rect 18512 23468 18564 23520
rect 19340 23468 19392 23520
rect 19984 23468 20036 23520
rect 20720 23468 20772 23520
rect 23388 23536 23440 23588
rect 26056 23715 26108 23724
rect 26056 23681 26065 23715
rect 26065 23681 26099 23715
rect 26099 23681 26108 23715
rect 26056 23672 26108 23681
rect 25964 23604 26016 23656
rect 22192 23511 22244 23520
rect 22192 23477 22201 23511
rect 22201 23477 22235 23511
rect 22235 23477 22244 23511
rect 22192 23468 22244 23477
rect 23848 23511 23900 23520
rect 23848 23477 23857 23511
rect 23857 23477 23891 23511
rect 23891 23477 23900 23511
rect 23848 23468 23900 23477
rect 24032 23511 24084 23520
rect 24032 23477 24041 23511
rect 24041 23477 24075 23511
rect 24075 23477 24084 23511
rect 24032 23468 24084 23477
rect 25780 23468 25832 23520
rect 27804 23468 27856 23520
rect 27896 23468 27948 23520
rect 28724 23468 28776 23520
rect 29000 23468 29052 23520
rect 29460 23468 29512 23520
rect 30196 23715 30248 23724
rect 30196 23681 30205 23715
rect 30205 23681 30239 23715
rect 30239 23681 30248 23715
rect 30196 23672 30248 23681
rect 30288 23715 30340 23724
rect 30288 23681 30297 23715
rect 30297 23681 30331 23715
rect 30331 23681 30340 23715
rect 30288 23672 30340 23681
rect 30656 23672 30708 23724
rect 32588 23672 32640 23724
rect 30380 23536 30432 23588
rect 30564 23468 30616 23520
rect 32404 23511 32456 23520
rect 32404 23477 32413 23511
rect 32413 23477 32447 23511
rect 32447 23477 32456 23511
rect 32404 23468 32456 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 2044 23264 2096 23316
rect 3792 23264 3844 23316
rect 3884 23196 3936 23248
rect 2320 23103 2372 23112
rect 2320 23069 2329 23103
rect 2329 23069 2363 23103
rect 2363 23069 2372 23103
rect 2320 23060 2372 23069
rect 2780 23128 2832 23180
rect 5172 23264 5224 23316
rect 4436 23196 4488 23248
rect 4896 23196 4948 23248
rect 3148 23060 3200 23112
rect 4528 23128 4580 23180
rect 5356 23196 5408 23248
rect 2228 22992 2280 23044
rect 3976 23103 4028 23112
rect 3976 23069 3985 23103
rect 3985 23069 4019 23103
rect 4019 23069 4028 23103
rect 3976 23060 4028 23069
rect 3792 22992 3844 23044
rect 4620 23103 4672 23112
rect 4620 23069 4629 23103
rect 4629 23069 4663 23103
rect 4663 23069 4672 23103
rect 4620 23060 4672 23069
rect 4988 23060 5040 23112
rect 5264 23060 5316 23112
rect 5356 23103 5408 23112
rect 5356 23069 5365 23103
rect 5365 23069 5399 23103
rect 5399 23069 5408 23103
rect 5356 23060 5408 23069
rect 5908 23264 5960 23316
rect 6736 23264 6788 23316
rect 4804 22992 4856 23044
rect 6920 23196 6972 23248
rect 7196 23196 7248 23248
rect 7564 23264 7616 23316
rect 9680 23264 9732 23316
rect 11612 23264 11664 23316
rect 13820 23264 13872 23316
rect 7288 23128 7340 23180
rect 3148 22967 3200 22976
rect 3148 22933 3157 22967
rect 3157 22933 3191 22967
rect 3191 22933 3200 22967
rect 3148 22924 3200 22933
rect 3240 22924 3292 22976
rect 4896 22924 4948 22976
rect 5540 22924 5592 22976
rect 6092 23060 6144 23112
rect 6184 23060 6236 23112
rect 6552 23103 6604 23112
rect 6552 23069 6561 23103
rect 6561 23069 6595 23103
rect 6595 23069 6604 23103
rect 6552 23060 6604 23069
rect 6736 23103 6788 23112
rect 6736 23069 6745 23103
rect 6745 23069 6779 23103
rect 6779 23069 6788 23103
rect 6736 23060 6788 23069
rect 6828 23103 6880 23112
rect 6828 23069 6837 23103
rect 6837 23069 6871 23103
rect 6871 23069 6880 23103
rect 6828 23060 6880 23069
rect 6920 23103 6972 23112
rect 6920 23069 6929 23103
rect 6929 23069 6963 23103
rect 6963 23069 6972 23103
rect 6920 23060 6972 23069
rect 5908 22924 5960 22976
rect 6736 22924 6788 22976
rect 7564 23103 7616 23112
rect 7564 23069 7573 23103
rect 7573 23069 7607 23103
rect 7607 23069 7616 23103
rect 7564 23060 7616 23069
rect 7932 23128 7984 23180
rect 11796 23196 11848 23248
rect 14004 23196 14056 23248
rect 7840 23103 7892 23112
rect 7840 23069 7849 23103
rect 7849 23069 7883 23103
rect 7883 23069 7892 23103
rect 7840 23060 7892 23069
rect 8116 23103 8168 23112
rect 8116 23069 8125 23103
rect 8125 23069 8159 23103
rect 8159 23069 8168 23103
rect 8116 23060 8168 23069
rect 8208 23103 8260 23112
rect 8208 23069 8217 23103
rect 8217 23069 8251 23103
rect 8251 23069 8260 23103
rect 8208 23060 8260 23069
rect 10784 23103 10836 23112
rect 10784 23069 10793 23103
rect 10793 23069 10827 23103
rect 10827 23069 10836 23103
rect 10784 23060 10836 23069
rect 11060 23103 11112 23112
rect 11060 23069 11069 23103
rect 11069 23069 11103 23103
rect 11103 23069 11112 23103
rect 11060 23060 11112 23069
rect 11980 23060 12032 23112
rect 12808 23060 12860 23112
rect 7656 22924 7708 22976
rect 8300 22924 8352 22976
rect 11060 22924 11112 22976
rect 11244 22967 11296 22976
rect 11244 22933 11253 22967
rect 11253 22933 11287 22967
rect 11287 22933 11296 22967
rect 11244 22924 11296 22933
rect 11520 23035 11572 23044
rect 11520 23001 11529 23035
rect 11529 23001 11563 23035
rect 11563 23001 11572 23035
rect 11520 22992 11572 23001
rect 12072 22992 12124 23044
rect 11704 22967 11756 22976
rect 11704 22933 11713 22967
rect 11713 22933 11747 22967
rect 11747 22933 11756 22967
rect 11704 22924 11756 22933
rect 11888 22924 11940 22976
rect 12624 22924 12676 22976
rect 13452 23060 13504 23112
rect 16304 23264 16356 23316
rect 16580 23264 16632 23316
rect 17776 23307 17828 23316
rect 17776 23273 17785 23307
rect 17785 23273 17819 23307
rect 17819 23273 17828 23307
rect 17776 23264 17828 23273
rect 18052 23264 18104 23316
rect 16580 23128 16632 23180
rect 16856 23128 16908 23180
rect 17592 23128 17644 23180
rect 14004 22992 14056 23044
rect 14372 23103 14424 23112
rect 14372 23069 14381 23103
rect 14381 23069 14415 23103
rect 14415 23069 14424 23103
rect 14372 23060 14424 23069
rect 15016 23060 15068 23112
rect 15384 23060 15436 23112
rect 14556 22992 14608 23044
rect 15200 22992 15252 23044
rect 16396 23060 16448 23112
rect 18512 23171 18564 23180
rect 18512 23137 18521 23171
rect 18521 23137 18555 23171
rect 18555 23137 18564 23171
rect 18512 23128 18564 23137
rect 19708 23264 19760 23316
rect 20352 23264 20404 23316
rect 20720 23264 20772 23316
rect 21732 23307 21784 23316
rect 21732 23273 21741 23307
rect 21741 23273 21775 23307
rect 21775 23273 21784 23307
rect 21732 23264 21784 23273
rect 20812 23196 20864 23248
rect 20904 23196 20956 23248
rect 22560 23264 22612 23316
rect 22836 23264 22888 23316
rect 23572 23264 23624 23316
rect 24676 23307 24728 23316
rect 24676 23273 24685 23307
rect 24685 23273 24719 23307
rect 24719 23273 24728 23307
rect 24676 23264 24728 23273
rect 25044 23264 25096 23316
rect 25780 23307 25832 23316
rect 25780 23273 25789 23307
rect 25789 23273 25823 23307
rect 25823 23273 25832 23307
rect 25780 23264 25832 23273
rect 26240 23264 26292 23316
rect 26424 23307 26476 23316
rect 26424 23273 26433 23307
rect 26433 23273 26467 23307
rect 26467 23273 26476 23307
rect 26424 23264 26476 23273
rect 19524 23128 19576 23180
rect 19064 23060 19116 23112
rect 19156 23060 19208 23112
rect 22376 23128 22428 23180
rect 17592 23035 17644 23044
rect 17592 23001 17601 23035
rect 17601 23001 17635 23035
rect 17635 23001 17644 23035
rect 17592 22992 17644 23001
rect 17684 22992 17736 23044
rect 20260 23060 20312 23112
rect 21180 23060 21232 23112
rect 15660 22924 15712 22976
rect 16028 22924 16080 22976
rect 16396 22924 16448 22976
rect 16948 22924 17000 22976
rect 18236 22967 18288 22976
rect 18236 22933 18245 22967
rect 18245 22933 18279 22967
rect 18279 22933 18288 22967
rect 18236 22924 18288 22933
rect 18880 22967 18932 22976
rect 18880 22933 18889 22967
rect 18889 22933 18923 22967
rect 18923 22933 18932 22967
rect 18880 22924 18932 22933
rect 18972 22924 19024 22976
rect 20720 22992 20772 23044
rect 21824 23103 21876 23112
rect 21824 23069 21833 23103
rect 21833 23069 21867 23103
rect 21867 23069 21876 23103
rect 21824 23060 21876 23069
rect 22192 23060 22244 23112
rect 23296 23103 23348 23112
rect 23296 23069 23305 23103
rect 23305 23069 23339 23103
rect 23339 23069 23348 23103
rect 23296 23060 23348 23069
rect 25044 23128 25096 23180
rect 26056 23128 26108 23180
rect 26516 23171 26568 23180
rect 26516 23137 26525 23171
rect 26525 23137 26559 23171
rect 26559 23137 26568 23171
rect 26516 23128 26568 23137
rect 24492 23060 24544 23112
rect 19984 22924 20036 22976
rect 21916 22924 21968 22976
rect 22008 22967 22060 22976
rect 22008 22933 22017 22967
rect 22017 22933 22051 22967
rect 22051 22933 22060 22967
rect 22008 22924 22060 22933
rect 22100 22967 22152 22976
rect 22100 22933 22109 22967
rect 22109 22933 22143 22967
rect 22143 22933 22152 22967
rect 22100 22924 22152 22933
rect 22560 22992 22612 23044
rect 22652 23035 22704 23044
rect 22652 23001 22661 23035
rect 22661 23001 22695 23035
rect 22695 23001 22704 23035
rect 22652 22992 22704 23001
rect 24860 23060 24912 23112
rect 25504 23035 25556 23044
rect 25504 23001 25513 23035
rect 25513 23001 25547 23035
rect 25547 23001 25556 23035
rect 25504 22992 25556 23001
rect 25596 22992 25648 23044
rect 25964 23060 26016 23112
rect 26148 23060 26200 23112
rect 27160 23060 27212 23112
rect 32680 23264 32732 23316
rect 30656 23128 30708 23180
rect 28908 23103 28960 23112
rect 28908 23069 28917 23103
rect 28917 23069 28951 23103
rect 28951 23069 28960 23103
rect 28908 23060 28960 23069
rect 31760 23060 31812 23112
rect 26240 22992 26292 23044
rect 22744 22967 22796 22976
rect 22744 22933 22753 22967
rect 22753 22933 22787 22967
rect 22787 22933 22796 22967
rect 22744 22924 22796 22933
rect 22836 22924 22888 22976
rect 31484 22992 31536 23044
rect 29828 22924 29880 22976
rect 30104 22924 30156 22976
rect 32588 22924 32640 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 2320 22720 2372 22772
rect 2964 22720 3016 22772
rect 3056 22652 3108 22704
rect 3976 22695 4028 22704
rect 3976 22661 3985 22695
rect 3985 22661 4019 22695
rect 4019 22661 4028 22695
rect 3976 22652 4028 22661
rect 4436 22652 4488 22704
rect 1676 22627 1728 22636
rect 1676 22593 1710 22627
rect 1710 22593 1728 22627
rect 1676 22584 1728 22593
rect 2780 22584 2832 22636
rect 1400 22559 1452 22568
rect 1400 22525 1409 22559
rect 1409 22525 1443 22559
rect 1443 22525 1452 22559
rect 1400 22516 1452 22525
rect 3700 22516 3752 22568
rect 4804 22627 4856 22636
rect 4804 22593 4813 22627
rect 4813 22593 4847 22627
rect 4847 22593 4856 22627
rect 4804 22584 4856 22593
rect 4988 22627 5040 22636
rect 4988 22593 4997 22627
rect 4997 22593 5031 22627
rect 5031 22593 5040 22627
rect 4988 22584 5040 22593
rect 5080 22584 5132 22636
rect 2964 22448 3016 22500
rect 3792 22448 3844 22500
rect 4896 22516 4948 22568
rect 4712 22448 4764 22500
rect 4804 22448 4856 22500
rect 6092 22652 6144 22704
rect 6644 22720 6696 22772
rect 6736 22720 6788 22772
rect 7564 22720 7616 22772
rect 7840 22720 7892 22772
rect 9404 22720 9456 22772
rect 10692 22720 10744 22772
rect 11612 22720 11664 22772
rect 12348 22720 12400 22772
rect 12900 22720 12952 22772
rect 13360 22720 13412 22772
rect 13452 22720 13504 22772
rect 13820 22720 13872 22772
rect 18144 22720 18196 22772
rect 19156 22720 19208 22772
rect 19432 22720 19484 22772
rect 19616 22720 19668 22772
rect 20260 22720 20312 22772
rect 6552 22695 6604 22704
rect 6552 22661 6561 22695
rect 6561 22661 6595 22695
rect 6595 22661 6604 22695
rect 6552 22652 6604 22661
rect 5908 22584 5960 22636
rect 6276 22584 6328 22636
rect 5264 22380 5316 22432
rect 5356 22423 5408 22432
rect 5356 22389 5365 22423
rect 5365 22389 5399 22423
rect 5399 22389 5408 22423
rect 5356 22380 5408 22389
rect 6092 22448 6144 22500
rect 7196 22584 7248 22636
rect 7380 22584 7432 22636
rect 7840 22584 7892 22636
rect 9772 22652 9824 22704
rect 10508 22652 10560 22704
rect 8668 22584 8720 22636
rect 8852 22627 8904 22636
rect 8852 22593 8861 22627
rect 8861 22593 8895 22627
rect 8895 22593 8904 22627
rect 8852 22584 8904 22593
rect 8944 22627 8996 22636
rect 8944 22593 8977 22627
rect 8977 22593 8996 22627
rect 8944 22584 8996 22593
rect 9956 22516 10008 22568
rect 10232 22627 10284 22636
rect 10232 22593 10241 22627
rect 10241 22593 10275 22627
rect 10275 22593 10284 22627
rect 10232 22584 10284 22593
rect 11244 22584 11296 22636
rect 11888 22627 11940 22636
rect 11888 22593 11897 22627
rect 11897 22593 11931 22627
rect 11931 22593 11940 22627
rect 11888 22584 11940 22593
rect 12072 22627 12124 22636
rect 12072 22593 12081 22627
rect 12081 22593 12115 22627
rect 12115 22593 12124 22627
rect 12072 22584 12124 22593
rect 12256 22584 12308 22636
rect 13084 22652 13136 22704
rect 14280 22652 14332 22704
rect 20720 22720 20772 22772
rect 22468 22720 22520 22772
rect 23388 22720 23440 22772
rect 24768 22720 24820 22772
rect 25780 22720 25832 22772
rect 10968 22516 11020 22568
rect 11428 22516 11480 22568
rect 8944 22448 8996 22500
rect 9128 22491 9180 22500
rect 9128 22457 9137 22491
rect 9137 22457 9171 22491
rect 9171 22457 9180 22491
rect 9128 22448 9180 22457
rect 12624 22516 12676 22568
rect 13268 22516 13320 22568
rect 14372 22516 14424 22568
rect 12072 22448 12124 22500
rect 12256 22491 12308 22500
rect 12256 22457 12265 22491
rect 12265 22457 12299 22491
rect 12299 22457 12308 22491
rect 12256 22448 12308 22457
rect 12532 22448 12584 22500
rect 12900 22448 12952 22500
rect 14280 22448 14332 22500
rect 14556 22516 14608 22568
rect 20628 22652 20680 22704
rect 20996 22695 21048 22704
rect 20996 22661 21005 22695
rect 21005 22661 21039 22695
rect 21039 22661 21048 22695
rect 20996 22652 21048 22661
rect 27896 22652 27948 22704
rect 16488 22584 16540 22636
rect 17224 22584 17276 22636
rect 17500 22584 17552 22636
rect 17684 22584 17736 22636
rect 18696 22584 18748 22636
rect 16396 22516 16448 22568
rect 19340 22584 19392 22636
rect 19432 22627 19484 22636
rect 19432 22593 19441 22627
rect 19441 22593 19475 22627
rect 19475 22593 19484 22627
rect 19432 22584 19484 22593
rect 19524 22584 19576 22636
rect 18788 22448 18840 22500
rect 19616 22516 19668 22568
rect 19800 22627 19852 22636
rect 19800 22593 19809 22627
rect 19809 22593 19843 22627
rect 19843 22593 19852 22627
rect 19800 22584 19852 22593
rect 20168 22584 20220 22636
rect 7104 22380 7156 22432
rect 7196 22380 7248 22432
rect 8208 22380 8260 22432
rect 9680 22380 9732 22432
rect 9864 22380 9916 22432
rect 10784 22380 10836 22432
rect 11796 22423 11848 22432
rect 11796 22389 11805 22423
rect 11805 22389 11839 22423
rect 11839 22389 11848 22423
rect 11796 22380 11848 22389
rect 11980 22380 12032 22432
rect 12164 22380 12216 22432
rect 12716 22423 12768 22432
rect 12716 22389 12725 22423
rect 12725 22389 12759 22423
rect 12759 22389 12768 22423
rect 12716 22380 12768 22389
rect 12992 22380 13044 22432
rect 13360 22380 13412 22432
rect 14372 22380 14424 22432
rect 15476 22380 15528 22432
rect 16212 22423 16264 22432
rect 16212 22389 16221 22423
rect 16221 22389 16255 22423
rect 16255 22389 16264 22423
rect 16212 22380 16264 22389
rect 16396 22380 16448 22432
rect 17776 22423 17828 22432
rect 17776 22389 17785 22423
rect 17785 22389 17819 22423
rect 17819 22389 17828 22423
rect 17776 22380 17828 22389
rect 19524 22380 19576 22432
rect 19892 22559 19944 22568
rect 19892 22525 19901 22559
rect 19901 22525 19935 22559
rect 19935 22525 19944 22559
rect 19892 22516 19944 22525
rect 19984 22516 20036 22568
rect 20904 22516 20956 22568
rect 21180 22584 21232 22636
rect 22376 22584 22428 22636
rect 22744 22584 22796 22636
rect 25044 22627 25096 22636
rect 25044 22593 25053 22627
rect 25053 22593 25087 22627
rect 25087 22593 25096 22627
rect 25044 22584 25096 22593
rect 25228 22627 25280 22636
rect 25228 22593 25237 22627
rect 25237 22593 25271 22627
rect 25271 22593 25280 22627
rect 25228 22584 25280 22593
rect 27620 22627 27672 22636
rect 27620 22593 27629 22627
rect 27629 22593 27663 22627
rect 27663 22593 27672 22627
rect 27620 22584 27672 22593
rect 27988 22584 28040 22636
rect 29828 22584 29880 22636
rect 21640 22516 21692 22568
rect 20260 22423 20312 22432
rect 20260 22389 20269 22423
rect 20269 22389 20303 22423
rect 20303 22389 20312 22423
rect 20260 22380 20312 22389
rect 22560 22448 22612 22500
rect 20904 22423 20956 22432
rect 20904 22389 20913 22423
rect 20913 22389 20947 22423
rect 20947 22389 20956 22423
rect 20904 22380 20956 22389
rect 21272 22380 21324 22432
rect 22284 22423 22336 22432
rect 22284 22389 22293 22423
rect 22293 22389 22327 22423
rect 22327 22389 22336 22423
rect 22284 22380 22336 22389
rect 23020 22423 23072 22432
rect 23020 22389 23029 22423
rect 23029 22389 23063 22423
rect 23063 22389 23072 22423
rect 23020 22380 23072 22389
rect 27804 22423 27856 22432
rect 27804 22389 27813 22423
rect 27813 22389 27847 22423
rect 27847 22389 27856 22423
rect 27804 22380 27856 22389
rect 29828 22380 29880 22432
rect 30104 22627 30156 22636
rect 30104 22593 30113 22627
rect 30113 22593 30147 22627
rect 30147 22593 30156 22627
rect 30104 22584 30156 22593
rect 30932 22584 30984 22636
rect 32220 22627 32272 22636
rect 32220 22593 32229 22627
rect 32229 22593 32263 22627
rect 32263 22593 32272 22627
rect 32220 22584 32272 22593
rect 30380 22559 30432 22568
rect 30380 22525 30389 22559
rect 30389 22525 30423 22559
rect 30423 22525 30432 22559
rect 30380 22516 30432 22525
rect 31024 22380 31076 22432
rect 31760 22423 31812 22432
rect 31760 22389 31769 22423
rect 31769 22389 31803 22423
rect 31803 22389 31812 22423
rect 31760 22380 31812 22389
rect 32496 22380 32548 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 2228 22219 2280 22228
rect 2228 22185 2237 22219
rect 2237 22185 2271 22219
rect 2271 22185 2280 22219
rect 2228 22176 2280 22185
rect 4436 22176 4488 22228
rect 3148 22108 3200 22160
rect 2044 22015 2096 22024
rect 2044 21981 2053 22015
rect 2053 21981 2087 22015
rect 2087 21981 2096 22015
rect 2044 21972 2096 21981
rect 2688 21972 2740 22024
rect 3240 22040 3292 22092
rect 4712 22108 4764 22160
rect 3332 22015 3384 22024
rect 3332 21981 3341 22015
rect 3341 21981 3375 22015
rect 3375 21981 3384 22015
rect 3332 21972 3384 21981
rect 3884 22015 3936 22024
rect 3884 21981 3893 22015
rect 3893 21981 3927 22015
rect 3927 21981 3936 22015
rect 3884 21972 3936 21981
rect 3976 22015 4028 22024
rect 3976 21981 3985 22015
rect 3985 21981 4019 22015
rect 4019 21981 4028 22015
rect 3976 21972 4028 21981
rect 4528 21972 4580 22024
rect 4988 22176 5040 22228
rect 5540 22176 5592 22228
rect 5724 22176 5776 22228
rect 7840 22176 7892 22228
rect 8668 22176 8720 22228
rect 9404 22176 9456 22228
rect 12716 22176 12768 22228
rect 12808 22176 12860 22228
rect 13728 22176 13780 22228
rect 18972 22176 19024 22228
rect 20168 22176 20220 22228
rect 21180 22176 21232 22228
rect 22008 22176 22060 22228
rect 22652 22176 22704 22228
rect 23020 22176 23072 22228
rect 24952 22176 25004 22228
rect 5908 22151 5960 22160
rect 5908 22117 5917 22151
rect 5917 22117 5951 22151
rect 5951 22117 5960 22151
rect 5908 22108 5960 22117
rect 6920 22108 6972 22160
rect 3792 21904 3844 21956
rect 2320 21879 2372 21888
rect 2320 21845 2329 21879
rect 2329 21845 2363 21879
rect 2363 21845 2372 21879
rect 2320 21836 2372 21845
rect 2964 21836 3016 21888
rect 3056 21879 3108 21888
rect 3056 21845 3065 21879
rect 3065 21845 3099 21879
rect 3099 21845 3108 21879
rect 3056 21836 3108 21845
rect 3148 21879 3200 21888
rect 3148 21845 3157 21879
rect 3157 21845 3191 21879
rect 3191 21845 3200 21879
rect 3148 21836 3200 21845
rect 3332 21836 3384 21888
rect 3424 21836 3476 21888
rect 3700 21836 3752 21888
rect 4528 21836 4580 21888
rect 5264 21836 5316 21888
rect 5632 21972 5684 22024
rect 6000 22015 6052 22024
rect 6000 21981 6009 22015
rect 6009 21981 6043 22015
rect 6043 21981 6052 22015
rect 6000 21972 6052 21981
rect 6828 22015 6880 22024
rect 6828 21981 6837 22015
rect 6837 21981 6871 22015
rect 6871 21981 6880 22015
rect 6828 21972 6880 21981
rect 7196 22015 7248 22024
rect 7196 21981 7205 22015
rect 7205 21981 7239 22015
rect 7239 21981 7248 22015
rect 7196 21972 7248 21981
rect 8852 22108 8904 22160
rect 10140 22108 10192 22160
rect 8668 21972 8720 22024
rect 8944 22015 8996 22024
rect 8944 21981 8953 22015
rect 8953 21981 8987 22015
rect 8987 21981 8996 22015
rect 8944 21972 8996 21981
rect 11152 22083 11204 22092
rect 11152 22049 11161 22083
rect 11161 22049 11195 22083
rect 11195 22049 11204 22083
rect 11152 22040 11204 22049
rect 11980 22083 12032 22092
rect 11980 22049 11989 22083
rect 11989 22049 12023 22083
rect 12023 22049 12032 22083
rect 11980 22040 12032 22049
rect 12992 22108 13044 22160
rect 17132 22151 17184 22160
rect 17132 22117 17141 22151
rect 17141 22117 17175 22151
rect 17175 22117 17184 22151
rect 17132 22108 17184 22117
rect 9588 21972 9640 22024
rect 9680 21972 9732 22024
rect 9864 21972 9916 22024
rect 9956 21972 10008 22024
rect 5908 21904 5960 21956
rect 6092 21904 6144 21956
rect 9220 21904 9272 21956
rect 10876 22015 10928 22024
rect 10876 21981 10885 22015
rect 10885 21981 10919 22015
rect 10919 21981 10928 22015
rect 10876 21972 10928 21981
rect 11612 22015 11664 22024
rect 11612 21981 11621 22015
rect 11621 21981 11655 22015
rect 11655 21981 11664 22015
rect 11612 21972 11664 21981
rect 11888 21997 11897 22024
rect 11897 21997 11931 22024
rect 11931 21997 11940 22024
rect 11888 21972 11940 21997
rect 12164 21972 12216 22024
rect 12624 21972 12676 22024
rect 13636 22015 13688 22024
rect 13636 21981 13645 22015
rect 13645 21981 13679 22015
rect 13679 21981 13688 22015
rect 13636 21972 13688 21981
rect 14280 21972 14332 22024
rect 15752 22040 15804 22092
rect 18788 22040 18840 22092
rect 15660 21972 15712 22024
rect 17684 21972 17736 22024
rect 6184 21879 6236 21888
rect 6184 21845 6193 21879
rect 6193 21845 6227 21879
rect 6227 21845 6236 21879
rect 6184 21836 6236 21845
rect 8668 21836 8720 21888
rect 9312 21836 9364 21888
rect 9864 21879 9916 21888
rect 9864 21845 9873 21879
rect 9873 21845 9907 21879
rect 9907 21845 9916 21879
rect 9864 21836 9916 21845
rect 10692 21904 10744 21956
rect 10968 21904 11020 21956
rect 10508 21836 10560 21888
rect 11244 21879 11296 21888
rect 11244 21845 11253 21879
rect 11253 21845 11287 21879
rect 11287 21845 11296 21879
rect 11244 21836 11296 21845
rect 12348 21904 12400 21956
rect 13176 21904 13228 21956
rect 11520 21836 11572 21888
rect 12164 21836 12216 21888
rect 13820 21879 13872 21888
rect 13820 21845 13829 21879
rect 13829 21845 13863 21879
rect 13863 21845 13872 21879
rect 13820 21836 13872 21845
rect 15016 21947 15068 21956
rect 15016 21913 15025 21947
rect 15025 21913 15059 21947
rect 15059 21913 15068 21947
rect 15016 21904 15068 21913
rect 17592 21904 17644 21956
rect 19156 21972 19208 22024
rect 19616 22040 19668 22092
rect 19984 22108 20036 22160
rect 29828 22176 29880 22228
rect 30748 22176 30800 22228
rect 31484 22219 31536 22228
rect 31484 22185 31493 22219
rect 31493 22185 31527 22219
rect 31527 22185 31536 22219
rect 31484 22176 31536 22185
rect 20168 22040 20220 22092
rect 20260 22040 20312 22092
rect 20720 22040 20772 22092
rect 21180 22040 21232 22092
rect 21824 22040 21876 22092
rect 25412 22040 25464 22092
rect 25688 22040 25740 22092
rect 25872 22083 25924 22092
rect 25872 22049 25881 22083
rect 25881 22049 25915 22083
rect 25915 22049 25924 22083
rect 25872 22040 25924 22049
rect 32588 22040 32640 22092
rect 19892 21972 19944 22024
rect 20628 21972 20680 22024
rect 21364 21972 21416 22024
rect 17868 21904 17920 21956
rect 22192 22015 22244 22024
rect 22192 21981 22201 22015
rect 22201 21981 22235 22015
rect 22235 21981 22244 22015
rect 22192 21972 22244 21981
rect 22284 21972 22336 22024
rect 22560 21972 22612 22024
rect 23204 21972 23256 22024
rect 23940 22015 23992 22024
rect 23940 21981 23949 22015
rect 23949 21981 23983 22015
rect 23983 21981 23992 22015
rect 23940 21972 23992 21981
rect 25136 21972 25188 22024
rect 27068 21972 27120 22024
rect 30748 21972 30800 22024
rect 17684 21879 17736 21888
rect 17684 21845 17693 21879
rect 17693 21845 17727 21879
rect 17727 21845 17736 21879
rect 17684 21836 17736 21845
rect 17776 21836 17828 21888
rect 21364 21836 21416 21888
rect 22560 21836 22612 21888
rect 23112 21879 23164 21888
rect 23112 21845 23121 21879
rect 23121 21845 23155 21879
rect 23155 21845 23164 21879
rect 23112 21836 23164 21845
rect 23756 21947 23808 21956
rect 23756 21913 23765 21947
rect 23765 21913 23799 21947
rect 23799 21913 23808 21947
rect 23756 21904 23808 21913
rect 24400 21836 24452 21888
rect 25688 21904 25740 21956
rect 30748 21836 30800 21888
rect 31208 21947 31260 21956
rect 31208 21913 31217 21947
rect 31217 21913 31251 21947
rect 31251 21913 31260 21947
rect 31208 21904 31260 21913
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 2044 21632 2096 21684
rect 2964 21632 3016 21684
rect 2320 21564 2372 21616
rect 3516 21564 3568 21616
rect 3792 21632 3844 21684
rect 4436 21632 4488 21684
rect 5632 21632 5684 21684
rect 3976 21607 4028 21616
rect 3976 21573 3985 21607
rect 3985 21573 4019 21607
rect 4019 21573 4028 21607
rect 3976 21564 4028 21573
rect 6828 21632 6880 21684
rect 7932 21632 7984 21684
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 1492 21496 1544 21548
rect 2412 21360 2464 21412
rect 4068 21539 4120 21548
rect 4068 21505 4077 21539
rect 4077 21505 4111 21539
rect 4111 21505 4120 21539
rect 4068 21496 4120 21505
rect 3056 21428 3108 21480
rect 3976 21428 4028 21480
rect 4344 21539 4396 21548
rect 4344 21505 4353 21539
rect 4353 21505 4387 21539
rect 4387 21505 4396 21539
rect 4344 21496 4396 21505
rect 5264 21496 5316 21548
rect 6736 21607 6788 21616
rect 6736 21573 6745 21607
rect 6745 21573 6779 21607
rect 6779 21573 6788 21607
rect 6736 21564 6788 21573
rect 5724 21539 5776 21548
rect 5724 21505 5733 21539
rect 5733 21505 5767 21539
rect 5767 21505 5776 21539
rect 5724 21496 5776 21505
rect 5540 21428 5592 21480
rect 6460 21496 6512 21548
rect 8024 21564 8076 21616
rect 7012 21496 7064 21548
rect 7564 21496 7616 21548
rect 664 21292 716 21344
rect 1768 21292 1820 21344
rect 2688 21292 2740 21344
rect 5080 21360 5132 21412
rect 3516 21335 3568 21344
rect 3516 21301 3525 21335
rect 3525 21301 3559 21335
rect 3559 21301 3568 21335
rect 3516 21292 3568 21301
rect 3608 21292 3660 21344
rect 4068 21292 4120 21344
rect 4252 21335 4304 21344
rect 4252 21301 4261 21335
rect 4261 21301 4295 21335
rect 4295 21301 4304 21335
rect 4252 21292 4304 21301
rect 4712 21292 4764 21344
rect 5356 21292 5408 21344
rect 5448 21292 5500 21344
rect 6736 21428 6788 21480
rect 7840 21496 7892 21548
rect 9680 21564 9732 21616
rect 11060 21632 11112 21684
rect 11704 21632 11756 21684
rect 13268 21632 13320 21684
rect 13820 21632 13872 21684
rect 10508 21564 10560 21616
rect 9312 21539 9364 21548
rect 9312 21505 9321 21539
rect 9321 21505 9355 21539
rect 9355 21505 9364 21539
rect 9312 21496 9364 21505
rect 9588 21496 9640 21548
rect 10692 21496 10744 21548
rect 8576 21428 8628 21480
rect 5724 21360 5776 21412
rect 8760 21360 8812 21412
rect 9496 21360 9548 21412
rect 10416 21428 10468 21480
rect 10968 21539 11020 21548
rect 10968 21505 10977 21539
rect 10977 21505 11011 21539
rect 11011 21505 11020 21539
rect 10968 21496 11020 21505
rect 11612 21496 11664 21548
rect 11796 21496 11848 21548
rect 12072 21496 12124 21548
rect 12900 21496 12952 21548
rect 12992 21539 13044 21548
rect 12992 21505 13001 21539
rect 13001 21505 13035 21539
rect 13035 21505 13044 21539
rect 12992 21496 13044 21505
rect 13268 21496 13320 21548
rect 13360 21539 13412 21548
rect 13360 21505 13369 21539
rect 13369 21505 13403 21539
rect 13403 21505 13412 21539
rect 13360 21496 13412 21505
rect 15476 21496 15528 21548
rect 15844 21496 15896 21548
rect 17776 21564 17828 21616
rect 18788 21564 18840 21616
rect 12624 21428 12676 21480
rect 11428 21360 11480 21412
rect 6368 21292 6420 21344
rect 7288 21292 7340 21344
rect 7564 21292 7616 21344
rect 8024 21292 8076 21344
rect 8208 21292 8260 21344
rect 9680 21292 9732 21344
rect 9864 21292 9916 21344
rect 10232 21335 10284 21344
rect 10232 21301 10241 21335
rect 10241 21301 10275 21335
rect 10275 21301 10284 21335
rect 10232 21292 10284 21301
rect 11796 21292 11848 21344
rect 11980 21360 12032 21412
rect 13728 21428 13780 21480
rect 15200 21428 15252 21480
rect 12716 21292 12768 21344
rect 13176 21292 13228 21344
rect 14924 21360 14976 21412
rect 17408 21496 17460 21548
rect 17132 21428 17184 21480
rect 17776 21471 17828 21480
rect 17776 21437 17785 21471
rect 17785 21437 17819 21471
rect 17819 21437 17828 21471
rect 17776 21428 17828 21437
rect 18052 21496 18104 21548
rect 18236 21539 18288 21548
rect 18236 21505 18245 21539
rect 18245 21505 18279 21539
rect 18279 21505 18288 21539
rect 18236 21496 18288 21505
rect 18512 21496 18564 21548
rect 19340 21632 19392 21684
rect 19800 21632 19852 21684
rect 19156 21496 19208 21548
rect 19248 21539 19300 21548
rect 19248 21505 19257 21539
rect 19257 21505 19291 21539
rect 19291 21505 19300 21539
rect 19248 21496 19300 21505
rect 19340 21496 19392 21548
rect 19524 21539 19576 21548
rect 19524 21505 19533 21539
rect 19533 21505 19567 21539
rect 19567 21505 19576 21539
rect 19524 21496 19576 21505
rect 19892 21496 19944 21548
rect 20352 21632 20404 21684
rect 23848 21632 23900 21684
rect 20260 21564 20312 21616
rect 20812 21564 20864 21616
rect 23112 21564 23164 21616
rect 27620 21675 27672 21684
rect 27620 21641 27629 21675
rect 27629 21641 27663 21675
rect 27663 21641 27672 21675
rect 27620 21632 27672 21641
rect 27804 21632 27856 21684
rect 27988 21632 28040 21684
rect 29552 21632 29604 21684
rect 32220 21632 32272 21684
rect 18420 21428 18472 21480
rect 19432 21471 19484 21480
rect 19432 21437 19441 21471
rect 19441 21437 19475 21471
rect 19475 21437 19484 21471
rect 19432 21428 19484 21437
rect 20720 21471 20772 21480
rect 20720 21437 20729 21471
rect 20729 21437 20763 21471
rect 20763 21437 20772 21471
rect 20720 21428 20772 21437
rect 13636 21292 13688 21344
rect 14280 21292 14332 21344
rect 14740 21292 14792 21344
rect 16856 21335 16908 21344
rect 16856 21301 16865 21335
rect 16865 21301 16899 21335
rect 16899 21301 16908 21335
rect 16856 21292 16908 21301
rect 17408 21335 17460 21344
rect 17408 21301 17417 21335
rect 17417 21301 17451 21335
rect 17451 21301 17460 21335
rect 17408 21292 17460 21301
rect 17684 21335 17736 21344
rect 17684 21301 17693 21335
rect 17693 21301 17727 21335
rect 17727 21301 17736 21335
rect 17684 21292 17736 21301
rect 17776 21292 17828 21344
rect 18144 21335 18196 21344
rect 18144 21301 18153 21335
rect 18153 21301 18187 21335
rect 18187 21301 18196 21335
rect 18144 21292 18196 21301
rect 18420 21335 18472 21344
rect 18420 21301 18429 21335
rect 18429 21301 18463 21335
rect 18463 21301 18472 21335
rect 18420 21292 18472 21301
rect 19892 21360 19944 21412
rect 21180 21496 21232 21548
rect 24768 21539 24820 21548
rect 24768 21505 24777 21539
rect 24777 21505 24811 21539
rect 24811 21505 24820 21539
rect 24768 21496 24820 21505
rect 26976 21539 27028 21548
rect 26976 21505 26985 21539
rect 26985 21505 27019 21539
rect 27019 21505 27028 21539
rect 26976 21496 27028 21505
rect 27252 21539 27304 21548
rect 27252 21505 27261 21539
rect 27261 21505 27295 21539
rect 27295 21505 27304 21539
rect 27252 21496 27304 21505
rect 27528 21496 27580 21548
rect 30380 21564 30432 21616
rect 28356 21496 28408 21548
rect 28632 21496 28684 21548
rect 23480 21428 23532 21480
rect 24032 21471 24084 21480
rect 24032 21437 24041 21471
rect 24041 21437 24075 21471
rect 24075 21437 24084 21471
rect 24032 21428 24084 21437
rect 26516 21428 26568 21480
rect 27620 21428 27672 21480
rect 27988 21428 28040 21480
rect 24584 21360 24636 21412
rect 30288 21496 30340 21548
rect 31116 21564 31168 21616
rect 31300 21496 31352 21548
rect 32128 21496 32180 21548
rect 28816 21471 28868 21480
rect 28816 21437 28825 21471
rect 28825 21437 28859 21471
rect 28859 21437 28868 21471
rect 28816 21428 28868 21437
rect 19524 21335 19576 21344
rect 19524 21301 19533 21335
rect 19533 21301 19567 21335
rect 19567 21301 19576 21335
rect 19524 21292 19576 21301
rect 19800 21335 19852 21344
rect 19800 21301 19809 21335
rect 19809 21301 19843 21335
rect 19843 21301 19852 21335
rect 19800 21292 19852 21301
rect 20260 21335 20312 21344
rect 20260 21301 20269 21335
rect 20269 21301 20303 21335
rect 20303 21301 20312 21335
rect 20260 21292 20312 21301
rect 20812 21335 20864 21344
rect 20812 21301 20821 21335
rect 20821 21301 20855 21335
rect 20855 21301 20864 21335
rect 20812 21292 20864 21301
rect 23480 21292 23532 21344
rect 23848 21335 23900 21344
rect 23848 21301 23857 21335
rect 23857 21301 23891 21335
rect 23891 21301 23900 21335
rect 23848 21292 23900 21301
rect 24308 21292 24360 21344
rect 24400 21335 24452 21344
rect 24400 21301 24409 21335
rect 24409 21301 24443 21335
rect 24443 21301 24452 21335
rect 24400 21292 24452 21301
rect 24492 21335 24544 21344
rect 24492 21301 24501 21335
rect 24501 21301 24535 21335
rect 24535 21301 24544 21335
rect 24492 21292 24544 21301
rect 25504 21292 25556 21344
rect 25872 21292 25924 21344
rect 26608 21292 26660 21344
rect 27160 21292 27212 21344
rect 28172 21292 28224 21344
rect 28264 21335 28316 21344
rect 28264 21301 28273 21335
rect 28273 21301 28307 21335
rect 28307 21301 28316 21335
rect 28264 21292 28316 21301
rect 28724 21335 28776 21344
rect 28724 21301 28733 21335
rect 28733 21301 28767 21335
rect 28767 21301 28776 21335
rect 28724 21292 28776 21301
rect 32404 21335 32456 21344
rect 32404 21301 32413 21335
rect 32413 21301 32447 21335
rect 32447 21301 32456 21335
rect 32404 21292 32456 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 2228 21131 2280 21140
rect 2228 21097 2237 21131
rect 2237 21097 2271 21131
rect 2271 21097 2280 21131
rect 2228 21088 2280 21097
rect 3240 21088 3292 21140
rect 4436 21088 4488 21140
rect 4896 21088 4948 21140
rect 4988 21088 5040 21140
rect 6000 21088 6052 21140
rect 6092 21088 6144 21140
rect 1768 21020 1820 21072
rect 2412 21020 2464 21072
rect 2596 21020 2648 21072
rect 3148 21020 3200 21072
rect 4344 21020 4396 21072
rect 5540 21020 5592 21072
rect 3608 20952 3660 21004
rect 2044 20927 2096 20936
rect 2044 20893 2053 20927
rect 2053 20893 2087 20927
rect 2087 20893 2096 20927
rect 2044 20884 2096 20893
rect 2228 20884 2280 20936
rect 2412 20884 2464 20936
rect 3792 20884 3844 20936
rect 1676 20791 1728 20800
rect 1676 20757 1685 20791
rect 1685 20757 1719 20791
rect 1719 20757 1728 20791
rect 1676 20748 1728 20757
rect 3700 20816 3752 20868
rect 4988 20952 5040 21004
rect 5080 20952 5132 21004
rect 6460 21020 6512 21072
rect 7288 21020 7340 21072
rect 8208 21020 8260 21072
rect 8668 21088 8720 21140
rect 8944 21020 8996 21072
rect 9220 21088 9272 21140
rect 10508 21088 10560 21140
rect 11244 21088 11296 21140
rect 12716 21088 12768 21140
rect 12808 21131 12860 21140
rect 12808 21097 12817 21131
rect 12817 21097 12851 21131
rect 12851 21097 12860 21131
rect 12808 21088 12860 21097
rect 12992 21088 13044 21140
rect 13912 21088 13964 21140
rect 14740 21131 14792 21140
rect 14740 21097 14749 21131
rect 14749 21097 14783 21131
rect 14783 21097 14792 21131
rect 14740 21088 14792 21097
rect 15936 21088 15988 21140
rect 19800 21088 19852 21140
rect 20260 21088 20312 21140
rect 21180 21088 21232 21140
rect 21272 21088 21324 21140
rect 21548 21131 21600 21140
rect 21548 21097 21557 21131
rect 21557 21097 21591 21131
rect 21591 21097 21600 21131
rect 21548 21088 21600 21097
rect 22192 21088 22244 21140
rect 23480 21088 23532 21140
rect 24860 21088 24912 21140
rect 25320 21088 25372 21140
rect 25780 21131 25832 21140
rect 25780 21097 25789 21131
rect 25789 21097 25823 21131
rect 25823 21097 25832 21131
rect 25780 21088 25832 21097
rect 4252 20884 4304 20936
rect 4344 20927 4396 20936
rect 4344 20893 4353 20927
rect 4353 20893 4387 20927
rect 4387 20893 4396 20927
rect 4344 20884 4396 20893
rect 4712 20927 4764 20936
rect 4712 20893 4721 20927
rect 4721 20893 4755 20927
rect 4755 20893 4764 20927
rect 4712 20884 4764 20893
rect 5356 20884 5408 20936
rect 5448 20927 5500 20936
rect 5448 20893 5457 20927
rect 5457 20893 5491 20927
rect 5491 20893 5500 20927
rect 5448 20884 5500 20893
rect 5540 20884 5592 20936
rect 4896 20816 4948 20868
rect 6092 20927 6144 20936
rect 6092 20893 6101 20927
rect 6101 20893 6135 20927
rect 6135 20893 6144 20927
rect 6092 20884 6144 20893
rect 6368 20884 6420 20936
rect 8208 20927 8260 20936
rect 8208 20893 8217 20927
rect 8217 20893 8251 20927
rect 8251 20893 8260 20927
rect 8208 20884 8260 20893
rect 9220 20952 9272 21004
rect 10692 21020 10744 21072
rect 10416 20995 10468 21004
rect 10416 20961 10425 20995
rect 10425 20961 10459 20995
rect 10459 20961 10468 20995
rect 10416 20952 10468 20961
rect 10508 20952 10560 21004
rect 11704 20952 11756 21004
rect 5908 20859 5960 20868
rect 5908 20825 5917 20859
rect 5917 20825 5951 20859
rect 5951 20825 5960 20859
rect 5908 20816 5960 20825
rect 6000 20859 6052 20868
rect 6000 20825 6009 20859
rect 6009 20825 6043 20859
rect 6043 20825 6052 20859
rect 6000 20816 6052 20825
rect 2964 20748 3016 20800
rect 3148 20791 3200 20800
rect 3148 20757 3157 20791
rect 3157 20757 3191 20791
rect 3191 20757 3200 20791
rect 3148 20748 3200 20757
rect 3240 20791 3292 20800
rect 3240 20757 3249 20791
rect 3249 20757 3283 20791
rect 3283 20757 3292 20791
rect 3240 20748 3292 20757
rect 3424 20791 3476 20800
rect 3424 20757 3433 20791
rect 3433 20757 3467 20791
rect 3467 20757 3476 20791
rect 3424 20748 3476 20757
rect 3792 20791 3844 20800
rect 3792 20757 3801 20791
rect 3801 20757 3835 20791
rect 3835 20757 3844 20791
rect 3792 20748 3844 20757
rect 5264 20748 5316 20800
rect 5724 20748 5776 20800
rect 7840 20816 7892 20868
rect 7932 20816 7984 20868
rect 6276 20791 6328 20800
rect 6276 20757 6285 20791
rect 6285 20757 6319 20791
rect 6319 20757 6328 20791
rect 6276 20748 6328 20757
rect 6368 20748 6420 20800
rect 7380 20748 7432 20800
rect 8760 20816 8812 20868
rect 9220 20816 9272 20868
rect 12164 20952 12216 21004
rect 13360 21020 13412 21072
rect 12624 20952 12676 21004
rect 12808 20952 12860 21004
rect 14556 20952 14608 21004
rect 15476 21020 15528 21072
rect 9864 20816 9916 20868
rect 11980 20884 12032 20936
rect 12900 20927 12952 20936
rect 12900 20893 12909 20927
rect 12909 20893 12943 20927
rect 12943 20893 12952 20927
rect 12900 20884 12952 20893
rect 13360 20884 13412 20936
rect 13912 20884 13964 20936
rect 14464 20927 14516 20936
rect 14464 20893 14473 20927
rect 14473 20893 14507 20927
rect 14507 20893 14516 20927
rect 14464 20884 14516 20893
rect 14648 20927 14700 20936
rect 14648 20893 14657 20927
rect 14657 20893 14691 20927
rect 14691 20893 14700 20927
rect 14648 20884 14700 20893
rect 15936 20952 15988 21004
rect 16488 20952 16540 21004
rect 18420 20952 18472 21004
rect 13636 20816 13688 20868
rect 13820 20816 13872 20868
rect 18512 20884 18564 20936
rect 19708 20884 19760 20936
rect 20812 20952 20864 21004
rect 21180 20952 21232 21004
rect 22376 21020 22428 21072
rect 24308 21020 24360 21072
rect 26976 21088 27028 21140
rect 27068 21088 27120 21140
rect 27528 21088 27580 21140
rect 31300 21131 31352 21140
rect 31300 21097 31309 21131
rect 31309 21097 31343 21131
rect 31343 21097 31352 21131
rect 31300 21088 31352 21097
rect 22560 20952 22612 21004
rect 26424 21020 26476 21072
rect 27436 21020 27488 21072
rect 30748 21020 30800 21072
rect 30840 21020 30892 21072
rect 31024 21020 31076 21072
rect 30472 20952 30524 21004
rect 23112 20884 23164 20936
rect 24768 20884 24820 20936
rect 24860 20884 24912 20936
rect 25872 20927 25924 20936
rect 25872 20893 25881 20927
rect 25881 20893 25915 20927
rect 25915 20893 25924 20927
rect 25872 20884 25924 20893
rect 25964 20884 26016 20936
rect 26424 20884 26476 20936
rect 27436 20927 27488 20936
rect 27436 20893 27445 20927
rect 27445 20893 27479 20927
rect 27479 20893 27488 20927
rect 27436 20884 27488 20893
rect 28356 20884 28408 20936
rect 28816 20884 28868 20936
rect 30748 20927 30800 20936
rect 30748 20893 30757 20927
rect 30757 20893 30791 20927
rect 30791 20893 30800 20927
rect 30748 20884 30800 20893
rect 32220 20995 32272 21004
rect 32220 20961 32229 20995
rect 32229 20961 32263 20995
rect 32263 20961 32272 20995
rect 32220 20952 32272 20961
rect 31852 20884 31904 20936
rect 10232 20748 10284 20800
rect 11704 20748 11756 20800
rect 12072 20748 12124 20800
rect 14188 20748 14240 20800
rect 14464 20748 14516 20800
rect 15384 20748 15436 20800
rect 16120 20748 16172 20800
rect 18144 20748 18196 20800
rect 19432 20748 19484 20800
rect 20444 20748 20496 20800
rect 21548 20859 21600 20868
rect 21548 20825 21557 20859
rect 21557 20825 21591 20859
rect 21591 20825 21600 20859
rect 21548 20816 21600 20825
rect 21640 20816 21692 20868
rect 28724 20816 28776 20868
rect 31024 20859 31076 20868
rect 31024 20825 31033 20859
rect 31033 20825 31067 20859
rect 31067 20825 31076 20859
rect 31024 20816 31076 20825
rect 31208 20816 31260 20868
rect 24216 20748 24268 20800
rect 26608 20748 26660 20800
rect 30012 20748 30064 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 1676 20544 1728 20596
rect 3148 20544 3200 20596
rect 3240 20544 3292 20596
rect 3884 20544 3936 20596
rect 1768 20451 1820 20460
rect 1768 20417 1777 20451
rect 1777 20417 1811 20451
rect 1811 20417 1820 20451
rect 1768 20408 1820 20417
rect 3056 20476 3108 20528
rect 3516 20476 3568 20528
rect 3240 20408 3292 20460
rect 2320 20383 2372 20392
rect 2320 20349 2329 20383
rect 2329 20349 2363 20383
rect 2363 20349 2372 20383
rect 2320 20340 2372 20349
rect 2596 20340 2648 20392
rect 2688 20315 2740 20324
rect 2688 20281 2697 20315
rect 2697 20281 2731 20315
rect 2731 20281 2740 20315
rect 2688 20272 2740 20281
rect 3148 20272 3200 20324
rect 4436 20451 4488 20460
rect 4436 20417 4445 20451
rect 4445 20417 4479 20451
rect 4479 20417 4488 20451
rect 4436 20408 4488 20417
rect 4804 20476 4856 20528
rect 4068 20340 4120 20392
rect 2780 20204 2832 20256
rect 5448 20451 5500 20460
rect 5448 20417 5457 20451
rect 5457 20417 5491 20451
rect 5491 20417 5500 20451
rect 5448 20408 5500 20417
rect 6368 20476 6420 20528
rect 6920 20476 6972 20528
rect 5632 20408 5684 20460
rect 8208 20519 8260 20528
rect 8208 20485 8217 20519
rect 8217 20485 8251 20519
rect 8251 20485 8260 20519
rect 8208 20476 8260 20485
rect 8300 20451 8352 20460
rect 8300 20417 8309 20451
rect 8309 20417 8343 20451
rect 8343 20417 8352 20451
rect 8300 20408 8352 20417
rect 9772 20544 9824 20596
rect 10508 20544 10560 20596
rect 12440 20544 12492 20596
rect 10416 20408 10468 20460
rect 5356 20272 5408 20324
rect 3332 20204 3384 20256
rect 3792 20204 3844 20256
rect 5448 20204 5500 20256
rect 8852 20340 8904 20392
rect 6276 20272 6328 20324
rect 10508 20272 10560 20324
rect 6368 20204 6420 20256
rect 8852 20204 8904 20256
rect 9220 20204 9272 20256
rect 9864 20204 9916 20256
rect 10876 20340 10928 20392
rect 11428 20476 11480 20528
rect 13360 20544 13412 20596
rect 11704 20451 11756 20460
rect 11704 20417 11713 20451
rect 11713 20417 11747 20451
rect 11747 20417 11756 20451
rect 11704 20408 11756 20417
rect 11796 20451 11848 20460
rect 11796 20417 11805 20451
rect 11805 20417 11839 20451
rect 11839 20417 11848 20451
rect 11796 20408 11848 20417
rect 12256 20451 12308 20460
rect 12256 20417 12265 20451
rect 12265 20417 12299 20451
rect 12299 20417 12308 20451
rect 12256 20408 12308 20417
rect 15108 20544 15160 20596
rect 15752 20544 15804 20596
rect 14464 20476 14516 20528
rect 15200 20476 15252 20528
rect 16488 20544 16540 20596
rect 17040 20544 17092 20596
rect 16028 20476 16080 20528
rect 11428 20340 11480 20392
rect 12716 20340 12768 20392
rect 14648 20408 14700 20460
rect 15568 20408 15620 20460
rect 16488 20408 16540 20460
rect 16764 20408 16816 20460
rect 16948 20451 17000 20460
rect 16948 20417 16957 20451
rect 16957 20417 16991 20451
rect 16991 20417 17000 20451
rect 16948 20408 17000 20417
rect 17224 20408 17276 20460
rect 19340 20408 19392 20460
rect 19984 20451 20036 20460
rect 19984 20417 19993 20451
rect 19993 20417 20027 20451
rect 20027 20417 20036 20451
rect 19984 20408 20036 20417
rect 20260 20451 20312 20460
rect 20260 20417 20269 20451
rect 20269 20417 20303 20451
rect 20303 20417 20312 20451
rect 20260 20408 20312 20417
rect 20904 20476 20956 20528
rect 23940 20476 23992 20528
rect 30748 20544 30800 20596
rect 20720 20408 20772 20460
rect 21088 20451 21140 20460
rect 21088 20417 21097 20451
rect 21097 20417 21131 20451
rect 21131 20417 21140 20451
rect 21088 20408 21140 20417
rect 21640 20408 21692 20460
rect 22560 20451 22612 20460
rect 22560 20417 22569 20451
rect 22569 20417 22603 20451
rect 22603 20417 22612 20451
rect 22560 20408 22612 20417
rect 23296 20408 23348 20460
rect 30840 20519 30892 20528
rect 30840 20485 30849 20519
rect 30849 20485 30883 20519
rect 30883 20485 30892 20519
rect 30840 20476 30892 20485
rect 30932 20519 30984 20528
rect 30932 20485 30941 20519
rect 30941 20485 30975 20519
rect 30975 20485 30984 20519
rect 30932 20476 30984 20485
rect 14004 20383 14056 20392
rect 14004 20349 14013 20383
rect 14013 20349 14047 20383
rect 14047 20349 14056 20383
rect 14004 20340 14056 20349
rect 11152 20272 11204 20324
rect 11612 20272 11664 20324
rect 11704 20272 11756 20324
rect 11244 20204 11296 20256
rect 12440 20272 12492 20324
rect 12532 20315 12584 20324
rect 12532 20281 12541 20315
rect 12541 20281 12575 20315
rect 12575 20281 12584 20315
rect 12532 20272 12584 20281
rect 13636 20272 13688 20324
rect 14464 20340 14516 20392
rect 14740 20340 14792 20392
rect 14924 20340 14976 20392
rect 16304 20340 16356 20392
rect 13084 20204 13136 20256
rect 16764 20272 16816 20324
rect 17132 20315 17184 20324
rect 17132 20281 17141 20315
rect 17141 20281 17175 20315
rect 17175 20281 17184 20315
rect 17132 20272 17184 20281
rect 18328 20340 18380 20392
rect 19800 20340 19852 20392
rect 19892 20272 19944 20324
rect 22284 20340 22336 20392
rect 23020 20340 23072 20392
rect 24032 20340 24084 20392
rect 28724 20408 28776 20460
rect 30196 20408 30248 20460
rect 30380 20408 30432 20460
rect 30748 20408 30800 20460
rect 31760 20408 31812 20460
rect 26424 20340 26476 20392
rect 29736 20340 29788 20392
rect 21456 20272 21508 20324
rect 21640 20272 21692 20324
rect 14004 20247 14056 20256
rect 14004 20213 14013 20247
rect 14013 20213 14047 20247
rect 14047 20213 14056 20247
rect 14004 20204 14056 20213
rect 15384 20204 15436 20256
rect 15660 20247 15712 20256
rect 15660 20213 15669 20247
rect 15669 20213 15703 20247
rect 15703 20213 15712 20247
rect 15660 20204 15712 20213
rect 17776 20247 17828 20256
rect 17776 20213 17785 20247
rect 17785 20213 17819 20247
rect 17819 20213 17828 20247
rect 17776 20204 17828 20213
rect 19156 20204 19208 20256
rect 20352 20204 20404 20256
rect 20720 20204 20772 20256
rect 23020 20204 23072 20256
rect 24584 20272 24636 20324
rect 29184 20272 29236 20324
rect 29828 20272 29880 20324
rect 30104 20383 30156 20392
rect 30104 20349 30113 20383
rect 30113 20349 30147 20383
rect 30147 20349 30156 20383
rect 30104 20340 30156 20349
rect 32128 20340 32180 20392
rect 32496 20340 32548 20392
rect 24492 20204 24544 20256
rect 26884 20204 26936 20256
rect 27436 20204 27488 20256
rect 29460 20204 29512 20256
rect 29736 20204 29788 20256
rect 30012 20247 30064 20256
rect 30012 20213 30021 20247
rect 30021 20213 30055 20247
rect 30055 20213 30064 20247
rect 30012 20204 30064 20213
rect 30104 20204 30156 20256
rect 31208 20247 31260 20256
rect 31208 20213 31217 20247
rect 31217 20213 31251 20247
rect 31251 20213 31260 20247
rect 31208 20204 31260 20213
rect 32404 20247 32456 20256
rect 32404 20213 32413 20247
rect 32413 20213 32447 20247
rect 32447 20213 32456 20247
rect 32404 20204 32456 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 3976 20000 4028 20052
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 2964 19932 3016 19984
rect 3884 19932 3936 19984
rect 4896 20000 4948 20052
rect 8208 20043 8260 20052
rect 8208 20009 8217 20043
rect 8217 20009 8251 20043
rect 8251 20009 8260 20043
rect 8208 20000 8260 20009
rect 9404 20043 9456 20052
rect 9404 20009 9413 20043
rect 9413 20009 9447 20043
rect 9447 20009 9456 20043
rect 9404 20000 9456 20009
rect 12808 20000 12860 20052
rect 13636 20000 13688 20052
rect 2596 19796 2648 19848
rect 1676 19771 1728 19780
rect 1676 19737 1710 19771
rect 1710 19737 1728 19771
rect 1676 19728 1728 19737
rect 2320 19728 2372 19780
rect 3148 19839 3200 19848
rect 3148 19805 3157 19839
rect 3157 19805 3191 19839
rect 3191 19805 3200 19839
rect 3148 19796 3200 19805
rect 3240 19839 3292 19848
rect 3240 19805 3249 19839
rect 3249 19805 3283 19839
rect 3283 19805 3292 19839
rect 3240 19796 3292 19805
rect 5448 19932 5500 19984
rect 6276 19932 6328 19984
rect 6552 19932 6604 19984
rect 4896 19796 4948 19848
rect 7196 19864 7248 19916
rect 5356 19839 5408 19848
rect 5356 19805 5365 19839
rect 5365 19805 5399 19839
rect 5399 19805 5408 19839
rect 5356 19796 5408 19805
rect 5724 19796 5776 19848
rect 2412 19660 2464 19712
rect 4068 19728 4120 19780
rect 4804 19728 4856 19780
rect 5448 19728 5500 19780
rect 6368 19839 6420 19848
rect 6368 19805 6377 19839
rect 6377 19805 6411 19839
rect 6411 19805 6420 19839
rect 6368 19796 6420 19805
rect 6460 19839 6512 19848
rect 6460 19805 6469 19839
rect 6469 19805 6503 19839
rect 6503 19805 6512 19839
rect 6460 19796 6512 19805
rect 7564 19932 7616 19984
rect 14004 20000 14056 20052
rect 14648 20043 14700 20052
rect 14648 20009 14657 20043
rect 14657 20009 14691 20043
rect 14691 20009 14700 20043
rect 14648 20000 14700 20009
rect 16028 20000 16080 20052
rect 16488 20043 16540 20052
rect 16488 20009 16497 20043
rect 16497 20009 16531 20043
rect 16531 20009 16540 20043
rect 16488 20000 16540 20009
rect 17224 20000 17276 20052
rect 19616 20000 19668 20052
rect 20260 20000 20312 20052
rect 20720 20043 20772 20052
rect 20720 20009 20729 20043
rect 20729 20009 20763 20043
rect 20763 20009 20772 20043
rect 20720 20000 20772 20009
rect 20904 20043 20956 20052
rect 20904 20009 20913 20043
rect 20913 20009 20947 20043
rect 20947 20009 20956 20043
rect 20904 20000 20956 20009
rect 23664 20000 23716 20052
rect 24768 20043 24820 20052
rect 24768 20009 24777 20043
rect 24777 20009 24811 20043
rect 24811 20009 24820 20043
rect 24768 20000 24820 20009
rect 26056 20043 26108 20052
rect 26056 20009 26065 20043
rect 26065 20009 26099 20043
rect 26099 20009 26108 20043
rect 26056 20000 26108 20009
rect 26424 20000 26476 20052
rect 26700 20000 26752 20052
rect 26792 20043 26844 20052
rect 26792 20009 26801 20043
rect 26801 20009 26835 20043
rect 26835 20009 26844 20043
rect 26792 20000 26844 20009
rect 27896 20043 27948 20052
rect 27896 20009 27905 20043
rect 27905 20009 27939 20043
rect 27939 20009 27948 20043
rect 27896 20000 27948 20009
rect 29000 20000 29052 20052
rect 8116 19864 8168 19916
rect 7380 19839 7432 19848
rect 7380 19805 7389 19839
rect 7389 19805 7423 19839
rect 7423 19805 7432 19839
rect 7380 19796 7432 19805
rect 6000 19660 6052 19712
rect 8668 19796 8720 19848
rect 8944 19839 8996 19848
rect 8944 19805 8953 19839
rect 8953 19805 8987 19839
rect 8987 19805 8996 19839
rect 8944 19796 8996 19805
rect 9680 19864 9732 19916
rect 10232 19907 10284 19916
rect 10232 19873 10241 19907
rect 10241 19873 10275 19907
rect 10275 19873 10284 19907
rect 10232 19864 10284 19873
rect 11152 19864 11204 19916
rect 12072 19864 12124 19916
rect 12348 19864 12400 19916
rect 14464 19907 14516 19916
rect 14464 19873 14473 19907
rect 14473 19873 14507 19907
rect 14507 19873 14516 19907
rect 14464 19864 14516 19873
rect 6460 19660 6512 19712
rect 7380 19660 7432 19712
rect 7564 19703 7616 19712
rect 7564 19669 7573 19703
rect 7573 19669 7607 19703
rect 7607 19669 7616 19703
rect 7564 19660 7616 19669
rect 8760 19728 8812 19780
rect 9404 19660 9456 19712
rect 9588 19703 9640 19712
rect 9588 19669 9597 19703
rect 9597 19669 9631 19703
rect 9631 19669 9640 19703
rect 9588 19660 9640 19669
rect 9772 19728 9824 19780
rect 9956 19660 10008 19712
rect 10508 19815 10560 19848
rect 10508 19796 10517 19815
rect 10517 19796 10551 19815
rect 10551 19796 10560 19815
rect 11888 19796 11940 19848
rect 13360 19796 13412 19848
rect 13820 19796 13872 19848
rect 14188 19796 14240 19848
rect 14924 19796 14976 19848
rect 17040 19932 17092 19984
rect 15660 19864 15712 19916
rect 16488 19796 16540 19848
rect 16672 19839 16724 19848
rect 16672 19805 16681 19839
rect 16681 19805 16715 19839
rect 16715 19805 16724 19839
rect 16672 19796 16724 19805
rect 16764 19839 16816 19848
rect 16764 19805 16773 19839
rect 16773 19805 16807 19839
rect 16807 19805 16816 19839
rect 16764 19796 16816 19805
rect 19432 19864 19484 19916
rect 19892 19864 19944 19916
rect 19984 19796 20036 19848
rect 11796 19728 11848 19780
rect 12532 19728 12584 19780
rect 22192 19864 22244 19916
rect 23112 19864 23164 19916
rect 24492 19907 24544 19916
rect 24492 19873 24501 19907
rect 24501 19873 24535 19907
rect 24535 19873 24544 19907
rect 24492 19864 24544 19873
rect 24584 19864 24636 19916
rect 24952 19864 25004 19916
rect 25228 19864 25280 19916
rect 20996 19796 21048 19848
rect 21088 19839 21140 19848
rect 21088 19805 21097 19839
rect 21097 19805 21131 19839
rect 21131 19805 21140 19839
rect 21088 19796 21140 19805
rect 24124 19796 24176 19848
rect 25780 19839 25832 19848
rect 25780 19805 25789 19839
rect 25789 19805 25823 19839
rect 25823 19805 25832 19839
rect 25780 19796 25832 19805
rect 26056 19839 26108 19848
rect 26056 19805 26065 19839
rect 26065 19805 26099 19839
rect 26099 19805 26108 19839
rect 26056 19796 26108 19805
rect 26240 19907 26292 19916
rect 26240 19873 26249 19907
rect 26249 19873 26283 19907
rect 26283 19873 26292 19907
rect 26240 19864 26292 19873
rect 26700 19907 26752 19916
rect 26700 19873 26709 19907
rect 26709 19873 26743 19907
rect 26743 19873 26752 19907
rect 26700 19864 26752 19873
rect 26884 19932 26936 19984
rect 30564 20043 30616 20052
rect 30564 20009 30573 20043
rect 30573 20009 30607 20043
rect 30607 20009 30616 20043
rect 30564 20000 30616 20009
rect 30932 20000 30984 20052
rect 32496 20043 32548 20052
rect 32496 20009 32505 20043
rect 32505 20009 32539 20043
rect 32539 20009 32548 20043
rect 32496 20000 32548 20009
rect 28172 19864 28224 19916
rect 26424 19796 26476 19848
rect 10692 19660 10744 19712
rect 11980 19660 12032 19712
rect 12716 19660 12768 19712
rect 13268 19660 13320 19712
rect 13728 19660 13780 19712
rect 14004 19660 14056 19712
rect 14096 19660 14148 19712
rect 14188 19660 14240 19712
rect 14556 19660 14608 19712
rect 14648 19660 14700 19712
rect 21180 19728 21232 19780
rect 16672 19660 16724 19712
rect 17776 19660 17828 19712
rect 19892 19660 19944 19712
rect 25228 19660 25280 19712
rect 25320 19660 25372 19712
rect 26056 19660 26108 19712
rect 27988 19839 28040 19848
rect 27988 19805 27997 19839
rect 27997 19805 28031 19839
rect 28031 19805 28040 19839
rect 27988 19796 28040 19805
rect 28816 19796 28868 19848
rect 28080 19728 28132 19780
rect 28632 19771 28684 19780
rect 28632 19737 28641 19771
rect 28641 19737 28675 19771
rect 28675 19737 28684 19771
rect 28632 19728 28684 19737
rect 29184 19728 29236 19780
rect 29368 19796 29420 19848
rect 30380 19796 30432 19848
rect 31116 19839 31168 19848
rect 31116 19805 31125 19839
rect 31125 19805 31159 19839
rect 31159 19805 31168 19839
rect 31116 19796 31168 19805
rect 31208 19796 31260 19848
rect 29000 19660 29052 19712
rect 30104 19660 30156 19712
rect 30564 19660 30616 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 1676 19456 1728 19508
rect 2780 19456 2832 19508
rect 3792 19456 3844 19508
rect 4344 19456 4396 19508
rect 7380 19456 7432 19508
rect 7656 19456 7708 19508
rect 10508 19456 10560 19508
rect 1308 19320 1360 19372
rect 4068 19363 4120 19372
rect 4068 19329 4077 19363
rect 4077 19329 4111 19363
rect 4111 19329 4120 19363
rect 4068 19320 4120 19329
rect 4620 19388 4672 19440
rect 7472 19388 7524 19440
rect 8116 19388 8168 19440
rect 8576 19388 8628 19440
rect 8760 19388 8812 19440
rect 9680 19388 9732 19440
rect 9956 19388 10008 19440
rect 10876 19388 10928 19440
rect 11152 19388 11204 19440
rect 12808 19456 12860 19508
rect 13268 19456 13320 19508
rect 13360 19456 13412 19508
rect 13820 19456 13872 19508
rect 14924 19456 14976 19508
rect 16212 19499 16264 19508
rect 16212 19465 16221 19499
rect 16221 19465 16255 19499
rect 16255 19465 16264 19499
rect 16212 19456 16264 19465
rect 16488 19456 16540 19508
rect 17592 19456 17644 19508
rect 18972 19456 19024 19508
rect 23940 19456 23992 19508
rect 14648 19388 14700 19440
rect 5080 19320 5132 19372
rect 3976 19252 4028 19304
rect 3608 19184 3660 19236
rect 1216 19116 1268 19168
rect 3148 19116 3200 19168
rect 4068 19116 4120 19168
rect 4804 19116 4856 19168
rect 6000 19252 6052 19304
rect 7564 19252 7616 19304
rect 7932 19252 7984 19304
rect 10232 19320 10284 19372
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 12072 19320 12124 19372
rect 12532 19320 12584 19372
rect 11152 19252 11204 19304
rect 11520 19252 11572 19304
rect 7472 19184 7524 19236
rect 9956 19184 10008 19236
rect 11980 19252 12032 19304
rect 13268 19252 13320 19304
rect 14188 19320 14240 19372
rect 13912 19252 13964 19304
rect 15016 19431 15068 19440
rect 15016 19397 15025 19431
rect 15025 19397 15059 19431
rect 15059 19397 15068 19431
rect 15016 19388 15068 19397
rect 15200 19363 15252 19396
rect 15200 19344 15209 19363
rect 15209 19344 15243 19363
rect 15243 19344 15252 19363
rect 15752 19431 15804 19440
rect 15752 19397 15768 19431
rect 15768 19397 15802 19431
rect 15802 19397 15804 19431
rect 15752 19388 15804 19397
rect 20168 19388 20220 19440
rect 20352 19388 20404 19440
rect 15292 19363 15344 19372
rect 15292 19329 15317 19363
rect 15317 19329 15344 19363
rect 15292 19320 15344 19329
rect 6552 19116 6604 19168
rect 8484 19116 8536 19168
rect 12072 19184 12124 19236
rect 13084 19184 13136 19236
rect 14188 19184 14240 19236
rect 10968 19116 11020 19168
rect 11980 19116 12032 19168
rect 12624 19116 12676 19168
rect 13820 19116 13872 19168
rect 14832 19184 14884 19236
rect 16028 19363 16080 19372
rect 16028 19329 16037 19363
rect 16037 19329 16071 19363
rect 16071 19329 16080 19363
rect 16028 19320 16080 19329
rect 17684 19320 17736 19372
rect 18052 19320 18104 19372
rect 19984 19363 20036 19372
rect 19984 19329 19993 19363
rect 19993 19329 20027 19363
rect 20027 19329 20036 19363
rect 19984 19320 20036 19329
rect 20444 19320 20496 19372
rect 22560 19320 22612 19372
rect 23020 19320 23072 19372
rect 16580 19252 16632 19304
rect 20168 19252 20220 19304
rect 20812 19252 20864 19304
rect 24492 19320 24544 19372
rect 25044 19388 25096 19440
rect 25228 19388 25280 19440
rect 28172 19456 28224 19508
rect 29368 19499 29420 19508
rect 29368 19465 29377 19499
rect 29377 19465 29411 19499
rect 29411 19465 29420 19499
rect 29368 19456 29420 19465
rect 30380 19456 30432 19508
rect 26884 19388 26936 19440
rect 28724 19388 28776 19440
rect 24768 19320 24820 19372
rect 25044 19252 25096 19304
rect 25780 19363 25832 19372
rect 25780 19329 25789 19363
rect 25789 19329 25823 19363
rect 25823 19329 25832 19363
rect 25780 19320 25832 19329
rect 25964 19320 26016 19372
rect 26056 19320 26108 19372
rect 26240 19320 26292 19372
rect 26424 19363 26476 19372
rect 26424 19329 26433 19363
rect 26433 19329 26467 19363
rect 26467 19329 26476 19363
rect 26424 19320 26476 19329
rect 26792 19320 26844 19372
rect 28080 19320 28132 19372
rect 27528 19252 27580 19304
rect 29000 19320 29052 19372
rect 29460 19388 29512 19440
rect 30472 19388 30524 19440
rect 31024 19456 31076 19508
rect 32404 19499 32456 19508
rect 32404 19465 32413 19499
rect 32413 19465 32447 19499
rect 32447 19465 32456 19499
rect 32404 19456 32456 19465
rect 29184 19363 29236 19372
rect 29184 19329 29193 19363
rect 29193 19329 29227 19363
rect 29227 19329 29236 19363
rect 29184 19320 29236 19329
rect 29644 19320 29696 19372
rect 14464 19159 14516 19168
rect 14464 19125 14473 19159
rect 14473 19125 14507 19159
rect 14507 19125 14516 19159
rect 15108 19159 15160 19168
rect 14464 19116 14516 19125
rect 15108 19125 15117 19159
rect 15117 19125 15151 19159
rect 15151 19125 15160 19159
rect 15108 19116 15160 19125
rect 15200 19116 15252 19168
rect 17776 19184 17828 19236
rect 16120 19116 16172 19168
rect 17040 19116 17092 19168
rect 18880 19184 18932 19236
rect 19616 19184 19668 19236
rect 20076 19184 20128 19236
rect 19892 19116 19944 19168
rect 20168 19159 20220 19168
rect 20168 19125 20177 19159
rect 20177 19125 20211 19159
rect 20211 19125 20220 19159
rect 20168 19116 20220 19125
rect 20444 19184 20496 19236
rect 20996 19184 21048 19236
rect 22376 19116 22428 19168
rect 22744 19116 22796 19168
rect 23572 19116 23624 19168
rect 23940 19159 23992 19168
rect 23940 19125 23949 19159
rect 23949 19125 23983 19159
rect 23983 19125 23992 19159
rect 23940 19116 23992 19125
rect 24400 19159 24452 19168
rect 24400 19125 24409 19159
rect 24409 19125 24443 19159
rect 24443 19125 24452 19159
rect 24400 19116 24452 19125
rect 25872 19159 25924 19168
rect 25872 19125 25881 19159
rect 25881 19125 25915 19159
rect 25915 19125 25924 19159
rect 25872 19116 25924 19125
rect 26240 19116 26292 19168
rect 28632 19184 28684 19236
rect 29000 19184 29052 19236
rect 30564 19363 30616 19372
rect 30564 19329 30573 19363
rect 30573 19329 30607 19363
rect 30607 19329 30616 19363
rect 30564 19320 30616 19329
rect 30748 19320 30800 19372
rect 32220 19363 32272 19372
rect 32220 19329 32229 19363
rect 32229 19329 32263 19363
rect 32263 19329 32272 19363
rect 32220 19320 32272 19329
rect 27896 19116 27948 19168
rect 29368 19116 29420 19168
rect 29828 19116 29880 19168
rect 31208 19159 31260 19168
rect 31208 19125 31217 19159
rect 31217 19125 31251 19159
rect 31251 19125 31260 19159
rect 31208 19116 31260 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 2044 18912 2096 18964
rect 7472 18912 7524 18964
rect 7656 18912 7708 18964
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 1308 18708 1360 18760
rect 3332 18751 3384 18760
rect 3332 18717 3341 18751
rect 3341 18717 3375 18751
rect 3375 18717 3384 18751
rect 3332 18708 3384 18717
rect 3424 18751 3476 18760
rect 3424 18717 3433 18751
rect 3433 18717 3467 18751
rect 3467 18717 3476 18751
rect 3424 18708 3476 18717
rect 4068 18708 4120 18760
rect 4344 18776 4396 18828
rect 4712 18776 4764 18828
rect 5080 18776 5132 18828
rect 4804 18708 4856 18760
rect 5448 18708 5500 18760
rect 6184 18776 6236 18828
rect 6092 18751 6144 18760
rect 6092 18717 6101 18751
rect 6101 18717 6135 18751
rect 6135 18717 6144 18751
rect 6092 18708 6144 18717
rect 6736 18776 6788 18828
rect 8208 18776 8260 18828
rect 10048 18844 10100 18896
rect 10232 18955 10284 18964
rect 10232 18921 10241 18955
rect 10241 18921 10275 18955
rect 10275 18921 10284 18955
rect 10232 18912 10284 18921
rect 10508 18955 10560 18964
rect 10508 18921 10517 18955
rect 10517 18921 10551 18955
rect 10551 18921 10560 18955
rect 10508 18912 10560 18921
rect 11152 18912 11204 18964
rect 11888 18912 11940 18964
rect 10600 18844 10652 18896
rect 12072 18955 12124 18964
rect 12072 18921 12081 18955
rect 12081 18921 12115 18955
rect 12115 18921 12124 18955
rect 12072 18912 12124 18921
rect 12624 18955 12676 18964
rect 12624 18921 12633 18955
rect 12633 18921 12667 18955
rect 12667 18921 12676 18955
rect 12624 18912 12676 18921
rect 13268 18912 13320 18964
rect 14096 18912 14148 18964
rect 14464 18912 14516 18964
rect 15016 18912 15068 18964
rect 16488 18912 16540 18964
rect 16764 18912 16816 18964
rect 1676 18683 1728 18692
rect 1676 18649 1710 18683
rect 1710 18649 1728 18683
rect 1676 18640 1728 18649
rect 5724 18640 5776 18692
rect 7012 18751 7064 18760
rect 7012 18717 7021 18751
rect 7021 18717 7055 18751
rect 7055 18717 7064 18751
rect 7012 18708 7064 18717
rect 6736 18640 6788 18692
rect 3332 18572 3384 18624
rect 3608 18615 3660 18624
rect 3608 18581 3617 18615
rect 3617 18581 3651 18615
rect 3651 18581 3660 18615
rect 3608 18572 3660 18581
rect 3792 18615 3844 18624
rect 3792 18581 3801 18615
rect 3801 18581 3835 18615
rect 3835 18581 3844 18615
rect 3792 18572 3844 18581
rect 5356 18572 5408 18624
rect 7472 18751 7524 18760
rect 7472 18717 7481 18751
rect 7481 18717 7515 18751
rect 7515 18717 7524 18751
rect 7472 18708 7524 18717
rect 7932 18751 7984 18760
rect 7932 18717 7941 18751
rect 7941 18717 7975 18751
rect 7975 18717 7984 18751
rect 7932 18708 7984 18717
rect 8944 18708 8996 18760
rect 12532 18844 12584 18896
rect 9496 18751 9548 18760
rect 9496 18717 9505 18751
rect 9505 18717 9539 18751
rect 9539 18717 9548 18751
rect 9496 18708 9548 18717
rect 9680 18708 9732 18760
rect 10324 18751 10376 18760
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 8760 18640 8812 18692
rect 9220 18683 9272 18692
rect 9220 18649 9229 18683
rect 9229 18649 9263 18683
rect 9263 18649 9272 18683
rect 9220 18640 9272 18649
rect 9956 18640 10008 18692
rect 7472 18572 7524 18624
rect 7656 18615 7708 18624
rect 7656 18581 7665 18615
rect 7665 18581 7699 18615
rect 7699 18581 7708 18615
rect 7656 18572 7708 18581
rect 7748 18572 7800 18624
rect 12072 18776 12124 18828
rect 13268 18776 13320 18828
rect 11244 18708 11296 18760
rect 11060 18640 11112 18692
rect 12256 18708 12308 18760
rect 12624 18708 12676 18760
rect 12808 18751 12860 18760
rect 12808 18717 12817 18751
rect 12817 18717 12851 18751
rect 12851 18717 12860 18751
rect 12808 18708 12860 18717
rect 16580 18844 16632 18896
rect 14280 18776 14332 18828
rect 16304 18776 16356 18828
rect 14188 18751 14240 18760
rect 14188 18717 14197 18751
rect 14197 18717 14231 18751
rect 14231 18717 14240 18751
rect 14188 18708 14240 18717
rect 17500 18844 17552 18896
rect 17776 18912 17828 18964
rect 18696 18912 18748 18964
rect 21272 18955 21324 18964
rect 21272 18921 21281 18955
rect 21281 18921 21315 18955
rect 21315 18921 21324 18955
rect 21272 18912 21324 18921
rect 21916 18912 21968 18964
rect 11888 18572 11940 18624
rect 12624 18572 12676 18624
rect 14648 18683 14700 18692
rect 14648 18649 14657 18683
rect 14657 18649 14691 18683
rect 14691 18649 14700 18683
rect 14648 18640 14700 18649
rect 13728 18572 13780 18624
rect 22468 18955 22520 18964
rect 22468 18921 22477 18955
rect 22477 18921 22511 18955
rect 22511 18921 22520 18955
rect 22468 18912 22520 18921
rect 22652 18912 22704 18964
rect 22928 18912 22980 18964
rect 23388 18912 23440 18964
rect 22744 18844 22796 18896
rect 24124 18955 24176 18964
rect 24124 18921 24133 18955
rect 24133 18921 24167 18955
rect 24167 18921 24176 18955
rect 24124 18912 24176 18921
rect 24308 18912 24360 18964
rect 25872 18912 25924 18964
rect 26148 18912 26200 18964
rect 29828 18912 29880 18964
rect 30196 18912 30248 18964
rect 30288 18912 30340 18964
rect 31852 18912 31904 18964
rect 17500 18751 17552 18760
rect 17500 18717 17509 18751
rect 17509 18717 17543 18751
rect 17543 18717 17552 18751
rect 17500 18708 17552 18717
rect 17776 18751 17828 18760
rect 17776 18717 17785 18751
rect 17785 18717 17819 18751
rect 17819 18717 17828 18751
rect 17776 18708 17828 18717
rect 16764 18615 16816 18624
rect 16764 18581 16773 18615
rect 16773 18581 16807 18615
rect 16807 18581 16816 18615
rect 16764 18572 16816 18581
rect 17132 18572 17184 18624
rect 17500 18572 17552 18624
rect 18052 18572 18104 18624
rect 19248 18683 19300 18692
rect 19248 18649 19257 18683
rect 19257 18649 19291 18683
rect 19291 18649 19300 18683
rect 19248 18640 19300 18649
rect 19340 18640 19392 18692
rect 19892 18708 19944 18760
rect 20996 18708 21048 18760
rect 21456 18708 21508 18760
rect 20352 18640 20404 18692
rect 20536 18640 20588 18692
rect 21732 18819 21784 18828
rect 21732 18785 21741 18819
rect 21741 18785 21775 18819
rect 21775 18785 21784 18819
rect 21732 18776 21784 18785
rect 21824 18751 21876 18760
rect 21824 18717 21833 18751
rect 21833 18717 21867 18751
rect 21867 18717 21876 18751
rect 21824 18708 21876 18717
rect 20720 18572 20772 18624
rect 22468 18708 22520 18760
rect 23480 18776 23532 18828
rect 27528 18776 27580 18828
rect 30656 18776 30708 18828
rect 23112 18708 23164 18760
rect 22928 18640 22980 18692
rect 23848 18751 23900 18760
rect 23848 18717 23857 18751
rect 23857 18717 23891 18751
rect 23891 18717 23900 18751
rect 23848 18708 23900 18717
rect 23480 18683 23532 18692
rect 23480 18649 23489 18683
rect 23489 18649 23523 18683
rect 23523 18649 23532 18683
rect 23480 18640 23532 18649
rect 23572 18640 23624 18692
rect 25136 18751 25188 18760
rect 25136 18717 25145 18751
rect 25145 18717 25179 18751
rect 25179 18717 25188 18751
rect 25136 18708 25188 18717
rect 29000 18708 29052 18760
rect 29184 18708 29236 18760
rect 30104 18640 30156 18692
rect 28172 18572 28224 18624
rect 29184 18615 29236 18624
rect 29184 18581 29193 18615
rect 29193 18581 29227 18615
rect 29227 18581 29236 18615
rect 29184 18572 29236 18581
rect 30932 18708 30984 18760
rect 31208 18708 31260 18760
rect 31392 18572 31444 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 2596 18368 2648 18420
rect 3516 18411 3568 18420
rect 3516 18377 3525 18411
rect 3525 18377 3559 18411
rect 3559 18377 3568 18411
rect 3516 18368 3568 18377
rect 2872 18343 2924 18352
rect 2872 18309 2881 18343
rect 2881 18309 2915 18343
rect 2915 18309 2924 18343
rect 2872 18300 2924 18309
rect 4620 18368 4672 18420
rect 7932 18368 7984 18420
rect 8116 18368 8168 18420
rect 2688 18275 2740 18284
rect 2688 18241 2697 18275
rect 2697 18241 2731 18275
rect 2731 18241 2740 18275
rect 2688 18232 2740 18241
rect 3056 18232 3108 18284
rect 3332 18275 3384 18284
rect 3332 18241 3341 18275
rect 3341 18241 3375 18275
rect 3375 18241 3384 18275
rect 3332 18232 3384 18241
rect 3700 18232 3752 18284
rect 4344 18275 4396 18284
rect 4344 18241 4353 18275
rect 4353 18241 4387 18275
rect 4387 18241 4396 18275
rect 4344 18232 4396 18241
rect 4620 18232 4672 18284
rect 4896 18232 4948 18284
rect 3516 18164 3568 18216
rect 4712 18164 4764 18216
rect 5356 18300 5408 18352
rect 6460 18300 6512 18352
rect 8944 18368 8996 18420
rect 9864 18368 9916 18420
rect 11704 18368 11756 18420
rect 11888 18368 11940 18420
rect 12164 18411 12216 18420
rect 12164 18377 12173 18411
rect 12173 18377 12207 18411
rect 12207 18377 12216 18411
rect 12164 18368 12216 18377
rect 12440 18368 12492 18420
rect 12716 18368 12768 18420
rect 12900 18368 12952 18420
rect 14280 18368 14332 18420
rect 15292 18368 15344 18420
rect 17224 18368 17276 18420
rect 17316 18368 17368 18420
rect 20260 18368 20312 18420
rect 5632 18232 5684 18284
rect 6276 18164 6328 18216
rect 6552 18164 6604 18216
rect 7748 18275 7800 18284
rect 7748 18241 7757 18275
rect 7757 18241 7791 18275
rect 7791 18241 7800 18275
rect 7748 18232 7800 18241
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 7932 18164 7984 18216
rect 8116 18164 8168 18216
rect 7012 18096 7064 18148
rect 7472 18096 7524 18148
rect 3608 18028 3660 18080
rect 3700 18028 3752 18080
rect 6092 18028 6144 18080
rect 7840 18096 7892 18148
rect 9404 18232 9456 18284
rect 10876 18300 10928 18352
rect 11520 18232 11572 18284
rect 11796 18232 11848 18284
rect 11888 18232 11940 18284
rect 12164 18232 12216 18284
rect 8668 18164 8720 18216
rect 11244 18164 11296 18216
rect 12256 18164 12308 18216
rect 12532 18164 12584 18216
rect 16120 18300 16172 18352
rect 16856 18300 16908 18352
rect 14740 18232 14792 18284
rect 14832 18275 14884 18284
rect 14832 18241 14841 18275
rect 14841 18241 14875 18275
rect 14875 18241 14884 18275
rect 14832 18232 14884 18241
rect 15476 18232 15528 18284
rect 15660 18232 15712 18284
rect 17224 18275 17276 18284
rect 17224 18241 17233 18275
rect 17233 18241 17267 18275
rect 17267 18241 17276 18275
rect 17224 18232 17276 18241
rect 18604 18300 18656 18352
rect 18788 18232 18840 18284
rect 14648 18207 14700 18216
rect 14648 18173 14657 18207
rect 14657 18173 14691 18207
rect 14691 18173 14700 18207
rect 14648 18164 14700 18173
rect 16764 18164 16816 18216
rect 10508 18096 10560 18148
rect 11520 18096 11572 18148
rect 12348 18096 12400 18148
rect 17776 18164 17828 18216
rect 8760 18028 8812 18080
rect 10600 18028 10652 18080
rect 17500 18096 17552 18148
rect 18972 18275 19024 18284
rect 18972 18241 18981 18275
rect 18981 18241 19015 18275
rect 19015 18241 19024 18275
rect 18972 18232 19024 18241
rect 19892 18300 19944 18352
rect 21456 18368 21508 18420
rect 21824 18368 21876 18420
rect 23848 18411 23900 18420
rect 23848 18377 23857 18411
rect 23857 18377 23891 18411
rect 23891 18377 23900 18411
rect 23848 18368 23900 18377
rect 28908 18368 28960 18420
rect 30472 18411 30524 18420
rect 30472 18377 30481 18411
rect 30481 18377 30515 18411
rect 30515 18377 30524 18411
rect 30472 18368 30524 18377
rect 32220 18368 32272 18420
rect 21180 18300 21232 18352
rect 22744 18300 22796 18352
rect 19524 18232 19576 18284
rect 20076 18232 20128 18284
rect 20260 18232 20312 18284
rect 23480 18275 23532 18284
rect 23480 18241 23489 18275
rect 23489 18241 23523 18275
rect 23523 18241 23532 18275
rect 23480 18232 23532 18241
rect 26148 18232 26200 18284
rect 27528 18232 27580 18284
rect 27712 18232 27764 18284
rect 27896 18275 27948 18284
rect 27896 18241 27905 18275
rect 27905 18241 27939 18275
rect 27939 18241 27948 18275
rect 27896 18232 27948 18241
rect 21456 18096 21508 18148
rect 22192 18096 22244 18148
rect 28264 18232 28316 18284
rect 29276 18164 29328 18216
rect 30288 18275 30340 18284
rect 30288 18241 30297 18275
rect 30297 18241 30331 18275
rect 30331 18241 30340 18275
rect 30288 18232 30340 18241
rect 30656 18232 30708 18284
rect 31392 18232 31444 18284
rect 13360 18028 13412 18080
rect 14464 18028 14516 18080
rect 15016 18028 15068 18080
rect 15200 18071 15252 18080
rect 15200 18037 15209 18071
rect 15209 18037 15243 18071
rect 15243 18037 15252 18071
rect 15200 18028 15252 18037
rect 18052 18028 18104 18080
rect 18696 18071 18748 18080
rect 18696 18037 18705 18071
rect 18705 18037 18739 18071
rect 18739 18037 18748 18071
rect 18696 18028 18748 18037
rect 19524 18028 19576 18080
rect 19984 18028 20036 18080
rect 20628 18028 20680 18080
rect 20996 18028 21048 18080
rect 22376 18028 22428 18080
rect 25412 18028 25464 18080
rect 26700 18028 26752 18080
rect 27896 18071 27948 18080
rect 27896 18037 27905 18071
rect 27905 18037 27939 18071
rect 27939 18037 27948 18071
rect 27896 18028 27948 18037
rect 29644 18028 29696 18080
rect 32404 18071 32456 18080
rect 32404 18037 32413 18071
rect 32413 18037 32447 18071
rect 32447 18037 32456 18071
rect 32404 18028 32456 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 2688 17867 2740 17876
rect 2688 17833 2697 17867
rect 2697 17833 2731 17867
rect 2731 17833 2740 17867
rect 2688 17824 2740 17833
rect 5356 17824 5408 17876
rect 7840 17824 7892 17876
rect 11152 17824 11204 17876
rect 11428 17824 11480 17876
rect 11612 17824 11664 17876
rect 12072 17824 12124 17876
rect 12440 17867 12492 17876
rect 12440 17833 12449 17867
rect 12449 17833 12483 17867
rect 12483 17833 12492 17867
rect 12440 17824 12492 17833
rect 12716 17824 12768 17876
rect 13084 17824 13136 17876
rect 5448 17756 5500 17808
rect 6368 17756 6420 17808
rect 3700 17688 3752 17740
rect 3148 17663 3200 17672
rect 3148 17629 3157 17663
rect 3157 17629 3191 17663
rect 3191 17629 3200 17663
rect 3148 17620 3200 17629
rect 3424 17663 3476 17672
rect 3424 17629 3433 17663
rect 3433 17629 3467 17663
rect 3467 17629 3476 17663
rect 3424 17620 3476 17629
rect 3700 17552 3752 17604
rect 4160 17663 4212 17672
rect 4160 17629 4169 17663
rect 4169 17629 4203 17663
rect 4203 17629 4212 17663
rect 4160 17620 4212 17629
rect 4620 17620 4672 17672
rect 4988 17688 5040 17740
rect 7288 17688 7340 17740
rect 7656 17756 7708 17808
rect 8024 17756 8076 17808
rect 8760 17756 8812 17808
rect 10508 17756 10560 17808
rect 10876 17756 10928 17808
rect 11980 17756 12032 17808
rect 9680 17688 9732 17740
rect 11612 17688 11664 17740
rect 12532 17756 12584 17808
rect 12992 17756 13044 17808
rect 12348 17688 12400 17740
rect 14648 17867 14700 17876
rect 14648 17833 14657 17867
rect 14657 17833 14691 17867
rect 14691 17833 14700 17867
rect 14648 17824 14700 17833
rect 14740 17756 14792 17808
rect 14832 17799 14884 17808
rect 14832 17765 14841 17799
rect 14841 17765 14875 17799
rect 14875 17765 14884 17799
rect 14832 17756 14884 17765
rect 4896 17620 4948 17672
rect 5540 17663 5592 17672
rect 5540 17629 5549 17663
rect 5549 17629 5583 17663
rect 5583 17629 5592 17663
rect 5540 17620 5592 17629
rect 6460 17620 6512 17672
rect 6552 17620 6604 17672
rect 7840 17620 7892 17672
rect 8576 17620 8628 17672
rect 10416 17620 10468 17672
rect 10508 17663 10560 17672
rect 10508 17629 10517 17663
rect 10517 17629 10551 17663
rect 10551 17629 10560 17663
rect 10508 17620 10560 17629
rect 11796 17620 11848 17672
rect 4252 17595 4304 17604
rect 4252 17561 4261 17595
rect 4261 17561 4295 17595
rect 4295 17561 4304 17595
rect 4252 17552 4304 17561
rect 2688 17484 2740 17536
rect 3148 17484 3200 17536
rect 3240 17527 3292 17536
rect 3240 17493 3249 17527
rect 3249 17493 3283 17527
rect 3283 17493 3292 17527
rect 3240 17484 3292 17493
rect 4620 17527 4672 17536
rect 4620 17493 4629 17527
rect 4629 17493 4663 17527
rect 4663 17493 4672 17527
rect 4620 17484 4672 17493
rect 7196 17552 7248 17604
rect 5356 17527 5408 17536
rect 5356 17493 5365 17527
rect 5365 17493 5399 17527
rect 5399 17493 5408 17527
rect 5356 17484 5408 17493
rect 5632 17527 5684 17536
rect 5632 17493 5641 17527
rect 5641 17493 5675 17527
rect 5675 17493 5684 17527
rect 5632 17484 5684 17493
rect 6460 17484 6512 17536
rect 9128 17484 9180 17536
rect 10232 17527 10284 17536
rect 10232 17493 10241 17527
rect 10241 17493 10275 17527
rect 10275 17493 10284 17527
rect 10232 17484 10284 17493
rect 10324 17527 10376 17536
rect 10324 17493 10333 17527
rect 10333 17493 10367 17527
rect 10367 17493 10376 17527
rect 10324 17484 10376 17493
rect 12716 17663 12768 17672
rect 12716 17629 12725 17663
rect 12725 17629 12759 17663
rect 12759 17629 12768 17663
rect 12716 17620 12768 17629
rect 12348 17484 12400 17536
rect 12808 17552 12860 17604
rect 13268 17663 13320 17672
rect 13268 17629 13277 17663
rect 13277 17629 13311 17663
rect 13311 17629 13320 17663
rect 13268 17620 13320 17629
rect 14280 17663 14332 17672
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 14280 17620 14332 17629
rect 14464 17731 14516 17740
rect 14464 17697 14473 17731
rect 14473 17697 14507 17731
rect 14507 17697 14516 17731
rect 14464 17688 14516 17697
rect 15200 17824 15252 17876
rect 17316 17867 17368 17876
rect 17316 17833 17325 17867
rect 17325 17833 17359 17867
rect 17359 17833 17368 17867
rect 17316 17824 17368 17833
rect 18052 17824 18104 17876
rect 15292 17756 15344 17808
rect 20260 17824 20312 17876
rect 22192 17824 22244 17876
rect 22652 17824 22704 17876
rect 23480 17824 23532 17876
rect 16304 17688 16356 17740
rect 17224 17688 17276 17740
rect 13360 17484 13412 17536
rect 13912 17595 13964 17604
rect 13912 17561 13921 17595
rect 13921 17561 13955 17595
rect 13955 17561 13964 17595
rect 13912 17552 13964 17561
rect 14188 17552 14240 17604
rect 14740 17552 14792 17604
rect 15200 17620 15252 17672
rect 16856 17620 16908 17672
rect 19432 17620 19484 17672
rect 19892 17620 19944 17672
rect 24308 17756 24360 17808
rect 26700 17824 26752 17876
rect 26516 17756 26568 17808
rect 20628 17688 20680 17740
rect 21916 17731 21968 17740
rect 21916 17697 21925 17731
rect 21925 17697 21959 17731
rect 21959 17697 21968 17731
rect 21916 17688 21968 17697
rect 22284 17688 22336 17740
rect 22652 17688 22704 17740
rect 26148 17731 26200 17740
rect 26148 17697 26157 17731
rect 26157 17697 26191 17731
rect 26191 17697 26200 17731
rect 26148 17688 26200 17697
rect 26240 17688 26292 17740
rect 20536 17552 20588 17604
rect 20628 17595 20680 17604
rect 20628 17561 20637 17595
rect 20637 17561 20671 17595
rect 20671 17561 20680 17595
rect 20628 17552 20680 17561
rect 15476 17484 15528 17536
rect 16120 17484 16172 17536
rect 16672 17484 16724 17536
rect 18052 17484 18104 17536
rect 19892 17484 19944 17536
rect 19984 17484 20036 17536
rect 21548 17620 21600 17672
rect 21824 17595 21876 17604
rect 21824 17561 21833 17595
rect 21833 17561 21867 17595
rect 21867 17561 21876 17595
rect 21824 17552 21876 17561
rect 22468 17620 22520 17672
rect 23204 17663 23256 17672
rect 23204 17629 23213 17663
rect 23213 17629 23247 17663
rect 23247 17629 23256 17663
rect 23204 17620 23256 17629
rect 22192 17484 22244 17536
rect 24400 17595 24452 17604
rect 24400 17561 24409 17595
rect 24409 17561 24443 17595
rect 24443 17561 24452 17595
rect 24400 17552 24452 17561
rect 25136 17620 25188 17672
rect 26148 17552 26200 17604
rect 27804 17824 27856 17876
rect 31024 17824 31076 17876
rect 31392 17824 31444 17876
rect 32220 17731 32272 17740
rect 32220 17697 32229 17731
rect 32229 17697 32263 17731
rect 32263 17697 32272 17731
rect 32220 17688 32272 17697
rect 27160 17620 27212 17672
rect 28448 17620 28500 17672
rect 28908 17663 28960 17672
rect 28908 17629 28917 17663
rect 28917 17629 28951 17663
rect 28951 17629 28960 17663
rect 28908 17620 28960 17629
rect 30380 17620 30432 17672
rect 30932 17663 30984 17672
rect 30932 17629 30941 17663
rect 30941 17629 30975 17663
rect 30975 17629 30984 17663
rect 30932 17620 30984 17629
rect 31024 17620 31076 17672
rect 25964 17484 26016 17536
rect 26700 17527 26752 17536
rect 26700 17493 26709 17527
rect 26709 17493 26743 17527
rect 26743 17493 26752 17527
rect 26700 17484 26752 17493
rect 30472 17552 30524 17604
rect 27068 17484 27120 17536
rect 28632 17484 28684 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 3240 17280 3292 17332
rect 3976 17212 4028 17264
rect 4160 17212 4212 17264
rect 4712 17212 4764 17264
rect 5540 17280 5592 17332
rect 6552 17280 6604 17332
rect 2688 17187 2740 17196
rect 2688 17153 2697 17187
rect 2697 17153 2731 17187
rect 2731 17153 2740 17187
rect 2688 17144 2740 17153
rect 3884 17144 3936 17196
rect 4252 17187 4304 17196
rect 4252 17153 4261 17187
rect 4261 17153 4295 17187
rect 4295 17153 4304 17187
rect 4252 17144 4304 17153
rect 4620 17187 4672 17196
rect 4620 17153 4629 17187
rect 4629 17153 4663 17187
rect 4663 17153 4672 17187
rect 4620 17144 4672 17153
rect 4804 17144 4856 17196
rect 6460 17212 6512 17264
rect 7196 17280 7248 17332
rect 7288 17280 7340 17332
rect 5724 17144 5776 17196
rect 6368 17187 6420 17196
rect 6368 17153 6377 17187
rect 6377 17153 6411 17187
rect 6411 17153 6420 17187
rect 6368 17144 6420 17153
rect 7380 17255 7432 17264
rect 7380 17221 7389 17255
rect 7389 17221 7423 17255
rect 7423 17221 7432 17255
rect 7380 17212 7432 17221
rect 6644 17187 6696 17196
rect 6644 17153 6653 17187
rect 6653 17153 6687 17187
rect 6687 17153 6696 17187
rect 6644 17144 6696 17153
rect 6920 17187 6972 17196
rect 6920 17153 6929 17187
rect 6929 17153 6963 17187
rect 6963 17153 6972 17187
rect 6920 17144 6972 17153
rect 7656 17280 7708 17332
rect 2688 17008 2740 17060
rect 3884 17008 3936 17060
rect 4988 17008 5040 17060
rect 3148 16940 3200 16992
rect 3700 16940 3752 16992
rect 7288 17008 7340 17060
rect 7656 17144 7708 17196
rect 8024 17280 8076 17332
rect 8208 17144 8260 17196
rect 9128 17144 9180 17196
rect 8668 17076 8720 17128
rect 9864 17212 9916 17264
rect 10324 17280 10376 17332
rect 11060 17280 11112 17332
rect 11796 17280 11848 17332
rect 12624 17280 12676 17332
rect 12716 17280 12768 17332
rect 15016 17280 15068 17332
rect 15292 17280 15344 17332
rect 15660 17280 15712 17332
rect 17776 17280 17828 17332
rect 17868 17280 17920 17332
rect 24400 17280 24452 17332
rect 10140 17255 10192 17264
rect 10140 17221 10149 17255
rect 10149 17221 10183 17255
rect 10183 17221 10192 17255
rect 10140 17212 10192 17221
rect 10416 17187 10468 17196
rect 10416 17153 10425 17187
rect 10425 17153 10459 17187
rect 10459 17153 10468 17187
rect 10416 17144 10468 17153
rect 10508 17144 10560 17196
rect 11060 17187 11112 17196
rect 11060 17153 11069 17187
rect 11069 17153 11103 17187
rect 11103 17153 11112 17187
rect 11060 17144 11112 17153
rect 11244 17144 11296 17196
rect 12164 17212 12216 17264
rect 12348 17212 12400 17264
rect 9864 17076 9916 17128
rect 10232 17076 10284 17128
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 11980 17187 12032 17196
rect 11980 17153 11989 17187
rect 11989 17153 12023 17187
rect 12023 17153 12032 17187
rect 11980 17144 12032 17153
rect 13820 17144 13872 17196
rect 14464 17144 14516 17196
rect 15936 17212 15988 17264
rect 16396 17212 16448 17264
rect 17960 17212 18012 17264
rect 18052 17212 18104 17264
rect 22008 17212 22060 17264
rect 22560 17255 22612 17264
rect 16580 17144 16632 17196
rect 17592 17144 17644 17196
rect 19616 17144 19668 17196
rect 22560 17221 22569 17255
rect 22569 17221 22603 17255
rect 22603 17221 22612 17255
rect 22560 17212 22612 17221
rect 23848 17212 23900 17264
rect 6552 16940 6604 16992
rect 7472 16940 7524 16992
rect 7656 16940 7708 16992
rect 12164 17076 12216 17128
rect 8208 16940 8260 16992
rect 8392 16940 8444 16992
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 10876 16983 10928 16992
rect 10876 16949 10885 16983
rect 10885 16949 10919 16983
rect 10919 16949 10928 16983
rect 10876 16940 10928 16949
rect 14832 17119 14884 17128
rect 14832 17085 14841 17119
rect 14841 17085 14875 17119
rect 14875 17085 14884 17119
rect 14832 17076 14884 17085
rect 14924 17076 14976 17128
rect 17868 17076 17920 17128
rect 18236 17076 18288 17128
rect 20260 17076 20312 17128
rect 20628 17076 20680 17128
rect 23204 17144 23256 17196
rect 24216 17187 24268 17196
rect 24216 17153 24225 17187
rect 24225 17153 24259 17187
rect 24259 17153 24268 17187
rect 24216 17144 24268 17153
rect 24308 17144 24360 17196
rect 25780 17187 25832 17196
rect 25780 17153 25789 17187
rect 25789 17153 25823 17187
rect 25823 17153 25832 17187
rect 25780 17144 25832 17153
rect 26148 17144 26200 17196
rect 26884 17144 26936 17196
rect 27252 17280 27304 17332
rect 30932 17280 30984 17332
rect 23480 17076 23532 17128
rect 27528 17144 27580 17196
rect 28448 17187 28500 17196
rect 28448 17153 28457 17187
rect 28457 17153 28491 17187
rect 28491 17153 28500 17187
rect 28448 17144 28500 17153
rect 28540 17144 28592 17196
rect 30656 17144 30708 17196
rect 31576 17144 31628 17196
rect 27712 17119 27764 17128
rect 27712 17085 27721 17119
rect 27721 17085 27755 17119
rect 27755 17085 27764 17119
rect 27712 17076 27764 17085
rect 27804 17076 27856 17128
rect 13912 17008 13964 17060
rect 16856 17008 16908 17060
rect 18144 17008 18196 17060
rect 22284 17008 22336 17060
rect 24124 17008 24176 17060
rect 32312 17144 32364 17196
rect 12164 16983 12216 16992
rect 12164 16949 12173 16983
rect 12173 16949 12207 16983
rect 12207 16949 12216 16983
rect 12164 16940 12216 16949
rect 12256 16983 12308 16992
rect 12256 16949 12265 16983
rect 12265 16949 12299 16983
rect 12299 16949 12308 16983
rect 12256 16940 12308 16949
rect 12716 16983 12768 16992
rect 12716 16949 12725 16983
rect 12725 16949 12759 16983
rect 12759 16949 12768 16983
rect 12716 16940 12768 16949
rect 12808 16940 12860 16992
rect 14004 16940 14056 16992
rect 14188 16940 14240 16992
rect 16028 16940 16080 16992
rect 16948 16940 17000 16992
rect 17776 16940 17828 16992
rect 23112 16983 23164 16992
rect 23112 16949 23121 16983
rect 23121 16949 23155 16983
rect 23155 16949 23164 16983
rect 23112 16940 23164 16949
rect 23848 16940 23900 16992
rect 24216 16940 24268 16992
rect 24676 16940 24728 16992
rect 28080 16983 28132 16992
rect 28080 16949 28089 16983
rect 28089 16949 28123 16983
rect 28123 16949 28132 16983
rect 28080 16940 28132 16949
rect 32404 17051 32456 17060
rect 32404 17017 32413 17051
rect 32413 17017 32447 17051
rect 32447 17017 32456 17051
rect 32404 17008 32456 17017
rect 30288 16940 30340 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 3240 16736 3292 16788
rect 3516 16736 3568 16788
rect 7472 16736 7524 16788
rect 8024 16779 8076 16788
rect 8024 16745 8033 16779
rect 8033 16745 8067 16779
rect 8067 16745 8076 16779
rect 8024 16736 8076 16745
rect 8484 16736 8536 16788
rect 10416 16736 10468 16788
rect 10692 16736 10744 16788
rect 11796 16736 11848 16788
rect 12164 16736 12216 16788
rect 13176 16736 13228 16788
rect 14004 16736 14056 16788
rect 15660 16736 15712 16788
rect 15936 16736 15988 16788
rect 16028 16779 16080 16788
rect 16028 16745 16037 16779
rect 16037 16745 16071 16779
rect 16071 16745 16080 16779
rect 16028 16736 16080 16745
rect 16488 16779 16540 16788
rect 16488 16745 16497 16779
rect 16497 16745 16531 16779
rect 16531 16745 16540 16779
rect 16488 16736 16540 16745
rect 16580 16736 16632 16788
rect 480 16668 532 16720
rect 3608 16600 3660 16652
rect 848 16532 900 16584
rect 2688 16575 2740 16584
rect 2688 16541 2697 16575
rect 2697 16541 2731 16575
rect 2731 16541 2740 16575
rect 2688 16532 2740 16541
rect 2964 16575 3016 16584
rect 2964 16541 2973 16575
rect 2973 16541 3007 16575
rect 3007 16541 3016 16575
rect 2964 16532 3016 16541
rect 3056 16575 3108 16584
rect 3056 16541 3065 16575
rect 3065 16541 3099 16575
rect 3099 16541 3108 16575
rect 3056 16532 3108 16541
rect 2412 16464 2464 16516
rect 2596 16464 2648 16516
rect 1584 16439 1636 16448
rect 1584 16405 1593 16439
rect 1593 16405 1627 16439
rect 1627 16405 1636 16439
rect 1584 16396 1636 16405
rect 2228 16396 2280 16448
rect 3240 16439 3292 16448
rect 3240 16405 3249 16439
rect 3249 16405 3283 16439
rect 3283 16405 3292 16439
rect 3240 16396 3292 16405
rect 4436 16668 4488 16720
rect 6000 16668 6052 16720
rect 9772 16668 9824 16720
rect 11980 16668 12032 16720
rect 4528 16600 4580 16652
rect 4988 16600 5040 16652
rect 4620 16575 4672 16584
rect 4620 16541 4629 16575
rect 4629 16541 4663 16575
rect 4663 16541 4672 16575
rect 4620 16532 4672 16541
rect 5172 16532 5224 16584
rect 5356 16575 5408 16584
rect 5356 16541 5365 16575
rect 5365 16541 5399 16575
rect 5399 16541 5408 16575
rect 5356 16532 5408 16541
rect 5540 16575 5592 16584
rect 5540 16541 5549 16575
rect 5549 16541 5583 16575
rect 5583 16541 5592 16575
rect 5540 16532 5592 16541
rect 5724 16575 5776 16584
rect 5724 16541 5733 16575
rect 5733 16541 5767 16575
rect 5767 16541 5776 16575
rect 5724 16532 5776 16541
rect 6092 16532 6144 16584
rect 7472 16532 7524 16584
rect 4528 16507 4580 16516
rect 4528 16473 4537 16507
rect 4537 16473 4571 16507
rect 4571 16473 4580 16507
rect 4528 16464 4580 16473
rect 5632 16507 5684 16516
rect 5632 16473 5641 16507
rect 5641 16473 5675 16507
rect 5675 16473 5684 16507
rect 5632 16464 5684 16473
rect 8300 16643 8352 16652
rect 8300 16609 8309 16643
rect 8309 16609 8343 16643
rect 8343 16609 8352 16643
rect 8300 16600 8352 16609
rect 8392 16575 8444 16584
rect 8392 16541 8401 16575
rect 8401 16541 8435 16575
rect 8435 16541 8444 16575
rect 8392 16532 8444 16541
rect 9864 16600 9916 16652
rect 14832 16668 14884 16720
rect 15016 16668 15068 16720
rect 15384 16668 15436 16720
rect 9956 16464 10008 16516
rect 11704 16464 11756 16516
rect 11980 16532 12032 16584
rect 12808 16575 12860 16584
rect 12808 16541 12817 16575
rect 12817 16541 12851 16575
rect 12851 16541 12860 16575
rect 12808 16532 12860 16541
rect 12992 16575 13044 16584
rect 12992 16541 13001 16575
rect 13001 16541 13035 16575
rect 13035 16541 13044 16575
rect 12992 16532 13044 16541
rect 13452 16575 13504 16584
rect 13452 16541 13461 16575
rect 13461 16541 13495 16575
rect 13495 16541 13504 16575
rect 13452 16532 13504 16541
rect 14372 16532 14424 16584
rect 4712 16396 4764 16448
rect 4804 16396 4856 16448
rect 6092 16396 6144 16448
rect 9496 16396 9548 16448
rect 9864 16396 9916 16448
rect 11152 16396 11204 16448
rect 12440 16396 12492 16448
rect 15108 16532 15160 16584
rect 15200 16575 15252 16584
rect 15200 16541 15209 16575
rect 15209 16541 15243 16575
rect 15243 16541 15252 16575
rect 15200 16532 15252 16541
rect 16948 16668 17000 16720
rect 17868 16736 17920 16788
rect 18788 16736 18840 16788
rect 16028 16600 16080 16652
rect 15016 16507 15068 16516
rect 15016 16473 15025 16507
rect 15025 16473 15059 16507
rect 15059 16473 15068 16507
rect 15016 16464 15068 16473
rect 15476 16507 15528 16516
rect 15476 16473 15485 16507
rect 15485 16473 15519 16507
rect 15519 16473 15528 16507
rect 15476 16464 15528 16473
rect 16304 16464 16356 16516
rect 16396 16507 16448 16516
rect 16396 16473 16405 16507
rect 16405 16473 16439 16507
rect 16439 16473 16448 16507
rect 16396 16464 16448 16473
rect 16580 16600 16632 16652
rect 16672 16575 16724 16584
rect 16672 16541 16681 16575
rect 16681 16541 16715 16575
rect 16715 16541 16724 16575
rect 16672 16532 16724 16541
rect 17316 16643 17368 16652
rect 17316 16609 17325 16643
rect 17325 16609 17359 16643
rect 17359 16609 17368 16643
rect 17316 16600 17368 16609
rect 18420 16600 18472 16652
rect 20260 16668 20312 16720
rect 22284 16736 22336 16788
rect 23848 16736 23900 16788
rect 25412 16779 25464 16788
rect 25412 16745 25421 16779
rect 25421 16745 25455 16779
rect 25455 16745 25464 16779
rect 25412 16736 25464 16745
rect 25780 16736 25832 16788
rect 27160 16736 27212 16788
rect 28080 16779 28132 16788
rect 28080 16745 28089 16779
rect 28089 16745 28123 16779
rect 28123 16745 28132 16779
rect 28080 16736 28132 16745
rect 28540 16736 28592 16788
rect 28724 16779 28776 16788
rect 28724 16745 28733 16779
rect 28733 16745 28767 16779
rect 28767 16745 28776 16779
rect 28724 16736 28776 16745
rect 21640 16668 21692 16720
rect 24492 16668 24544 16720
rect 22468 16600 22520 16652
rect 23388 16600 23440 16652
rect 23664 16600 23716 16652
rect 17500 16532 17552 16584
rect 17960 16575 18012 16584
rect 17960 16541 17969 16575
rect 17969 16541 18003 16575
rect 18003 16541 18012 16575
rect 17960 16532 18012 16541
rect 18052 16575 18104 16584
rect 18052 16541 18061 16575
rect 18061 16541 18095 16575
rect 18095 16541 18104 16575
rect 18052 16532 18104 16541
rect 12900 16396 12952 16448
rect 15660 16396 15712 16448
rect 15936 16439 15988 16448
rect 15936 16405 15945 16439
rect 15945 16405 15979 16439
rect 15979 16405 15988 16439
rect 15936 16396 15988 16405
rect 17132 16507 17184 16516
rect 17132 16473 17141 16507
rect 17141 16473 17175 16507
rect 17175 16473 17184 16507
rect 17132 16464 17184 16473
rect 17500 16396 17552 16448
rect 18420 16507 18472 16516
rect 18420 16473 18429 16507
rect 18429 16473 18463 16507
rect 18463 16473 18472 16507
rect 18420 16464 18472 16473
rect 18696 16575 18748 16584
rect 18696 16541 18705 16575
rect 18705 16541 18739 16575
rect 18739 16541 18748 16575
rect 18696 16532 18748 16541
rect 20996 16532 21048 16584
rect 23572 16532 23624 16584
rect 27620 16668 27672 16720
rect 29368 16736 29420 16788
rect 31576 16779 31628 16788
rect 31576 16745 31585 16779
rect 31585 16745 31619 16779
rect 31619 16745 31628 16779
rect 31576 16736 31628 16745
rect 26884 16600 26936 16652
rect 27160 16600 27212 16652
rect 27528 16600 27580 16652
rect 27804 16600 27856 16652
rect 28080 16600 28132 16652
rect 28908 16600 28960 16652
rect 32312 16643 32364 16652
rect 32312 16609 32321 16643
rect 32321 16609 32355 16643
rect 32355 16609 32364 16643
rect 32312 16600 32364 16609
rect 26700 16532 26752 16584
rect 18328 16439 18380 16448
rect 18328 16405 18337 16439
rect 18337 16405 18371 16439
rect 18371 16405 18380 16439
rect 18328 16396 18380 16405
rect 18880 16439 18932 16448
rect 18880 16405 18889 16439
rect 18889 16405 18923 16439
rect 18923 16405 18932 16439
rect 18880 16396 18932 16405
rect 19984 16396 20036 16448
rect 20536 16464 20588 16516
rect 22284 16464 22336 16516
rect 24860 16464 24912 16516
rect 25136 16464 25188 16516
rect 25412 16464 25464 16516
rect 28264 16532 28316 16584
rect 30288 16532 30340 16584
rect 29460 16464 29512 16516
rect 30932 16464 30984 16516
rect 28264 16396 28316 16448
rect 28632 16396 28684 16448
rect 29368 16439 29420 16448
rect 29368 16405 29377 16439
rect 29377 16405 29411 16439
rect 29411 16405 29420 16439
rect 29368 16396 29420 16405
rect 30380 16396 30432 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 2964 16192 3016 16244
rect 4436 16192 4488 16244
rect 4528 16192 4580 16244
rect 7012 16192 7064 16244
rect 9128 16192 9180 16244
rect 9864 16192 9916 16244
rect 10140 16192 10192 16244
rect 2688 16056 2740 16108
rect 2964 16099 3016 16108
rect 2964 16065 2973 16099
rect 2973 16065 3007 16099
rect 3007 16065 3016 16099
rect 2964 16056 3016 16065
rect 4344 16099 4396 16108
rect 4344 16065 4353 16099
rect 4353 16065 4387 16099
rect 4387 16065 4396 16099
rect 4344 16056 4396 16065
rect 5172 16056 5224 16108
rect 5816 16124 5868 16176
rect 6920 16124 6972 16176
rect 8484 16167 8536 16176
rect 8484 16133 8493 16167
rect 8493 16133 8527 16167
rect 8527 16133 8536 16167
rect 8484 16124 8536 16133
rect 9496 16124 9548 16176
rect 12532 16167 12584 16176
rect 12532 16133 12541 16167
rect 12541 16133 12575 16167
rect 12575 16133 12584 16167
rect 12532 16124 12584 16133
rect 12808 16192 12860 16244
rect 13084 16192 13136 16244
rect 16672 16192 16724 16244
rect 14280 16124 14332 16176
rect 6184 16056 6236 16108
rect 6736 16056 6788 16108
rect 3148 15988 3200 16040
rect 5908 15988 5960 16040
rect 7012 16099 7064 16108
rect 7012 16065 7021 16099
rect 7021 16065 7055 16099
rect 7055 16065 7064 16099
rect 7012 16056 7064 16065
rect 8668 16099 8720 16108
rect 8668 16065 8677 16099
rect 8677 16065 8711 16099
rect 8711 16065 8720 16099
rect 8668 16056 8720 16065
rect 8852 16099 8904 16108
rect 8852 16065 8861 16099
rect 8861 16065 8895 16099
rect 8895 16065 8904 16099
rect 8852 16056 8904 16065
rect 9036 16056 9088 16108
rect 10784 16099 10836 16108
rect 10784 16065 10793 16099
rect 10793 16065 10827 16099
rect 10827 16065 10836 16099
rect 10784 16056 10836 16065
rect 10968 16099 11020 16108
rect 10968 16065 10977 16099
rect 10977 16065 11011 16099
rect 11011 16065 11020 16099
rect 10968 16056 11020 16065
rect 12164 16056 12216 16108
rect 12808 16099 12860 16108
rect 12808 16065 12817 16099
rect 12817 16065 12851 16099
rect 12851 16065 12860 16099
rect 12808 16056 12860 16065
rect 15016 16056 15068 16108
rect 15384 16056 15436 16108
rect 16396 16124 16448 16176
rect 19340 16192 19392 16244
rect 16948 16124 17000 16176
rect 19156 16124 19208 16176
rect 19708 16124 19760 16176
rect 19984 16167 20036 16176
rect 19984 16133 19993 16167
rect 19993 16133 20027 16167
rect 20027 16133 20036 16167
rect 19984 16124 20036 16133
rect 22836 16167 22888 16176
rect 22836 16133 22845 16167
rect 22845 16133 22879 16167
rect 22879 16133 22888 16167
rect 22836 16124 22888 16133
rect 23480 16235 23532 16244
rect 23480 16201 23489 16235
rect 23489 16201 23523 16235
rect 23523 16201 23532 16235
rect 23480 16192 23532 16201
rect 27528 16192 27580 16244
rect 30196 16235 30248 16244
rect 30196 16201 30205 16235
rect 30205 16201 30239 16235
rect 30239 16201 30248 16235
rect 30196 16192 30248 16201
rect 30564 16192 30616 16244
rect 31760 16192 31812 16244
rect 30748 16124 30800 16176
rect 11152 15988 11204 16040
rect 11612 15988 11664 16040
rect 12624 15988 12676 16040
rect 13176 15988 13228 16040
rect 17684 16056 17736 16108
rect 18328 16056 18380 16108
rect 20536 16099 20588 16108
rect 20536 16065 20545 16099
rect 20545 16065 20579 16099
rect 20579 16065 20588 16099
rect 20536 16056 20588 16065
rect 20720 16099 20772 16108
rect 20720 16065 20729 16099
rect 20729 16065 20763 16099
rect 20763 16065 20772 16099
rect 20720 16056 20772 16065
rect 20904 16056 20956 16108
rect 1124 15920 1176 15972
rect 3608 15852 3660 15904
rect 4712 15963 4764 15972
rect 4712 15929 4721 15963
rect 4721 15929 4755 15963
rect 4755 15929 4764 15963
rect 4712 15920 4764 15929
rect 6000 15920 6052 15972
rect 6276 15920 6328 15972
rect 8300 15920 8352 15972
rect 5816 15852 5868 15904
rect 6184 15852 6236 15904
rect 12440 15920 12492 15972
rect 12900 15920 12952 15972
rect 14004 15920 14056 15972
rect 16304 15988 16356 16040
rect 18788 15988 18840 16040
rect 19708 15988 19760 16040
rect 22928 16031 22980 16040
rect 22928 15997 22937 16031
rect 22937 15997 22971 16031
rect 22971 15997 22980 16031
rect 22928 15988 22980 15997
rect 8852 15852 8904 15904
rect 10324 15852 10376 15904
rect 10692 15895 10744 15904
rect 10692 15861 10701 15895
rect 10701 15861 10735 15895
rect 10735 15861 10744 15895
rect 10692 15852 10744 15861
rect 11152 15895 11204 15904
rect 11152 15861 11161 15895
rect 11161 15861 11195 15895
rect 11195 15861 11204 15895
rect 11152 15852 11204 15861
rect 11796 15852 11848 15904
rect 13912 15852 13964 15904
rect 15752 15963 15804 15972
rect 15752 15929 15761 15963
rect 15761 15929 15795 15963
rect 15795 15929 15804 15963
rect 15752 15920 15804 15929
rect 15936 15920 15988 15972
rect 24308 16056 24360 16108
rect 23388 15988 23440 16040
rect 24860 16056 24912 16108
rect 25780 16056 25832 16108
rect 26424 16099 26476 16108
rect 26424 16065 26433 16099
rect 26433 16065 26467 16099
rect 26467 16065 26476 16099
rect 26424 16056 26476 16065
rect 29644 16056 29696 16108
rect 30012 16099 30064 16108
rect 30012 16065 30021 16099
rect 30021 16065 30055 16099
rect 30055 16065 30064 16099
rect 30012 16056 30064 16065
rect 30196 16056 30248 16108
rect 30564 16099 30616 16108
rect 30564 16065 30573 16099
rect 30573 16065 30607 16099
rect 30607 16065 30616 16099
rect 30564 16056 30616 16065
rect 26332 15988 26384 16040
rect 29276 15988 29328 16040
rect 29828 16031 29880 16040
rect 29828 15997 29837 16031
rect 29837 15997 29871 16031
rect 29871 15997 29880 16031
rect 29828 15988 29880 15997
rect 26792 15963 26844 15972
rect 26792 15929 26801 15963
rect 26801 15929 26835 15963
rect 26835 15929 26844 15963
rect 26792 15920 26844 15929
rect 30564 15920 30616 15972
rect 30840 16099 30892 16108
rect 30840 16065 30849 16099
rect 30849 16065 30883 16099
rect 30883 16065 30892 16099
rect 30840 16056 30892 16065
rect 32220 16099 32272 16108
rect 32220 16065 32229 16099
rect 32229 16065 32263 16099
rect 32263 16065 32272 16099
rect 32220 16056 32272 16065
rect 17040 15852 17092 15904
rect 18144 15852 18196 15904
rect 18696 15852 18748 15904
rect 19892 15852 19944 15904
rect 20444 15852 20496 15904
rect 21180 15852 21232 15904
rect 21272 15852 21324 15904
rect 21916 15852 21968 15904
rect 22468 15852 22520 15904
rect 23296 15895 23348 15904
rect 23296 15861 23305 15895
rect 23305 15861 23339 15895
rect 23339 15861 23348 15895
rect 23296 15852 23348 15861
rect 23480 15852 23532 15904
rect 23848 15852 23900 15904
rect 25504 15895 25556 15904
rect 25504 15861 25513 15895
rect 25513 15861 25547 15895
rect 25547 15861 25556 15895
rect 25504 15852 25556 15861
rect 26700 15852 26752 15904
rect 29460 15852 29512 15904
rect 30472 15852 30524 15904
rect 31208 15895 31260 15904
rect 31208 15861 31217 15895
rect 31217 15861 31251 15895
rect 31251 15861 31260 15895
rect 31208 15852 31260 15861
rect 32404 15895 32456 15904
rect 32404 15861 32413 15895
rect 32413 15861 32447 15895
rect 32447 15861 32456 15895
rect 32404 15852 32456 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 3884 15648 3936 15700
rect 5540 15648 5592 15700
rect 6000 15648 6052 15700
rect 6276 15648 6328 15700
rect 6552 15580 6604 15632
rect 6736 15691 6788 15700
rect 6736 15657 6745 15691
rect 6745 15657 6779 15691
rect 6779 15657 6788 15691
rect 6736 15648 6788 15657
rect 7840 15648 7892 15700
rect 12808 15648 12860 15700
rect 14924 15648 14976 15700
rect 15108 15648 15160 15700
rect 15200 15691 15252 15700
rect 15200 15657 15209 15691
rect 15209 15657 15243 15691
rect 15243 15657 15252 15691
rect 15200 15648 15252 15657
rect 15292 15648 15344 15700
rect 16764 15691 16816 15700
rect 16764 15657 16773 15691
rect 16773 15657 16807 15691
rect 16807 15657 16816 15691
rect 16764 15648 16816 15657
rect 18144 15648 18196 15700
rect 18512 15648 18564 15700
rect 20444 15648 20496 15700
rect 21824 15648 21876 15700
rect 22468 15691 22520 15700
rect 22468 15657 22477 15691
rect 22477 15657 22511 15691
rect 22511 15657 22520 15691
rect 22468 15648 22520 15657
rect 23020 15691 23072 15700
rect 23020 15657 23029 15691
rect 23029 15657 23063 15691
rect 23063 15657 23072 15691
rect 23020 15648 23072 15657
rect 27528 15648 27580 15700
rect 29460 15648 29512 15700
rect 30196 15691 30248 15700
rect 30196 15657 30205 15691
rect 30205 15657 30239 15691
rect 30239 15657 30248 15691
rect 30196 15648 30248 15657
rect 30564 15691 30616 15700
rect 30564 15657 30573 15691
rect 30573 15657 30607 15691
rect 30607 15657 30616 15691
rect 30564 15648 30616 15657
rect 32220 15648 32272 15700
rect 9128 15580 9180 15632
rect 9312 15580 9364 15632
rect 10232 15623 10284 15632
rect 10232 15589 10241 15623
rect 10241 15589 10275 15623
rect 10275 15589 10284 15623
rect 10232 15580 10284 15589
rect 10416 15580 10468 15632
rect 3792 15512 3844 15564
rect 6184 15512 6236 15564
rect 3884 15487 3936 15496
rect 3884 15453 3893 15487
rect 3893 15453 3927 15487
rect 3927 15453 3936 15487
rect 3884 15444 3936 15453
rect 4528 15444 4580 15496
rect 5264 15487 5316 15496
rect 5264 15453 5273 15487
rect 5273 15453 5307 15487
rect 5307 15453 5316 15487
rect 5264 15444 5316 15453
rect 5632 15444 5684 15496
rect 6552 15487 6604 15496
rect 6552 15453 6561 15487
rect 6561 15453 6595 15487
rect 6595 15453 6604 15487
rect 6552 15444 6604 15453
rect 7656 15512 7708 15564
rect 10508 15512 10560 15564
rect 6736 15444 6788 15496
rect 8300 15444 8352 15496
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 10048 15487 10100 15496
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 10600 15444 10652 15496
rect 10784 15487 10836 15496
rect 10784 15453 10793 15487
rect 10793 15453 10827 15487
rect 10827 15453 10836 15487
rect 10784 15444 10836 15453
rect 2504 15376 2556 15428
rect 7380 15376 7432 15428
rect 7472 15376 7524 15428
rect 15384 15580 15436 15632
rect 12348 15512 12400 15564
rect 13912 15512 13964 15564
rect 14004 15512 14056 15564
rect 16212 15580 16264 15632
rect 18880 15580 18932 15632
rect 21640 15580 21692 15632
rect 15660 15512 15712 15564
rect 17960 15512 18012 15564
rect 22284 15580 22336 15632
rect 22192 15555 22244 15564
rect 22192 15521 22201 15555
rect 22201 15521 22235 15555
rect 22235 15521 22244 15555
rect 22192 15512 22244 15521
rect 22928 15512 22980 15564
rect 23572 15512 23624 15564
rect 27068 15555 27120 15564
rect 27068 15521 27077 15555
rect 27077 15521 27111 15555
rect 27111 15521 27120 15555
rect 27068 15512 27120 15521
rect 12164 15444 12216 15496
rect 12440 15444 12492 15496
rect 12808 15376 12860 15428
rect 13084 15376 13136 15428
rect 13544 15419 13596 15428
rect 13544 15385 13553 15419
rect 13553 15385 13587 15419
rect 13587 15385 13596 15419
rect 13544 15376 13596 15385
rect 15016 15487 15068 15496
rect 15016 15453 15025 15487
rect 15025 15453 15059 15487
rect 15059 15453 15068 15487
rect 15016 15444 15068 15453
rect 15384 15444 15436 15496
rect 16120 15444 16172 15496
rect 18788 15444 18840 15496
rect 20444 15444 20496 15496
rect 22008 15444 22060 15496
rect 4068 15308 4120 15360
rect 8392 15308 8444 15360
rect 8484 15308 8536 15360
rect 9312 15308 9364 15360
rect 9772 15308 9824 15360
rect 10324 15308 10376 15360
rect 10784 15308 10836 15360
rect 10876 15308 10928 15360
rect 14188 15308 14240 15360
rect 17224 15376 17276 15428
rect 15844 15308 15896 15360
rect 19340 15376 19392 15428
rect 19616 15376 19668 15428
rect 19708 15308 19760 15360
rect 21824 15376 21876 15428
rect 23204 15444 23256 15496
rect 24952 15444 25004 15496
rect 25504 15487 25556 15496
rect 25504 15453 25513 15487
rect 25513 15453 25547 15487
rect 25547 15453 25556 15487
rect 25504 15444 25556 15453
rect 22468 15376 22520 15428
rect 22652 15419 22704 15428
rect 22652 15385 22661 15419
rect 22661 15385 22695 15419
rect 22695 15385 22704 15419
rect 22652 15376 22704 15385
rect 22928 15376 22980 15428
rect 20260 15308 20312 15360
rect 20536 15308 20588 15360
rect 20812 15308 20864 15360
rect 27344 15444 27396 15496
rect 27528 15444 27580 15496
rect 28816 15444 28868 15496
rect 29828 15555 29880 15564
rect 29828 15521 29837 15555
rect 29837 15521 29871 15555
rect 29871 15521 29880 15555
rect 29828 15512 29880 15521
rect 30656 15512 30708 15564
rect 26976 15419 27028 15428
rect 26976 15385 26985 15419
rect 26985 15385 27019 15419
rect 27019 15385 27028 15419
rect 26976 15376 27028 15385
rect 27436 15376 27488 15428
rect 28540 15376 28592 15428
rect 29276 15376 29328 15428
rect 29460 15376 29512 15428
rect 29736 15376 29788 15428
rect 31208 15444 31260 15496
rect 30012 15376 30064 15428
rect 23480 15351 23532 15360
rect 23480 15317 23489 15351
rect 23489 15317 23523 15351
rect 23523 15317 23532 15351
rect 23480 15308 23532 15317
rect 25872 15308 25924 15360
rect 28172 15308 28224 15360
rect 28448 15308 28500 15360
rect 30564 15308 30616 15360
rect 30932 15308 30984 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 3056 15104 3108 15156
rect 3884 15147 3936 15156
rect 3884 15113 3893 15147
rect 3893 15113 3927 15147
rect 3927 15113 3936 15147
rect 3884 15104 3936 15113
rect 6736 15104 6788 15156
rect 7012 15104 7064 15156
rect 2228 15011 2280 15020
rect 2228 14977 2237 15011
rect 2237 14977 2271 15011
rect 2271 14977 2280 15011
rect 2228 14968 2280 14977
rect 2412 15011 2464 15020
rect 2412 14977 2421 15011
rect 2421 14977 2455 15011
rect 2455 14977 2464 15011
rect 2412 14968 2464 14977
rect 2964 15011 3016 15020
rect 2964 14977 2973 15011
rect 2973 14977 3007 15011
rect 3007 14977 3016 15011
rect 2964 14968 3016 14977
rect 3148 15011 3200 15020
rect 3148 14977 3157 15011
rect 3157 14977 3191 15011
rect 3191 14977 3200 15011
rect 3148 14968 3200 14977
rect 3792 14968 3844 15020
rect 4712 15036 4764 15088
rect 4620 15011 4672 15020
rect 4620 14977 4629 15011
rect 4629 14977 4663 15011
rect 4663 14977 4672 15011
rect 4620 14968 4672 14977
rect 4804 14968 4856 15020
rect 5448 15036 5500 15088
rect 7380 15036 7432 15088
rect 8852 15104 8904 15156
rect 10968 15104 11020 15156
rect 12164 15104 12216 15156
rect 8760 15036 8812 15088
rect 3976 14900 4028 14952
rect 4712 14900 4764 14952
rect 4988 14900 5040 14952
rect 7472 14968 7524 15020
rect 8116 14968 8168 15020
rect 8300 15011 8352 15020
rect 8300 14977 8309 15011
rect 8309 14977 8343 15011
rect 8343 14977 8352 15011
rect 8300 14968 8352 14977
rect 8392 15011 8444 15020
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 8484 14968 8536 15020
rect 8852 14968 8904 15020
rect 5540 14900 5592 14952
rect 5724 14900 5776 14952
rect 6368 14943 6420 14952
rect 6368 14909 6377 14943
rect 6377 14909 6411 14943
rect 6411 14909 6420 14943
rect 6368 14900 6420 14909
rect 7012 14900 7064 14952
rect 8024 14900 8076 14952
rect 9312 14968 9364 15020
rect 10048 15079 10100 15088
rect 10048 15045 10057 15079
rect 10057 15045 10091 15079
rect 10091 15045 10100 15079
rect 10048 15036 10100 15045
rect 11244 15036 11296 15088
rect 13544 15079 13596 15088
rect 13544 15045 13553 15079
rect 13553 15045 13587 15079
rect 13587 15045 13596 15079
rect 13544 15036 13596 15045
rect 14096 15036 14148 15088
rect 14372 15036 14424 15088
rect 9588 14968 9640 15020
rect 10324 15011 10376 15020
rect 10324 14977 10333 15011
rect 10333 14977 10367 15011
rect 10367 14977 10376 15011
rect 10324 14968 10376 14977
rect 10784 15011 10836 15020
rect 10784 14977 10793 15011
rect 10793 14977 10827 15011
rect 10827 14977 10836 15011
rect 10784 14968 10836 14977
rect 10968 14968 11020 15020
rect 11152 14968 11204 15020
rect 11796 14968 11848 15020
rect 11888 14968 11940 15020
rect 13728 15011 13780 15020
rect 8668 14832 8720 14884
rect 3792 14764 3844 14816
rect 3976 14764 4028 14816
rect 4528 14764 4580 14816
rect 4896 14764 4948 14816
rect 5080 14807 5132 14816
rect 5080 14773 5089 14807
rect 5089 14773 5123 14807
rect 5123 14773 5132 14807
rect 5080 14764 5132 14773
rect 7656 14764 7708 14816
rect 7748 14807 7800 14816
rect 7748 14773 7757 14807
rect 7757 14773 7791 14807
rect 7791 14773 7800 14807
rect 7748 14764 7800 14773
rect 8024 14764 8076 14816
rect 8852 14807 8904 14816
rect 8852 14773 8861 14807
rect 8861 14773 8895 14807
rect 8895 14773 8904 14807
rect 8852 14764 8904 14773
rect 11060 14832 11112 14884
rect 12256 14900 12308 14952
rect 13728 14977 13737 15011
rect 13737 14977 13771 15011
rect 13771 14977 13780 15011
rect 13728 14968 13780 14977
rect 14280 15011 14332 15020
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14280 14968 14332 14977
rect 15844 15104 15896 15156
rect 16396 15104 16448 15156
rect 16764 15104 16816 15156
rect 17776 15104 17828 15156
rect 20628 15104 20680 15156
rect 22468 15104 22520 15156
rect 12440 14900 12492 14952
rect 13268 14900 13320 14952
rect 9588 14764 9640 14816
rect 9864 14807 9916 14816
rect 9864 14773 9873 14807
rect 9873 14773 9907 14807
rect 9907 14773 9916 14807
rect 9864 14764 9916 14773
rect 10048 14807 10100 14816
rect 10048 14773 10057 14807
rect 10057 14773 10091 14807
rect 10091 14773 10100 14807
rect 10048 14764 10100 14773
rect 10692 14764 10744 14816
rect 10876 14807 10928 14816
rect 10876 14773 10885 14807
rect 10885 14773 10919 14807
rect 10919 14773 10928 14807
rect 10876 14764 10928 14773
rect 13176 14832 13228 14884
rect 13452 14832 13504 14884
rect 13636 14832 13688 14884
rect 17132 14900 17184 14952
rect 12072 14807 12124 14816
rect 12072 14773 12081 14807
rect 12081 14773 12115 14807
rect 12115 14773 12124 14807
rect 12072 14764 12124 14773
rect 13268 14764 13320 14816
rect 13544 14764 13596 14816
rect 14924 14832 14976 14884
rect 17684 15011 17736 15020
rect 17684 14977 17693 15011
rect 17693 14977 17727 15011
rect 17727 14977 17736 15011
rect 17684 14968 17736 14977
rect 17776 15011 17828 15020
rect 17776 14977 17785 15011
rect 17785 14977 17819 15011
rect 17819 14977 17828 15011
rect 17776 14968 17828 14977
rect 18236 14968 18288 15020
rect 18420 15011 18472 15020
rect 18420 14977 18429 15011
rect 18429 14977 18463 15011
rect 18463 14977 18472 15011
rect 18420 14968 18472 14977
rect 18880 15011 18932 15020
rect 18880 14977 18889 15011
rect 18889 14977 18923 15011
rect 18923 14977 18932 15011
rect 18880 14968 18932 14977
rect 19616 14968 19668 15020
rect 20444 15036 20496 15088
rect 21640 15036 21692 15088
rect 23388 15079 23440 15088
rect 23388 15045 23397 15079
rect 23397 15045 23431 15079
rect 23431 15045 23440 15079
rect 23388 15036 23440 15045
rect 23756 15104 23808 15156
rect 26056 15147 26108 15156
rect 26056 15113 26065 15147
rect 26065 15113 26099 15147
rect 26099 15113 26108 15147
rect 26056 15104 26108 15113
rect 29552 15104 29604 15156
rect 30196 15104 30248 15156
rect 32404 15147 32456 15156
rect 32404 15113 32413 15147
rect 32413 15113 32447 15147
rect 32447 15113 32456 15147
rect 32404 15104 32456 15113
rect 30380 15036 30432 15088
rect 31208 15036 31260 15088
rect 22100 14968 22152 15020
rect 23572 14968 23624 15020
rect 23664 15011 23716 15020
rect 23664 14977 23673 15011
rect 23673 14977 23707 15011
rect 23707 14977 23716 15011
rect 23664 14968 23716 14977
rect 23756 14968 23808 15020
rect 24676 14968 24728 15020
rect 28080 15011 28132 15020
rect 28080 14977 28089 15011
rect 28089 14977 28123 15011
rect 28123 14977 28132 15011
rect 28080 14968 28132 14977
rect 30840 14968 30892 15020
rect 31024 15011 31076 15020
rect 31024 14977 31033 15011
rect 31033 14977 31067 15011
rect 31067 14977 31076 15011
rect 31024 14968 31076 14977
rect 32220 15011 32272 15020
rect 32220 14977 32229 15011
rect 32229 14977 32263 15011
rect 32263 14977 32272 15011
rect 32220 14968 32272 14977
rect 14648 14764 14700 14816
rect 15292 14764 15344 14816
rect 16212 14764 16264 14816
rect 16672 14764 16724 14816
rect 16948 14764 17000 14816
rect 17040 14807 17092 14816
rect 17040 14773 17049 14807
rect 17049 14773 17083 14807
rect 17083 14773 17092 14807
rect 17040 14764 17092 14773
rect 17132 14764 17184 14816
rect 17684 14832 17736 14884
rect 17776 14832 17828 14884
rect 18788 14875 18840 14884
rect 18788 14841 18797 14875
rect 18797 14841 18831 14875
rect 18831 14841 18840 14875
rect 18788 14832 18840 14841
rect 18880 14832 18932 14884
rect 22928 14900 22980 14952
rect 23296 14900 23348 14952
rect 24952 14900 25004 14952
rect 26056 14900 26108 14952
rect 30380 14900 30432 14952
rect 19156 14875 19208 14884
rect 19156 14841 19165 14875
rect 19165 14841 19199 14875
rect 19199 14841 19208 14875
rect 19156 14832 19208 14841
rect 18420 14807 18472 14816
rect 18420 14773 18429 14807
rect 18429 14773 18463 14807
rect 18463 14773 18472 14807
rect 18420 14764 18472 14773
rect 18512 14764 18564 14816
rect 24676 14832 24728 14884
rect 19616 14764 19668 14816
rect 20076 14764 20128 14816
rect 21272 14764 21324 14816
rect 23204 14764 23256 14816
rect 23848 14764 23900 14816
rect 24492 14764 24544 14816
rect 24860 14764 24912 14816
rect 25596 14764 25648 14816
rect 29000 14764 29052 14816
rect 29736 14764 29788 14816
rect 30472 14764 30524 14816
rect 30656 14764 30708 14816
rect 30840 14807 30892 14816
rect 30840 14773 30849 14807
rect 30849 14773 30883 14807
rect 30883 14773 30892 14807
rect 30840 14764 30892 14773
rect 31392 14764 31444 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 1492 14560 1544 14612
rect 3884 14560 3936 14612
rect 4068 14603 4120 14612
rect 4068 14569 4077 14603
rect 4077 14569 4111 14603
rect 4111 14569 4120 14603
rect 4068 14560 4120 14569
rect 4712 14560 4764 14612
rect 5540 14560 5592 14612
rect 5724 14603 5776 14612
rect 5724 14569 5733 14603
rect 5733 14569 5767 14603
rect 5767 14569 5776 14603
rect 5724 14560 5776 14569
rect 3240 14424 3292 14476
rect 848 14356 900 14408
rect 3976 14356 4028 14408
rect 6644 14560 6696 14612
rect 7380 14603 7432 14612
rect 7380 14569 7389 14603
rect 7389 14569 7423 14603
rect 7423 14569 7432 14603
rect 7380 14560 7432 14569
rect 8300 14560 8352 14612
rect 9128 14560 9180 14612
rect 11244 14603 11296 14612
rect 11244 14569 11253 14603
rect 11253 14569 11287 14603
rect 11287 14569 11296 14603
rect 11244 14560 11296 14569
rect 11612 14603 11664 14612
rect 11612 14569 11621 14603
rect 11621 14569 11655 14603
rect 11655 14569 11664 14603
rect 11612 14560 11664 14569
rect 11704 14560 11756 14612
rect 4620 14424 4672 14476
rect 4804 14356 4856 14408
rect 5908 14424 5960 14476
rect 6828 14492 6880 14544
rect 8944 14492 8996 14544
rect 9496 14492 9548 14544
rect 9680 14492 9732 14544
rect 7288 14424 7340 14476
rect 7748 14424 7800 14476
rect 7932 14467 7984 14476
rect 7932 14433 7941 14467
rect 7941 14433 7975 14467
rect 7975 14433 7984 14467
rect 7932 14424 7984 14433
rect 8392 14424 8444 14476
rect 9956 14424 10008 14476
rect 10600 14492 10652 14544
rect 11152 14492 11204 14544
rect 4988 14288 5040 14340
rect 5080 14288 5132 14340
rect 5816 14399 5868 14408
rect 5816 14365 5825 14399
rect 5825 14365 5859 14399
rect 5859 14365 5868 14399
rect 5816 14356 5868 14365
rect 6460 14356 6512 14408
rect 6552 14356 6604 14408
rect 6736 14399 6788 14408
rect 6736 14365 6745 14399
rect 6745 14365 6779 14399
rect 6779 14365 6788 14399
rect 6736 14356 6788 14365
rect 7012 14356 7064 14408
rect 7656 14399 7708 14408
rect 7656 14365 7665 14399
rect 7665 14365 7699 14399
rect 7699 14365 7708 14399
rect 7656 14356 7708 14365
rect 8300 14356 8352 14408
rect 9312 14356 9364 14408
rect 9772 14356 9824 14408
rect 10876 14424 10928 14476
rect 11336 14492 11388 14544
rect 11704 14467 11756 14476
rect 11704 14433 11713 14467
rect 11713 14433 11747 14467
rect 11747 14433 11756 14467
rect 11704 14424 11756 14433
rect 12440 14560 12492 14612
rect 13084 14560 13136 14612
rect 15016 14560 15068 14612
rect 11980 14492 12032 14544
rect 12624 14492 12676 14544
rect 14648 14492 14700 14544
rect 16120 14492 16172 14544
rect 16488 14603 16540 14612
rect 16488 14569 16497 14603
rect 16497 14569 16531 14603
rect 16531 14569 16540 14603
rect 16488 14560 16540 14569
rect 16672 14560 16724 14612
rect 16764 14603 16816 14612
rect 16764 14569 16773 14603
rect 16773 14569 16807 14603
rect 16807 14569 16816 14603
rect 16764 14560 16816 14569
rect 17592 14560 17644 14612
rect 18512 14560 18564 14612
rect 18880 14560 18932 14612
rect 19524 14560 19576 14612
rect 6000 14288 6052 14340
rect 6184 14288 6236 14340
rect 7288 14288 7340 14340
rect 8852 14288 8904 14340
rect 10232 14399 10284 14408
rect 10232 14365 10241 14399
rect 10241 14365 10275 14399
rect 10275 14365 10284 14399
rect 10232 14356 10284 14365
rect 9956 14331 10008 14340
rect 9956 14297 9965 14331
rect 9965 14297 9999 14331
rect 9999 14297 10008 14331
rect 9956 14288 10008 14297
rect 5540 14220 5592 14272
rect 5816 14220 5868 14272
rect 6828 14220 6880 14272
rect 7472 14220 7524 14272
rect 11796 14356 11848 14408
rect 11888 14399 11940 14408
rect 11888 14365 11897 14399
rect 11897 14365 11931 14399
rect 11931 14365 11940 14399
rect 11888 14356 11940 14365
rect 10600 14288 10652 14340
rect 10968 14288 11020 14340
rect 10416 14263 10468 14272
rect 10416 14229 10425 14263
rect 10425 14229 10459 14263
rect 10459 14229 10468 14263
rect 10416 14220 10468 14229
rect 11520 14288 11572 14340
rect 11704 14288 11756 14340
rect 12256 14424 12308 14476
rect 12072 14356 12124 14408
rect 12256 14288 12308 14340
rect 13084 14356 13136 14408
rect 13268 14356 13320 14408
rect 12624 14288 12676 14340
rect 14096 14356 14148 14408
rect 11336 14220 11388 14272
rect 14648 14288 14700 14340
rect 15384 14331 15436 14340
rect 15384 14297 15393 14331
rect 15393 14297 15427 14331
rect 15427 14297 15436 14331
rect 15384 14288 15436 14297
rect 15568 14331 15620 14340
rect 15568 14297 15577 14331
rect 15577 14297 15611 14331
rect 15611 14297 15620 14331
rect 15568 14288 15620 14297
rect 16212 14356 16264 14408
rect 19984 14535 20036 14544
rect 19984 14501 19993 14535
rect 19993 14501 20027 14535
rect 20027 14501 20036 14535
rect 19984 14492 20036 14501
rect 20812 14560 20864 14612
rect 17040 14424 17092 14476
rect 16396 14399 16448 14408
rect 16396 14365 16405 14399
rect 16405 14365 16439 14399
rect 16439 14365 16448 14399
rect 16396 14356 16448 14365
rect 16488 14399 16540 14408
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 16948 14356 17000 14408
rect 17776 14424 17828 14476
rect 18788 14356 18840 14408
rect 15200 14220 15252 14272
rect 16028 14220 16080 14272
rect 17684 14263 17736 14272
rect 17684 14229 17693 14263
rect 17693 14229 17727 14263
rect 17727 14229 17736 14263
rect 17684 14220 17736 14229
rect 18236 14288 18288 14340
rect 19340 14288 19392 14340
rect 19708 14356 19760 14408
rect 19800 14399 19852 14408
rect 19800 14365 19809 14399
rect 19809 14365 19843 14399
rect 19843 14365 19852 14399
rect 19800 14356 19852 14365
rect 20076 14399 20128 14408
rect 20076 14365 20085 14399
rect 20085 14365 20119 14399
rect 20119 14365 20128 14399
rect 20076 14356 20128 14365
rect 20720 14492 20772 14544
rect 24308 14560 24360 14612
rect 24768 14560 24820 14612
rect 27068 14560 27120 14612
rect 27528 14560 27580 14612
rect 30288 14603 30340 14612
rect 30288 14569 30297 14603
rect 30297 14569 30331 14603
rect 30331 14569 30340 14603
rect 30288 14560 30340 14569
rect 30564 14560 30616 14612
rect 27804 14492 27856 14544
rect 30012 14492 30064 14544
rect 30748 14560 30800 14612
rect 30932 14560 30984 14612
rect 20352 14356 20404 14408
rect 23296 14356 23348 14408
rect 24492 14424 24544 14476
rect 25228 14424 25280 14476
rect 19248 14220 19300 14272
rect 21456 14331 21508 14340
rect 21456 14297 21465 14331
rect 21465 14297 21499 14331
rect 21499 14297 21508 14331
rect 21456 14288 21508 14297
rect 21640 14331 21692 14340
rect 21640 14297 21649 14331
rect 21649 14297 21683 14331
rect 21683 14297 21692 14331
rect 21640 14288 21692 14297
rect 20536 14220 20588 14272
rect 22560 14288 22612 14340
rect 22928 14288 22980 14340
rect 23204 14288 23256 14340
rect 24768 14399 24820 14408
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 24492 14263 24544 14272
rect 24492 14229 24501 14263
rect 24501 14229 24535 14263
rect 24535 14229 24544 14263
rect 24492 14220 24544 14229
rect 25228 14331 25280 14340
rect 25228 14297 25237 14331
rect 25237 14297 25271 14331
rect 25271 14297 25280 14331
rect 25228 14288 25280 14297
rect 25596 14288 25648 14340
rect 25964 14288 26016 14340
rect 26240 14288 26292 14340
rect 26976 14356 27028 14408
rect 27068 14356 27120 14408
rect 27436 14356 27488 14408
rect 27620 14424 27672 14476
rect 27988 14356 28040 14408
rect 29000 14467 29052 14476
rect 29000 14433 29009 14467
rect 29009 14433 29043 14467
rect 29043 14433 29052 14467
rect 29000 14424 29052 14433
rect 29828 14424 29880 14476
rect 29184 14356 29236 14408
rect 31760 14424 31812 14476
rect 27620 14288 27672 14340
rect 27712 14288 27764 14340
rect 28816 14331 28868 14340
rect 28816 14297 28825 14331
rect 28825 14297 28859 14331
rect 28859 14297 28868 14331
rect 28816 14288 28868 14297
rect 26608 14220 26660 14272
rect 27436 14220 27488 14272
rect 29828 14220 29880 14272
rect 30932 14399 30984 14408
rect 30932 14365 30941 14399
rect 30941 14365 30975 14399
rect 30975 14365 30984 14399
rect 30932 14356 30984 14365
rect 31392 14399 31444 14408
rect 31392 14365 31401 14399
rect 31401 14365 31435 14399
rect 31435 14365 31444 14399
rect 31392 14356 31444 14365
rect 31668 14399 31720 14408
rect 31668 14365 31677 14399
rect 31677 14365 31711 14399
rect 31711 14365 31720 14399
rect 31668 14356 31720 14365
rect 30288 14220 30340 14272
rect 31024 14220 31076 14272
rect 31852 14220 31904 14272
rect 32128 14220 32180 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 4620 14016 4672 14068
rect 4712 14016 4764 14068
rect 5724 14016 5776 14068
rect 6000 14059 6052 14068
rect 6000 14025 6009 14059
rect 6009 14025 6043 14059
rect 6043 14025 6052 14059
rect 6000 14016 6052 14025
rect 7288 14059 7340 14068
rect 7288 14025 7297 14059
rect 7297 14025 7331 14059
rect 7331 14025 7340 14059
rect 7288 14016 7340 14025
rect 3148 13880 3200 13932
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 3700 13880 3752 13932
rect 3884 13880 3936 13932
rect 5540 13991 5592 14000
rect 5540 13957 5549 13991
rect 5549 13957 5583 13991
rect 5583 13957 5592 13991
rect 5540 13948 5592 13957
rect 8208 14016 8260 14068
rect 4988 13880 5040 13932
rect 5356 13880 5408 13932
rect 5724 13880 5776 13932
rect 7748 13991 7800 14000
rect 7748 13957 7757 13991
rect 7757 13957 7791 13991
rect 7791 13957 7800 13991
rect 7748 13948 7800 13957
rect 8392 13948 8444 14000
rect 8576 13880 8628 13932
rect 8668 13923 8720 13932
rect 8668 13889 8677 13923
rect 8677 13889 8711 13923
rect 8711 13889 8720 13923
rect 8668 13880 8720 13889
rect 3976 13812 4028 13864
rect 4896 13812 4948 13864
rect 5632 13855 5684 13864
rect 5632 13821 5641 13855
rect 5641 13821 5675 13855
rect 5675 13821 5684 13855
rect 5632 13812 5684 13821
rect 6000 13812 6052 13864
rect 6368 13812 6420 13864
rect 2688 13744 2740 13796
rect 7196 13855 7248 13864
rect 7196 13821 7205 13855
rect 7205 13821 7239 13855
rect 7239 13821 7248 13855
rect 7196 13812 7248 13821
rect 7380 13812 7432 13864
rect 7656 13812 7708 13864
rect 7012 13744 7064 13796
rect 8668 13744 8720 13796
rect 2504 13719 2556 13728
rect 2504 13685 2513 13719
rect 2513 13685 2547 13719
rect 2547 13685 2556 13719
rect 2504 13676 2556 13685
rect 3700 13676 3752 13728
rect 4252 13719 4304 13728
rect 4252 13685 4261 13719
rect 4261 13685 4295 13719
rect 4295 13685 4304 13719
rect 4252 13676 4304 13685
rect 4712 13676 4764 13728
rect 6644 13676 6696 13728
rect 7472 13719 7524 13728
rect 7472 13685 7481 13719
rect 7481 13685 7515 13719
rect 7515 13685 7524 13719
rect 7472 13676 7524 13685
rect 8484 13719 8536 13728
rect 8484 13685 8493 13719
rect 8493 13685 8527 13719
rect 8527 13685 8536 13719
rect 8484 13676 8536 13685
rect 8852 13676 8904 13728
rect 9036 13719 9088 13728
rect 9036 13685 9045 13719
rect 9045 13685 9079 13719
rect 9079 13685 9088 13719
rect 9036 13676 9088 13685
rect 9312 14016 9364 14068
rect 10232 14016 10284 14068
rect 10416 14016 10468 14068
rect 11244 14016 11296 14068
rect 11336 14059 11388 14068
rect 11336 14025 11345 14059
rect 11345 14025 11379 14059
rect 11379 14025 11388 14059
rect 11336 14016 11388 14025
rect 11520 14016 11572 14068
rect 12256 14016 12308 14068
rect 12532 14016 12584 14068
rect 13176 14059 13228 14068
rect 13176 14025 13185 14059
rect 13185 14025 13219 14059
rect 13219 14025 13228 14059
rect 13176 14016 13228 14025
rect 13452 14059 13504 14068
rect 13452 14025 13461 14059
rect 13461 14025 13495 14059
rect 13495 14025 13504 14059
rect 13452 14016 13504 14025
rect 13636 14016 13688 14068
rect 9312 13923 9364 13932
rect 9312 13889 9321 13923
rect 9321 13889 9355 13923
rect 9355 13889 9364 13923
rect 9312 13880 9364 13889
rect 9588 13880 9640 13932
rect 9864 13923 9916 13932
rect 9864 13889 9873 13923
rect 9873 13889 9907 13923
rect 9907 13889 9916 13923
rect 9864 13880 9916 13889
rect 10140 13880 10192 13932
rect 10876 13880 10928 13932
rect 11704 13923 11756 13932
rect 11704 13889 11713 13923
rect 11713 13889 11747 13923
rect 11747 13889 11756 13923
rect 11704 13880 11756 13889
rect 11980 13991 12032 14000
rect 11980 13957 11989 13991
rect 11989 13957 12023 13991
rect 12023 13957 12032 13991
rect 11980 13948 12032 13957
rect 14924 14016 14976 14068
rect 20812 14016 20864 14068
rect 21088 14059 21140 14068
rect 21088 14025 21097 14059
rect 21097 14025 21131 14059
rect 21131 14025 21140 14059
rect 21088 14016 21140 14025
rect 12440 13880 12492 13932
rect 12532 13880 12584 13932
rect 12808 13880 12860 13932
rect 9496 13812 9548 13864
rect 11060 13812 11112 13864
rect 11520 13812 11572 13864
rect 12164 13855 12216 13864
rect 11336 13744 11388 13796
rect 11428 13744 11480 13796
rect 11704 13744 11756 13796
rect 12164 13821 12173 13855
rect 12173 13821 12207 13855
rect 12207 13821 12216 13855
rect 12164 13812 12216 13821
rect 13176 13880 13228 13932
rect 13728 13923 13780 13932
rect 13728 13889 13737 13923
rect 13737 13889 13771 13923
rect 13771 13889 13780 13923
rect 13728 13880 13780 13889
rect 14556 13880 14608 13932
rect 16304 13948 16356 14000
rect 13452 13812 13504 13864
rect 12808 13744 12860 13796
rect 14280 13744 14332 13796
rect 15016 13855 15068 13864
rect 15016 13821 15025 13855
rect 15025 13821 15059 13855
rect 15059 13821 15068 13855
rect 15016 13812 15068 13821
rect 15936 13880 15988 13932
rect 16212 13880 16264 13932
rect 16672 13880 16724 13932
rect 19892 13948 19944 14000
rect 20536 13948 20588 14000
rect 18696 13923 18748 13932
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 18788 13880 18840 13932
rect 18972 13880 19024 13932
rect 20444 13880 20496 13932
rect 21088 13880 21140 13932
rect 21272 13880 21324 13932
rect 21364 13923 21416 13932
rect 21364 13889 21373 13923
rect 21373 13889 21407 13923
rect 21407 13889 21416 13923
rect 21364 13880 21416 13889
rect 21456 13923 21508 13932
rect 21456 13889 21465 13923
rect 21465 13889 21499 13923
rect 21499 13889 21508 13923
rect 21456 13880 21508 13889
rect 21732 13880 21784 13932
rect 22376 13948 22428 14000
rect 23204 13948 23256 14000
rect 23572 13948 23624 14000
rect 23940 13948 23992 14000
rect 15292 13744 15344 13796
rect 10048 13719 10100 13728
rect 10048 13685 10057 13719
rect 10057 13685 10091 13719
rect 10091 13685 10100 13719
rect 10048 13676 10100 13685
rect 10140 13719 10192 13728
rect 10140 13685 10149 13719
rect 10149 13685 10183 13719
rect 10183 13685 10192 13719
rect 10140 13676 10192 13685
rect 10600 13676 10652 13728
rect 14740 13676 14792 13728
rect 14924 13719 14976 13728
rect 14924 13685 14933 13719
rect 14933 13685 14967 13719
rect 14967 13685 14976 13719
rect 14924 13676 14976 13685
rect 16028 13812 16080 13864
rect 20720 13812 20772 13864
rect 22100 13812 22152 13864
rect 15844 13744 15896 13796
rect 16304 13744 16356 13796
rect 18236 13744 18288 13796
rect 18328 13719 18380 13728
rect 18328 13685 18337 13719
rect 18337 13685 18371 13719
rect 18371 13685 18380 13719
rect 18328 13676 18380 13685
rect 20352 13744 20404 13796
rect 21640 13787 21692 13796
rect 21640 13753 21649 13787
rect 21649 13753 21683 13787
rect 21683 13753 21692 13787
rect 21640 13744 21692 13753
rect 22468 13880 22520 13932
rect 22652 13855 22704 13864
rect 22652 13821 22661 13855
rect 22661 13821 22695 13855
rect 22695 13821 22704 13855
rect 22652 13812 22704 13821
rect 23112 13812 23164 13864
rect 23940 13855 23992 13864
rect 23940 13821 23949 13855
rect 23949 13821 23983 13855
rect 23983 13821 23992 13855
rect 23940 13812 23992 13821
rect 25228 14016 25280 14068
rect 26424 13948 26476 14000
rect 26792 13948 26844 14000
rect 26976 14016 27028 14068
rect 28816 14016 28868 14068
rect 30932 14016 30984 14068
rect 32220 14016 32272 14068
rect 32404 14059 32456 14068
rect 32404 14025 32413 14059
rect 32413 14025 32447 14059
rect 32447 14025 32456 14059
rect 32404 14016 32456 14025
rect 24216 13880 24268 13932
rect 26240 13880 26292 13932
rect 26608 13923 26660 13932
rect 26608 13889 26617 13923
rect 26617 13889 26651 13923
rect 26651 13889 26660 13923
rect 26608 13880 26660 13889
rect 26516 13855 26568 13864
rect 26516 13821 26525 13855
rect 26525 13821 26559 13855
rect 26559 13821 26568 13855
rect 26516 13812 26568 13821
rect 22928 13787 22980 13796
rect 22928 13753 22937 13787
rect 22937 13753 22971 13787
rect 22971 13753 22980 13787
rect 22928 13744 22980 13753
rect 24584 13744 24636 13796
rect 20076 13676 20128 13728
rect 20536 13676 20588 13728
rect 20720 13719 20772 13728
rect 20720 13685 20729 13719
rect 20729 13685 20763 13719
rect 20763 13685 20772 13719
rect 20720 13676 20772 13685
rect 21824 13719 21876 13728
rect 21824 13685 21833 13719
rect 21833 13685 21867 13719
rect 21867 13685 21876 13719
rect 21824 13676 21876 13685
rect 22284 13719 22336 13728
rect 22284 13685 22293 13719
rect 22293 13685 22327 13719
rect 22327 13685 22336 13719
rect 22284 13676 22336 13685
rect 22468 13719 22520 13728
rect 22468 13685 22477 13719
rect 22477 13685 22511 13719
rect 22511 13685 22520 13719
rect 22468 13676 22520 13685
rect 22560 13719 22612 13728
rect 22560 13685 22569 13719
rect 22569 13685 22603 13719
rect 22603 13685 22612 13719
rect 22560 13676 22612 13685
rect 24124 13719 24176 13728
rect 24124 13685 24133 13719
rect 24133 13685 24167 13719
rect 24167 13685 24176 13719
rect 24124 13676 24176 13685
rect 26240 13676 26292 13728
rect 26700 13676 26752 13728
rect 26884 13880 26936 13932
rect 27436 13948 27488 14000
rect 27252 13923 27304 13932
rect 27252 13889 27261 13923
rect 27261 13889 27295 13923
rect 27295 13889 27304 13923
rect 27252 13880 27304 13889
rect 27804 13948 27856 14000
rect 27436 13812 27488 13864
rect 29276 13812 29328 13864
rect 29828 13923 29880 13932
rect 29828 13889 29837 13923
rect 29837 13889 29871 13923
rect 29871 13889 29880 13923
rect 29828 13880 29880 13889
rect 30288 13880 30340 13932
rect 31760 13880 31812 13932
rect 32128 13880 32180 13932
rect 26976 13744 27028 13796
rect 28264 13744 28316 13796
rect 28448 13744 28500 13796
rect 29184 13744 29236 13796
rect 30012 13812 30064 13864
rect 30564 13855 30616 13864
rect 30564 13821 30573 13855
rect 30573 13821 30607 13855
rect 30607 13821 30616 13855
rect 30564 13812 30616 13821
rect 26884 13676 26936 13728
rect 27160 13719 27212 13728
rect 27160 13685 27169 13719
rect 27169 13685 27203 13719
rect 27203 13685 27212 13719
rect 27160 13676 27212 13685
rect 27436 13719 27488 13728
rect 27436 13685 27445 13719
rect 27445 13685 27479 13719
rect 27479 13685 27488 13719
rect 27436 13676 27488 13685
rect 27712 13719 27764 13728
rect 27712 13685 27721 13719
rect 27721 13685 27755 13719
rect 27755 13685 27764 13719
rect 27712 13676 27764 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 3240 13472 3292 13524
rect 3976 13472 4028 13524
rect 4528 13472 4580 13524
rect 572 13404 624 13456
rect 3424 13404 3476 13456
rect 2780 13336 2832 13388
rect 4712 13404 4764 13456
rect 4988 13404 5040 13456
rect 6368 13404 6420 13456
rect 2504 13311 2556 13320
rect 2504 13277 2513 13311
rect 2513 13277 2547 13311
rect 2547 13277 2556 13311
rect 2504 13268 2556 13277
rect 2872 13268 2924 13320
rect 3700 13268 3752 13320
rect 2964 13200 3016 13252
rect 3976 13311 4028 13320
rect 3976 13277 3985 13311
rect 3985 13277 4019 13311
rect 4019 13277 4028 13311
rect 3976 13268 4028 13277
rect 4436 13336 4488 13388
rect 7840 13472 7892 13524
rect 8760 13472 8812 13524
rect 9588 13515 9640 13524
rect 9588 13481 9597 13515
rect 9597 13481 9631 13515
rect 9631 13481 9640 13515
rect 9588 13472 9640 13481
rect 9772 13472 9824 13524
rect 10232 13472 10284 13524
rect 11244 13515 11296 13524
rect 11244 13481 11253 13515
rect 11253 13481 11287 13515
rect 11287 13481 11296 13515
rect 11244 13472 11296 13481
rect 11428 13472 11480 13524
rect 12072 13472 12124 13524
rect 12440 13472 12492 13524
rect 7288 13447 7340 13456
rect 7288 13413 7312 13447
rect 7312 13413 7340 13447
rect 7288 13404 7340 13413
rect 7748 13404 7800 13456
rect 7472 13379 7524 13388
rect 7472 13345 7481 13379
rect 7481 13345 7515 13379
rect 7515 13345 7524 13379
rect 7472 13336 7524 13345
rect 7656 13336 7708 13388
rect 12532 13404 12584 13456
rect 13636 13472 13688 13524
rect 14556 13472 14608 13524
rect 17776 13472 17828 13524
rect 4344 13268 4396 13320
rect 4620 13311 4672 13320
rect 4620 13277 4629 13311
rect 4629 13277 4663 13311
rect 4663 13277 4672 13311
rect 4620 13268 4672 13277
rect 3700 13132 3752 13184
rect 4344 13175 4396 13184
rect 4344 13141 4353 13175
rect 4353 13141 4387 13175
rect 4387 13141 4396 13175
rect 4344 13132 4396 13141
rect 4896 13200 4948 13252
rect 4620 13132 4672 13184
rect 5448 13132 5500 13184
rect 5816 13311 5868 13320
rect 5816 13277 5825 13311
rect 5825 13277 5859 13311
rect 5859 13277 5868 13311
rect 5816 13268 5868 13277
rect 5908 13268 5960 13320
rect 6276 13268 6328 13320
rect 5632 13200 5684 13252
rect 8484 13268 8536 13320
rect 10140 13336 10192 13388
rect 7380 13200 7432 13252
rect 7656 13200 7708 13252
rect 7840 13243 7892 13252
rect 7840 13209 7849 13243
rect 7849 13209 7883 13243
rect 7883 13209 7892 13243
rect 7840 13200 7892 13209
rect 6184 13132 6236 13184
rect 6736 13132 6788 13184
rect 8852 13200 8904 13252
rect 9864 13268 9916 13320
rect 12808 13336 12860 13388
rect 12992 13336 13044 13388
rect 13084 13379 13136 13388
rect 13084 13345 13093 13379
rect 13093 13345 13127 13379
rect 13127 13345 13136 13379
rect 13084 13336 13136 13345
rect 11704 13268 11756 13320
rect 11888 13268 11940 13320
rect 12256 13268 12308 13320
rect 10140 13200 10192 13252
rect 10968 13200 11020 13252
rect 8208 13132 8260 13184
rect 10876 13132 10928 13184
rect 13084 13200 13136 13252
rect 13544 13336 13596 13388
rect 13268 13311 13320 13320
rect 13268 13277 13277 13311
rect 13277 13277 13311 13311
rect 13311 13277 13320 13311
rect 13268 13268 13320 13277
rect 14740 13268 14792 13320
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 15844 13268 15896 13320
rect 17224 13268 17276 13320
rect 14096 13243 14148 13252
rect 14096 13209 14105 13243
rect 14105 13209 14139 13243
rect 14139 13209 14148 13243
rect 14096 13200 14148 13209
rect 15936 13200 15988 13252
rect 16672 13200 16724 13252
rect 17592 13200 17644 13252
rect 18696 13472 18748 13524
rect 20076 13472 20128 13524
rect 18604 13404 18656 13456
rect 22560 13472 22612 13524
rect 22928 13472 22980 13524
rect 28356 13472 28408 13524
rect 28632 13472 28684 13524
rect 30380 13472 30432 13524
rect 31760 13472 31812 13524
rect 18972 13268 19024 13320
rect 19524 13268 19576 13320
rect 19800 13268 19852 13320
rect 21272 13404 21324 13456
rect 21640 13404 21692 13456
rect 22376 13404 22428 13456
rect 25780 13404 25832 13456
rect 20352 13336 20404 13388
rect 20536 13200 20588 13252
rect 20812 13268 20864 13320
rect 13452 13175 13504 13184
rect 13452 13141 13461 13175
rect 13461 13141 13495 13175
rect 13495 13141 13504 13175
rect 13452 13132 13504 13141
rect 13912 13132 13964 13184
rect 14372 13132 14424 13184
rect 14924 13132 14976 13184
rect 18696 13132 18748 13184
rect 21364 13268 21416 13320
rect 21732 13336 21784 13388
rect 24860 13336 24912 13388
rect 24124 13268 24176 13320
rect 24400 13311 24452 13320
rect 24400 13277 24409 13311
rect 24409 13277 24443 13311
rect 24443 13277 24452 13311
rect 24400 13268 24452 13277
rect 21272 13200 21324 13252
rect 21548 13132 21600 13184
rect 22376 13200 22428 13252
rect 26056 13200 26108 13252
rect 23112 13132 23164 13184
rect 24584 13132 24636 13184
rect 27804 13311 27856 13320
rect 27804 13277 27813 13311
rect 27813 13277 27847 13311
rect 27847 13277 27856 13311
rect 27804 13268 27856 13277
rect 29460 13404 29512 13456
rect 29920 13404 29972 13456
rect 28448 13268 28500 13320
rect 28540 13311 28592 13320
rect 28540 13277 28549 13311
rect 28549 13277 28583 13311
rect 28583 13277 28592 13311
rect 28540 13268 28592 13277
rect 30564 13336 30616 13388
rect 32220 13379 32272 13388
rect 32220 13345 32229 13379
rect 32229 13345 32263 13379
rect 32263 13345 32272 13379
rect 32220 13336 32272 13345
rect 28908 13311 28960 13320
rect 28908 13277 28917 13311
rect 28917 13277 28951 13311
rect 28951 13277 28960 13311
rect 28908 13268 28960 13277
rect 30288 13268 30340 13320
rect 30932 13311 30984 13320
rect 30932 13277 30941 13311
rect 30941 13277 30975 13311
rect 30975 13277 30984 13311
rect 30932 13268 30984 13277
rect 31208 13311 31260 13320
rect 31208 13277 31217 13311
rect 31217 13277 31251 13311
rect 31251 13277 31260 13311
rect 31208 13268 31260 13277
rect 29736 13200 29788 13252
rect 30104 13200 30156 13252
rect 30656 13200 30708 13252
rect 30840 13200 30892 13252
rect 27712 13132 27764 13184
rect 28448 13132 28500 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 2504 12928 2556 12980
rect 6092 12928 6144 12980
rect 6460 12928 6512 12980
rect 6736 12928 6788 12980
rect 3240 12835 3292 12844
rect 3240 12801 3249 12835
rect 3249 12801 3283 12835
rect 3283 12801 3292 12835
rect 3240 12792 3292 12801
rect 3608 12835 3660 12844
rect 3608 12801 3617 12835
rect 3617 12801 3651 12835
rect 3651 12801 3660 12835
rect 3608 12792 3660 12801
rect 3792 12835 3844 12844
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 3884 12792 3936 12844
rect 4528 12792 4580 12844
rect 3148 12656 3200 12708
rect 3240 12656 3292 12708
rect 5264 12835 5316 12844
rect 5264 12801 5273 12835
rect 5273 12801 5307 12835
rect 5307 12801 5316 12835
rect 5264 12792 5316 12801
rect 5080 12699 5132 12708
rect 5080 12665 5089 12699
rect 5089 12665 5123 12699
rect 5123 12665 5132 12699
rect 5080 12656 5132 12665
rect 3792 12588 3844 12640
rect 5264 12588 5316 12640
rect 5724 12860 5776 12912
rect 8208 12928 8260 12980
rect 5908 12835 5960 12844
rect 5908 12801 5917 12835
rect 5917 12801 5951 12835
rect 5951 12801 5960 12835
rect 5908 12792 5960 12801
rect 7656 12860 7708 12912
rect 14096 12928 14148 12980
rect 15476 12928 15528 12980
rect 6552 12835 6604 12844
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 7012 12792 7064 12844
rect 7288 12792 7340 12844
rect 8576 12792 8628 12844
rect 8760 12792 8812 12844
rect 10416 12860 10468 12912
rect 12532 12860 12584 12912
rect 15660 12903 15712 12912
rect 15660 12869 15669 12903
rect 15669 12869 15703 12903
rect 15703 12869 15712 12903
rect 15660 12860 15712 12869
rect 16764 12903 16816 12912
rect 8944 12835 8996 12844
rect 8944 12801 8953 12835
rect 8953 12801 8987 12835
rect 8987 12801 8996 12835
rect 8944 12792 8996 12801
rect 9496 12835 9548 12844
rect 9496 12801 9505 12835
rect 9505 12801 9539 12835
rect 9539 12801 9548 12835
rect 9496 12792 9548 12801
rect 9864 12792 9916 12844
rect 10048 12792 10100 12844
rect 11428 12792 11480 12844
rect 11796 12835 11848 12844
rect 11796 12801 11805 12835
rect 11805 12801 11839 12835
rect 11839 12801 11848 12835
rect 11796 12792 11848 12801
rect 11888 12792 11940 12844
rect 11980 12792 12032 12844
rect 12348 12835 12400 12844
rect 12348 12801 12357 12835
rect 12357 12801 12391 12835
rect 12391 12801 12400 12835
rect 12348 12792 12400 12801
rect 15108 12792 15160 12844
rect 15292 12792 15344 12844
rect 15384 12792 15436 12844
rect 6184 12724 6236 12776
rect 6276 12724 6328 12776
rect 6552 12656 6604 12708
rect 6828 12656 6880 12708
rect 7104 12767 7156 12776
rect 7104 12733 7113 12767
rect 7113 12733 7147 12767
rect 7147 12733 7156 12767
rect 7104 12724 7156 12733
rect 9312 12724 9364 12776
rect 10876 12724 10928 12776
rect 11244 12767 11296 12776
rect 11244 12733 11253 12767
rect 11253 12733 11287 12767
rect 11287 12733 11296 12767
rect 11244 12724 11296 12733
rect 12440 12724 12492 12776
rect 12532 12724 12584 12776
rect 12992 12724 13044 12776
rect 14924 12724 14976 12776
rect 16764 12869 16773 12903
rect 16773 12869 16807 12903
rect 16807 12869 16816 12903
rect 16764 12860 16816 12869
rect 20536 12928 20588 12980
rect 22744 12928 22796 12980
rect 23756 12928 23808 12980
rect 23940 12928 23992 12980
rect 15936 12835 15988 12844
rect 15936 12801 15945 12835
rect 15945 12801 15979 12835
rect 15979 12801 15988 12835
rect 15936 12792 15988 12801
rect 16028 12792 16080 12844
rect 16488 12792 16540 12844
rect 16396 12724 16448 12776
rect 8760 12656 8812 12708
rect 7012 12588 7064 12640
rect 7932 12588 7984 12640
rect 9128 12631 9180 12640
rect 9128 12597 9137 12631
rect 9137 12597 9171 12631
rect 9171 12597 9180 12631
rect 9128 12588 9180 12597
rect 9312 12631 9364 12640
rect 9312 12597 9321 12631
rect 9321 12597 9355 12631
rect 9355 12597 9364 12631
rect 9312 12588 9364 12597
rect 9496 12588 9548 12640
rect 9772 12656 9824 12708
rect 10600 12656 10652 12708
rect 10048 12588 10100 12640
rect 10876 12631 10928 12640
rect 10876 12597 10885 12631
rect 10885 12597 10919 12631
rect 10919 12597 10928 12631
rect 10876 12588 10928 12597
rect 11152 12631 11204 12640
rect 11152 12597 11161 12631
rect 11161 12597 11195 12631
rect 11195 12597 11204 12631
rect 11152 12588 11204 12597
rect 12072 12588 12124 12640
rect 12532 12588 12584 12640
rect 14832 12656 14884 12708
rect 16948 12724 17000 12776
rect 13728 12588 13780 12640
rect 15200 12588 15252 12640
rect 15476 12588 15528 12640
rect 15660 12588 15712 12640
rect 16212 12631 16264 12640
rect 16212 12597 16221 12631
rect 16221 12597 16255 12631
rect 16255 12597 16264 12631
rect 16212 12588 16264 12597
rect 16304 12588 16356 12640
rect 17316 12835 17368 12844
rect 17316 12801 17325 12835
rect 17325 12801 17359 12835
rect 17359 12801 17368 12835
rect 17316 12792 17368 12801
rect 18512 12792 18564 12844
rect 18696 12835 18748 12844
rect 18696 12801 18705 12835
rect 18705 12801 18739 12835
rect 18739 12801 18748 12835
rect 18696 12792 18748 12801
rect 20076 12835 20128 12844
rect 20076 12801 20085 12835
rect 20085 12801 20119 12835
rect 20119 12801 20128 12835
rect 20076 12792 20128 12801
rect 21088 12860 21140 12912
rect 17960 12724 18012 12776
rect 18788 12724 18840 12776
rect 21640 12724 21692 12776
rect 22100 12792 22152 12844
rect 22192 12835 22244 12844
rect 22192 12801 22201 12835
rect 22201 12801 22235 12835
rect 22235 12801 22244 12835
rect 22192 12792 22244 12801
rect 22468 12792 22520 12844
rect 23940 12792 23992 12844
rect 24400 12928 24452 12980
rect 24676 12928 24728 12980
rect 21916 12724 21968 12776
rect 22652 12724 22704 12776
rect 23204 12724 23256 12776
rect 17592 12656 17644 12708
rect 17776 12656 17828 12708
rect 22468 12656 22520 12708
rect 17316 12588 17368 12640
rect 18788 12588 18840 12640
rect 18880 12588 18932 12640
rect 21640 12588 21692 12640
rect 22836 12588 22888 12640
rect 23664 12724 23716 12776
rect 26148 12860 26200 12912
rect 28908 12928 28960 12980
rect 29552 12928 29604 12980
rect 30104 12928 30156 12980
rect 31668 12928 31720 12980
rect 28080 12860 28132 12912
rect 28172 12903 28224 12912
rect 28172 12869 28181 12903
rect 28181 12869 28215 12903
rect 28215 12869 28224 12903
rect 28172 12860 28224 12869
rect 30564 12860 30616 12912
rect 24768 12835 24820 12844
rect 24768 12801 24777 12835
rect 24777 12801 24811 12835
rect 24811 12801 24820 12835
rect 24768 12792 24820 12801
rect 24860 12835 24912 12844
rect 24860 12801 24869 12835
rect 24869 12801 24903 12835
rect 24903 12801 24912 12835
rect 24860 12792 24912 12801
rect 26056 12835 26108 12844
rect 26056 12801 26065 12835
rect 26065 12801 26099 12835
rect 26099 12801 26108 12835
rect 26056 12792 26108 12801
rect 27160 12835 27212 12844
rect 27160 12801 27169 12835
rect 27169 12801 27203 12835
rect 27203 12801 27212 12835
rect 27160 12792 27212 12801
rect 27436 12835 27488 12844
rect 27436 12801 27445 12835
rect 27445 12801 27479 12835
rect 27479 12801 27488 12835
rect 27436 12792 27488 12801
rect 24676 12656 24728 12708
rect 26884 12724 26936 12776
rect 27252 12767 27304 12776
rect 27252 12733 27261 12767
rect 27261 12733 27295 12767
rect 27295 12733 27304 12767
rect 27252 12724 27304 12733
rect 30288 12835 30340 12844
rect 30288 12801 30297 12835
rect 30297 12801 30331 12835
rect 30331 12801 30340 12835
rect 30288 12792 30340 12801
rect 30656 12792 30708 12844
rect 31208 12792 31260 12844
rect 28632 12724 28684 12776
rect 32496 12835 32548 12844
rect 32496 12801 32505 12835
rect 32505 12801 32539 12835
rect 32539 12801 32548 12835
rect 32496 12792 32548 12801
rect 23756 12631 23808 12640
rect 23756 12597 23765 12631
rect 23765 12597 23799 12631
rect 23799 12597 23808 12631
rect 23756 12588 23808 12597
rect 24124 12588 24176 12640
rect 24400 12588 24452 12640
rect 25044 12631 25096 12640
rect 25044 12597 25053 12631
rect 25053 12597 25087 12631
rect 25087 12597 25096 12631
rect 25044 12588 25096 12597
rect 25780 12631 25832 12640
rect 25780 12597 25789 12631
rect 25789 12597 25823 12631
rect 25823 12597 25832 12631
rect 25780 12588 25832 12597
rect 26608 12588 26660 12640
rect 30932 12588 30984 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 3056 12427 3108 12436
rect 3056 12393 3065 12427
rect 3065 12393 3099 12427
rect 3099 12393 3108 12427
rect 3056 12384 3108 12393
rect 2780 12248 2832 12300
rect 3792 12316 3844 12368
rect 4988 12384 5040 12436
rect 6368 12384 6420 12436
rect 6828 12384 6880 12436
rect 6920 12384 6972 12436
rect 7932 12384 7984 12436
rect 9312 12384 9364 12436
rect 3056 12248 3108 12300
rect 2872 12223 2924 12232
rect 2872 12189 2881 12223
rect 2881 12189 2915 12223
rect 2915 12189 2924 12223
rect 2872 12180 2924 12189
rect 3424 12180 3476 12232
rect 3700 12180 3752 12232
rect 2228 12087 2280 12096
rect 2228 12053 2237 12087
rect 2237 12053 2271 12087
rect 2271 12053 2280 12087
rect 2228 12044 2280 12053
rect 2780 12155 2832 12164
rect 2780 12121 2789 12155
rect 2789 12121 2823 12155
rect 2823 12121 2832 12155
rect 4068 12180 4120 12232
rect 5080 12316 5132 12368
rect 4988 12223 5040 12232
rect 4988 12189 4997 12223
rect 4997 12189 5031 12223
rect 5031 12189 5040 12223
rect 4988 12180 5040 12189
rect 5080 12223 5132 12232
rect 5080 12189 5113 12223
rect 5113 12189 5132 12223
rect 5080 12180 5132 12189
rect 2780 12112 2832 12121
rect 2964 12044 3016 12096
rect 3516 12044 3568 12096
rect 5816 12316 5868 12368
rect 11428 12384 11480 12436
rect 15844 12384 15896 12436
rect 16396 12427 16448 12436
rect 16396 12393 16405 12427
rect 16405 12393 16439 12427
rect 16439 12393 16448 12427
rect 16396 12384 16448 12393
rect 16672 12384 16724 12436
rect 6092 12248 6144 12300
rect 5724 12180 5776 12232
rect 6552 12248 6604 12300
rect 8576 12248 8628 12300
rect 11796 12316 11848 12368
rect 12532 12316 12584 12368
rect 13084 12316 13136 12368
rect 20076 12384 20128 12436
rect 20536 12384 20588 12436
rect 21456 12384 21508 12436
rect 21916 12427 21968 12436
rect 21916 12393 21925 12427
rect 21925 12393 21959 12427
rect 21959 12393 21968 12427
rect 21916 12384 21968 12393
rect 22100 12384 22152 12436
rect 23296 12384 23348 12436
rect 23664 12427 23716 12436
rect 23664 12393 23673 12427
rect 23673 12393 23707 12427
rect 23707 12393 23716 12427
rect 23664 12384 23716 12393
rect 24400 12427 24452 12436
rect 24400 12393 24409 12427
rect 24409 12393 24443 12427
rect 24443 12393 24452 12427
rect 24400 12384 24452 12393
rect 24952 12427 25004 12436
rect 24952 12393 24961 12427
rect 24961 12393 24995 12427
rect 24995 12393 25004 12427
rect 24952 12384 25004 12393
rect 17224 12359 17276 12368
rect 17224 12325 17233 12359
rect 17233 12325 17267 12359
rect 17267 12325 17276 12359
rect 17224 12316 17276 12325
rect 18788 12316 18840 12368
rect 10232 12248 10284 12300
rect 6644 12180 6696 12232
rect 7012 12180 7064 12232
rect 7288 12180 7340 12232
rect 7472 12180 7524 12232
rect 9128 12223 9180 12232
rect 9128 12189 9144 12223
rect 9144 12189 9178 12223
rect 9178 12189 9180 12223
rect 9128 12180 9180 12189
rect 9312 12223 9364 12232
rect 9312 12189 9321 12223
rect 9321 12189 9355 12223
rect 9355 12189 9364 12223
rect 9312 12180 9364 12189
rect 9680 12180 9732 12232
rect 6552 12155 6604 12164
rect 6552 12121 6561 12155
rect 6561 12121 6595 12155
rect 6595 12121 6604 12155
rect 6552 12112 6604 12121
rect 7840 12155 7892 12164
rect 7840 12121 7849 12155
rect 7849 12121 7883 12155
rect 7883 12121 7892 12155
rect 7840 12112 7892 12121
rect 7932 12112 7984 12164
rect 11428 12180 11480 12232
rect 11704 12291 11756 12300
rect 11704 12257 11713 12291
rect 11713 12257 11747 12291
rect 11747 12257 11756 12291
rect 11704 12248 11756 12257
rect 12072 12248 12124 12300
rect 12808 12248 12860 12300
rect 16028 12248 16080 12300
rect 16764 12248 16816 12300
rect 10508 12112 10560 12164
rect 10784 12112 10836 12164
rect 10876 12112 10928 12164
rect 13084 12180 13136 12232
rect 13820 12180 13872 12232
rect 17592 12180 17644 12232
rect 21272 12248 21324 12300
rect 6920 12044 6972 12096
rect 8760 12044 8812 12096
rect 9404 12044 9456 12096
rect 9680 12044 9732 12096
rect 11888 12044 11940 12096
rect 12164 12044 12216 12096
rect 17132 12112 17184 12164
rect 21456 12180 21508 12232
rect 21640 12248 21692 12300
rect 22100 12223 22152 12232
rect 22100 12189 22109 12223
rect 22109 12189 22143 12223
rect 22143 12189 22152 12223
rect 22100 12180 22152 12189
rect 22744 12180 22796 12232
rect 23940 12316 23992 12368
rect 23020 12248 23072 12300
rect 23204 12248 23256 12300
rect 23756 12248 23808 12300
rect 24768 12316 24820 12368
rect 25320 12316 25372 12368
rect 25596 12427 25648 12436
rect 25596 12393 25605 12427
rect 25605 12393 25639 12427
rect 25639 12393 25648 12427
rect 25596 12384 25648 12393
rect 26608 12384 26660 12436
rect 26884 12427 26936 12436
rect 26884 12393 26893 12427
rect 26893 12393 26927 12427
rect 26927 12393 26936 12427
rect 26884 12384 26936 12393
rect 27160 12384 27212 12436
rect 27804 12384 27856 12436
rect 28080 12384 28132 12436
rect 29460 12384 29512 12436
rect 25504 12316 25556 12368
rect 25780 12316 25832 12368
rect 24584 12180 24636 12232
rect 24860 12180 24912 12232
rect 16580 12044 16632 12096
rect 19340 12112 19392 12164
rect 19432 12155 19484 12164
rect 19432 12121 19441 12155
rect 19441 12121 19475 12155
rect 19475 12121 19484 12155
rect 19432 12112 19484 12121
rect 19616 12155 19668 12164
rect 19616 12121 19625 12155
rect 19625 12121 19659 12155
rect 19659 12121 19668 12155
rect 19616 12112 19668 12121
rect 20996 12112 21048 12164
rect 21640 12112 21692 12164
rect 21824 12155 21876 12164
rect 21824 12121 21833 12155
rect 21833 12121 21867 12155
rect 21867 12121 21876 12155
rect 21824 12112 21876 12121
rect 22376 12155 22428 12164
rect 22376 12121 22385 12155
rect 22385 12121 22419 12155
rect 22419 12121 22428 12155
rect 22376 12112 22428 12121
rect 23480 12112 23532 12164
rect 25964 12248 26016 12300
rect 26148 12180 26200 12232
rect 28908 12316 28960 12368
rect 27160 12248 27212 12300
rect 28264 12248 28316 12300
rect 28540 12248 28592 12300
rect 29920 12291 29972 12300
rect 29920 12257 29929 12291
rect 29929 12257 29963 12291
rect 29963 12257 29972 12291
rect 29920 12248 29972 12257
rect 25964 12112 26016 12164
rect 26608 12112 26660 12164
rect 27804 12112 27856 12164
rect 18512 12044 18564 12096
rect 19064 12044 19116 12096
rect 19524 12044 19576 12096
rect 22192 12044 22244 12096
rect 22744 12044 22796 12096
rect 30932 12223 30984 12232
rect 30932 12189 30941 12223
rect 30941 12189 30975 12223
rect 30975 12189 30984 12223
rect 30932 12180 30984 12189
rect 32220 12223 32272 12232
rect 32220 12189 32229 12223
rect 32229 12189 32263 12223
rect 32263 12189 32272 12223
rect 32220 12180 32272 12189
rect 30380 12112 30432 12164
rect 30840 12112 30892 12164
rect 31208 12155 31260 12164
rect 31208 12121 31217 12155
rect 31217 12121 31251 12155
rect 31251 12121 31260 12155
rect 31208 12112 31260 12121
rect 28448 12044 28500 12096
rect 30472 12087 30524 12096
rect 30472 12053 30481 12087
rect 30481 12053 30515 12087
rect 30515 12053 30524 12087
rect 30472 12044 30524 12053
rect 30656 12044 30708 12096
rect 31484 12087 31536 12096
rect 31484 12053 31493 12087
rect 31493 12053 31527 12087
rect 31527 12053 31536 12087
rect 31484 12044 31536 12053
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 3516 11840 3568 11892
rect 2136 11704 2188 11756
rect 3332 11704 3384 11756
rect 3516 11747 3568 11756
rect 3516 11713 3525 11747
rect 3525 11713 3559 11747
rect 3559 11713 3568 11747
rect 3516 11704 3568 11713
rect 3608 11704 3660 11756
rect 4344 11840 4396 11892
rect 4436 11747 4488 11756
rect 4436 11713 4445 11747
rect 4445 11713 4479 11747
rect 4479 11713 4488 11747
rect 4436 11704 4488 11713
rect 5356 11840 5408 11892
rect 5632 11840 5684 11892
rect 5724 11840 5776 11892
rect 7012 11883 7064 11892
rect 3424 11636 3476 11688
rect 6460 11772 6512 11824
rect 7012 11849 7021 11883
rect 7021 11849 7055 11883
rect 7055 11849 7064 11883
rect 7012 11840 7064 11849
rect 7840 11840 7892 11892
rect 7196 11772 7248 11824
rect 7656 11772 7708 11824
rect 4804 11704 4856 11756
rect 5356 11704 5408 11756
rect 5632 11704 5684 11756
rect 6276 11704 6328 11756
rect 7012 11704 7064 11756
rect 1860 11568 1912 11620
rect 3056 11568 3108 11620
rect 3148 11568 3200 11620
rect 2504 11500 2556 11552
rect 2780 11500 2832 11552
rect 2964 11543 3016 11552
rect 2964 11509 2973 11543
rect 2973 11509 3007 11543
rect 3007 11509 3016 11543
rect 2964 11500 3016 11509
rect 3332 11543 3384 11552
rect 3332 11509 3341 11543
rect 3341 11509 3375 11543
rect 3375 11509 3384 11543
rect 3332 11500 3384 11509
rect 3516 11568 3568 11620
rect 5908 11568 5960 11620
rect 4068 11500 4120 11552
rect 5080 11500 5132 11552
rect 6000 11543 6052 11552
rect 6000 11509 6009 11543
rect 6009 11509 6043 11543
rect 6043 11509 6052 11543
rect 6000 11500 6052 11509
rect 6460 11568 6512 11620
rect 7196 11568 7248 11620
rect 9956 11840 10008 11892
rect 10232 11840 10284 11892
rect 10508 11772 10560 11824
rect 9588 11704 9640 11756
rect 10048 11704 10100 11756
rect 10416 11704 10468 11756
rect 9680 11636 9732 11688
rect 9956 11636 10008 11688
rect 10968 11840 11020 11892
rect 11152 11883 11204 11892
rect 11152 11849 11161 11883
rect 11161 11849 11195 11883
rect 11195 11849 11204 11883
rect 11152 11840 11204 11849
rect 12808 11840 12860 11892
rect 13728 11840 13780 11892
rect 11428 11704 11480 11756
rect 11796 11747 11848 11756
rect 11796 11713 11805 11747
rect 11805 11713 11839 11747
rect 11839 11713 11848 11747
rect 11796 11704 11848 11713
rect 12256 11704 12308 11756
rect 12348 11747 12400 11756
rect 12348 11713 12357 11747
rect 12357 11713 12391 11747
rect 12391 11713 12400 11747
rect 12348 11704 12400 11713
rect 12624 11772 12676 11824
rect 13084 11704 13136 11756
rect 14096 11772 14148 11824
rect 14556 11772 14608 11824
rect 15108 11840 15160 11892
rect 13360 11704 13412 11756
rect 14832 11747 14884 11756
rect 14832 11713 14841 11747
rect 14841 11713 14875 11747
rect 14875 11713 14884 11747
rect 14832 11704 14884 11713
rect 15016 11747 15068 11756
rect 15016 11713 15025 11747
rect 15025 11713 15059 11747
rect 15059 11713 15068 11747
rect 15016 11704 15068 11713
rect 15476 11772 15528 11824
rect 16120 11772 16172 11824
rect 17132 11883 17184 11892
rect 17132 11849 17141 11883
rect 17141 11849 17175 11883
rect 17175 11849 17184 11883
rect 17132 11840 17184 11849
rect 17500 11883 17552 11892
rect 17500 11849 17509 11883
rect 17509 11849 17543 11883
rect 17543 11849 17552 11883
rect 17500 11840 17552 11849
rect 17960 11883 18012 11892
rect 17960 11849 17969 11883
rect 17969 11849 18003 11883
rect 18003 11849 18012 11883
rect 17960 11840 18012 11849
rect 16396 11704 16448 11756
rect 11612 11679 11664 11688
rect 11612 11645 11621 11679
rect 11621 11645 11655 11679
rect 11655 11645 11664 11679
rect 11612 11636 11664 11645
rect 12072 11636 12124 11688
rect 12992 11679 13044 11688
rect 12992 11645 13001 11679
rect 13001 11645 13035 11679
rect 13035 11645 13044 11679
rect 12992 11636 13044 11645
rect 15476 11636 15528 11688
rect 16304 11636 16356 11688
rect 17040 11704 17092 11756
rect 17868 11772 17920 11824
rect 18328 11772 18380 11824
rect 17224 11636 17276 11688
rect 18512 11704 18564 11756
rect 19064 11883 19116 11892
rect 19064 11849 19073 11883
rect 19073 11849 19107 11883
rect 19107 11849 19116 11883
rect 19064 11840 19116 11849
rect 20720 11883 20772 11892
rect 20720 11849 20729 11883
rect 20729 11849 20763 11883
rect 20763 11849 20772 11883
rect 20720 11840 20772 11849
rect 21364 11840 21416 11892
rect 21548 11840 21600 11892
rect 24124 11815 24176 11824
rect 24124 11781 24133 11815
rect 24133 11781 24167 11815
rect 24167 11781 24176 11815
rect 24124 11772 24176 11781
rect 24860 11840 24912 11892
rect 29184 11840 29236 11892
rect 32220 11840 32272 11892
rect 25596 11772 25648 11824
rect 27160 11772 27212 11824
rect 28540 11772 28592 11824
rect 17868 11636 17920 11688
rect 17960 11636 18012 11688
rect 10692 11568 10744 11620
rect 6552 11500 6604 11552
rect 6736 11543 6788 11552
rect 6736 11509 6745 11543
rect 6745 11509 6779 11543
rect 6779 11509 6788 11543
rect 6736 11500 6788 11509
rect 7288 11500 7340 11552
rect 7840 11500 7892 11552
rect 8024 11500 8076 11552
rect 8208 11500 8260 11552
rect 8668 11543 8720 11552
rect 8668 11509 8677 11543
rect 8677 11509 8711 11543
rect 8711 11509 8720 11543
rect 8668 11500 8720 11509
rect 9128 11500 9180 11552
rect 9680 11500 9732 11552
rect 9956 11500 10008 11552
rect 10416 11543 10468 11552
rect 10416 11509 10425 11543
rect 10425 11509 10459 11543
rect 10459 11509 10468 11543
rect 10416 11500 10468 11509
rect 10508 11500 10560 11552
rect 11152 11500 11204 11552
rect 11244 11500 11296 11552
rect 11888 11500 11940 11552
rect 12256 11568 12308 11620
rect 17316 11568 17368 11620
rect 17408 11568 17460 11620
rect 20352 11747 20404 11756
rect 20352 11713 20361 11747
rect 20361 11713 20395 11747
rect 20395 11713 20404 11747
rect 20352 11704 20404 11713
rect 20536 11747 20588 11756
rect 20536 11713 20545 11747
rect 20545 11713 20579 11747
rect 20579 11713 20588 11747
rect 20536 11704 20588 11713
rect 20628 11704 20680 11756
rect 25044 11704 25096 11756
rect 25320 11704 25372 11756
rect 25780 11704 25832 11756
rect 28080 11704 28132 11756
rect 28632 11747 28684 11756
rect 28632 11713 28641 11747
rect 28641 11713 28675 11747
rect 28675 11713 28684 11747
rect 28632 11704 28684 11713
rect 28724 11747 28776 11756
rect 28724 11713 28733 11747
rect 28733 11713 28767 11747
rect 28767 11713 28776 11747
rect 28724 11704 28776 11713
rect 29368 11772 29420 11824
rect 31484 11772 31536 11824
rect 32220 11747 32272 11756
rect 32220 11713 32229 11747
rect 32229 11713 32263 11747
rect 32263 11713 32272 11747
rect 32220 11704 32272 11713
rect 19340 11636 19392 11688
rect 21640 11636 21692 11688
rect 22376 11636 22428 11688
rect 22744 11636 22796 11688
rect 30564 11679 30616 11688
rect 30564 11645 30573 11679
rect 30573 11645 30607 11679
rect 30607 11645 30616 11679
rect 30564 11636 30616 11645
rect 12164 11543 12216 11552
rect 12164 11509 12173 11543
rect 12173 11509 12207 11543
rect 12207 11509 12216 11543
rect 12164 11500 12216 11509
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 13360 11543 13412 11552
rect 13360 11509 13369 11543
rect 13369 11509 13403 11543
rect 13403 11509 13412 11543
rect 13360 11500 13412 11509
rect 14280 11543 14332 11552
rect 14280 11509 14289 11543
rect 14289 11509 14323 11543
rect 14323 11509 14332 11543
rect 14280 11500 14332 11509
rect 14740 11543 14792 11552
rect 14740 11509 14749 11543
rect 14749 11509 14783 11543
rect 14783 11509 14792 11543
rect 14740 11500 14792 11509
rect 15476 11500 15528 11552
rect 16488 11500 16540 11552
rect 16764 11543 16816 11552
rect 16764 11509 16773 11543
rect 16773 11509 16807 11543
rect 16807 11509 16816 11543
rect 16764 11500 16816 11509
rect 16856 11500 16908 11552
rect 18604 11543 18656 11552
rect 18604 11509 18613 11543
rect 18613 11509 18647 11543
rect 18647 11509 18656 11543
rect 18604 11500 18656 11509
rect 18696 11543 18748 11552
rect 18696 11509 18705 11543
rect 18705 11509 18739 11543
rect 18739 11509 18748 11543
rect 18696 11500 18748 11509
rect 18788 11500 18840 11552
rect 20536 11500 20588 11552
rect 22008 11568 22060 11620
rect 23296 11568 23348 11620
rect 25964 11568 26016 11620
rect 21364 11500 21416 11552
rect 23480 11500 23532 11552
rect 24032 11500 24084 11552
rect 24492 11500 24544 11552
rect 24768 11500 24820 11552
rect 26792 11500 26844 11552
rect 28448 11543 28500 11552
rect 28448 11509 28457 11543
rect 28457 11509 28491 11543
rect 28491 11509 28500 11543
rect 28448 11500 28500 11509
rect 29092 11500 29144 11552
rect 30472 11568 30524 11620
rect 30012 11543 30064 11552
rect 30012 11509 30021 11543
rect 30021 11509 30055 11543
rect 30055 11509 30064 11543
rect 30012 11500 30064 11509
rect 32404 11611 32456 11620
rect 32404 11577 32413 11611
rect 32413 11577 32447 11611
rect 32447 11577 32456 11611
rect 32404 11568 32456 11577
rect 30840 11500 30892 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 1676 11296 1728 11348
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 2504 11160 2556 11212
rect 3608 11296 3660 11348
rect 2872 11228 2924 11280
rect 3424 11228 3476 11280
rect 6276 11296 6328 11348
rect 6368 11296 6420 11348
rect 6828 11296 6880 11348
rect 2136 11135 2188 11144
rect 2136 11101 2145 11135
rect 2145 11101 2179 11135
rect 2179 11101 2188 11135
rect 2136 11092 2188 11101
rect 2228 11135 2280 11144
rect 2228 11101 2237 11135
rect 2237 11101 2271 11135
rect 2271 11101 2280 11135
rect 2228 11092 2280 11101
rect 4252 11160 4304 11212
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 3332 11092 3384 11144
rect 2688 11024 2740 11076
rect 3516 11092 3568 11144
rect 4160 11135 4212 11144
rect 4160 11101 4169 11135
rect 4169 11101 4203 11135
rect 4203 11101 4212 11135
rect 4160 11092 4212 11101
rect 4620 11092 4672 11144
rect 6552 11228 6604 11280
rect 2504 10999 2556 11008
rect 2504 10965 2513 10999
rect 2513 10965 2547 10999
rect 2547 10965 2556 10999
rect 2504 10956 2556 10965
rect 3056 10956 3108 11008
rect 3700 11024 3752 11076
rect 4252 11024 4304 11076
rect 3976 10956 4028 11008
rect 4436 11067 4488 11076
rect 4436 11033 4445 11067
rect 4445 11033 4479 11067
rect 4479 11033 4488 11067
rect 4436 11024 4488 11033
rect 5632 11092 5684 11144
rect 5264 11067 5316 11076
rect 5264 11033 5273 11067
rect 5273 11033 5307 11067
rect 5307 11033 5316 11067
rect 5264 11024 5316 11033
rect 4528 10956 4580 11008
rect 4712 10956 4764 11008
rect 4896 10956 4948 11008
rect 5172 10956 5224 11008
rect 5816 11024 5868 11076
rect 5724 10956 5776 11008
rect 6368 11135 6420 11144
rect 6368 11101 6377 11135
rect 6377 11101 6411 11135
rect 6411 11101 6420 11135
rect 6368 11092 6420 11101
rect 6644 11024 6696 11076
rect 7196 11296 7248 11348
rect 9680 11296 9732 11348
rect 7748 11228 7800 11280
rect 7012 11092 7064 11144
rect 7288 11160 7340 11212
rect 7472 11160 7524 11212
rect 10416 11296 10468 11348
rect 11428 11296 11480 11348
rect 11888 11339 11940 11348
rect 11888 11305 11897 11339
rect 11897 11305 11931 11339
rect 11931 11305 11940 11339
rect 11888 11296 11940 11305
rect 12900 11296 12952 11348
rect 13544 11296 13596 11348
rect 15568 11296 15620 11348
rect 16396 11296 16448 11348
rect 19524 11296 19576 11348
rect 19984 11296 20036 11348
rect 20444 11339 20496 11348
rect 20444 11305 20453 11339
rect 20453 11305 20487 11339
rect 20487 11305 20496 11339
rect 20444 11296 20496 11305
rect 20812 11296 20864 11348
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 7472 11067 7524 11076
rect 7472 11033 7481 11067
rect 7481 11033 7515 11067
rect 7515 11033 7524 11067
rect 7472 11024 7524 11033
rect 7748 11135 7800 11144
rect 7748 11101 7757 11135
rect 7757 11101 7791 11135
rect 7791 11101 7800 11135
rect 7748 11092 7800 11101
rect 8944 11160 8996 11212
rect 7288 10956 7340 11008
rect 7932 10956 7984 11008
rect 8116 11067 8168 11076
rect 8116 11033 8125 11067
rect 8125 11033 8159 11067
rect 8159 11033 8168 11067
rect 8116 11024 8168 11033
rect 8576 11135 8628 11144
rect 8576 11101 8585 11135
rect 8585 11101 8619 11135
rect 8619 11101 8628 11135
rect 8576 11092 8628 11101
rect 8760 11092 8812 11144
rect 9312 11092 9364 11144
rect 10692 11203 10744 11212
rect 10692 11169 10701 11203
rect 10701 11169 10735 11203
rect 10735 11169 10744 11203
rect 10692 11160 10744 11169
rect 14832 11228 14884 11280
rect 14096 11160 14148 11212
rect 14280 11160 14332 11212
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 10508 11135 10560 11144
rect 10508 11101 10517 11135
rect 10517 11101 10551 11135
rect 10551 11101 10560 11135
rect 10508 11092 10560 11101
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 10876 11135 10928 11144
rect 10876 11101 10885 11135
rect 10885 11101 10919 11135
rect 10919 11101 10928 11135
rect 10876 11092 10928 11101
rect 14464 11135 14516 11144
rect 14464 11101 14473 11135
rect 14473 11101 14507 11135
rect 14507 11101 14516 11135
rect 14464 11092 14516 11101
rect 8392 10999 8444 11008
rect 8392 10965 8401 10999
rect 8401 10965 8435 10999
rect 8435 10965 8444 10999
rect 8392 10956 8444 10965
rect 9128 10956 9180 11008
rect 12164 11024 12216 11076
rect 14832 11092 14884 11144
rect 15476 11228 15528 11280
rect 15936 11228 15988 11280
rect 17316 11228 17368 11280
rect 20444 11160 20496 11212
rect 20536 11203 20588 11212
rect 20536 11169 20545 11203
rect 20545 11169 20579 11203
rect 20579 11169 20588 11203
rect 20536 11160 20588 11169
rect 15752 11092 15804 11144
rect 15844 11092 15896 11144
rect 16488 11135 16540 11144
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 16488 11092 16540 11101
rect 16948 11092 17000 11144
rect 17500 11092 17552 11144
rect 18604 11092 18656 11144
rect 11980 10956 12032 11008
rect 12072 10956 12124 11008
rect 15016 10956 15068 11008
rect 15476 10956 15528 11008
rect 15660 10999 15712 11008
rect 15660 10965 15669 10999
rect 15669 10965 15703 10999
rect 15703 10965 15712 10999
rect 15660 10956 15712 10965
rect 17316 11024 17368 11076
rect 18696 11024 18748 11076
rect 19892 11024 19944 11076
rect 20720 11135 20772 11144
rect 20720 11101 20729 11135
rect 20729 11101 20763 11135
rect 20763 11101 20772 11135
rect 20720 11092 20772 11101
rect 22928 11296 22980 11348
rect 23664 11296 23716 11348
rect 23940 11296 23992 11348
rect 25504 11296 25556 11348
rect 26240 11339 26292 11348
rect 26240 11305 26249 11339
rect 26249 11305 26283 11339
rect 26283 11305 26292 11339
rect 26240 11296 26292 11305
rect 26792 11339 26844 11348
rect 26792 11305 26801 11339
rect 26801 11305 26835 11339
rect 26835 11305 26844 11339
rect 26792 11296 26844 11305
rect 28080 11339 28132 11348
rect 28080 11305 28089 11339
rect 28089 11305 28123 11339
rect 28123 11305 28132 11339
rect 28080 11296 28132 11305
rect 32128 11296 32180 11348
rect 22008 11228 22060 11280
rect 22468 11228 22520 11280
rect 21180 11160 21232 11212
rect 25964 11228 26016 11280
rect 22192 11135 22244 11144
rect 22192 11101 22201 11135
rect 22201 11101 22235 11135
rect 22235 11101 22244 11135
rect 22192 11092 22244 11101
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 23112 11092 23164 11144
rect 22284 11024 22336 11076
rect 22560 10956 22612 11008
rect 23296 11024 23348 11076
rect 24216 11092 24268 11144
rect 25688 11135 25740 11144
rect 25688 11101 25697 11135
rect 25697 11101 25731 11135
rect 25731 11101 25740 11135
rect 25688 11092 25740 11101
rect 26332 11228 26384 11280
rect 28632 11228 28684 11280
rect 27344 11160 27396 11212
rect 28264 11160 28316 11212
rect 28448 11160 28500 11212
rect 24032 10999 24084 11008
rect 24032 10965 24041 10999
rect 24041 10965 24075 10999
rect 24075 10965 24084 10999
rect 24032 10956 24084 10965
rect 25412 11024 25464 11076
rect 26608 11092 26660 11144
rect 26792 11135 26844 11144
rect 26792 11101 26801 11135
rect 26801 11101 26835 11135
rect 26835 11101 26844 11135
rect 26792 11092 26844 11101
rect 28540 11092 28592 11144
rect 30196 11135 30248 11144
rect 30196 11101 30205 11135
rect 30205 11101 30239 11135
rect 30239 11101 30248 11135
rect 30196 11092 30248 11101
rect 30380 11135 30432 11144
rect 30380 11101 30389 11135
rect 30389 11101 30423 11135
rect 30423 11101 30432 11135
rect 30380 11092 30432 11101
rect 30564 11135 30616 11144
rect 30564 11101 30573 11135
rect 30573 11101 30607 11135
rect 30607 11101 30616 11135
rect 30564 11092 30616 11101
rect 30840 11135 30892 11144
rect 30840 11101 30849 11135
rect 30849 11101 30883 11135
rect 30883 11101 30892 11135
rect 30840 11092 30892 11101
rect 26976 11024 27028 11076
rect 26608 10956 26660 11008
rect 27436 10956 27488 11008
rect 27804 11024 27856 11076
rect 31208 11024 31260 11076
rect 28264 10956 28316 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 3608 10752 3660 10804
rect 4436 10752 4488 10804
rect 4620 10752 4672 10804
rect 3976 10684 4028 10736
rect 4988 10752 5040 10804
rect 5724 10752 5776 10804
rect 5632 10684 5684 10736
rect 5908 10752 5960 10804
rect 6920 10795 6972 10804
rect 6920 10761 6929 10795
rect 6929 10761 6963 10795
rect 6963 10761 6972 10795
rect 6920 10752 6972 10761
rect 7472 10795 7524 10804
rect 7472 10761 7481 10795
rect 7481 10761 7515 10795
rect 7515 10761 7524 10795
rect 7472 10752 7524 10761
rect 9036 10752 9088 10804
rect 3148 10616 3200 10668
rect 3700 10616 3752 10668
rect 4344 10659 4396 10668
rect 4344 10625 4353 10659
rect 4353 10625 4387 10659
rect 4387 10625 4396 10659
rect 4344 10616 4396 10625
rect 4620 10616 4672 10668
rect 3148 10480 3200 10532
rect 4436 10480 4488 10532
rect 4896 10659 4948 10668
rect 4896 10625 4905 10659
rect 4905 10625 4939 10659
rect 4939 10625 4948 10659
rect 4896 10616 4948 10625
rect 5356 10616 5408 10668
rect 5080 10548 5132 10600
rect 6000 10663 6052 10668
rect 6000 10629 6009 10663
rect 6009 10629 6043 10663
rect 6043 10629 6052 10663
rect 6000 10616 6052 10629
rect 6644 10659 6696 10668
rect 6644 10625 6653 10659
rect 6653 10625 6687 10659
rect 6687 10625 6696 10659
rect 6644 10616 6696 10625
rect 6736 10659 6788 10668
rect 6736 10625 6769 10659
rect 6769 10625 6788 10659
rect 6736 10616 6788 10625
rect 6552 10548 6604 10600
rect 7104 10591 7156 10600
rect 7104 10557 7113 10591
rect 7113 10557 7147 10591
rect 7147 10557 7156 10591
rect 7104 10548 7156 10557
rect 4528 10412 4580 10464
rect 5172 10455 5224 10464
rect 5172 10421 5181 10455
rect 5181 10421 5215 10455
rect 5215 10421 5224 10455
rect 5172 10412 5224 10421
rect 5540 10412 5592 10464
rect 6920 10480 6972 10532
rect 7564 10727 7616 10736
rect 7564 10693 7573 10727
rect 7573 10693 7607 10727
rect 7607 10693 7616 10727
rect 7564 10684 7616 10693
rect 9312 10684 9364 10736
rect 11612 10684 11664 10736
rect 12716 10752 12768 10804
rect 12256 10684 12308 10736
rect 14004 10684 14056 10736
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 7748 10659 7800 10668
rect 7748 10625 7757 10659
rect 7757 10625 7791 10659
rect 7791 10625 7800 10659
rect 7748 10616 7800 10625
rect 9956 10616 10008 10668
rect 10140 10616 10192 10668
rect 10968 10616 11020 10668
rect 11428 10616 11480 10668
rect 11704 10659 11756 10668
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 11980 10659 12032 10668
rect 11980 10625 11989 10659
rect 11989 10625 12023 10659
rect 12023 10625 12032 10659
rect 11980 10616 12032 10625
rect 7656 10548 7708 10600
rect 8392 10548 8444 10600
rect 9588 10548 9640 10600
rect 12716 10591 12768 10600
rect 12716 10557 12725 10591
rect 12725 10557 12759 10591
rect 12759 10557 12768 10591
rect 12716 10548 12768 10557
rect 13084 10616 13136 10668
rect 12808 10480 12860 10532
rect 14556 10659 14608 10668
rect 14556 10625 14565 10659
rect 14565 10625 14599 10659
rect 14599 10625 14608 10659
rect 14556 10616 14608 10625
rect 14372 10591 14424 10600
rect 14372 10557 14381 10591
rect 14381 10557 14415 10591
rect 14415 10557 14424 10591
rect 14372 10548 14424 10557
rect 5816 10412 5868 10464
rect 6092 10412 6144 10464
rect 6276 10412 6328 10464
rect 7380 10412 7432 10464
rect 9404 10412 9456 10464
rect 9680 10412 9732 10464
rect 11428 10412 11480 10464
rect 11704 10412 11756 10464
rect 12164 10455 12216 10464
rect 12164 10421 12173 10455
rect 12173 10421 12207 10455
rect 12207 10421 12216 10455
rect 12164 10412 12216 10421
rect 12256 10412 12308 10464
rect 15936 10684 15988 10736
rect 15200 10616 15252 10668
rect 16212 10616 16264 10668
rect 16764 10616 16816 10668
rect 17408 10616 17460 10668
rect 17592 10659 17644 10668
rect 17592 10625 17601 10659
rect 17601 10625 17635 10659
rect 17635 10625 17644 10659
rect 17592 10616 17644 10625
rect 18420 10684 18472 10736
rect 18880 10684 18932 10736
rect 19432 10795 19484 10804
rect 19432 10761 19441 10795
rect 19441 10761 19475 10795
rect 19475 10761 19484 10795
rect 19432 10752 19484 10761
rect 20352 10752 20404 10804
rect 20536 10752 20588 10804
rect 20720 10752 20772 10804
rect 22100 10752 22152 10804
rect 22192 10795 22244 10804
rect 22192 10761 22201 10795
rect 22201 10761 22235 10795
rect 22235 10761 22244 10795
rect 22192 10752 22244 10761
rect 18788 10616 18840 10668
rect 13084 10412 13136 10464
rect 15476 10412 15528 10464
rect 15568 10412 15620 10464
rect 16120 10480 16172 10532
rect 18144 10548 18196 10600
rect 19064 10591 19116 10600
rect 19064 10557 19073 10591
rect 19073 10557 19107 10591
rect 19107 10557 19116 10591
rect 19064 10548 19116 10557
rect 19340 10616 19392 10668
rect 18052 10480 18104 10532
rect 18420 10480 18472 10532
rect 21088 10727 21140 10736
rect 21088 10693 21097 10727
rect 21097 10693 21131 10727
rect 21131 10693 21140 10727
rect 21088 10684 21140 10693
rect 20536 10659 20588 10668
rect 20536 10625 20545 10659
rect 20545 10625 20579 10659
rect 20579 10625 20588 10659
rect 20536 10616 20588 10625
rect 20904 10591 20956 10600
rect 20904 10557 20913 10591
rect 20913 10557 20947 10591
rect 20947 10557 20956 10591
rect 20904 10548 20956 10557
rect 21364 10616 21416 10668
rect 22560 10684 22612 10736
rect 23572 10684 23624 10736
rect 23940 10727 23992 10736
rect 23940 10693 23949 10727
rect 23949 10693 23983 10727
rect 23983 10693 23992 10727
rect 23940 10684 23992 10693
rect 26792 10752 26844 10804
rect 27068 10752 27120 10804
rect 27988 10795 28040 10804
rect 27988 10761 27997 10795
rect 27997 10761 28031 10795
rect 28031 10761 28040 10795
rect 27988 10752 28040 10761
rect 28356 10752 28408 10804
rect 30564 10752 30616 10804
rect 21824 10659 21876 10668
rect 21824 10625 21833 10659
rect 21833 10625 21867 10659
rect 21867 10625 21876 10659
rect 21824 10616 21876 10625
rect 22008 10659 22060 10668
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 22100 10616 22152 10668
rect 22652 10659 22704 10668
rect 22652 10625 22661 10659
rect 22661 10625 22695 10659
rect 22695 10625 22704 10659
rect 22652 10616 22704 10625
rect 22928 10659 22980 10668
rect 22928 10625 22937 10659
rect 22937 10625 22971 10659
rect 22971 10625 22980 10659
rect 22928 10616 22980 10625
rect 22192 10548 22244 10600
rect 22284 10548 22336 10600
rect 23572 10591 23624 10600
rect 23572 10557 23581 10591
rect 23581 10557 23615 10591
rect 23615 10557 23624 10591
rect 23572 10548 23624 10557
rect 16304 10455 16356 10464
rect 16304 10421 16313 10455
rect 16313 10421 16347 10455
rect 16347 10421 16356 10455
rect 16304 10412 16356 10421
rect 16764 10455 16816 10464
rect 16764 10421 16773 10455
rect 16773 10421 16807 10455
rect 16807 10421 16816 10455
rect 16764 10412 16816 10421
rect 17500 10412 17552 10464
rect 17776 10455 17828 10464
rect 17776 10421 17785 10455
rect 17785 10421 17819 10455
rect 17819 10421 17828 10455
rect 17776 10412 17828 10421
rect 19248 10455 19300 10464
rect 19248 10421 19257 10455
rect 19257 10421 19291 10455
rect 19291 10421 19300 10455
rect 19248 10412 19300 10421
rect 19340 10412 19392 10464
rect 19892 10455 19944 10464
rect 19892 10421 19901 10455
rect 19901 10421 19935 10455
rect 19935 10421 19944 10455
rect 19892 10412 19944 10421
rect 20720 10480 20772 10532
rect 20352 10455 20404 10464
rect 20352 10421 20361 10455
rect 20361 10421 20395 10455
rect 20395 10421 20404 10455
rect 20352 10412 20404 10421
rect 20628 10412 20680 10464
rect 20904 10412 20956 10464
rect 21548 10480 21600 10532
rect 22560 10480 22612 10532
rect 21180 10412 21232 10464
rect 21824 10412 21876 10464
rect 23388 10480 23440 10532
rect 22928 10455 22980 10464
rect 22928 10421 22937 10455
rect 22937 10421 22971 10455
rect 22971 10421 22980 10455
rect 22928 10412 22980 10421
rect 23020 10412 23072 10464
rect 23480 10455 23532 10464
rect 23480 10421 23489 10455
rect 23489 10421 23523 10455
rect 23523 10421 23532 10455
rect 23480 10412 23532 10421
rect 24124 10659 24176 10668
rect 24124 10625 24133 10659
rect 24133 10625 24167 10659
rect 24167 10625 24176 10659
rect 24124 10616 24176 10625
rect 24308 10616 24360 10668
rect 24584 10616 24636 10668
rect 24952 10659 25004 10668
rect 24952 10625 24961 10659
rect 24961 10625 24995 10659
rect 24995 10625 25004 10659
rect 24952 10616 25004 10625
rect 26148 10684 26200 10736
rect 30196 10684 30248 10736
rect 24768 10591 24820 10600
rect 24768 10557 24777 10591
rect 24777 10557 24811 10591
rect 24811 10557 24820 10591
rect 24768 10548 24820 10557
rect 24860 10548 24912 10600
rect 25688 10548 25740 10600
rect 26792 10616 26844 10668
rect 25872 10548 25924 10600
rect 26976 10548 27028 10600
rect 27344 10659 27396 10668
rect 27344 10625 27353 10659
rect 27353 10625 27387 10659
rect 27387 10625 27396 10659
rect 27344 10616 27396 10625
rect 25320 10412 25372 10464
rect 25596 10455 25648 10464
rect 25596 10421 25605 10455
rect 25605 10421 25639 10455
rect 25639 10421 25648 10455
rect 25596 10412 25648 10421
rect 25964 10480 26016 10532
rect 26148 10412 26200 10464
rect 26240 10455 26292 10464
rect 26240 10421 26249 10455
rect 26249 10421 26283 10455
rect 26283 10421 26292 10455
rect 26240 10412 26292 10421
rect 26608 10412 26660 10464
rect 28264 10659 28316 10668
rect 28264 10625 28273 10659
rect 28273 10625 28307 10659
rect 28307 10625 28316 10659
rect 28264 10616 28316 10625
rect 29552 10548 29604 10600
rect 29736 10548 29788 10600
rect 30472 10659 30524 10668
rect 30472 10625 30481 10659
rect 30481 10625 30515 10659
rect 30515 10625 30524 10659
rect 31392 10684 31444 10736
rect 30472 10616 30524 10625
rect 31024 10659 31076 10668
rect 31024 10625 31033 10659
rect 31033 10625 31067 10659
rect 31067 10625 31076 10659
rect 31024 10616 31076 10625
rect 31484 10616 31536 10668
rect 32128 10548 32180 10600
rect 29736 10412 29788 10464
rect 30564 10412 30616 10464
rect 31576 10412 31628 10464
rect 32404 10455 32456 10464
rect 32404 10421 32413 10455
rect 32413 10421 32447 10455
rect 32447 10421 32456 10455
rect 32404 10412 32456 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 4068 10208 4120 10260
rect 3976 10140 4028 10192
rect 5356 10140 5408 10192
rect 5724 10208 5776 10260
rect 6092 10208 6144 10260
rect 6736 10208 6788 10260
rect 8116 10208 8168 10260
rect 9220 10208 9272 10260
rect 9588 10251 9640 10260
rect 9588 10217 9597 10251
rect 9597 10217 9631 10251
rect 9631 10217 9640 10251
rect 9588 10208 9640 10217
rect 10140 10208 10192 10260
rect 10416 10208 10468 10260
rect 12900 10208 12952 10260
rect 15476 10208 15528 10260
rect 15936 10208 15988 10260
rect 16028 10251 16080 10260
rect 16028 10217 16037 10251
rect 16037 10217 16071 10251
rect 16071 10217 16080 10251
rect 16028 10208 16080 10217
rect 16948 10251 17000 10260
rect 16948 10217 16957 10251
rect 16957 10217 16991 10251
rect 16991 10217 17000 10251
rect 16948 10208 17000 10217
rect 17408 10251 17460 10260
rect 17408 10217 17417 10251
rect 17417 10217 17451 10251
rect 17451 10217 17460 10251
rect 17408 10208 17460 10217
rect 17500 10208 17552 10260
rect 19800 10208 19852 10260
rect 20720 10208 20772 10260
rect 22284 10208 22336 10260
rect 4896 10072 4948 10124
rect 3608 10004 3660 10056
rect 3884 10004 3936 10056
rect 4160 10047 4212 10056
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 4252 10004 4304 10056
rect 5264 10004 5316 10056
rect 3976 9979 4028 9988
rect 3976 9945 3985 9979
rect 3985 9945 4019 9979
rect 4019 9945 4028 9979
rect 3976 9936 4028 9945
rect 3332 9868 3384 9920
rect 5080 9936 5132 9988
rect 5816 10004 5868 10056
rect 6644 10140 6696 10192
rect 6920 10140 6972 10192
rect 7748 10140 7800 10192
rect 6276 10047 6328 10056
rect 6276 10013 6285 10047
rect 6285 10013 6319 10047
rect 6319 10013 6328 10047
rect 6276 10004 6328 10013
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 4896 9868 4948 9920
rect 5448 9868 5500 9920
rect 5632 9868 5684 9920
rect 5816 9868 5868 9920
rect 7104 9936 7156 9988
rect 8484 10072 8536 10124
rect 12992 10140 13044 10192
rect 9496 10072 9548 10124
rect 7564 9911 7616 9920
rect 7564 9877 7573 9911
rect 7573 9877 7607 9911
rect 7607 9877 7616 9911
rect 7564 9868 7616 9877
rect 9680 10004 9732 10056
rect 9864 10047 9916 10056
rect 9864 10013 9873 10047
rect 9873 10013 9907 10047
rect 9907 10013 9916 10047
rect 9864 10004 9916 10013
rect 10600 10072 10652 10124
rect 10968 10072 11020 10124
rect 14556 10072 14608 10124
rect 9036 9936 9088 9988
rect 10048 9936 10100 9988
rect 10324 9936 10376 9988
rect 12440 10004 12492 10056
rect 12716 10004 12768 10056
rect 12900 10004 12952 10056
rect 13268 10004 13320 10056
rect 13820 9936 13872 9988
rect 15844 10047 15896 10056
rect 15844 10013 15853 10047
rect 15853 10013 15887 10047
rect 15887 10013 15896 10047
rect 15844 10004 15896 10013
rect 16396 10047 16448 10056
rect 16396 10013 16405 10047
rect 16405 10013 16439 10047
rect 16439 10013 16448 10047
rect 16396 10004 16448 10013
rect 16580 10004 16632 10056
rect 18052 10072 18104 10124
rect 19616 10115 19668 10124
rect 19616 10081 19625 10115
rect 19625 10081 19659 10115
rect 19659 10081 19668 10115
rect 19616 10072 19668 10081
rect 20076 10140 20128 10192
rect 20352 10140 20404 10192
rect 22192 10140 22244 10192
rect 23388 10208 23440 10260
rect 27712 10251 27764 10260
rect 27712 10217 27721 10251
rect 27721 10217 27755 10251
rect 27755 10217 27764 10251
rect 27712 10208 27764 10217
rect 29644 10251 29696 10260
rect 29644 10217 29653 10251
rect 29653 10217 29687 10251
rect 29687 10217 29696 10251
rect 29644 10208 29696 10217
rect 16028 9936 16080 9988
rect 16488 9936 16540 9988
rect 17132 9936 17184 9988
rect 19156 10004 19208 10056
rect 8852 9868 8904 9920
rect 10876 9868 10928 9920
rect 11244 9911 11296 9920
rect 11244 9877 11253 9911
rect 11253 9877 11287 9911
rect 11287 9877 11296 9911
rect 11244 9868 11296 9877
rect 16580 9911 16632 9920
rect 16580 9877 16589 9911
rect 16589 9877 16623 9911
rect 16623 9877 16632 9911
rect 16580 9868 16632 9877
rect 16672 9911 16724 9920
rect 16672 9877 16681 9911
rect 16681 9877 16715 9911
rect 16715 9877 16724 9911
rect 19340 9936 19392 9988
rect 19432 9979 19484 9988
rect 19432 9945 19441 9979
rect 19441 9945 19475 9979
rect 19475 9945 19484 9979
rect 19432 9936 19484 9945
rect 20352 10004 20404 10056
rect 20076 9936 20128 9988
rect 22652 10072 22704 10124
rect 22928 10072 22980 10124
rect 22560 10047 22612 10056
rect 22560 10013 22569 10047
rect 22569 10013 22603 10047
rect 22603 10013 22612 10047
rect 22560 10004 22612 10013
rect 22836 10004 22888 10056
rect 24216 10004 24268 10056
rect 24492 10115 24544 10124
rect 24492 10081 24501 10115
rect 24501 10081 24535 10115
rect 24535 10081 24544 10115
rect 24492 10072 24544 10081
rect 28356 10072 28408 10124
rect 28632 10140 28684 10192
rect 26516 10004 26568 10056
rect 27528 10047 27580 10056
rect 27528 10013 27537 10047
rect 27537 10013 27571 10047
rect 27571 10013 27580 10047
rect 27528 10004 27580 10013
rect 27988 10004 28040 10056
rect 30104 10004 30156 10056
rect 31484 10047 31536 10056
rect 31484 10013 31493 10047
rect 31493 10013 31527 10047
rect 31527 10013 31536 10047
rect 31484 10004 31536 10013
rect 31576 10047 31628 10056
rect 31576 10013 31585 10047
rect 31585 10013 31619 10047
rect 31619 10013 31628 10047
rect 31576 10004 31628 10013
rect 32496 10047 32548 10056
rect 32496 10013 32505 10047
rect 32505 10013 32539 10047
rect 32539 10013 32548 10047
rect 32496 10004 32548 10013
rect 24768 9936 24820 9988
rect 27160 9979 27212 9988
rect 27160 9945 27169 9979
rect 27169 9945 27203 9979
rect 27203 9945 27212 9979
rect 27160 9936 27212 9945
rect 29736 9936 29788 9988
rect 30472 9979 30524 9988
rect 30472 9945 30481 9979
rect 30481 9945 30515 9979
rect 30515 9945 30524 9979
rect 30472 9936 30524 9945
rect 30656 9936 30708 9988
rect 16672 9868 16724 9877
rect 18236 9868 18288 9920
rect 20444 9868 20496 9920
rect 24676 9868 24728 9920
rect 25964 9868 26016 9920
rect 27344 9911 27396 9920
rect 27344 9877 27353 9911
rect 27353 9877 27387 9911
rect 27387 9877 27396 9911
rect 27344 9868 27396 9877
rect 29920 9868 29972 9920
rect 30748 9911 30800 9920
rect 30748 9877 30757 9911
rect 30757 9877 30791 9911
rect 30791 9877 30800 9911
rect 30748 9868 30800 9877
rect 31852 9868 31904 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 2780 9528 2832 9580
rect 3884 9664 3936 9716
rect 4712 9664 4764 9716
rect 3608 9639 3660 9648
rect 3608 9605 3617 9639
rect 3617 9605 3651 9639
rect 3651 9605 3660 9639
rect 3608 9596 3660 9605
rect 3516 9571 3568 9580
rect 3516 9537 3525 9571
rect 3525 9537 3559 9571
rect 3559 9537 3568 9571
rect 3516 9528 3568 9537
rect 3424 9460 3476 9512
rect 3884 9528 3936 9580
rect 4068 9460 4120 9512
rect 4252 9460 4304 9512
rect 4804 9528 4856 9580
rect 5356 9664 5408 9716
rect 5724 9664 5776 9716
rect 5816 9596 5868 9648
rect 4712 9392 4764 9444
rect 5264 9392 5316 9444
rect 6000 9664 6052 9716
rect 6736 9664 6788 9716
rect 6276 9596 6328 9648
rect 9220 9664 9272 9716
rect 9312 9664 9364 9716
rect 10048 9664 10100 9716
rect 10968 9664 11020 9716
rect 7012 9528 7064 9580
rect 7288 9571 7340 9580
rect 7288 9537 7297 9571
rect 7297 9537 7331 9571
rect 7331 9537 7340 9571
rect 7288 9528 7340 9537
rect 8944 9596 8996 9648
rect 12532 9664 12584 9716
rect 15844 9664 15896 9716
rect 16488 9707 16540 9716
rect 16488 9673 16497 9707
rect 16497 9673 16531 9707
rect 16531 9673 16540 9707
rect 16488 9664 16540 9673
rect 7656 9528 7708 9580
rect 7932 9571 7984 9580
rect 7932 9537 7941 9571
rect 7941 9537 7975 9571
rect 7975 9537 7984 9571
rect 7932 9528 7984 9537
rect 3792 9324 3844 9376
rect 5172 9324 5224 9376
rect 5448 9324 5500 9376
rect 7288 9392 7340 9444
rect 7748 9392 7800 9444
rect 7932 9392 7984 9444
rect 8300 9392 8352 9444
rect 6092 9324 6144 9376
rect 6460 9324 6512 9376
rect 6644 9324 6696 9376
rect 7472 9367 7524 9376
rect 7472 9333 7481 9367
rect 7481 9333 7515 9367
rect 7515 9333 7524 9367
rect 7472 9324 7524 9333
rect 7564 9324 7616 9376
rect 9864 9528 9916 9580
rect 10048 9571 10100 9580
rect 10048 9537 10057 9571
rect 10057 9537 10091 9571
rect 10091 9537 10100 9571
rect 10048 9528 10100 9537
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 8944 9503 8996 9512
rect 8944 9469 8953 9503
rect 8953 9469 8987 9503
rect 8987 9469 8996 9503
rect 8944 9460 8996 9469
rect 9496 9460 9548 9512
rect 9588 9460 9640 9512
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 10968 9571 11020 9580
rect 10968 9537 10977 9571
rect 10977 9537 11011 9571
rect 11011 9537 11020 9571
rect 10968 9528 11020 9537
rect 12900 9596 12952 9648
rect 12992 9596 13044 9648
rect 14372 9596 14424 9648
rect 16672 9664 16724 9716
rect 19156 9664 19208 9716
rect 20536 9664 20588 9716
rect 10876 9460 10928 9512
rect 9128 9392 9180 9444
rect 9680 9324 9732 9376
rect 10508 9392 10560 9444
rect 11152 9392 11204 9444
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 13360 9571 13412 9580
rect 13360 9537 13369 9571
rect 13369 9537 13403 9571
rect 13403 9537 13412 9571
rect 13360 9528 13412 9537
rect 13176 9460 13228 9512
rect 12440 9392 12492 9444
rect 13728 9460 13780 9512
rect 15568 9528 15620 9580
rect 16028 9571 16080 9580
rect 16028 9537 16037 9571
rect 16037 9537 16071 9571
rect 16071 9537 16080 9571
rect 16028 9528 16080 9537
rect 16580 9528 16632 9580
rect 17868 9528 17920 9580
rect 18144 9528 18196 9580
rect 18236 9571 18288 9580
rect 18236 9537 18245 9571
rect 18245 9537 18279 9571
rect 18279 9537 18288 9571
rect 18236 9528 18288 9537
rect 18328 9528 18380 9580
rect 20260 9596 20312 9648
rect 19800 9528 19852 9580
rect 19984 9528 20036 9580
rect 20444 9528 20496 9580
rect 20904 9571 20956 9580
rect 20904 9537 20913 9571
rect 20913 9537 20947 9571
rect 20947 9537 20956 9571
rect 20904 9528 20956 9537
rect 16672 9460 16724 9512
rect 12992 9367 13044 9376
rect 12992 9333 13001 9367
rect 13001 9333 13035 9367
rect 13035 9333 13044 9367
rect 12992 9324 13044 9333
rect 17776 9392 17828 9444
rect 18972 9460 19024 9512
rect 21180 9528 21232 9580
rect 21456 9571 21508 9580
rect 21456 9537 21465 9571
rect 21465 9537 21499 9571
rect 21499 9537 21508 9571
rect 21456 9528 21508 9537
rect 21916 9571 21968 9580
rect 21916 9537 21925 9571
rect 21925 9537 21959 9571
rect 21959 9537 21968 9571
rect 21916 9528 21968 9537
rect 22192 9571 22244 9580
rect 22192 9537 22201 9571
rect 22201 9537 22235 9571
rect 22235 9537 22244 9571
rect 22192 9528 22244 9537
rect 23020 9571 23072 9580
rect 23020 9537 23029 9571
rect 23029 9537 23063 9571
rect 23063 9537 23072 9571
rect 23020 9528 23072 9537
rect 21548 9460 21600 9512
rect 22744 9460 22796 9512
rect 24308 9460 24360 9512
rect 14096 9324 14148 9376
rect 14832 9324 14884 9376
rect 16120 9324 16172 9376
rect 16580 9324 16632 9376
rect 18144 9367 18196 9376
rect 18144 9333 18153 9367
rect 18153 9333 18187 9367
rect 18187 9333 18196 9367
rect 18144 9324 18196 9333
rect 19340 9324 19392 9376
rect 19984 9392 20036 9444
rect 21732 9392 21784 9444
rect 20996 9324 21048 9376
rect 22008 9324 22060 9376
rect 22284 9324 22336 9376
rect 22560 9367 22612 9376
rect 22560 9333 22569 9367
rect 22569 9333 22603 9367
rect 22603 9333 22612 9367
rect 22560 9324 22612 9333
rect 24676 9460 24728 9512
rect 27344 9596 27396 9648
rect 29000 9596 29052 9648
rect 29736 9639 29788 9648
rect 29736 9605 29745 9639
rect 29745 9605 29779 9639
rect 29779 9605 29788 9639
rect 29736 9596 29788 9605
rect 30472 9664 30524 9716
rect 26240 9528 26292 9580
rect 29276 9528 29328 9580
rect 30656 9596 30708 9648
rect 27436 9460 27488 9512
rect 24492 9392 24544 9444
rect 25136 9392 25188 9444
rect 25688 9392 25740 9444
rect 27252 9392 27304 9444
rect 27344 9392 27396 9444
rect 27712 9392 27764 9444
rect 26332 9324 26384 9376
rect 26516 9367 26568 9376
rect 26516 9333 26525 9367
rect 26525 9333 26559 9367
rect 26559 9333 26568 9367
rect 26516 9324 26568 9333
rect 27068 9324 27120 9376
rect 28356 9324 28408 9376
rect 30840 9324 30892 9376
rect 31116 9324 31168 9376
rect 31484 9664 31536 9716
rect 31852 9528 31904 9580
rect 32496 9571 32548 9580
rect 32496 9537 32505 9571
rect 32505 9537 32539 9571
rect 32539 9537 32548 9571
rect 32496 9528 32548 9537
rect 32312 9435 32364 9444
rect 32312 9401 32321 9435
rect 32321 9401 32355 9435
rect 32355 9401 32364 9435
rect 32312 9392 32364 9401
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 4068 9120 4120 9172
rect 5080 9120 5132 9172
rect 5816 9120 5868 9172
rect 6460 9120 6512 9172
rect 6736 9120 6788 9172
rect 9036 9120 9088 9172
rect 5448 9052 5500 9104
rect 6000 9052 6052 9104
rect 7196 9052 7248 9104
rect 9220 9120 9272 9172
rect 11796 9120 11848 9172
rect 10140 9052 10192 9104
rect 12164 9052 12216 9104
rect 5264 8984 5316 9036
rect 2964 8916 3016 8968
rect 3884 8916 3936 8968
rect 4160 8916 4212 8968
rect 4436 8959 4488 8968
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 4528 8916 4580 8968
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 4804 8916 4856 8968
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 5724 8916 5776 8968
rect 6092 8916 6144 8968
rect 3516 8848 3568 8900
rect 4344 8891 4396 8900
rect 4344 8857 4353 8891
rect 4353 8857 4387 8891
rect 4387 8857 4396 8891
rect 4344 8848 4396 8857
rect 4896 8780 4948 8832
rect 5816 8891 5868 8900
rect 5816 8857 5825 8891
rect 5825 8857 5859 8891
rect 5859 8857 5868 8891
rect 5816 8848 5868 8857
rect 5908 8891 5960 8900
rect 5908 8857 5917 8891
rect 5917 8857 5951 8891
rect 5951 8857 5960 8891
rect 5908 8848 5960 8857
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 6920 8984 6972 9036
rect 6644 8959 6696 8968
rect 6644 8925 6653 8959
rect 6653 8925 6687 8959
rect 6687 8925 6696 8959
rect 6644 8916 6696 8925
rect 9772 8984 9824 9036
rect 10968 8984 11020 9036
rect 5448 8780 5500 8832
rect 6092 8780 6144 8832
rect 6644 8780 6696 8832
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 9496 8916 9548 8968
rect 9956 8916 10008 8968
rect 11336 8959 11388 8968
rect 11336 8925 11345 8959
rect 11345 8925 11379 8959
rect 11379 8925 11388 8959
rect 11336 8916 11388 8925
rect 11612 9027 11664 9036
rect 11612 8993 11621 9027
rect 11621 8993 11655 9027
rect 11655 8993 11664 9027
rect 11612 8984 11664 8993
rect 12256 8984 12308 9036
rect 12440 9052 12492 9104
rect 13728 9120 13780 9172
rect 14556 9163 14608 9172
rect 14556 9129 14565 9163
rect 14565 9129 14599 9163
rect 14599 9129 14608 9163
rect 14556 9120 14608 9129
rect 15936 9120 15988 9172
rect 16396 9120 16448 9172
rect 16856 9120 16908 9172
rect 17040 9120 17092 9172
rect 15108 9052 15160 9104
rect 18420 9120 18472 9172
rect 18604 9163 18656 9172
rect 18604 9129 18613 9163
rect 18613 9129 18647 9163
rect 18647 9129 18656 9163
rect 18604 9120 18656 9129
rect 18696 9120 18748 9172
rect 18144 9052 18196 9104
rect 21916 9163 21968 9172
rect 21916 9129 21925 9163
rect 21925 9129 21959 9163
rect 21959 9129 21968 9163
rect 21916 9120 21968 9129
rect 22008 9120 22060 9172
rect 22376 9120 22428 9172
rect 12532 8959 12584 8968
rect 12532 8925 12541 8959
rect 12541 8925 12575 8959
rect 12575 8925 12584 8959
rect 12532 8916 12584 8925
rect 12900 8916 12952 8968
rect 13360 8916 13412 8968
rect 14096 8959 14148 8968
rect 14096 8925 14105 8959
rect 14105 8925 14139 8959
rect 14139 8925 14148 8959
rect 14096 8916 14148 8925
rect 14372 8959 14424 8968
rect 14372 8925 14381 8959
rect 14381 8925 14415 8959
rect 14415 8925 14424 8959
rect 14372 8916 14424 8925
rect 8208 8848 8260 8900
rect 9036 8848 9088 8900
rect 9404 8891 9456 8900
rect 9404 8857 9413 8891
rect 9413 8857 9447 8891
rect 9447 8857 9456 8891
rect 9404 8848 9456 8857
rect 9680 8848 9732 8900
rect 10968 8848 11020 8900
rect 11428 8848 11480 8900
rect 7012 8780 7064 8832
rect 7656 8780 7708 8832
rect 7748 8823 7800 8832
rect 7748 8789 7757 8823
rect 7757 8789 7791 8823
rect 7791 8789 7800 8823
rect 7748 8780 7800 8789
rect 7840 8823 7892 8832
rect 7840 8789 7849 8823
rect 7849 8789 7883 8823
rect 7883 8789 7892 8823
rect 7840 8780 7892 8789
rect 9864 8780 9916 8832
rect 11152 8780 11204 8832
rect 12348 8848 12400 8900
rect 16672 8916 16724 8968
rect 16856 8916 16908 8968
rect 18512 9027 18564 9036
rect 18512 8993 18521 9027
rect 18521 8993 18555 9027
rect 18555 8993 18564 9027
rect 18512 8984 18564 8993
rect 12900 8780 12952 8832
rect 13176 8780 13228 8832
rect 17224 8848 17276 8900
rect 14832 8780 14884 8832
rect 16396 8780 16448 8832
rect 16856 8780 16908 8832
rect 17776 8891 17828 8900
rect 17776 8857 17785 8891
rect 17785 8857 17819 8891
rect 17819 8857 17828 8891
rect 17776 8848 17828 8857
rect 23388 8984 23440 9036
rect 25688 9120 25740 9172
rect 26056 9120 26108 9172
rect 25872 9052 25924 9104
rect 26608 9163 26660 9172
rect 26608 9129 26617 9163
rect 26617 9129 26651 9163
rect 26651 9129 26660 9163
rect 26608 9120 26660 9129
rect 26148 8984 26200 9036
rect 26516 9052 26568 9104
rect 27620 9120 27672 9172
rect 27252 9052 27304 9104
rect 28172 9120 28224 9172
rect 29276 9163 29328 9172
rect 29276 9129 29285 9163
rect 29285 9129 29319 9163
rect 29319 9129 29328 9163
rect 29276 9120 29328 9129
rect 32496 9163 32548 9172
rect 32496 9129 32505 9163
rect 32505 9129 32539 9163
rect 32539 9129 32548 9163
rect 32496 9120 32548 9129
rect 22008 8916 22060 8968
rect 22284 8916 22336 8968
rect 22560 8916 22612 8968
rect 25596 8916 25648 8968
rect 25688 8959 25740 8968
rect 25688 8925 25697 8959
rect 25697 8925 25731 8959
rect 25731 8925 25740 8959
rect 25688 8916 25740 8925
rect 25780 8959 25832 8968
rect 25780 8925 25789 8959
rect 25789 8925 25823 8959
rect 25823 8925 25832 8959
rect 25780 8916 25832 8925
rect 26792 8984 26844 9036
rect 26608 8916 26660 8968
rect 27528 8984 27580 9036
rect 27804 8984 27856 9036
rect 28816 8984 28868 9036
rect 18236 8780 18288 8832
rect 24584 8848 24636 8900
rect 24952 8780 25004 8832
rect 26148 8891 26200 8900
rect 26148 8857 26157 8891
rect 26157 8857 26191 8891
rect 26191 8857 26200 8891
rect 26148 8848 26200 8857
rect 27344 8848 27396 8900
rect 28356 8959 28408 8968
rect 28356 8925 28365 8959
rect 28365 8925 28399 8959
rect 28399 8925 28408 8959
rect 28356 8916 28408 8925
rect 29092 8959 29144 8968
rect 29092 8925 29101 8959
rect 29101 8925 29135 8959
rect 29135 8925 29144 8959
rect 29092 8916 29144 8925
rect 31116 8959 31168 8968
rect 31116 8925 31125 8959
rect 31125 8925 31159 8959
rect 31159 8925 31168 8959
rect 31116 8916 31168 8925
rect 30748 8848 30800 8900
rect 27160 8823 27212 8832
rect 27160 8789 27169 8823
rect 27169 8789 27203 8823
rect 27203 8789 27212 8823
rect 27160 8780 27212 8789
rect 27528 8780 27580 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 4436 8576 4488 8628
rect 4804 8576 4856 8628
rect 5908 8576 5960 8628
rect 6276 8576 6328 8628
rect 6828 8576 6880 8628
rect 7472 8576 7524 8628
rect 4160 8508 4212 8560
rect 3148 8440 3200 8492
rect 4620 8440 4672 8492
rect 5264 8483 5316 8492
rect 5264 8449 5273 8483
rect 5273 8449 5307 8483
rect 5307 8449 5316 8483
rect 5264 8440 5316 8449
rect 4988 8372 5040 8424
rect 5448 8551 5500 8560
rect 5448 8517 5457 8551
rect 5457 8517 5491 8551
rect 5491 8517 5500 8551
rect 5448 8508 5500 8517
rect 7380 8551 7432 8560
rect 7380 8517 7389 8551
rect 7389 8517 7423 8551
rect 7423 8517 7432 8551
rect 7380 8508 7432 8517
rect 8760 8576 8812 8628
rect 9220 8576 9272 8628
rect 5540 8483 5592 8492
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 5724 8440 5776 8492
rect 6000 8440 6052 8492
rect 4344 8304 4396 8356
rect 4712 8304 4764 8356
rect 7840 8440 7892 8492
rect 8208 8440 8260 8492
rect 7656 8372 7708 8424
rect 8852 8483 8904 8492
rect 8852 8449 8861 8483
rect 8861 8449 8895 8483
rect 8895 8449 8904 8483
rect 8852 8440 8904 8449
rect 9036 8440 9088 8492
rect 9312 8508 9364 8560
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 9680 8551 9732 8560
rect 9680 8517 9689 8551
rect 9689 8517 9723 8551
rect 9723 8517 9732 8551
rect 9680 8508 9732 8517
rect 11336 8619 11388 8628
rect 11336 8585 11345 8619
rect 11345 8585 11379 8619
rect 11379 8585 11388 8619
rect 11336 8576 11388 8585
rect 11704 8576 11756 8628
rect 11888 8619 11940 8628
rect 11888 8585 11897 8619
rect 11897 8585 11931 8619
rect 11931 8585 11940 8619
rect 11888 8576 11940 8585
rect 13728 8576 13780 8628
rect 14372 8576 14424 8628
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10324 8483 10376 8492
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 10324 8440 10376 8449
rect 10968 8551 11020 8560
rect 10968 8517 10977 8551
rect 10977 8517 11011 8551
rect 11011 8517 11020 8551
rect 10968 8508 11020 8517
rect 11060 8551 11112 8560
rect 11060 8517 11069 8551
rect 11069 8517 11103 8551
rect 11103 8517 11112 8551
rect 11060 8508 11112 8517
rect 16948 8576 17000 8628
rect 11152 8483 11204 8492
rect 11152 8449 11161 8483
rect 11161 8449 11195 8483
rect 11195 8449 11204 8483
rect 11152 8440 11204 8449
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 12256 8483 12308 8492
rect 12256 8449 12265 8483
rect 12265 8449 12299 8483
rect 12299 8449 12308 8483
rect 12256 8440 12308 8449
rect 12532 8440 12584 8492
rect 12900 8440 12952 8492
rect 12992 8440 13044 8492
rect 13176 8440 13228 8492
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 8392 8372 8444 8424
rect 8024 8304 8076 8356
rect 8852 8304 8904 8356
rect 9588 8372 9640 8424
rect 9956 8372 10008 8424
rect 9404 8304 9456 8356
rect 10876 8372 10928 8424
rect 13268 8372 13320 8424
rect 10508 8304 10560 8356
rect 11428 8304 11480 8356
rect 12348 8304 12400 8356
rect 12624 8304 12676 8356
rect 5816 8279 5868 8288
rect 5816 8245 5825 8279
rect 5825 8245 5859 8279
rect 5859 8245 5868 8279
rect 5816 8236 5868 8245
rect 5908 8236 5960 8288
rect 8116 8236 8168 8288
rect 8484 8279 8536 8288
rect 8484 8245 8493 8279
rect 8493 8245 8527 8279
rect 8527 8245 8536 8279
rect 8484 8236 8536 8245
rect 10876 8236 10928 8288
rect 11520 8279 11572 8288
rect 11520 8245 11529 8279
rect 11529 8245 11563 8279
rect 11563 8245 11572 8279
rect 11520 8236 11572 8245
rect 12164 8279 12216 8288
rect 12164 8245 12173 8279
rect 12173 8245 12207 8279
rect 12207 8245 12216 8279
rect 12164 8236 12216 8245
rect 12256 8236 12308 8288
rect 17408 8576 17460 8628
rect 19800 8576 19852 8628
rect 19892 8576 19944 8628
rect 13912 8440 13964 8492
rect 14096 8440 14148 8492
rect 15108 8483 15160 8492
rect 15108 8449 15117 8483
rect 15117 8449 15151 8483
rect 15151 8449 15160 8483
rect 15108 8440 15160 8449
rect 15200 8483 15252 8492
rect 15200 8449 15209 8483
rect 15209 8449 15243 8483
rect 15243 8449 15252 8483
rect 15200 8440 15252 8449
rect 15568 8440 15620 8492
rect 15752 8483 15804 8492
rect 15752 8449 15761 8483
rect 15761 8449 15795 8483
rect 15795 8449 15804 8483
rect 15752 8440 15804 8449
rect 15844 8440 15896 8492
rect 16672 8483 16724 8492
rect 16672 8449 16681 8483
rect 16681 8449 16715 8483
rect 16715 8449 16724 8483
rect 16672 8440 16724 8449
rect 19432 8508 19484 8560
rect 17132 8440 17184 8492
rect 17684 8483 17736 8492
rect 17684 8449 17693 8483
rect 17693 8449 17727 8483
rect 17727 8449 17736 8483
rect 17684 8440 17736 8449
rect 13728 8415 13780 8424
rect 13728 8381 13737 8415
rect 13737 8381 13771 8415
rect 13771 8381 13780 8415
rect 13728 8372 13780 8381
rect 15384 8347 15436 8356
rect 15384 8313 15393 8347
rect 15393 8313 15427 8347
rect 15427 8313 15436 8347
rect 15384 8304 15436 8313
rect 16580 8372 16632 8424
rect 19800 8440 19852 8492
rect 20904 8508 20956 8560
rect 23480 8551 23532 8560
rect 23480 8517 23489 8551
rect 23489 8517 23523 8551
rect 23523 8517 23532 8551
rect 23480 8508 23532 8517
rect 23572 8508 23624 8560
rect 24676 8619 24728 8628
rect 24676 8585 24685 8619
rect 24685 8585 24719 8619
rect 24719 8585 24728 8619
rect 24676 8576 24728 8585
rect 24768 8576 24820 8628
rect 29552 8576 29604 8628
rect 20996 8440 21048 8492
rect 27620 8508 27672 8560
rect 23940 8483 23992 8492
rect 23940 8449 23949 8483
rect 23949 8449 23983 8483
rect 23983 8449 23992 8483
rect 23940 8440 23992 8449
rect 20168 8372 20220 8424
rect 20904 8372 20956 8424
rect 24768 8440 24820 8492
rect 30012 8440 30064 8492
rect 30564 8508 30616 8560
rect 31852 8508 31904 8560
rect 32220 8483 32272 8492
rect 32220 8449 32229 8483
rect 32229 8449 32263 8483
rect 32263 8449 32272 8483
rect 32220 8440 32272 8449
rect 30104 8347 30156 8356
rect 30104 8313 30113 8347
rect 30113 8313 30147 8347
rect 30147 8313 30156 8347
rect 30104 8304 30156 8313
rect 32404 8347 32456 8356
rect 32404 8313 32413 8347
rect 32413 8313 32447 8347
rect 32447 8313 32456 8347
rect 32404 8304 32456 8313
rect 14924 8279 14976 8288
rect 14924 8245 14933 8279
rect 14933 8245 14967 8279
rect 14967 8245 14976 8279
rect 14924 8236 14976 8245
rect 15108 8236 15160 8288
rect 15292 8236 15344 8288
rect 15568 8236 15620 8288
rect 15936 8279 15988 8288
rect 15936 8245 15945 8279
rect 15945 8245 15979 8279
rect 15979 8245 15988 8279
rect 15936 8236 15988 8245
rect 16028 8236 16080 8288
rect 17500 8279 17552 8288
rect 17500 8245 17509 8279
rect 17509 8245 17543 8279
rect 17543 8245 17552 8279
rect 17500 8236 17552 8245
rect 19892 8236 19944 8288
rect 21824 8236 21876 8288
rect 22652 8236 22704 8288
rect 23756 8279 23808 8288
rect 23756 8245 23765 8279
rect 23765 8245 23799 8279
rect 23799 8245 23808 8279
rect 23756 8236 23808 8245
rect 24032 8236 24084 8288
rect 24308 8236 24360 8288
rect 27344 8236 27396 8288
rect 29920 8279 29972 8288
rect 29920 8245 29929 8279
rect 29929 8245 29963 8279
rect 29963 8245 29972 8279
rect 29920 8236 29972 8245
rect 31208 8279 31260 8288
rect 31208 8245 31217 8279
rect 31217 8245 31251 8279
rect 31251 8245 31260 8279
rect 31208 8236 31260 8245
rect 31300 8236 31352 8288
rect 31760 8236 31812 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 4804 8032 4856 8084
rect 7932 8032 7984 8084
rect 8852 8032 8904 8084
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 9036 8032 9088 8084
rect 10876 8032 10928 8084
rect 11520 8032 11572 8084
rect 11704 8075 11756 8084
rect 11704 8041 11713 8075
rect 11713 8041 11747 8075
rect 11747 8041 11756 8075
rect 11704 8032 11756 8041
rect 5264 7964 5316 8016
rect 5908 7964 5960 8016
rect 6000 7964 6052 8016
rect 7840 7964 7892 8016
rect 9312 7964 9364 8016
rect 10784 7964 10836 8016
rect 12256 7964 12308 8016
rect 12624 8032 12676 8084
rect 13636 8032 13688 8084
rect 14464 7964 14516 8016
rect 15844 8032 15896 8084
rect 16672 8075 16724 8084
rect 16672 8041 16681 8075
rect 16681 8041 16715 8075
rect 16715 8041 16724 8075
rect 16672 8032 16724 8041
rect 5632 7896 5684 7948
rect 6276 7828 6328 7880
rect 8116 7896 8168 7948
rect 6736 7828 6788 7880
rect 7104 7828 7156 7880
rect 8484 7828 8536 7880
rect 8944 7828 8996 7880
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 9588 7828 9640 7880
rect 6368 7803 6420 7812
rect 6368 7769 6377 7803
rect 6377 7769 6411 7803
rect 6411 7769 6420 7803
rect 6368 7760 6420 7769
rect 6920 7760 6972 7812
rect 10416 7828 10468 7880
rect 11612 7896 11664 7948
rect 13360 7896 13412 7948
rect 13636 7896 13688 7948
rect 14556 7939 14608 7948
rect 14556 7905 14565 7939
rect 14565 7905 14599 7939
rect 14599 7905 14608 7939
rect 14556 7896 14608 7905
rect 15752 7896 15804 7948
rect 16948 7964 17000 8016
rect 17132 8075 17184 8084
rect 17132 8041 17141 8075
rect 17141 8041 17175 8075
rect 17175 8041 17184 8075
rect 17132 8032 17184 8041
rect 17868 8032 17920 8084
rect 19984 8032 20036 8084
rect 20168 8032 20220 8084
rect 20996 8032 21048 8084
rect 21732 8075 21784 8084
rect 21732 8041 21741 8075
rect 21741 8041 21775 8075
rect 21775 8041 21784 8075
rect 21732 8032 21784 8041
rect 22836 8075 22888 8084
rect 22836 8041 22845 8075
rect 22845 8041 22879 8075
rect 22879 8041 22888 8075
rect 22836 8032 22888 8041
rect 25780 8075 25832 8084
rect 25780 8041 25789 8075
rect 25789 8041 25823 8075
rect 25823 8041 25832 8075
rect 25780 8032 25832 8041
rect 11796 7828 11848 7880
rect 12624 7828 12676 7880
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 14372 7828 14424 7880
rect 16212 7871 16264 7880
rect 16212 7837 16221 7871
rect 16221 7837 16255 7871
rect 16255 7837 16264 7871
rect 16212 7828 16264 7837
rect 9956 7760 10008 7812
rect 5540 7692 5592 7744
rect 6644 7692 6696 7744
rect 10968 7692 11020 7744
rect 13820 7692 13872 7744
rect 14096 7760 14148 7812
rect 14556 7760 14608 7812
rect 16304 7760 16356 7812
rect 15844 7692 15896 7744
rect 16396 7735 16448 7744
rect 16396 7701 16405 7735
rect 16405 7701 16439 7735
rect 16439 7701 16448 7735
rect 16396 7692 16448 7701
rect 17132 7896 17184 7948
rect 17960 7896 18012 7948
rect 19984 7896 20036 7948
rect 21640 7896 21692 7948
rect 17040 7828 17092 7880
rect 17224 7871 17276 7880
rect 17224 7837 17233 7871
rect 17233 7837 17267 7871
rect 17267 7837 17276 7871
rect 17224 7828 17276 7837
rect 17592 7760 17644 7812
rect 18512 7760 18564 7812
rect 19340 7760 19392 7812
rect 20168 7828 20220 7880
rect 20628 7828 20680 7880
rect 22560 7964 22612 8016
rect 31300 8032 31352 8084
rect 32220 8032 32272 8084
rect 21824 7939 21876 7948
rect 21824 7905 21833 7939
rect 21833 7905 21867 7939
rect 21867 7905 21876 7939
rect 21824 7896 21876 7905
rect 21824 7760 21876 7812
rect 21916 7692 21968 7744
rect 22744 7871 22796 7880
rect 22744 7837 22753 7871
rect 22753 7837 22787 7871
rect 22787 7837 22796 7871
rect 22744 7828 22796 7837
rect 25504 7896 25556 7948
rect 27160 7896 27212 7948
rect 26884 7828 26936 7880
rect 28816 7871 28868 7880
rect 28816 7837 28825 7871
rect 28825 7837 28859 7871
rect 28859 7837 28868 7871
rect 28816 7828 28868 7837
rect 29184 7871 29236 7880
rect 29184 7837 29193 7871
rect 29193 7837 29227 7871
rect 29227 7837 29236 7871
rect 29184 7828 29236 7837
rect 22928 7760 22980 7812
rect 29000 7803 29052 7812
rect 29000 7769 29009 7803
rect 29009 7769 29043 7803
rect 29043 7769 29052 7803
rect 29000 7760 29052 7769
rect 29552 7871 29604 7880
rect 29552 7837 29561 7871
rect 29561 7837 29595 7871
rect 29595 7837 29604 7871
rect 31116 7871 31168 7880
rect 29552 7828 29604 7837
rect 31116 7837 31125 7871
rect 31125 7837 31159 7871
rect 31159 7837 31168 7871
rect 31116 7828 31168 7837
rect 31208 7828 31260 7880
rect 23112 7692 23164 7744
rect 26056 7692 26108 7744
rect 30472 7692 30524 7744
rect 30748 7692 30800 7744
rect 30932 7735 30984 7744
rect 30932 7701 30941 7735
rect 30941 7701 30975 7735
rect 30975 7701 30984 7735
rect 30932 7692 30984 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 6368 7488 6420 7540
rect 6920 7531 6972 7540
rect 6920 7497 6929 7531
rect 6929 7497 6963 7531
rect 6963 7497 6972 7531
rect 6920 7488 6972 7497
rect 3976 7420 4028 7472
rect 4160 7463 4212 7472
rect 4160 7429 4169 7463
rect 4169 7429 4203 7463
rect 4203 7429 4212 7463
rect 4160 7420 4212 7429
rect 4252 7395 4304 7404
rect 4252 7361 4261 7395
rect 4261 7361 4295 7395
rect 4295 7361 4304 7395
rect 4252 7352 4304 7361
rect 6644 7463 6696 7472
rect 6644 7429 6653 7463
rect 6653 7429 6687 7463
rect 6687 7429 6696 7463
rect 6644 7420 6696 7429
rect 4712 7395 4764 7404
rect 4712 7361 4721 7395
rect 4721 7361 4755 7395
rect 4755 7361 4764 7395
rect 4712 7352 4764 7361
rect 4804 7395 4856 7404
rect 4804 7361 4813 7395
rect 4813 7361 4847 7395
rect 4847 7361 4856 7395
rect 4804 7352 4856 7361
rect 4988 7352 5040 7404
rect 5540 7352 5592 7404
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 6368 7395 6420 7404
rect 6368 7361 6377 7395
rect 6377 7361 6411 7395
rect 6411 7361 6420 7395
rect 6368 7352 6420 7361
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 7472 7463 7524 7472
rect 7472 7429 7481 7463
rect 7481 7429 7515 7463
rect 7515 7429 7524 7463
rect 7472 7420 7524 7429
rect 12992 7488 13044 7540
rect 13268 7488 13320 7540
rect 14372 7488 14424 7540
rect 16212 7488 16264 7540
rect 18788 7488 18840 7540
rect 5080 7259 5132 7268
rect 5080 7225 5089 7259
rect 5089 7225 5123 7259
rect 5123 7225 5132 7259
rect 5080 7216 5132 7225
rect 5908 7216 5960 7268
rect 6368 7216 6420 7268
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 7840 7352 7892 7404
rect 8116 7395 8168 7404
rect 8116 7361 8125 7395
rect 8125 7361 8159 7395
rect 8159 7361 8168 7395
rect 8116 7352 8168 7361
rect 8208 7395 8260 7404
rect 8208 7361 8217 7395
rect 8217 7361 8251 7395
rect 8251 7361 8260 7395
rect 8208 7352 8260 7361
rect 8484 7352 8536 7404
rect 8576 7395 8628 7404
rect 8576 7361 8585 7395
rect 8585 7361 8619 7395
rect 8619 7361 8628 7395
rect 8576 7352 8628 7361
rect 8852 7395 8904 7404
rect 8852 7361 8861 7395
rect 8861 7361 8895 7395
rect 8895 7361 8904 7395
rect 8852 7352 8904 7361
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 9036 7352 9088 7404
rect 9496 7395 9548 7404
rect 9496 7361 9505 7395
rect 9505 7361 9539 7395
rect 9539 7361 9548 7395
rect 9496 7352 9548 7361
rect 10508 7420 10560 7472
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 12532 7395 12584 7404
rect 12532 7361 12541 7395
rect 12541 7361 12575 7395
rect 12575 7361 12584 7395
rect 12532 7352 12584 7361
rect 13084 7352 13136 7404
rect 13360 7463 13412 7472
rect 13360 7429 13369 7463
rect 13369 7429 13403 7463
rect 13403 7429 13412 7463
rect 13360 7420 13412 7429
rect 14464 7420 14516 7472
rect 15476 7420 15528 7472
rect 17592 7420 17644 7472
rect 19340 7463 19392 7472
rect 19340 7429 19349 7463
rect 19349 7429 19383 7463
rect 19383 7429 19392 7463
rect 19340 7420 19392 7429
rect 23388 7488 23440 7540
rect 13544 7352 13596 7404
rect 13820 7352 13872 7404
rect 8944 7216 8996 7268
rect 9956 7284 10008 7336
rect 12624 7327 12676 7336
rect 12624 7293 12633 7327
rect 12633 7293 12667 7327
rect 12667 7293 12676 7327
rect 12624 7284 12676 7293
rect 9864 7216 9916 7268
rect 5540 7148 5592 7200
rect 6092 7148 6144 7200
rect 6828 7148 6880 7200
rect 7012 7148 7064 7200
rect 9036 7148 9088 7200
rect 10508 7148 10560 7200
rect 10692 7148 10744 7200
rect 10876 7148 10928 7200
rect 12624 7148 12676 7200
rect 13176 7216 13228 7268
rect 12992 7191 13044 7200
rect 12992 7157 13001 7191
rect 13001 7157 13035 7191
rect 13035 7157 13044 7191
rect 12992 7148 13044 7157
rect 13452 7284 13504 7336
rect 16580 7352 16632 7404
rect 23664 7352 23716 7404
rect 27620 7488 27672 7540
rect 29184 7488 29236 7540
rect 27896 7420 27948 7472
rect 28172 7420 28224 7472
rect 16396 7284 16448 7336
rect 20168 7284 20220 7336
rect 13912 7216 13964 7268
rect 14280 7216 14332 7268
rect 23848 7284 23900 7336
rect 24216 7284 24268 7336
rect 25964 7395 26016 7404
rect 25964 7361 25973 7395
rect 25973 7361 26007 7395
rect 26007 7361 26016 7395
rect 25964 7352 26016 7361
rect 32496 7352 32548 7404
rect 30932 7284 30984 7336
rect 32220 7284 32272 7336
rect 19248 7148 19300 7200
rect 22376 7148 22428 7200
rect 24124 7191 24176 7200
rect 24124 7157 24133 7191
rect 24133 7157 24167 7191
rect 24167 7157 24176 7191
rect 24124 7148 24176 7157
rect 26056 7191 26108 7200
rect 26056 7157 26065 7191
rect 26065 7157 26099 7191
rect 26099 7157 26108 7191
rect 26056 7148 26108 7157
rect 27804 7191 27856 7200
rect 27804 7157 27813 7191
rect 27813 7157 27847 7191
rect 27847 7157 27856 7191
rect 27804 7148 27856 7157
rect 30840 7148 30892 7200
rect 32312 7191 32364 7200
rect 32312 7157 32321 7191
rect 32321 7157 32355 7191
rect 32355 7157 32364 7191
rect 32312 7148 32364 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 4712 6987 4764 6996
rect 4712 6953 4721 6987
rect 4721 6953 4755 6987
rect 4755 6953 4764 6987
rect 4712 6944 4764 6953
rect 5080 6944 5132 6996
rect 3976 6876 4028 6928
rect 5448 6876 5500 6928
rect 7012 6876 7064 6928
rect 7656 6944 7708 6996
rect 7932 6944 7984 6996
rect 9496 6944 9548 6996
rect 9864 6944 9916 6996
rect 10692 6944 10744 6996
rect 11244 6944 11296 6996
rect 11428 6944 11480 6996
rect 13084 6944 13136 6996
rect 13636 6987 13688 6996
rect 13636 6953 13645 6987
rect 13645 6953 13679 6987
rect 13679 6953 13688 6987
rect 13636 6944 13688 6953
rect 11520 6876 11572 6928
rect 9588 6808 9640 6860
rect 7748 6740 7800 6792
rect 9312 6783 9364 6792
rect 9312 6749 9321 6783
rect 9321 6749 9355 6783
rect 9355 6749 9364 6783
rect 9312 6740 9364 6749
rect 9404 6783 9456 6792
rect 9404 6749 9413 6783
rect 9413 6749 9447 6783
rect 9447 6749 9456 6783
rect 9404 6740 9456 6749
rect 10600 6740 10652 6792
rect 10784 6740 10836 6792
rect 10968 6672 11020 6724
rect 11244 6740 11296 6792
rect 11520 6740 11572 6792
rect 11704 6851 11756 6860
rect 11704 6817 11713 6851
rect 11713 6817 11747 6851
rect 11747 6817 11756 6851
rect 13452 6876 13504 6928
rect 14832 6944 14884 6996
rect 11704 6808 11756 6817
rect 13360 6808 13412 6860
rect 15476 6944 15528 6996
rect 18512 6987 18564 6996
rect 18512 6953 18521 6987
rect 18521 6953 18555 6987
rect 18555 6953 18564 6987
rect 18512 6944 18564 6953
rect 20628 6944 20680 6996
rect 23204 6944 23256 6996
rect 9496 6604 9548 6656
rect 10876 6604 10928 6656
rect 11520 6604 11572 6656
rect 12992 6740 13044 6792
rect 11888 6672 11940 6724
rect 16580 6808 16632 6860
rect 18880 6876 18932 6928
rect 19248 6876 19300 6928
rect 32496 6987 32548 6996
rect 32496 6953 32505 6987
rect 32505 6953 32539 6987
rect 32539 6953 32548 6987
rect 32496 6944 32548 6953
rect 13912 6740 13964 6792
rect 15108 6740 15160 6792
rect 15200 6783 15252 6792
rect 15200 6749 15209 6783
rect 15209 6749 15243 6783
rect 15243 6749 15252 6783
rect 15200 6740 15252 6749
rect 16212 6783 16264 6792
rect 16212 6749 16221 6783
rect 16221 6749 16255 6783
rect 16255 6749 16264 6783
rect 16212 6740 16264 6749
rect 17776 6783 17828 6792
rect 17776 6749 17785 6783
rect 17785 6749 17819 6783
rect 17819 6749 17828 6783
rect 17776 6740 17828 6749
rect 17960 6740 18012 6792
rect 14464 6672 14516 6724
rect 12348 6604 12400 6656
rect 15476 6672 15528 6724
rect 15844 6672 15896 6724
rect 16028 6715 16080 6724
rect 16028 6681 16037 6715
rect 16037 6681 16071 6715
rect 16071 6681 16080 6715
rect 16028 6672 16080 6681
rect 17592 6715 17644 6724
rect 17592 6681 17601 6715
rect 17601 6681 17635 6715
rect 17635 6681 17644 6715
rect 17592 6672 17644 6681
rect 18696 6672 18748 6724
rect 15660 6647 15712 6656
rect 15660 6613 15669 6647
rect 15669 6613 15703 6647
rect 15703 6613 15712 6647
rect 15660 6604 15712 6613
rect 17684 6604 17736 6656
rect 18052 6647 18104 6656
rect 18052 6613 18061 6647
rect 18061 6613 18095 6647
rect 18095 6613 18104 6647
rect 18052 6604 18104 6613
rect 18420 6604 18472 6656
rect 19984 6740 20036 6792
rect 20076 6783 20128 6792
rect 20076 6749 20085 6783
rect 20085 6749 20119 6783
rect 20119 6749 20128 6783
rect 20076 6740 20128 6749
rect 20260 6851 20312 6860
rect 20260 6817 20269 6851
rect 20269 6817 20303 6851
rect 20303 6817 20312 6851
rect 20260 6808 20312 6817
rect 21640 6808 21692 6860
rect 22100 6808 22152 6860
rect 22376 6740 22428 6792
rect 22468 6783 22520 6792
rect 22468 6749 22477 6783
rect 22477 6749 22511 6783
rect 22511 6749 22520 6783
rect 22468 6740 22520 6749
rect 22560 6783 22612 6792
rect 22560 6749 22569 6783
rect 22569 6749 22603 6783
rect 22603 6749 22612 6783
rect 22560 6740 22612 6749
rect 24768 6851 24820 6860
rect 24768 6817 24777 6851
rect 24777 6817 24811 6851
rect 24811 6817 24820 6851
rect 24768 6808 24820 6817
rect 26148 6808 26200 6860
rect 29552 6808 29604 6860
rect 25320 6740 25372 6792
rect 26516 6783 26568 6792
rect 26516 6749 26525 6783
rect 26525 6749 26559 6783
rect 26559 6749 26568 6783
rect 26516 6740 26568 6749
rect 30104 6740 30156 6792
rect 30748 6783 30800 6792
rect 30748 6749 30757 6783
rect 30757 6749 30791 6783
rect 30791 6749 30800 6783
rect 30748 6740 30800 6749
rect 30840 6783 30892 6792
rect 30840 6749 30849 6783
rect 30849 6749 30883 6783
rect 30883 6749 30892 6783
rect 30840 6740 30892 6749
rect 18880 6672 18932 6724
rect 24584 6715 24636 6724
rect 24584 6681 24593 6715
rect 24593 6681 24627 6715
rect 24627 6681 24636 6715
rect 24584 6672 24636 6681
rect 29000 6672 29052 6724
rect 18972 6647 19024 6656
rect 18972 6613 18981 6647
rect 18981 6613 19015 6647
rect 19015 6613 19024 6647
rect 18972 6604 19024 6613
rect 20536 6647 20588 6656
rect 20536 6613 20545 6647
rect 20545 6613 20579 6647
rect 20579 6613 20588 6647
rect 20536 6604 20588 6613
rect 20628 6604 20680 6656
rect 22652 6604 22704 6656
rect 23572 6604 23624 6656
rect 27896 6604 27948 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 10140 6400 10192 6452
rect 14096 6400 14148 6452
rect 14188 6400 14240 6452
rect 14924 6400 14976 6452
rect 15752 6443 15804 6452
rect 15752 6409 15761 6443
rect 15761 6409 15795 6443
rect 15795 6409 15804 6443
rect 15752 6400 15804 6409
rect 18604 6443 18656 6452
rect 18604 6409 18613 6443
rect 18613 6409 18647 6443
rect 18647 6409 18656 6443
rect 18604 6400 18656 6409
rect 2596 6196 2648 6248
rect 10692 6264 10744 6316
rect 11520 6307 11572 6316
rect 11520 6273 11529 6307
rect 11529 6273 11563 6307
rect 11563 6273 11572 6307
rect 11520 6264 11572 6273
rect 13912 6264 13964 6316
rect 15108 6264 15160 6316
rect 15660 6264 15712 6316
rect 17132 6264 17184 6316
rect 17316 6307 17368 6316
rect 17316 6273 17325 6307
rect 17325 6273 17359 6307
rect 17359 6273 17368 6307
rect 17316 6264 17368 6273
rect 11428 6196 11480 6248
rect 15476 6196 15528 6248
rect 17224 6239 17276 6248
rect 17224 6205 17233 6239
rect 17233 6205 17267 6239
rect 17267 6205 17276 6239
rect 17224 6196 17276 6205
rect 10600 6128 10652 6180
rect 11244 6128 11296 6180
rect 17776 6264 17828 6316
rect 19708 6332 19760 6384
rect 19984 6332 20036 6384
rect 17684 6196 17736 6248
rect 18788 6196 18840 6248
rect 19248 6307 19300 6316
rect 19248 6273 19257 6307
rect 19257 6273 19291 6307
rect 19291 6273 19300 6307
rect 19248 6264 19300 6273
rect 19616 6264 19668 6316
rect 20720 6332 20772 6384
rect 21180 6332 21232 6384
rect 22560 6400 22612 6452
rect 23020 6400 23072 6452
rect 19524 6196 19576 6248
rect 20536 6264 20588 6316
rect 22376 6307 22428 6316
rect 22376 6273 22385 6307
rect 22385 6273 22419 6307
rect 22419 6273 22428 6307
rect 22376 6264 22428 6273
rect 22652 6332 22704 6384
rect 20628 6128 20680 6180
rect 11336 6060 11388 6112
rect 11704 6103 11756 6112
rect 11704 6069 11713 6103
rect 11713 6069 11747 6103
rect 11747 6069 11756 6103
rect 11704 6060 11756 6069
rect 11980 6060 12032 6112
rect 14004 6060 14056 6112
rect 15476 6060 15528 6112
rect 17500 6103 17552 6112
rect 17500 6069 17509 6103
rect 17509 6069 17543 6103
rect 17543 6069 17552 6103
rect 17500 6060 17552 6069
rect 17776 6103 17828 6112
rect 17776 6069 17785 6103
rect 17785 6069 17819 6103
rect 17819 6069 17828 6103
rect 17776 6060 17828 6069
rect 17868 6060 17920 6112
rect 18972 6103 19024 6112
rect 18972 6069 18981 6103
rect 18981 6069 19015 6103
rect 19015 6069 19024 6103
rect 18972 6060 19024 6069
rect 20076 6103 20128 6112
rect 20076 6069 20085 6103
rect 20085 6069 20119 6103
rect 20119 6069 20128 6103
rect 20076 6060 20128 6069
rect 20352 6103 20404 6112
rect 20352 6069 20361 6103
rect 20361 6069 20395 6103
rect 20395 6069 20404 6103
rect 20352 6060 20404 6069
rect 22100 6103 22152 6112
rect 22100 6069 22109 6103
rect 22109 6069 22143 6103
rect 22143 6069 22152 6103
rect 22100 6060 22152 6069
rect 23020 6196 23072 6248
rect 23204 6307 23256 6316
rect 23204 6273 23213 6307
rect 23213 6273 23247 6307
rect 23247 6273 23256 6307
rect 23204 6264 23256 6273
rect 26424 6400 26476 6452
rect 26976 6400 27028 6452
rect 31668 6400 31720 6452
rect 25044 6307 25096 6316
rect 25044 6273 25053 6307
rect 25053 6273 25087 6307
rect 25087 6273 25096 6307
rect 25044 6264 25096 6273
rect 25228 6264 25280 6316
rect 25780 6264 25832 6316
rect 25964 6307 26016 6316
rect 25964 6273 25973 6307
rect 25973 6273 26007 6307
rect 26007 6273 26016 6307
rect 25964 6264 26016 6273
rect 25504 6196 25556 6248
rect 26516 6264 26568 6316
rect 32220 6307 32272 6316
rect 32220 6273 32229 6307
rect 32229 6273 32263 6307
rect 32263 6273 32272 6307
rect 32220 6264 32272 6273
rect 23388 6060 23440 6112
rect 24308 6060 24360 6112
rect 25228 6103 25280 6112
rect 25228 6069 25237 6103
rect 25237 6069 25271 6103
rect 25271 6069 25280 6103
rect 25228 6060 25280 6069
rect 25320 6103 25372 6112
rect 25320 6069 25329 6103
rect 25329 6069 25363 6103
rect 25363 6069 25372 6103
rect 25320 6060 25372 6069
rect 25688 6103 25740 6112
rect 25688 6069 25697 6103
rect 25697 6069 25731 6103
rect 25731 6069 25740 6103
rect 25688 6060 25740 6069
rect 25964 6060 26016 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 8208 5856 8260 5908
rect 9404 5856 9456 5908
rect 8484 5788 8536 5840
rect 11060 5788 11112 5840
rect 11520 5788 11572 5840
rect 13268 5788 13320 5840
rect 14188 5856 14240 5908
rect 14464 5856 14516 5908
rect 15108 5788 15160 5840
rect 16672 5856 16724 5908
rect 18052 5856 18104 5908
rect 19064 5856 19116 5908
rect 20904 5856 20956 5908
rect 20996 5856 21048 5908
rect 22376 5856 22428 5908
rect 23020 5899 23072 5908
rect 23020 5865 23029 5899
rect 23029 5865 23063 5899
rect 23063 5865 23072 5899
rect 23020 5856 23072 5865
rect 24400 5856 24452 5908
rect 20352 5788 20404 5840
rect 23296 5788 23348 5840
rect 5356 5720 5408 5772
rect 5540 5652 5592 5704
rect 7104 5627 7156 5636
rect 7104 5593 7113 5627
rect 7113 5593 7147 5627
rect 7147 5593 7156 5627
rect 7104 5584 7156 5593
rect 7380 5695 7432 5704
rect 7380 5661 7389 5695
rect 7389 5661 7423 5695
rect 7423 5661 7432 5695
rect 7380 5652 7432 5661
rect 8668 5652 8720 5704
rect 9312 5720 9364 5772
rect 11612 5720 11664 5772
rect 12532 5720 12584 5772
rect 17132 5720 17184 5772
rect 17224 5720 17276 5772
rect 18972 5720 19024 5772
rect 25044 5788 25096 5840
rect 25228 5720 25280 5772
rect 9128 5652 9180 5704
rect 11244 5652 11296 5704
rect 12072 5652 12124 5704
rect 15292 5652 15344 5704
rect 18512 5695 18564 5704
rect 18512 5661 18521 5695
rect 18521 5661 18555 5695
rect 18555 5661 18564 5695
rect 18512 5652 18564 5661
rect 18788 5652 18840 5704
rect 20444 5652 20496 5704
rect 20996 5652 21048 5704
rect 23388 5695 23440 5704
rect 23388 5661 23397 5695
rect 23397 5661 23431 5695
rect 23431 5661 23440 5695
rect 23388 5652 23440 5661
rect 31760 5652 31812 5704
rect 11428 5584 11480 5636
rect 11612 5584 11664 5636
rect 13452 5584 13504 5636
rect 8300 5559 8352 5568
rect 8300 5525 8309 5559
rect 8309 5525 8343 5559
rect 8343 5525 8352 5559
rect 8300 5516 8352 5525
rect 8392 5559 8444 5568
rect 8392 5525 8401 5559
rect 8401 5525 8435 5559
rect 8435 5525 8444 5559
rect 8392 5516 8444 5525
rect 11888 5516 11940 5568
rect 13268 5516 13320 5568
rect 17040 5584 17092 5636
rect 14096 5516 14148 5568
rect 14464 5516 14516 5568
rect 16672 5516 16724 5568
rect 16764 5516 16816 5568
rect 17868 5584 17920 5636
rect 19616 5584 19668 5636
rect 23204 5627 23256 5636
rect 23204 5593 23213 5627
rect 23213 5593 23247 5627
rect 23247 5593 23256 5627
rect 23204 5584 23256 5593
rect 23480 5627 23532 5636
rect 23480 5593 23489 5627
rect 23489 5593 23523 5627
rect 23523 5593 23532 5627
rect 23480 5584 23532 5593
rect 17224 5516 17276 5568
rect 24584 5516 24636 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 1308 5312 1360 5364
rect 12072 5355 12124 5364
rect 12072 5321 12081 5355
rect 12081 5321 12115 5355
rect 12115 5321 12124 5355
rect 12072 5312 12124 5321
rect 8208 5287 8260 5296
rect 8208 5253 8217 5287
rect 8217 5253 8251 5287
rect 8251 5253 8260 5287
rect 8208 5244 8260 5253
rect 3240 5176 3292 5228
rect 8484 5219 8536 5228
rect 8484 5185 8493 5219
rect 8493 5185 8527 5219
rect 8527 5185 8536 5219
rect 8484 5176 8536 5185
rect 10968 5244 11020 5296
rect 21088 5312 21140 5364
rect 23204 5312 23256 5364
rect 14372 5244 14424 5296
rect 11888 5219 11940 5228
rect 11888 5185 11897 5219
rect 11897 5185 11931 5219
rect 11931 5185 11940 5219
rect 11888 5176 11940 5185
rect 8300 5108 8352 5160
rect 9588 5108 9640 5160
rect 11336 5108 11388 5160
rect 8024 5040 8076 5092
rect 8392 5015 8444 5024
rect 8392 4981 8401 5015
rect 8401 4981 8435 5015
rect 8435 4981 8444 5015
rect 8392 4972 8444 4981
rect 10048 5040 10100 5092
rect 14280 5176 14332 5228
rect 14464 5219 14516 5228
rect 14464 5185 14473 5219
rect 14473 5185 14507 5219
rect 14507 5185 14516 5219
rect 14464 5176 14516 5185
rect 16120 5244 16172 5296
rect 15016 5176 15068 5228
rect 18512 5176 18564 5228
rect 23572 5219 23624 5228
rect 23572 5185 23581 5219
rect 23581 5185 23615 5219
rect 23615 5185 23624 5219
rect 23572 5176 23624 5185
rect 23756 5219 23808 5228
rect 23756 5185 23765 5219
rect 23765 5185 23799 5219
rect 23799 5185 23808 5219
rect 23756 5176 23808 5185
rect 23940 5219 23992 5228
rect 23940 5185 23949 5219
rect 23949 5185 23983 5219
rect 23983 5185 23992 5219
rect 23940 5176 23992 5185
rect 24216 5176 24268 5228
rect 15752 5108 15804 5160
rect 16028 5108 16080 5160
rect 18144 5151 18196 5160
rect 18144 5117 18153 5151
rect 18153 5117 18187 5151
rect 18187 5117 18196 5151
rect 18144 5108 18196 5117
rect 24492 5219 24544 5228
rect 24492 5185 24501 5219
rect 24501 5185 24535 5219
rect 24535 5185 24544 5219
rect 24492 5176 24544 5185
rect 31576 5312 31628 5364
rect 30380 5244 30432 5296
rect 29828 5176 29880 5228
rect 25688 5151 25740 5160
rect 25688 5117 25697 5151
rect 25697 5117 25731 5151
rect 25731 5117 25740 5151
rect 25688 5108 25740 5117
rect 14648 5083 14700 5092
rect 14648 5049 14657 5083
rect 14657 5049 14691 5083
rect 14691 5049 14700 5083
rect 14648 5040 14700 5049
rect 14372 4972 14424 5024
rect 16212 4972 16264 5024
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 24124 5015 24176 5024
rect 24124 4981 24133 5015
rect 24133 4981 24167 5015
rect 24167 4981 24176 5015
rect 24124 4972 24176 4981
rect 24216 5015 24268 5024
rect 24216 4981 24225 5015
rect 24225 4981 24259 5015
rect 24259 4981 24268 5015
rect 24216 4972 24268 4981
rect 24768 4972 24820 5024
rect 24952 4972 25004 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 9588 4632 9640 4684
rect 9956 4607 10008 4616
rect 9956 4573 9965 4607
rect 9965 4573 9999 4607
rect 9999 4573 10008 4607
rect 9956 4564 10008 4573
rect 10968 4564 11020 4616
rect 14464 4768 14516 4820
rect 14648 4768 14700 4820
rect 14740 4811 14792 4820
rect 14740 4777 14749 4811
rect 14749 4777 14783 4811
rect 14783 4777 14792 4811
rect 14740 4768 14792 4777
rect 12624 4743 12676 4752
rect 12624 4709 12633 4743
rect 12633 4709 12667 4743
rect 12667 4709 12676 4743
rect 12624 4700 12676 4709
rect 14372 4700 14424 4752
rect 16120 4811 16172 4820
rect 16120 4777 16129 4811
rect 16129 4777 16163 4811
rect 16163 4777 16172 4811
rect 16120 4768 16172 4777
rect 16304 4811 16356 4820
rect 16304 4777 16313 4811
rect 16313 4777 16347 4811
rect 16347 4777 16356 4811
rect 16304 4768 16356 4777
rect 26240 4768 26292 4820
rect 22468 4700 22520 4752
rect 12808 4607 12860 4616
rect 12808 4573 12817 4607
rect 12817 4573 12851 4607
rect 12851 4573 12860 4607
rect 12808 4564 12860 4573
rect 15752 4632 15804 4684
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 14556 4564 14608 4573
rect 14648 4564 14700 4616
rect 16212 4564 16264 4616
rect 18144 4564 18196 4616
rect 19708 4564 19760 4616
rect 20812 4607 20864 4616
rect 20812 4573 20821 4607
rect 20821 4573 20855 4607
rect 20855 4573 20864 4607
rect 20812 4564 20864 4573
rect 21180 4607 21232 4616
rect 21180 4573 21189 4607
rect 21189 4573 21223 4607
rect 21223 4573 21232 4607
rect 21180 4564 21232 4573
rect 22192 4564 22244 4616
rect 23572 4607 23624 4616
rect 23572 4573 23581 4607
rect 23581 4573 23615 4607
rect 23615 4573 23624 4607
rect 23572 4564 23624 4573
rect 23756 4564 23808 4616
rect 24216 4607 24268 4616
rect 24216 4573 24225 4607
rect 24225 4573 24259 4607
rect 24259 4573 24268 4607
rect 24216 4564 24268 4573
rect 24584 4607 24636 4616
rect 24584 4573 24593 4607
rect 24593 4573 24627 4607
rect 24627 4573 24636 4607
rect 24584 4564 24636 4573
rect 24860 4607 24912 4616
rect 24860 4573 24869 4607
rect 24869 4573 24903 4607
rect 24903 4573 24912 4607
rect 24860 4564 24912 4573
rect 24952 4564 25004 4616
rect 20996 4539 21048 4548
rect 20996 4505 21005 4539
rect 21005 4505 21039 4539
rect 21039 4505 21048 4539
rect 20996 4496 21048 4505
rect 21088 4539 21140 4548
rect 21088 4505 21097 4539
rect 21097 4505 21131 4539
rect 21131 4505 21140 4539
rect 21088 4496 21140 4505
rect 18512 4428 18564 4480
rect 21364 4471 21416 4480
rect 21364 4437 21373 4471
rect 21373 4437 21407 4471
rect 21407 4437 21416 4471
rect 21364 4428 21416 4437
rect 26148 4496 26200 4548
rect 25688 4428 25740 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 1124 4224 1176 4276
rect 12808 4224 12860 4276
rect 19708 4224 19760 4276
rect 21180 4224 21232 4276
rect 23940 4224 23992 4276
rect 2412 4088 2464 4140
rect 16580 4088 16632 4140
rect 16764 4088 16816 4140
rect 18788 4088 18840 4140
rect 21916 4088 21968 4140
rect 22468 4131 22520 4140
rect 22468 4097 22502 4131
rect 22502 4097 22520 4131
rect 22468 4088 22520 4097
rect 24124 4131 24176 4140
rect 24124 4097 24158 4131
rect 24158 4097 24176 4131
rect 24124 4088 24176 4097
rect 24860 4088 24912 4140
rect 20904 4063 20956 4072
rect 20904 4029 20913 4063
rect 20913 4029 20947 4063
rect 20947 4029 20956 4063
rect 20904 4020 20956 4029
rect 25228 4020 25280 4072
rect 25872 4063 25924 4072
rect 25872 4029 25881 4063
rect 25881 4029 25915 4063
rect 25915 4029 25924 4063
rect 25872 4020 25924 4029
rect 17684 3884 17736 3936
rect 23572 3927 23624 3936
rect 23572 3893 23581 3927
rect 23581 3893 23615 3927
rect 23615 3893 23624 3927
rect 23572 3884 23624 3893
rect 31024 3952 31076 4004
rect 25228 3927 25280 3936
rect 25228 3893 25237 3927
rect 25237 3893 25271 3927
rect 25271 3893 25280 3927
rect 25228 3884 25280 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 10232 3680 10284 3732
rect 31392 3680 31444 3732
rect 16764 3655 16816 3664
rect 16764 3621 16773 3655
rect 16773 3621 16807 3655
rect 16807 3621 16816 3655
rect 16764 3612 16816 3621
rect 18788 3655 18840 3664
rect 18788 3621 18797 3655
rect 18797 3621 18831 3655
rect 18831 3621 18840 3655
rect 18788 3612 18840 3621
rect 16488 3544 16540 3596
rect 17684 3544 17736 3596
rect 18236 3519 18288 3528
rect 18236 3485 18245 3519
rect 18245 3485 18279 3519
rect 18279 3485 18288 3519
rect 18236 3476 18288 3485
rect 18512 3519 18564 3528
rect 18512 3485 18521 3519
rect 18521 3485 18555 3519
rect 18555 3485 18564 3519
rect 18512 3476 18564 3485
rect 21916 3587 21968 3596
rect 21916 3553 21925 3587
rect 21925 3553 21959 3587
rect 21959 3553 21968 3587
rect 21916 3544 21968 3553
rect 21088 3476 21140 3528
rect 21364 3476 21416 3528
rect 20996 3408 21048 3460
rect 20904 3340 20956 3392
rect 21364 3340 21416 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 16580 3136 16632 3188
rect 28448 3136 28500 3188
rect 5816 3068 5868 3120
rect 28080 3068 28132 3120
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 17684 2388 17736 2440
rect 19708 2431 19760 2440
rect 19708 2397 19717 2431
rect 19717 2397 19751 2431
rect 19751 2397 19760 2431
rect 19708 2388 19760 2397
rect 21364 2431 21416 2440
rect 21364 2397 21373 2431
rect 21373 2397 21407 2431
rect 21407 2397 21416 2431
rect 21364 2388 21416 2397
rect 23572 2388 23624 2440
rect 25688 2388 25740 2440
rect 25872 2431 25924 2440
rect 25872 2397 25881 2431
rect 25881 2397 25915 2431
rect 25915 2397 25924 2431
rect 25872 2388 25924 2397
rect 29644 2388 29696 2440
rect 17408 2252 17460 2304
rect 19340 2252 19392 2304
rect 21272 2252 21324 2304
rect 22560 2252 22612 2304
rect 24492 2252 24544 2304
rect 25780 2252 25832 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 16762 33200 16818 34000
rect 18694 33200 18750 34000
rect 21270 33200 21326 34000
rect 23202 33200 23258 34000
rect 25134 33200 25190 34000
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 16776 31414 16804 33200
rect 18708 31482 18736 33200
rect 21284 31482 21312 33200
rect 18696 31476 18748 31482
rect 18696 31418 18748 31424
rect 21272 31476 21324 31482
rect 21272 31418 21324 31424
rect 23216 31414 23244 33200
rect 25148 31482 25176 33200
rect 25136 31476 25188 31482
rect 25136 31418 25188 31424
rect 16764 31408 16816 31414
rect 16764 31350 16816 31356
rect 23204 31408 23256 31414
rect 23204 31350 23256 31356
rect 17132 31340 17184 31346
rect 17132 31282 17184 31288
rect 19340 31340 19392 31346
rect 19340 31282 19392 31288
rect 21916 31340 21968 31346
rect 21916 31282 21968 31288
rect 23664 31340 23716 31346
rect 23664 31282 23716 31288
rect 25320 31340 25372 31346
rect 25320 31282 25372 31288
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 13726 30832 13782 30841
rect 13452 30796 13504 30802
rect 13726 30767 13782 30776
rect 13452 30738 13504 30744
rect 1308 30592 1360 30598
rect 1308 30534 1360 30540
rect 1122 30288 1178 30297
rect 1122 30223 1178 30232
rect 940 30048 992 30054
rect 940 29990 992 29996
rect 848 25900 900 25906
rect 848 25842 900 25848
rect 860 25809 888 25842
rect 846 25800 902 25809
rect 846 25735 902 25744
rect 386 24712 442 24721
rect 386 24647 442 24656
rect 400 7993 428 24647
rect 848 24200 900 24206
rect 754 24168 810 24177
rect 848 24142 900 24148
rect 754 24103 810 24112
rect 478 23216 534 23225
rect 478 23151 534 23160
rect 492 16726 520 23151
rect 664 21344 716 21350
rect 664 21286 716 21292
rect 570 20904 626 20913
rect 570 20839 626 20848
rect 480 16720 532 16726
rect 480 16662 532 16668
rect 584 13462 612 20839
rect 676 14113 704 21286
rect 662 14104 718 14113
rect 662 14039 718 14048
rect 572 13456 624 13462
rect 572 13398 624 13404
rect 768 10826 796 24103
rect 860 24041 888 24142
rect 846 24032 902 24041
rect 846 23967 902 23976
rect 952 23746 980 29990
rect 1032 29776 1084 29782
rect 1032 29718 1084 29724
rect 860 23718 980 23746
rect 860 18873 888 23718
rect 940 23656 992 23662
rect 940 23598 992 23604
rect 846 18864 902 18873
rect 846 18799 902 18808
rect 952 17649 980 23598
rect 1044 20777 1072 29718
rect 1030 20768 1086 20777
rect 1030 20703 1086 20712
rect 938 17640 994 17649
rect 938 17575 994 17584
rect 848 16584 900 16590
rect 846 16552 848 16561
rect 900 16552 902 16561
rect 846 16487 902 16496
rect 1136 15978 1164 30223
rect 1216 29844 1268 29850
rect 1216 29786 1268 29792
rect 1228 19174 1256 29786
rect 1320 23662 1348 30534
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 6826 30424 6882 30433
rect 6092 30388 6144 30394
rect 6826 30359 6882 30368
rect 6092 30330 6144 30336
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 5632 29708 5684 29714
rect 5632 29650 5684 29656
rect 3240 29640 3292 29646
rect 3240 29582 3292 29588
rect 2780 29232 2832 29238
rect 2780 29174 2832 29180
rect 1400 29164 1452 29170
rect 1400 29106 1452 29112
rect 1412 28665 1440 29106
rect 2228 29096 2280 29102
rect 2792 29050 2820 29174
rect 3056 29164 3108 29170
rect 3056 29106 3108 29112
rect 2228 29038 2280 29044
rect 1676 28960 1728 28966
rect 1676 28902 1728 28908
rect 1398 28656 1454 28665
rect 1398 28591 1454 28600
rect 1688 28558 1716 28902
rect 1400 28552 1452 28558
rect 1400 28494 1452 28500
rect 1676 28552 1728 28558
rect 1676 28494 1728 28500
rect 1412 28014 1440 28494
rect 1676 28076 1728 28082
rect 1676 28018 1728 28024
rect 1400 28008 1452 28014
rect 1400 27950 1452 27956
rect 1490 27976 1546 27985
rect 1412 26382 1440 27950
rect 1490 27911 1546 27920
rect 1504 27470 1532 27911
rect 1688 27674 1716 28018
rect 1676 27668 1728 27674
rect 1676 27610 1728 27616
rect 2240 27606 2268 29038
rect 2700 29022 2820 29050
rect 2872 29028 2924 29034
rect 2504 28552 2556 28558
rect 2504 28494 2556 28500
rect 2320 28416 2372 28422
rect 2320 28358 2372 28364
rect 2228 27600 2280 27606
rect 2228 27542 2280 27548
rect 1492 27464 1544 27470
rect 1492 27406 1544 27412
rect 2332 26994 2360 28358
rect 2516 27538 2544 28494
rect 2700 28422 2728 29022
rect 2872 28970 2924 28976
rect 2884 28762 2912 28970
rect 2964 28960 3016 28966
rect 2964 28902 3016 28908
rect 2872 28756 2924 28762
rect 2872 28698 2924 28704
rect 2688 28416 2740 28422
rect 2688 28358 2740 28364
rect 2884 27538 2912 28698
rect 2976 28490 3004 28902
rect 2964 28484 3016 28490
rect 2964 28426 3016 28432
rect 2976 28014 3004 28426
rect 2964 28008 3016 28014
rect 2964 27950 3016 27956
rect 2976 27606 3004 27950
rect 2964 27600 3016 27606
rect 2964 27542 3016 27548
rect 2504 27532 2556 27538
rect 2504 27474 2556 27480
rect 2872 27532 2924 27538
rect 2872 27474 2924 27480
rect 3068 27470 3096 29106
rect 3148 28960 3200 28966
rect 3148 28902 3200 28908
rect 3160 28626 3188 28902
rect 3148 28620 3200 28626
rect 3148 28562 3200 28568
rect 3160 28082 3188 28562
rect 3252 28218 3280 29582
rect 3332 29504 3384 29510
rect 3332 29446 3384 29452
rect 3424 29504 3476 29510
rect 3424 29446 3476 29452
rect 5264 29504 5316 29510
rect 5264 29446 5316 29452
rect 3344 28558 3372 29446
rect 3436 29238 3464 29446
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 3516 29300 3568 29306
rect 3516 29242 3568 29248
rect 3424 29232 3476 29238
rect 3424 29174 3476 29180
rect 3332 28552 3384 28558
rect 3332 28494 3384 28500
rect 3332 28416 3384 28422
rect 3330 28384 3332 28393
rect 3384 28384 3386 28393
rect 3330 28319 3386 28328
rect 3240 28212 3292 28218
rect 3240 28154 3292 28160
rect 3332 28144 3384 28150
rect 3332 28086 3384 28092
rect 3148 28076 3200 28082
rect 3148 28018 3200 28024
rect 3056 27464 3108 27470
rect 3056 27406 3108 27412
rect 3068 27130 3096 27406
rect 3160 27402 3188 28018
rect 3240 28008 3292 28014
rect 3240 27950 3292 27956
rect 3148 27396 3200 27402
rect 3148 27338 3200 27344
rect 3252 27334 3280 27950
rect 3344 27538 3372 28086
rect 3332 27532 3384 27538
rect 3332 27474 3384 27480
rect 3240 27328 3292 27334
rect 3240 27270 3292 27276
rect 3056 27124 3108 27130
rect 3056 27066 3108 27072
rect 2780 27056 2832 27062
rect 2780 26998 2832 27004
rect 2320 26988 2372 26994
rect 2320 26930 2372 26936
rect 2596 26920 2648 26926
rect 2594 26888 2596 26897
rect 2648 26888 2650 26897
rect 2594 26823 2650 26832
rect 1400 26376 1452 26382
rect 1400 26318 1452 26324
rect 1412 25294 1440 26318
rect 2792 26314 2820 26998
rect 3252 26994 3280 27270
rect 2872 26988 2924 26994
rect 2872 26930 2924 26936
rect 3240 26988 3292 26994
rect 3240 26930 3292 26936
rect 2884 26450 2912 26930
rect 3056 26920 3108 26926
rect 3108 26868 3188 26874
rect 3056 26862 3188 26868
rect 2964 26852 3016 26858
rect 3068 26846 3188 26862
rect 2964 26794 3016 26800
rect 2872 26444 2924 26450
rect 2872 26386 2924 26392
rect 1676 26308 1728 26314
rect 1676 26250 1728 26256
rect 2780 26308 2832 26314
rect 2780 26250 2832 26256
rect 1688 26042 1716 26250
rect 1676 26036 1728 26042
rect 1676 25978 1728 25984
rect 2792 25906 2820 26250
rect 2884 26042 2912 26386
rect 2976 26382 3004 26794
rect 3160 26790 3188 26846
rect 3148 26784 3200 26790
rect 3148 26726 3200 26732
rect 2964 26376 3016 26382
rect 2964 26318 3016 26324
rect 2872 26036 2924 26042
rect 2872 25978 2924 25984
rect 2976 25974 3004 26318
rect 3160 26246 3188 26726
rect 3148 26240 3200 26246
rect 3148 26182 3200 26188
rect 2964 25968 3016 25974
rect 2964 25910 3016 25916
rect 3160 25906 3188 26182
rect 3344 25906 3372 27474
rect 3424 27328 3476 27334
rect 3424 27270 3476 27276
rect 2780 25900 2832 25906
rect 2780 25842 2832 25848
rect 3148 25900 3200 25906
rect 3148 25842 3200 25848
rect 3332 25900 3384 25906
rect 3332 25842 3384 25848
rect 2134 25800 2190 25809
rect 3436 25786 3464 27270
rect 3528 27130 3556 29242
rect 4344 29164 4396 29170
rect 4172 29124 4344 29152
rect 3792 28960 3844 28966
rect 3698 28928 3754 28937
rect 3792 28902 3844 28908
rect 3884 28960 3936 28966
rect 4172 28948 4200 29124
rect 4344 29106 4396 29112
rect 4712 29164 4764 29170
rect 4712 29106 4764 29112
rect 4620 29096 4672 29102
rect 4620 29038 4672 29044
rect 3884 28902 3936 28908
rect 4080 28920 4200 28948
rect 4250 29008 4306 29017
rect 4250 28943 4252 28952
rect 3698 28863 3754 28872
rect 3712 28490 3740 28863
rect 3700 28484 3752 28490
rect 3700 28426 3752 28432
rect 3804 28150 3832 28902
rect 3792 28144 3844 28150
rect 3792 28086 3844 28092
rect 3608 27872 3660 27878
rect 3608 27814 3660 27820
rect 3516 27124 3568 27130
rect 3516 27066 3568 27072
rect 3528 26994 3556 27066
rect 3516 26988 3568 26994
rect 3516 26930 3568 26936
rect 3516 26784 3568 26790
rect 3516 26726 3568 26732
rect 2134 25735 2190 25744
rect 3252 25758 3464 25786
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 1308 23656 1360 23662
rect 1308 23598 1360 23604
rect 1412 22574 1440 25230
rect 1676 25220 1728 25226
rect 1676 25162 1728 25168
rect 1688 24410 1716 25162
rect 1766 25120 1822 25129
rect 1766 25055 1822 25064
rect 1676 24404 1728 24410
rect 1676 24346 1728 24352
rect 1676 22636 1728 22642
rect 1676 22578 1728 22584
rect 1400 22568 1452 22574
rect 1400 22510 1452 22516
rect 1412 21593 1440 22510
rect 1688 22094 1716 22578
rect 1596 22066 1716 22094
rect 1398 21584 1454 21593
rect 1398 21519 1400 21528
rect 1452 21519 1454 21528
rect 1492 21548 1544 21554
rect 1400 21490 1452 21496
rect 1492 21490 1544 21496
rect 1412 19922 1440 21490
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1308 19372 1360 19378
rect 1308 19314 1360 19320
rect 1216 19168 1268 19174
rect 1320 19145 1348 19314
rect 1216 19110 1268 19116
rect 1306 19136 1362 19145
rect 1306 19071 1362 19080
rect 1412 18834 1440 19858
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1308 18760 1360 18766
rect 1308 18702 1360 18708
rect 1124 15972 1176 15978
rect 1124 15914 1176 15920
rect 1122 15464 1178 15473
rect 1122 15399 1178 15408
rect 846 14512 902 14521
rect 846 14447 902 14456
rect 860 14414 888 14447
rect 848 14408 900 14414
rect 848 14350 900 14356
rect 938 10840 994 10849
rect 768 10798 938 10826
rect 938 10775 994 10784
rect 386 7984 442 7993
rect 386 7919 442 7928
rect 1136 4282 1164 15399
rect 1320 5370 1348 18702
rect 1504 14618 1532 21490
rect 1596 16454 1624 22066
rect 1780 21350 1808 25055
rect 2044 24812 2096 24818
rect 2044 24754 2096 24760
rect 1860 24200 1912 24206
rect 1860 24142 1912 24148
rect 1872 23798 1900 24142
rect 1860 23792 1912 23798
rect 1860 23734 1912 23740
rect 2056 23322 2084 24754
rect 2148 24410 2176 25735
rect 3056 25288 3108 25294
rect 3056 25230 3108 25236
rect 3148 25288 3200 25294
rect 3148 25230 3200 25236
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2884 24886 2912 25094
rect 2688 24880 2740 24886
rect 2688 24822 2740 24828
rect 2872 24880 2924 24886
rect 2872 24822 2924 24828
rect 2320 24812 2372 24818
rect 2320 24754 2372 24760
rect 2412 24812 2464 24818
rect 2412 24754 2464 24760
rect 2136 24404 2188 24410
rect 2136 24346 2188 24352
rect 2228 23724 2280 23730
rect 2228 23666 2280 23672
rect 2044 23316 2096 23322
rect 2044 23258 2096 23264
rect 2240 23050 2268 23666
rect 2332 23594 2360 24754
rect 2424 23866 2452 24754
rect 2596 24608 2648 24614
rect 2596 24550 2648 24556
rect 2608 24206 2636 24550
rect 2700 24342 2728 24822
rect 2688 24336 2740 24342
rect 2688 24278 2740 24284
rect 2700 24206 2728 24278
rect 2596 24200 2648 24206
rect 2596 24142 2648 24148
rect 2688 24200 2740 24206
rect 2688 24142 2740 24148
rect 2780 24132 2832 24138
rect 2884 24120 2912 24822
rect 2832 24092 2912 24120
rect 2780 24074 2832 24080
rect 3068 23866 3096 25230
rect 3160 24682 3188 25230
rect 3148 24676 3200 24682
rect 3148 24618 3200 24624
rect 3160 24274 3188 24618
rect 3148 24268 3200 24274
rect 3148 24210 3200 24216
rect 2412 23860 2464 23866
rect 2412 23802 2464 23808
rect 2964 23860 3016 23866
rect 2964 23802 3016 23808
rect 3056 23860 3108 23866
rect 3056 23802 3108 23808
rect 2872 23724 2924 23730
rect 2872 23666 2924 23672
rect 2412 23656 2464 23662
rect 2412 23598 2464 23604
rect 2320 23588 2372 23594
rect 2320 23530 2372 23536
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 2228 23044 2280 23050
rect 2228 22986 2280 22992
rect 2240 22234 2268 22986
rect 2332 22778 2360 23054
rect 2320 22772 2372 22778
rect 2320 22714 2372 22720
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 2424 22094 2452 23598
rect 2780 23588 2832 23594
rect 2780 23530 2832 23536
rect 2792 23186 2820 23530
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 2792 22642 2820 23122
rect 2780 22636 2832 22642
rect 2780 22578 2832 22584
rect 2240 22066 2452 22094
rect 2044 22024 2096 22030
rect 2044 21966 2096 21972
rect 2056 21690 2084 21966
rect 2044 21684 2096 21690
rect 2044 21626 2096 21632
rect 1768 21344 1820 21350
rect 1768 21286 1820 21292
rect 2240 21146 2268 22066
rect 2688 22024 2740 22030
rect 2688 21966 2740 21972
rect 2320 21888 2372 21894
rect 2320 21830 2372 21836
rect 2332 21622 2360 21830
rect 2700 21706 2728 21966
rect 2700 21678 2820 21706
rect 2320 21616 2372 21622
rect 2320 21558 2372 21564
rect 2228 21140 2280 21146
rect 2228 21082 2280 21088
rect 1768 21072 1820 21078
rect 1768 21014 1820 21020
rect 1676 20800 1728 20806
rect 1676 20742 1728 20748
rect 1688 20602 1716 20742
rect 1676 20596 1728 20602
rect 1676 20538 1728 20544
rect 1780 20466 1808 21014
rect 2240 20942 2268 21082
rect 2044 20936 2096 20942
rect 2044 20878 2096 20884
rect 2228 20936 2280 20942
rect 2228 20878 2280 20884
rect 2332 20890 2360 21558
rect 2412 21412 2464 21418
rect 2412 21354 2464 21360
rect 2424 21078 2452 21354
rect 2688 21344 2740 21350
rect 2688 21286 2740 21292
rect 2412 21072 2464 21078
rect 2412 21014 2464 21020
rect 2596 21072 2648 21078
rect 2596 21014 2648 21020
rect 2412 20936 2464 20942
rect 2332 20884 2412 20890
rect 2332 20878 2464 20884
rect 1768 20460 1820 20466
rect 1768 20402 1820 20408
rect 1676 19780 1728 19786
rect 1676 19722 1728 19728
rect 1688 19514 1716 19722
rect 1858 19680 1914 19689
rect 1858 19615 1914 19624
rect 1676 19508 1728 19514
rect 1676 19450 1728 19456
rect 1676 18692 1728 18698
rect 1676 18634 1728 18640
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 1688 11354 1716 18634
rect 1872 11626 1900 19615
rect 2056 18970 2084 20878
rect 2332 20862 2452 20878
rect 2226 20632 2282 20641
rect 2226 20567 2282 20576
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 2240 16538 2268 20567
rect 2332 20398 2360 20862
rect 2608 20398 2636 21014
rect 2320 20392 2372 20398
rect 2320 20334 2372 20340
rect 2596 20392 2648 20398
rect 2596 20334 2648 20340
rect 2332 19786 2360 20334
rect 2608 19854 2636 20334
rect 2700 20330 2728 21286
rect 2688 20324 2740 20330
rect 2688 20266 2740 20272
rect 2792 20262 2820 21678
rect 2884 20788 2912 23666
rect 2976 22778 3004 23802
rect 2964 22772 3016 22778
rect 2964 22714 3016 22720
rect 2976 22506 3004 22714
rect 3068 22710 3096 23802
rect 3252 23644 3280 25758
rect 3332 25152 3384 25158
rect 3332 25094 3384 25100
rect 3424 25152 3476 25158
rect 3424 25094 3476 25100
rect 3344 24274 3372 25094
rect 3436 24410 3464 25094
rect 3528 24954 3556 26726
rect 3620 25378 3648 27814
rect 3700 27600 3752 27606
rect 3698 27568 3700 27577
rect 3752 27568 3754 27577
rect 3698 27503 3754 27512
rect 3896 27402 3924 28902
rect 4080 28762 4108 28920
rect 4304 28943 4306 28952
rect 4252 28902 4304 28908
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4068 28756 4120 28762
rect 3988 28716 4068 28744
rect 3884 27396 3936 27402
rect 3884 27338 3936 27344
rect 3792 26988 3844 26994
rect 3792 26930 3844 26936
rect 3884 26988 3936 26994
rect 3884 26930 3936 26936
rect 3804 26586 3832 26930
rect 3792 26580 3844 26586
rect 3792 26522 3844 26528
rect 3700 26512 3752 26518
rect 3700 26454 3752 26460
rect 3712 26314 3740 26454
rect 3700 26308 3752 26314
rect 3700 26250 3752 26256
rect 3700 25900 3752 25906
rect 3700 25842 3752 25848
rect 3712 25702 3740 25842
rect 3700 25696 3752 25702
rect 3700 25638 3752 25644
rect 3896 25498 3924 26930
rect 3988 26926 4016 28716
rect 4068 28698 4120 28704
rect 4344 28756 4396 28762
rect 4344 28698 4396 28704
rect 4356 28558 4384 28698
rect 4632 28694 4660 29038
rect 4620 28688 4672 28694
rect 4620 28630 4672 28636
rect 4252 28552 4304 28558
rect 4252 28494 4304 28500
rect 4344 28552 4396 28558
rect 4344 28494 4396 28500
rect 4068 28416 4120 28422
rect 4068 28358 4120 28364
rect 4080 27946 4108 28358
rect 4264 28082 4292 28494
rect 4356 28150 4384 28494
rect 4528 28416 4580 28422
rect 4528 28358 4580 28364
rect 4620 28416 4672 28422
rect 4620 28358 4672 28364
rect 4344 28144 4396 28150
rect 4344 28086 4396 28092
rect 4252 28076 4304 28082
rect 4252 28018 4304 28024
rect 4068 27940 4120 27946
rect 4540 27928 4568 28358
rect 4632 28121 4660 28358
rect 4618 28112 4674 28121
rect 4618 28047 4674 28056
rect 4620 27940 4672 27946
rect 4540 27900 4620 27928
rect 4068 27882 4120 27888
rect 4620 27882 4672 27888
rect 4080 27606 4108 27882
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4068 27600 4120 27606
rect 4068 27542 4120 27548
rect 4632 27538 4660 27882
rect 4620 27532 4672 27538
rect 4620 27474 4672 27480
rect 4252 27464 4304 27470
rect 4252 27406 4304 27412
rect 3976 26920 4028 26926
rect 3976 26862 4028 26868
rect 4068 26852 4120 26858
rect 4068 26794 4120 26800
rect 3976 26512 4028 26518
rect 3976 26454 4028 26460
rect 3988 26246 4016 26454
rect 4080 26450 4108 26794
rect 4264 26790 4292 27406
rect 4724 27130 4752 29106
rect 4896 28960 4948 28966
rect 4896 28902 4948 28908
rect 4988 28960 5040 28966
rect 4988 28902 5040 28908
rect 4908 28762 4936 28902
rect 4896 28756 4948 28762
rect 4896 28698 4948 28704
rect 5000 28626 5028 28902
rect 4804 28620 4856 28626
rect 4804 28562 4856 28568
rect 4988 28620 5040 28626
rect 4988 28562 5040 28568
rect 4816 28150 4844 28562
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4804 28144 4856 28150
rect 4804 28086 4856 28092
rect 4816 27674 4844 28086
rect 5276 28064 5304 29446
rect 5448 28960 5500 28966
rect 5448 28902 5500 28908
rect 5356 28688 5408 28694
rect 5356 28630 5408 28636
rect 5368 28218 5396 28630
rect 5356 28212 5408 28218
rect 5356 28154 5408 28160
rect 5460 28082 5488 28902
rect 4908 28036 5304 28064
rect 5448 28076 5500 28082
rect 4804 27668 4856 27674
rect 4804 27610 4856 27616
rect 4908 27316 4936 28036
rect 5448 28018 5500 28024
rect 4988 27940 5040 27946
rect 4988 27882 5040 27888
rect 5000 27606 5028 27882
rect 5172 27668 5224 27674
rect 5172 27610 5224 27616
rect 4988 27600 5040 27606
rect 4988 27542 5040 27548
rect 5184 27418 5212 27610
rect 5460 27520 5488 28018
rect 5644 27606 5672 29650
rect 5908 28960 5960 28966
rect 5908 28902 5960 28908
rect 5816 28756 5868 28762
rect 5816 28698 5868 28704
rect 5828 28626 5856 28698
rect 5920 28626 5948 28902
rect 5816 28620 5868 28626
rect 5816 28562 5868 28568
rect 5908 28620 5960 28626
rect 5908 28562 5960 28568
rect 6000 28552 6052 28558
rect 6000 28494 6052 28500
rect 5724 28484 5776 28490
rect 5724 28426 5776 28432
rect 5632 27600 5684 27606
rect 5632 27542 5684 27548
rect 5460 27492 5512 27520
rect 5000 27402 5212 27418
rect 4988 27396 5212 27402
rect 5040 27390 5212 27396
rect 5484 27418 5512 27492
rect 5484 27402 5580 27418
rect 5484 27396 5592 27402
rect 5484 27390 5540 27396
rect 4988 27338 5040 27344
rect 5540 27338 5592 27344
rect 4816 27288 4936 27316
rect 5080 27328 5132 27334
rect 4712 27124 4764 27130
rect 4712 27066 4764 27072
rect 4710 27024 4766 27033
rect 4710 26959 4712 26968
rect 4764 26959 4766 26968
rect 4712 26930 4764 26936
rect 4620 26920 4672 26926
rect 4620 26862 4672 26868
rect 4252 26784 4304 26790
rect 4252 26726 4304 26732
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4160 26580 4212 26586
rect 4160 26522 4212 26528
rect 4068 26444 4120 26450
rect 4068 26386 4120 26392
rect 3976 26240 4028 26246
rect 3976 26182 4028 26188
rect 4172 25906 4200 26522
rect 4528 26444 4580 26450
rect 4528 26386 4580 26392
rect 4540 25906 4568 26386
rect 4632 26382 4660 26862
rect 4816 26790 4844 27288
rect 5132 27288 5488 27316
rect 5552 27305 5580 27338
rect 5632 27328 5684 27334
rect 5080 27270 5132 27276
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 5354 27160 5410 27169
rect 5080 27124 5132 27130
rect 5354 27095 5410 27104
rect 5080 27066 5132 27072
rect 4896 26988 4948 26994
rect 4896 26930 4948 26936
rect 4712 26784 4764 26790
rect 4712 26726 4764 26732
rect 4804 26784 4856 26790
rect 4804 26726 4856 26732
rect 4724 26382 4752 26726
rect 4908 26586 4936 26930
rect 4896 26580 4948 26586
rect 4896 26522 4948 26528
rect 5092 26518 5120 27066
rect 5080 26512 5132 26518
rect 5080 26454 5132 26460
rect 5368 26450 5396 27095
rect 5356 26444 5408 26450
rect 5356 26386 5408 26392
rect 4620 26376 4672 26382
rect 4620 26318 4672 26324
rect 4712 26376 4764 26382
rect 4712 26318 4764 26324
rect 5264 26376 5316 26382
rect 5264 26318 5316 26324
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4986 25936 5042 25945
rect 4160 25900 4212 25906
rect 4160 25842 4212 25848
rect 4528 25900 4580 25906
rect 4986 25871 4988 25880
rect 4528 25842 4580 25848
rect 5040 25871 5042 25880
rect 5080 25900 5132 25906
rect 4988 25842 5040 25848
rect 5080 25842 5132 25848
rect 5172 25900 5224 25906
rect 5172 25842 5224 25848
rect 4068 25696 4120 25702
rect 5092 25673 5120 25842
rect 5184 25702 5212 25842
rect 5276 25770 5304 26318
rect 5354 26208 5410 26217
rect 5354 26143 5410 26152
rect 5264 25764 5316 25770
rect 5264 25706 5316 25712
rect 5172 25696 5224 25702
rect 4068 25638 4120 25644
rect 5078 25664 5134 25673
rect 3884 25492 3936 25498
rect 3884 25434 3936 25440
rect 3620 25350 3924 25378
rect 3608 25288 3660 25294
rect 3608 25230 3660 25236
rect 3516 24948 3568 24954
rect 3516 24890 3568 24896
rect 3620 24682 3648 25230
rect 3792 24812 3844 24818
rect 3792 24754 3844 24760
rect 3608 24676 3660 24682
rect 3608 24618 3660 24624
rect 3700 24608 3752 24614
rect 3700 24550 3752 24556
rect 3712 24410 3740 24550
rect 3424 24404 3476 24410
rect 3424 24346 3476 24352
rect 3700 24404 3752 24410
rect 3700 24346 3752 24352
rect 3332 24268 3384 24274
rect 3332 24210 3384 24216
rect 3436 24070 3464 24346
rect 3332 24064 3384 24070
rect 3332 24006 3384 24012
rect 3424 24064 3476 24070
rect 3424 24006 3476 24012
rect 3344 23798 3372 24006
rect 3332 23792 3384 23798
rect 3332 23734 3384 23740
rect 3146 23624 3202 23633
rect 3252 23616 3372 23644
rect 3146 23559 3202 23568
rect 3160 23118 3188 23559
rect 3148 23112 3200 23118
rect 3148 23054 3200 23060
rect 3148 22976 3200 22982
rect 3148 22918 3200 22924
rect 3240 22976 3292 22982
rect 3240 22918 3292 22924
rect 3056 22704 3108 22710
rect 3056 22646 3108 22652
rect 3160 22545 3188 22918
rect 3146 22536 3202 22545
rect 2964 22500 3016 22506
rect 3146 22471 3202 22480
rect 2964 22442 3016 22448
rect 3148 22160 3200 22166
rect 3148 22102 3200 22108
rect 3160 21978 3188 22102
rect 3252 22098 3280 22918
rect 3240 22092 3292 22098
rect 3240 22034 3292 22040
rect 3344 22030 3372 23616
rect 3436 23594 3464 24006
rect 3514 23624 3570 23633
rect 3424 23588 3476 23594
rect 3514 23559 3570 23568
rect 3424 23530 3476 23536
rect 3332 22024 3384 22030
rect 3160 21950 3280 21978
rect 3332 21966 3384 21972
rect 2964 21888 3016 21894
rect 2964 21830 3016 21836
rect 3056 21888 3108 21894
rect 3056 21830 3108 21836
rect 3148 21888 3200 21894
rect 3148 21830 3200 21836
rect 2976 21690 3004 21830
rect 2964 21684 3016 21690
rect 2964 21626 3016 21632
rect 3068 21486 3096 21830
rect 3056 21480 3108 21486
rect 3056 21422 3108 21428
rect 2964 20800 3016 20806
rect 2884 20760 2964 20788
rect 2964 20742 3016 20748
rect 2780 20256 2832 20262
rect 2780 20198 2832 20204
rect 2976 19990 3004 20742
rect 3068 20534 3096 21422
rect 3160 21078 3188 21830
rect 3252 21146 3280 21950
rect 3332 21888 3384 21894
rect 3332 21830 3384 21836
rect 3424 21888 3476 21894
rect 3424 21830 3476 21836
rect 3240 21140 3292 21146
rect 3240 21082 3292 21088
rect 3148 21072 3200 21078
rect 3148 21014 3200 21020
rect 3148 20800 3200 20806
rect 3148 20742 3200 20748
rect 3240 20800 3292 20806
rect 3240 20742 3292 20748
rect 3160 20602 3188 20742
rect 3252 20602 3280 20742
rect 3148 20596 3200 20602
rect 3148 20538 3200 20544
rect 3240 20596 3292 20602
rect 3240 20538 3292 20544
rect 3056 20528 3108 20534
rect 3056 20470 3108 20476
rect 3160 20330 3188 20538
rect 3252 20466 3280 20538
rect 3344 20505 3372 21830
rect 3436 21049 3464 21830
rect 3528 21729 3556 23559
rect 3804 23322 3832 24754
rect 3896 23769 3924 25350
rect 3976 24948 4028 24954
rect 3976 24890 4028 24896
rect 3988 24274 4016 24890
rect 4080 24818 4108 25638
rect 5172 25638 5224 25644
rect 4214 25596 4522 25605
rect 5078 25599 5134 25608
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4620 25424 4672 25430
rect 4620 25366 4672 25372
rect 4344 25356 4396 25362
rect 4344 25298 4396 25304
rect 4160 25288 4212 25294
rect 4160 25230 4212 25236
rect 4068 24812 4120 24818
rect 4068 24754 4120 24760
rect 4172 24750 4200 25230
rect 4356 24857 4384 25298
rect 4342 24848 4398 24857
rect 4342 24783 4398 24792
rect 4356 24750 4384 24783
rect 4160 24744 4212 24750
rect 4160 24686 4212 24692
rect 4344 24744 4396 24750
rect 4344 24686 4396 24692
rect 4068 24676 4120 24682
rect 4068 24618 4120 24624
rect 3976 24268 4028 24274
rect 3976 24210 4028 24216
rect 3988 23866 4016 24210
rect 3976 23860 4028 23866
rect 3976 23802 4028 23808
rect 3882 23760 3938 23769
rect 4080 23730 4108 24618
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4344 24404 4396 24410
rect 4344 24346 4396 24352
rect 4160 24336 4212 24342
rect 4160 24278 4212 24284
rect 3882 23695 3938 23704
rect 4068 23724 4120 23730
rect 4068 23666 4120 23672
rect 4172 23594 4200 24278
rect 4356 23798 4384 24346
rect 4632 23798 4660 25366
rect 5264 25288 5316 25294
rect 5264 25230 5316 25236
rect 4712 25220 4764 25226
rect 4712 25162 4764 25168
rect 4724 24410 4752 25162
rect 4804 25152 4856 25158
rect 4804 25094 4856 25100
rect 4712 24404 4764 24410
rect 4712 24346 4764 24352
rect 4816 24138 4844 25094
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5276 24954 5304 25230
rect 5264 24948 5316 24954
rect 5264 24890 5316 24896
rect 5368 24410 5396 26143
rect 5356 24404 5408 24410
rect 5356 24346 5408 24352
rect 5262 24304 5318 24313
rect 5460 24290 5488 27288
rect 5538 27296 5594 27305
rect 5632 27270 5684 27276
rect 5538 27231 5594 27240
rect 5644 27169 5672 27270
rect 5630 27160 5686 27169
rect 5630 27095 5686 27104
rect 5632 26988 5684 26994
rect 5552 26948 5632 26976
rect 5552 26586 5580 26948
rect 5632 26930 5684 26936
rect 5540 26580 5592 26586
rect 5540 26522 5592 26528
rect 5552 26489 5580 26522
rect 5538 26480 5594 26489
rect 5538 26415 5594 26424
rect 5540 26376 5592 26382
rect 5736 26330 5764 28426
rect 6012 27946 6040 28494
rect 6000 27940 6052 27946
rect 6000 27882 6052 27888
rect 5816 27872 5868 27878
rect 5816 27814 5868 27820
rect 5828 27614 5856 27814
rect 5828 27586 5948 27614
rect 5920 27520 5948 27586
rect 5540 26318 5592 26324
rect 5552 25974 5580 26318
rect 5644 26302 5764 26330
rect 5828 27492 5948 27520
rect 5644 26246 5672 26302
rect 5632 26240 5684 26246
rect 5724 26240 5776 26246
rect 5632 26182 5684 26188
rect 5722 26208 5724 26217
rect 5776 26208 5778 26217
rect 5722 26143 5778 26152
rect 5632 26036 5684 26042
rect 5632 25978 5684 25984
rect 5540 25968 5592 25974
rect 5540 25910 5592 25916
rect 5644 25226 5672 25978
rect 5828 25922 5856 27492
rect 6104 26874 6132 30330
rect 6736 29028 6788 29034
rect 6736 28970 6788 28976
rect 6644 28620 6696 28626
rect 6644 28562 6696 28568
rect 6656 28422 6684 28562
rect 6748 28558 6776 28970
rect 6736 28552 6788 28558
rect 6736 28494 6788 28500
rect 6644 28416 6696 28422
rect 6748 28393 6776 28494
rect 6644 28358 6696 28364
rect 6734 28384 6790 28393
rect 6656 28218 6684 28358
rect 6734 28319 6790 28328
rect 6644 28212 6696 28218
rect 6644 28154 6696 28160
rect 6184 28076 6236 28082
rect 6184 28018 6236 28024
rect 6460 28076 6512 28082
rect 6644 28076 6696 28082
rect 6512 28036 6592 28064
rect 6460 28018 6512 28024
rect 6196 27062 6224 28018
rect 6564 27606 6592 28036
rect 6644 28018 6696 28024
rect 6552 27600 6604 27606
rect 6552 27542 6604 27548
rect 6368 27464 6420 27470
rect 6368 27406 6420 27412
rect 6276 27328 6328 27334
rect 6276 27270 6328 27276
rect 6184 27056 6236 27062
rect 6184 26998 6236 27004
rect 6104 26846 6224 26874
rect 5908 26784 5960 26790
rect 5908 26726 5960 26732
rect 6000 26784 6052 26790
rect 6000 26726 6052 26732
rect 5920 26081 5948 26726
rect 5906 26072 5962 26081
rect 5906 26007 5962 26016
rect 5736 25894 5856 25922
rect 5908 25900 5960 25906
rect 5632 25220 5684 25226
rect 5552 25180 5632 25208
rect 5552 24886 5580 25180
rect 5632 25162 5684 25168
rect 5540 24880 5592 24886
rect 5540 24822 5592 24828
rect 5262 24239 5318 24248
rect 5368 24262 5488 24290
rect 4804 24132 4856 24138
rect 4804 24074 4856 24080
rect 4344 23792 4396 23798
rect 4344 23734 4396 23740
rect 4620 23792 4672 23798
rect 4620 23734 4672 23740
rect 4712 23792 4764 23798
rect 4712 23734 4764 23740
rect 4356 23662 4384 23734
rect 4344 23656 4396 23662
rect 4344 23598 4396 23604
rect 4160 23588 4212 23594
rect 4160 23530 4212 23536
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3792 23316 3844 23322
rect 3792 23258 3844 23264
rect 3804 23202 3832 23258
rect 3712 23174 3832 23202
rect 3884 23248 3936 23254
rect 3884 23190 3936 23196
rect 4436 23248 4488 23254
rect 4436 23190 4488 23196
rect 3712 22574 3740 23174
rect 3792 23044 3844 23050
rect 3792 22986 3844 22992
rect 3700 22568 3752 22574
rect 3700 22510 3752 22516
rect 3804 22506 3832 22986
rect 3792 22500 3844 22506
rect 3792 22442 3844 22448
rect 3896 22030 3924 23190
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 3988 22710 4016 23054
rect 4448 22710 4476 23190
rect 4528 23180 4580 23186
rect 4528 23122 4580 23128
rect 4540 22964 4568 23122
rect 4632 23118 4660 23734
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 4540 22936 4660 22964
rect 3976 22704 4028 22710
rect 3976 22646 4028 22652
rect 4436 22704 4488 22710
rect 4436 22646 4488 22652
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4436 22228 4488 22234
rect 4436 22170 4488 22176
rect 3884 22024 3936 22030
rect 3884 21966 3936 21972
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 4342 21992 4398 22001
rect 3792 21956 3844 21962
rect 3792 21898 3844 21904
rect 3700 21888 3752 21894
rect 3700 21830 3752 21836
rect 3514 21720 3570 21729
rect 3514 21655 3570 21664
rect 3516 21616 3568 21622
rect 3568 21576 3648 21604
rect 3516 21558 3568 21564
rect 3620 21350 3648 21576
rect 3516 21344 3568 21350
rect 3516 21286 3568 21292
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 3422 21040 3478 21049
rect 3422 20975 3478 20984
rect 3424 20800 3476 20806
rect 3424 20742 3476 20748
rect 3330 20496 3386 20505
rect 3240 20460 3292 20466
rect 3330 20431 3386 20440
rect 3240 20402 3292 20408
rect 3148 20324 3200 20330
rect 3148 20266 3200 20272
rect 2964 19984 3016 19990
rect 2964 19926 3016 19932
rect 3160 19854 3188 20266
rect 3252 19854 3280 20402
rect 3332 20256 3384 20262
rect 3332 20198 3384 20204
rect 2596 19848 2648 19854
rect 2502 19816 2558 19825
rect 2320 19780 2372 19786
rect 2596 19790 2648 19796
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3240 19848 3292 19854
rect 3240 19790 3292 19796
rect 2502 19751 2558 19760
rect 2320 19722 2372 19728
rect 2412 19712 2464 19718
rect 2412 19654 2464 19660
rect 2424 16674 2452 19654
rect 2148 16510 2268 16538
rect 2332 16646 2452 16674
rect 2042 16280 2098 16289
rect 2042 16215 2098 16224
rect 2056 13138 2084 16215
rect 2148 13410 2176 16510
rect 2228 16448 2280 16454
rect 2228 16390 2280 16396
rect 2240 15026 2268 16390
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 2332 13433 2360 16646
rect 2412 16516 2464 16522
rect 2412 16458 2464 16464
rect 2424 15026 2452 16458
rect 2516 15434 2544 19751
rect 2870 19544 2926 19553
rect 2780 19508 2832 19514
rect 2870 19479 2926 19488
rect 2780 19450 2832 19456
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2608 16522 2636 18362
rect 2688 18284 2740 18290
rect 2688 18226 2740 18232
rect 2700 17882 2728 18226
rect 2688 17876 2740 17882
rect 2688 17818 2740 17824
rect 2700 17542 2728 17818
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2686 17232 2742 17241
rect 2686 17167 2688 17176
rect 2740 17167 2742 17176
rect 2688 17138 2740 17144
rect 2688 17060 2740 17066
rect 2688 17002 2740 17008
rect 2700 16590 2728 17002
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2700 16114 2728 16526
rect 2792 16266 2820 19450
rect 2884 18358 2912 19479
rect 3148 19168 3200 19174
rect 3148 19110 3200 19116
rect 2872 18352 2924 18358
rect 2872 18294 2924 18300
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 3068 16590 3096 18226
rect 3160 17678 3188 19110
rect 3344 18766 3372 20198
rect 3436 18766 3464 20742
rect 3528 20534 3556 21286
rect 3620 21010 3648 21286
rect 3608 21004 3660 21010
rect 3608 20946 3660 20952
rect 3712 20874 3740 21830
rect 3804 21690 3832 21898
rect 3792 21684 3844 21690
rect 3792 21626 3844 21632
rect 3790 21448 3846 21457
rect 3790 21383 3846 21392
rect 3804 20942 3832 21383
rect 3792 20936 3844 20942
rect 3792 20878 3844 20884
rect 3700 20868 3752 20874
rect 3700 20810 3752 20816
rect 3516 20528 3568 20534
rect 3516 20470 3568 20476
rect 3608 19236 3660 19242
rect 3608 19178 3660 19184
rect 3332 18760 3384 18766
rect 3332 18702 3384 18708
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3514 18728 3570 18737
rect 3514 18663 3570 18672
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3344 18290 3372 18566
rect 3528 18426 3556 18663
rect 3620 18630 3648 19178
rect 3608 18624 3660 18630
rect 3608 18566 3660 18572
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3332 18284 3384 18290
rect 3332 18226 3384 18232
rect 3148 17672 3200 17678
rect 3148 17614 3200 17620
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 3160 17241 3188 17478
rect 3252 17338 3280 17478
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 3146 17232 3202 17241
rect 3146 17167 3202 17176
rect 3160 16998 3188 17167
rect 3148 16992 3200 16998
rect 3148 16934 3200 16940
rect 3252 16794 3280 17274
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 2792 16238 2912 16266
rect 2976 16250 3004 16526
rect 3240 16448 3292 16454
rect 3054 16416 3110 16425
rect 3240 16390 3292 16396
rect 3054 16351 3110 16360
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 2778 16008 2834 16017
rect 2778 15943 2834 15952
rect 2504 15428 2556 15434
rect 2504 15370 2556 15376
rect 2502 15328 2558 15337
rect 2502 15263 2558 15272
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 2516 13920 2544 15263
rect 2792 15178 2820 15943
rect 2424 13892 2544 13920
rect 2608 15150 2820 15178
rect 2318 13424 2374 13433
rect 2148 13382 2268 13410
rect 2056 13110 2176 13138
rect 2148 12434 2176 13110
rect 2056 12406 2176 12434
rect 1860 11620 1912 11626
rect 1860 11562 1912 11568
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10985 1440 11086
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1308 5364 1360 5370
rect 1308 5306 1360 5312
rect 2056 5137 2084 12406
rect 2240 12186 2268 13382
rect 2318 13359 2374 13368
rect 2424 12434 2452 13892
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2516 13326 2544 13670
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2516 12986 2544 13262
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2148 12158 2268 12186
rect 2332 12406 2452 12434
rect 2148 11762 2176 12158
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2148 11150 2176 11698
rect 2240 11150 2268 12038
rect 2136 11144 2188 11150
rect 2228 11144 2280 11150
rect 2136 11086 2188 11092
rect 2226 11112 2228 11121
rect 2280 11112 2282 11121
rect 2226 11047 2282 11056
rect 2332 5681 2360 12406
rect 2608 11778 2636 15150
rect 2688 13796 2740 13802
rect 2688 13738 2740 13744
rect 2424 11750 2636 11778
rect 2318 5672 2374 5681
rect 2318 5607 2374 5616
rect 2042 5128 2098 5137
rect 2042 5063 2098 5072
rect 1124 4276 1176 4282
rect 1124 4218 1176 4224
rect 2424 4146 2452 11750
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 11218 2544 11494
rect 2700 11370 2728 13738
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2792 12306 2820 13330
rect 2884 13326 2912 16238
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 2964 16108 3016 16114
rect 2964 16050 3016 16056
rect 2976 15026 3004 16050
rect 3068 15473 3096 16351
rect 3148 16040 3200 16046
rect 3252 16017 3280 16390
rect 3148 15982 3200 15988
rect 3238 16008 3294 16017
rect 3054 15464 3110 15473
rect 3054 15399 3110 15408
rect 3054 15192 3110 15201
rect 3054 15127 3056 15136
rect 3108 15127 3110 15136
rect 3056 15098 3108 15104
rect 3160 15026 3188 15982
rect 3238 15943 3294 15952
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 3054 13832 3110 13841
rect 3054 13767 3110 13776
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2964 13252 3016 13258
rect 2964 13194 3016 13200
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2872 12232 2924 12238
rect 2976 12209 3004 13194
rect 3068 12442 3096 13767
rect 3160 13297 3188 13874
rect 3252 13530 3280 14418
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 3146 13288 3202 13297
rect 3146 13223 3202 13232
rect 3146 13152 3202 13161
rect 3146 13087 3202 13096
rect 3160 12714 3188 13087
rect 3252 12850 3280 13466
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3240 12708 3292 12714
rect 3240 12650 3292 12656
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 2872 12174 2924 12180
rect 2962 12200 3018 12209
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2792 11558 2820 12106
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2884 11370 2912 12174
rect 2962 12135 3018 12144
rect 2964 12096 3016 12102
rect 3068 12084 3096 12242
rect 3016 12056 3096 12084
rect 2964 12038 3016 12044
rect 2976 11558 3004 12038
rect 3056 11620 3108 11626
rect 3056 11562 3108 11568
rect 3148 11620 3200 11626
rect 3148 11562 3200 11568
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2608 11342 2728 11370
rect 2792 11342 2912 11370
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2504 11008 2556 11014
rect 2504 10950 2556 10956
rect 2516 9081 2544 10950
rect 2502 9072 2558 9081
rect 2502 9007 2558 9016
rect 2608 6254 2636 11342
rect 2688 11076 2740 11082
rect 2792 11064 2820 11342
rect 2872 11280 2924 11286
rect 2870 11248 2872 11257
rect 2924 11248 2926 11257
rect 2870 11183 2926 11192
rect 2872 11144 2924 11150
rect 2740 11036 2820 11064
rect 2870 11112 2872 11121
rect 2924 11112 2926 11121
rect 2870 11047 2926 11056
rect 2688 11018 2740 11024
rect 2792 9586 2820 11036
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2976 8974 3004 11494
rect 3068 11014 3096 11562
rect 3056 11008 3108 11014
rect 3056 10950 3108 10956
rect 3160 10674 3188 11562
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3148 10532 3200 10538
rect 3148 10474 3200 10480
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 3160 8498 3188 10474
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 3252 5234 3280 12650
rect 3344 11762 3372 18226
rect 3528 18222 3556 18362
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3620 18086 3648 18566
rect 3712 18290 3740 20810
rect 3792 20800 3844 20806
rect 3790 20768 3792 20777
rect 3844 20768 3846 20777
rect 3790 20703 3846 20712
rect 3896 20602 3924 21966
rect 3988 21622 4016 21966
rect 4342 21927 4398 21936
rect 4066 21856 4122 21865
rect 4066 21791 4122 21800
rect 3976 21616 4028 21622
rect 3976 21558 4028 21564
rect 4080 21554 4108 21791
rect 4356 21554 4384 21927
rect 4448 21690 4476 22170
rect 4526 22128 4582 22137
rect 4526 22063 4582 22072
rect 4540 22030 4568 22063
rect 4528 22024 4580 22030
rect 4528 21966 4580 21972
rect 4528 21888 4580 21894
rect 4526 21856 4528 21865
rect 4580 21856 4582 21865
rect 4526 21791 4582 21800
rect 4436 21684 4488 21690
rect 4436 21626 4488 21632
rect 4068 21548 4120 21554
rect 4068 21490 4120 21496
rect 4344 21548 4396 21554
rect 4344 21490 4396 21496
rect 3976 21480 4028 21486
rect 3976 21422 4028 21428
rect 4250 21448 4306 21457
rect 3884 20596 3936 20602
rect 3884 20538 3936 20544
rect 3790 20496 3846 20505
rect 3790 20431 3846 20440
rect 3804 20262 3832 20431
rect 3792 20256 3844 20262
rect 3792 20198 3844 20204
rect 3804 19514 3832 20198
rect 3988 20058 4016 21422
rect 4250 21383 4306 21392
rect 4264 21350 4292 21383
rect 4068 21344 4120 21350
rect 4068 21286 4120 21292
rect 4252 21344 4304 21350
rect 4252 21286 4304 21292
rect 4080 20398 4108 21286
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4436 21140 4488 21146
rect 4436 21082 4488 21088
rect 4344 21072 4396 21078
rect 4250 21040 4306 21049
rect 4344 21014 4396 21020
rect 4250 20975 4306 20984
rect 4264 20942 4292 20975
rect 4356 20942 4384 21014
rect 4252 20936 4304 20942
rect 4252 20878 4304 20884
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 4264 20244 4292 20878
rect 4448 20466 4476 21082
rect 4436 20460 4488 20466
rect 4436 20402 4488 20408
rect 4080 20216 4292 20244
rect 3976 20052 4028 20058
rect 4080 20040 4108 20216
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4080 20012 4200 20040
rect 3976 19994 4028 20000
rect 3884 19984 3936 19990
rect 3884 19926 3936 19932
rect 3792 19508 3844 19514
rect 3792 19450 3844 19456
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 3608 18080 3660 18086
rect 3608 18022 3660 18028
rect 3700 18080 3752 18086
rect 3700 18022 3752 18028
rect 3422 17912 3478 17921
rect 3422 17847 3478 17856
rect 3436 17678 3464 17847
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3620 17184 3648 18022
rect 3712 17746 3740 18022
rect 3700 17740 3752 17746
rect 3700 17682 3752 17688
rect 3700 17604 3752 17610
rect 3700 17546 3752 17552
rect 3436 17156 3648 17184
rect 3436 13818 3464 17156
rect 3712 17082 3740 17546
rect 3620 17054 3740 17082
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3528 13938 3556 16730
rect 3620 16658 3648 17054
rect 3700 16992 3752 16998
rect 3700 16934 3752 16940
rect 3608 16652 3660 16658
rect 3608 16594 3660 16600
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3620 13818 3648 15846
rect 3712 13938 3740 16934
rect 3804 15570 3832 18566
rect 3896 17202 3924 19926
rect 4068 19780 4120 19786
rect 3988 19740 4068 19768
rect 3988 19310 4016 19740
rect 4068 19722 4120 19728
rect 4066 19680 4122 19689
rect 4066 19615 4122 19624
rect 4080 19378 4108 19615
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3988 17270 4016 19246
rect 4172 19224 4200 20012
rect 4344 19508 4396 19514
rect 4344 19450 4396 19456
rect 4356 19334 4384 19450
rect 4632 19446 4660 22936
rect 4724 22506 4752 23734
rect 4816 23662 4844 24074
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5276 23848 5304 24239
rect 5092 23820 5304 23848
rect 4804 23656 4856 23662
rect 4804 23598 4856 23604
rect 5092 23526 5120 23820
rect 5368 23730 5396 24262
rect 5448 24200 5500 24206
rect 5448 24142 5500 24148
rect 5460 23866 5488 24142
rect 5552 24138 5580 24822
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 5644 24342 5672 24754
rect 5632 24336 5684 24342
rect 5632 24278 5684 24284
rect 5540 24132 5592 24138
rect 5540 24074 5592 24080
rect 5736 24041 5764 25894
rect 5908 25842 5960 25848
rect 5816 25832 5868 25838
rect 5816 25774 5868 25780
rect 5828 25294 5856 25774
rect 5920 25673 5948 25842
rect 5906 25664 5962 25673
rect 5906 25599 5962 25608
rect 5816 25288 5868 25294
rect 5816 25230 5868 25236
rect 5828 25158 5856 25230
rect 5816 25152 5868 25158
rect 5816 25094 5868 25100
rect 5828 24818 5856 25094
rect 6012 24954 6040 26726
rect 6196 26625 6224 26846
rect 6182 26616 6238 26625
rect 6182 26551 6238 26560
rect 6196 26518 6224 26551
rect 6184 26512 6236 26518
rect 6184 26454 6236 26460
rect 6184 26376 6236 26382
rect 6184 26318 6236 26324
rect 6196 26246 6224 26318
rect 6184 26240 6236 26246
rect 6090 26208 6146 26217
rect 6184 26182 6236 26188
rect 6090 26143 6146 26152
rect 6104 25906 6132 26143
rect 6092 25900 6144 25906
rect 6092 25842 6144 25848
rect 6104 25430 6132 25842
rect 6196 25498 6224 26182
rect 6184 25492 6236 25498
rect 6184 25434 6236 25440
rect 6092 25424 6144 25430
rect 6092 25366 6144 25372
rect 6196 25294 6224 25434
rect 6184 25288 6236 25294
rect 6184 25230 6236 25236
rect 6000 24948 6052 24954
rect 6000 24890 6052 24896
rect 5816 24812 5868 24818
rect 5816 24754 5868 24760
rect 6092 24812 6144 24818
rect 6092 24754 6144 24760
rect 6184 24812 6236 24818
rect 6184 24754 6236 24760
rect 5908 24676 5960 24682
rect 5908 24618 5960 24624
rect 6000 24676 6052 24682
rect 6000 24618 6052 24624
rect 5920 24290 5948 24618
rect 5828 24262 5948 24290
rect 5722 24032 5778 24041
rect 5722 23967 5778 23976
rect 5448 23860 5500 23866
rect 5448 23802 5500 23808
rect 5172 23724 5224 23730
rect 5172 23666 5224 23672
rect 5356 23724 5408 23730
rect 5356 23666 5408 23672
rect 4896 23520 4948 23526
rect 4896 23462 4948 23468
rect 5080 23520 5132 23526
rect 5080 23462 5132 23468
rect 4908 23254 4936 23462
rect 5184 23322 5212 23666
rect 5264 23656 5316 23662
rect 5316 23604 5488 23610
rect 5264 23598 5488 23604
rect 5276 23582 5488 23598
rect 5460 23526 5488 23582
rect 5356 23520 5408 23526
rect 5356 23462 5408 23468
rect 5448 23520 5500 23526
rect 5724 23520 5776 23526
rect 5448 23462 5500 23468
rect 5538 23488 5594 23497
rect 5172 23316 5224 23322
rect 5172 23258 5224 23264
rect 5368 23254 5396 23462
rect 4896 23248 4948 23254
rect 5356 23248 5408 23254
rect 4896 23190 4948 23196
rect 4986 23216 5042 23225
rect 5356 23190 5408 23196
rect 4986 23151 5042 23160
rect 5000 23118 5028 23151
rect 5368 23118 5396 23190
rect 4988 23112 5040 23118
rect 4894 23080 4950 23089
rect 4804 23044 4856 23050
rect 4988 23054 5040 23060
rect 5264 23112 5316 23118
rect 5264 23054 5316 23060
rect 5356 23112 5408 23118
rect 5356 23054 5408 23060
rect 4894 23015 4950 23024
rect 4804 22986 4856 22992
rect 4816 22642 4844 22986
rect 4908 22982 4936 23015
rect 4896 22976 4948 22982
rect 4896 22918 4948 22924
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5276 22794 5304 23054
rect 5368 22953 5396 23054
rect 5354 22944 5410 22953
rect 5354 22879 5410 22888
rect 5354 22808 5410 22817
rect 5276 22766 5354 22794
rect 5354 22743 5410 22752
rect 4804 22636 4856 22642
rect 4804 22578 4856 22584
rect 4988 22636 5040 22642
rect 4988 22578 5040 22584
rect 5080 22636 5132 22642
rect 5080 22578 5132 22584
rect 4816 22506 4844 22578
rect 4896 22568 4948 22574
rect 4896 22510 4948 22516
rect 4712 22500 4764 22506
rect 4712 22442 4764 22448
rect 4804 22500 4856 22506
rect 4804 22442 4856 22448
rect 4710 22264 4766 22273
rect 4710 22199 4766 22208
rect 4724 22166 4752 22199
rect 4712 22160 4764 22166
rect 4712 22102 4764 22108
rect 4712 21344 4764 21350
rect 4712 21286 4764 21292
rect 4724 20942 4752 21286
rect 4712 20936 4764 20942
rect 4712 20878 4764 20884
rect 4724 20641 4752 20878
rect 4710 20632 4766 20641
rect 4710 20567 4766 20576
rect 4724 20346 4752 20567
rect 4816 20534 4844 22442
rect 4908 22216 4936 22510
rect 5000 22409 5028 22578
rect 5092 22545 5120 22578
rect 5078 22536 5134 22545
rect 5078 22471 5134 22480
rect 5368 22438 5396 22743
rect 5264 22432 5316 22438
rect 4986 22400 5042 22409
rect 5264 22374 5316 22380
rect 5356 22432 5408 22438
rect 5356 22374 5408 22380
rect 4986 22335 5042 22344
rect 4988 22228 5040 22234
rect 4908 22188 4988 22216
rect 4988 22170 5040 22176
rect 5276 22094 5304 22374
rect 5276 22066 5396 22094
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5276 21554 5304 21830
rect 5264 21548 5316 21554
rect 5264 21490 5316 21496
rect 5368 21457 5396 22066
rect 5460 21978 5488 23462
rect 5724 23462 5776 23468
rect 5538 23423 5594 23432
rect 5552 23066 5580 23423
rect 5552 23038 5672 23066
rect 5540 22976 5592 22982
rect 5540 22918 5592 22924
rect 5552 22234 5580 22918
rect 5540 22228 5592 22234
rect 5540 22170 5592 22176
rect 5644 22030 5672 23038
rect 5736 22545 5764 23462
rect 5722 22536 5778 22545
rect 5722 22471 5778 22480
rect 5724 22228 5776 22234
rect 5724 22170 5776 22176
rect 5632 22024 5684 22030
rect 5538 21992 5594 22001
rect 5460 21950 5538 21978
rect 5632 21966 5684 21972
rect 5538 21927 5594 21936
rect 5632 21684 5684 21690
rect 5632 21626 5684 21632
rect 5540 21480 5592 21486
rect 5354 21448 5410 21457
rect 5080 21412 5132 21418
rect 5540 21422 5592 21428
rect 5354 21383 5410 21392
rect 5080 21354 5132 21360
rect 4894 21176 4950 21185
rect 4894 21111 4896 21120
rect 4948 21111 4950 21120
rect 4988 21140 5040 21146
rect 4896 21082 4948 21088
rect 4988 21082 5040 21088
rect 4908 20874 4936 21082
rect 5000 21010 5028 21082
rect 5092 21010 5120 21354
rect 5356 21344 5408 21350
rect 5356 21286 5408 21292
rect 5448 21344 5500 21350
rect 5552 21332 5580 21422
rect 5644 21400 5672 21626
rect 5736 21554 5764 22170
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5724 21412 5776 21418
rect 5644 21372 5724 21400
rect 5724 21354 5776 21360
rect 5552 21304 5672 21332
rect 5448 21286 5500 21292
rect 4988 21004 5040 21010
rect 4988 20946 5040 20952
rect 5080 21004 5132 21010
rect 5080 20946 5132 20952
rect 5368 20942 5396 21286
rect 5460 20942 5488 21286
rect 5540 21072 5592 21078
rect 5540 21014 5592 21020
rect 5552 20942 5580 21014
rect 5356 20936 5408 20942
rect 5448 20936 5500 20942
rect 5356 20878 5408 20884
rect 5446 20904 5448 20913
rect 5540 20936 5592 20942
rect 5500 20904 5502 20913
rect 4896 20868 4948 20874
rect 4896 20810 4948 20816
rect 5264 20800 5316 20806
rect 5264 20742 5316 20748
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4804 20528 4856 20534
rect 4804 20470 4856 20476
rect 4802 20360 4858 20369
rect 4724 20318 4802 20346
rect 4802 20295 4858 20304
rect 4896 20052 4948 20058
rect 4896 19994 4948 20000
rect 4908 19854 4936 19994
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4804 19780 4856 19786
rect 4724 19740 4804 19768
rect 4724 19553 4752 19740
rect 4804 19722 4856 19728
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4710 19544 4766 19553
rect 4874 19547 5182 19556
rect 4710 19479 4766 19488
rect 4620 19440 4672 19446
rect 4620 19382 4672 19388
rect 5080 19372 5132 19378
rect 4356 19306 4752 19334
rect 5080 19314 5132 19320
rect 4172 19196 4660 19224
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 4080 18766 4108 19110
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4344 18828 4396 18834
rect 4344 18770 4396 18776
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 3976 17264 4028 17270
rect 3976 17206 4028 17212
rect 3884 17196 3936 17202
rect 3884 17138 3936 17144
rect 4080 17116 4108 18702
rect 4356 18290 4384 18770
rect 4632 18426 4660 19196
rect 4724 18834 4752 19306
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4816 18766 4844 19110
rect 5092 18834 5120 19314
rect 5080 18828 5132 18834
rect 5080 18770 5132 18776
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4620 18420 4672 18426
rect 4816 18408 4844 18702
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4816 18380 5028 18408
rect 4620 18362 4672 18368
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4896 18284 4948 18290
rect 4896 18226 4948 18232
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17762 4660 18226
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4540 17734 4660 17762
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4172 17270 4200 17614
rect 4252 17604 4304 17610
rect 4252 17546 4304 17552
rect 4160 17264 4212 17270
rect 4160 17206 4212 17212
rect 4264 17202 4292 17546
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 3882 17096 3938 17105
rect 3882 17031 3884 17040
rect 3936 17031 3938 17040
rect 3988 17088 4108 17116
rect 3884 17002 3936 17008
rect 3882 16552 3938 16561
rect 3882 16487 3938 16496
rect 3896 15706 3924 16487
rect 3884 15700 3936 15706
rect 3884 15642 3936 15648
rect 3882 15600 3938 15609
rect 3792 15564 3844 15570
rect 3882 15535 3938 15544
rect 3792 15506 3844 15512
rect 3896 15502 3924 15535
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 3884 15156 3936 15162
rect 3884 15098 3936 15104
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3804 14822 3832 14962
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3804 14385 3832 14758
rect 3896 14618 3924 15098
rect 3988 14958 4016 17088
rect 4540 16980 4568 17734
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4632 17542 4660 17614
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4632 17202 4660 17478
rect 4724 17270 4752 18158
rect 4802 17776 4858 17785
rect 4802 17711 4858 17720
rect 4712 17264 4764 17270
rect 4712 17206 4764 17212
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 4540 16952 4660 16980
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16776 4660 16952
rect 4540 16748 4660 16776
rect 4436 16720 4488 16726
rect 4436 16662 4488 16668
rect 4342 16552 4398 16561
rect 4342 16487 4398 16496
rect 4356 16114 4384 16487
rect 4448 16250 4476 16662
rect 4540 16658 4568 16748
rect 4724 16674 4752 17206
rect 4816 17202 4844 17711
rect 4908 17678 4936 18226
rect 5000 17746 5028 18380
rect 4988 17740 5040 17746
rect 4988 17682 5040 17688
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 5170 17096 5226 17105
rect 4988 17060 5040 17066
rect 5170 17031 5226 17040
rect 4988 17002 5040 17008
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 4632 16646 4752 16674
rect 5000 16658 5028 17002
rect 4988 16652 5040 16658
rect 4632 16590 4660 16646
rect 4988 16594 5040 16600
rect 5184 16590 5212 17031
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 4528 16516 4580 16522
rect 4528 16458 4580 16464
rect 4540 16250 4568 16458
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4528 16244 4580 16250
rect 4528 16186 4580 16192
rect 4448 16130 4476 16186
rect 4344 16108 4396 16114
rect 4448 16102 4660 16130
rect 4344 16050 4396 16056
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4434 15600 4490 15609
rect 4434 15535 4490 15544
rect 4068 15360 4120 15366
rect 4448 15337 4476 15535
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 4068 15302 4120 15308
rect 4434 15328 4490 15337
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 3882 14512 3938 14521
rect 3882 14447 3938 14456
rect 3790 14376 3846 14385
rect 3790 14311 3846 14320
rect 3896 13938 3924 14447
rect 3988 14414 4016 14758
rect 4080 14618 4108 15302
rect 4434 15263 4490 15272
rect 4540 14822 4568 15438
rect 4632 15026 4660 16102
rect 4724 15978 4752 16390
rect 4712 15972 4764 15978
rect 4712 15914 4764 15920
rect 4724 15094 4752 15914
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 4816 15026 4844 16390
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 5184 15881 5212 16050
rect 5170 15872 5226 15881
rect 5170 15807 5226 15816
rect 5276 15502 5304 20742
rect 5368 20330 5396 20878
rect 5540 20878 5592 20884
rect 5446 20839 5502 20848
rect 5448 20460 5500 20466
rect 5448 20402 5500 20408
rect 5356 20324 5408 20330
rect 5356 20266 5408 20272
rect 5460 20262 5488 20402
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 5460 19990 5488 20198
rect 5448 19984 5500 19990
rect 5448 19926 5500 19932
rect 5356 19848 5408 19854
rect 5356 19790 5408 19796
rect 5368 19428 5396 19790
rect 5460 19786 5488 19926
rect 5448 19780 5500 19786
rect 5448 19722 5500 19728
rect 5368 19400 5414 19428
rect 5386 19292 5414 19400
rect 5368 19264 5414 19292
rect 5368 18737 5396 19264
rect 5552 19224 5580 20878
rect 5644 20466 5672 21304
rect 5724 20800 5776 20806
rect 5724 20742 5776 20748
rect 5736 20505 5764 20742
rect 5722 20496 5778 20505
rect 5632 20460 5684 20466
rect 5722 20431 5778 20440
rect 5632 20402 5684 20408
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5460 19196 5580 19224
rect 5460 18766 5488 19196
rect 5538 19136 5594 19145
rect 5538 19071 5594 19080
rect 5448 18760 5500 18766
rect 5354 18728 5410 18737
rect 5448 18702 5500 18708
rect 5354 18663 5410 18672
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5368 18358 5396 18566
rect 5356 18352 5408 18358
rect 5356 18294 5408 18300
rect 5460 18204 5488 18702
rect 5368 18176 5488 18204
rect 5368 17882 5396 18176
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 5448 17808 5500 17814
rect 5448 17750 5500 17756
rect 5356 17536 5408 17542
rect 5356 17478 5408 17484
rect 5368 16590 5396 17478
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4620 15020 4672 15026
rect 4620 14962 4672 14968
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3700 13932 3752 13938
rect 3700 13874 3752 13880
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3976 13864 4028 13870
rect 3436 13790 3556 13818
rect 3620 13790 3924 13818
rect 3976 13806 4028 13812
rect 3424 13456 3476 13462
rect 3424 13398 3476 13404
rect 3436 12238 3464 13398
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3528 12186 3556 13790
rect 3700 13728 3752 13734
rect 3700 13670 3752 13676
rect 3712 13326 3740 13670
rect 3700 13320 3752 13326
rect 3752 13280 3832 13308
rect 3700 13262 3752 13268
rect 3700 13184 3752 13190
rect 3700 13126 3752 13132
rect 3606 12880 3662 12889
rect 3606 12815 3608 12824
rect 3660 12815 3662 12824
rect 3608 12786 3660 12792
rect 3712 12238 3740 13126
rect 3804 13025 3832 13280
rect 3790 13016 3846 13025
rect 3790 12951 3846 12960
rect 3896 12850 3924 13790
rect 3988 13530 4016 13806
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 3988 13326 4016 13466
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3804 12646 3832 12786
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 4080 12434 4108 14554
rect 4632 14482 4660 14962
rect 4712 14952 4764 14958
rect 4988 14952 5040 14958
rect 4764 14900 4844 14906
rect 4712 14894 4844 14900
rect 4988 14894 5040 14900
rect 4724 14878 4844 14894
rect 4710 14648 4766 14657
rect 4710 14583 4712 14592
rect 4764 14583 4766 14592
rect 4712 14554 4764 14560
rect 4816 14498 4844 14878
rect 4896 14816 4948 14822
rect 4894 14784 4896 14793
rect 4948 14784 4950 14793
rect 4894 14719 4950 14728
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4724 14470 4844 14498
rect 4250 14376 4306 14385
rect 4250 14311 4306 14320
rect 4264 13734 4292 14311
rect 4724 14074 4752 14470
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4252 13728 4304 13734
rect 4252 13670 4304 13676
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4434 13424 4490 13433
rect 4434 13359 4436 13368
rect 4488 13359 4490 13368
rect 4436 13330 4488 13336
rect 4344 13320 4396 13326
rect 4342 13288 4344 13297
rect 4396 13288 4398 13297
rect 4342 13223 4398 13232
rect 4356 13190 4384 13223
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4540 12850 4568 13466
rect 4632 13326 4660 14010
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4724 13462 4752 13670
rect 4816 13569 4844 14350
rect 5000 14346 5028 14894
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 5092 14346 5120 14758
rect 4988 14340 5040 14346
rect 4988 14282 5040 14288
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 4896 13864 4948 13870
rect 4894 13832 4896 13841
rect 4948 13832 4950 13841
rect 4894 13767 4950 13776
rect 4802 13560 4858 13569
rect 4802 13495 4858 13504
rect 5000 13462 5028 13874
rect 4712 13456 4764 13462
rect 4988 13456 5040 13462
rect 4764 13416 4844 13444
rect 4712 13398 4764 13404
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4080 12406 4200 12434
rect 3792 12368 3844 12374
rect 3792 12310 3844 12316
rect 3700 12232 3752 12238
rect 3528 12158 3648 12186
rect 3700 12174 3752 12180
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3528 11898 3556 12038
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3528 11762 3556 11834
rect 3620 11762 3648 12158
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 3344 11150 3372 11494
rect 3436 11286 3464 11630
rect 3516 11620 3568 11626
rect 3516 11562 3568 11568
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3528 11150 3556 11562
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3344 9926 3372 11086
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3344 9466 3372 9862
rect 3528 9586 3556 11086
rect 3620 10810 3648 11290
rect 3712 11082 3740 12174
rect 3700 11076 3752 11082
rect 3700 11018 3752 11024
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3620 9654 3648 9998
rect 3608 9648 3660 9654
rect 3608 9590 3660 9596
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3424 9512 3476 9518
rect 3344 9460 3424 9466
rect 3344 9454 3476 9460
rect 3344 9438 3464 9454
rect 3528 8906 3556 9522
rect 3712 9466 3740 10610
rect 3804 10044 3832 12310
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4080 11558 4108 12174
rect 4172 11665 4200 12406
rect 4342 11928 4398 11937
rect 4342 11863 4344 11872
rect 4396 11863 4398 11872
rect 4344 11834 4396 11840
rect 4436 11756 4488 11762
rect 4632 11744 4660 13126
rect 4710 13016 4766 13025
rect 4710 12951 4766 12960
rect 4488 11716 4660 11744
rect 4724 11744 4752 12951
rect 4816 11880 4844 13416
rect 4988 13398 5040 13404
rect 4894 13288 4950 13297
rect 4894 13223 4896 13232
rect 4948 13223 4950 13232
rect 4896 13194 4948 13200
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5276 12850 5304 15438
rect 5368 13938 5396 16526
rect 5460 15094 5488 17750
rect 5552 17678 5580 19071
rect 5736 18698 5764 19790
rect 5724 18692 5776 18698
rect 5724 18634 5776 18640
rect 5630 18456 5686 18465
rect 5630 18391 5686 18400
rect 5644 18290 5672 18391
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5552 16590 5580 17274
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5644 16522 5672 17478
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 5736 16590 5764 17138
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 5632 16516 5684 16522
rect 5632 16458 5684 16464
rect 5538 16416 5594 16425
rect 5538 16351 5594 16360
rect 5552 15706 5580 16351
rect 5644 15745 5672 16458
rect 5828 16182 5856 24262
rect 6012 24206 6040 24618
rect 6104 24206 6132 24754
rect 6196 24410 6224 24754
rect 6184 24404 6236 24410
rect 6184 24346 6236 24352
rect 6000 24200 6052 24206
rect 5906 24168 5962 24177
rect 6000 24142 6052 24148
rect 6092 24200 6144 24206
rect 6092 24142 6144 24148
rect 5906 24103 5962 24112
rect 5920 23866 5948 24103
rect 6184 24064 6236 24070
rect 5998 24032 6054 24041
rect 6184 24006 6236 24012
rect 5998 23967 6054 23976
rect 5908 23860 5960 23866
rect 5908 23802 5960 23808
rect 5920 23730 5948 23802
rect 5908 23724 5960 23730
rect 5908 23666 5960 23672
rect 5906 23488 5962 23497
rect 5906 23423 5962 23432
rect 5920 23322 5948 23423
rect 5908 23316 5960 23322
rect 5908 23258 5960 23264
rect 5906 23080 5962 23089
rect 5906 23015 5962 23024
rect 5920 22982 5948 23015
rect 5908 22976 5960 22982
rect 5908 22918 5960 22924
rect 5908 22636 5960 22642
rect 5908 22578 5960 22584
rect 5920 22273 5948 22578
rect 5906 22264 5962 22273
rect 5906 22199 5962 22208
rect 5908 22160 5960 22166
rect 5906 22128 5908 22137
rect 5960 22128 5962 22137
rect 5906 22063 5962 22072
rect 5920 21962 5948 22063
rect 6012 22030 6040 23967
rect 6090 23352 6146 23361
rect 6090 23287 6146 23296
rect 6104 23118 6132 23287
rect 6196 23118 6224 24006
rect 6092 23112 6144 23118
rect 6092 23054 6144 23060
rect 6184 23112 6236 23118
rect 6184 23054 6236 23060
rect 6090 22808 6146 22817
rect 6090 22743 6146 22752
rect 6104 22710 6132 22743
rect 6092 22704 6144 22710
rect 6092 22646 6144 22652
rect 6288 22642 6316 27270
rect 6380 26897 6408 27406
rect 6460 27396 6512 27402
rect 6460 27338 6512 27344
rect 6472 27130 6500 27338
rect 6460 27124 6512 27130
rect 6460 27066 6512 27072
rect 6564 26994 6592 27542
rect 6656 27130 6684 28018
rect 6734 27704 6790 27713
rect 6734 27639 6790 27648
rect 6644 27124 6696 27130
rect 6644 27066 6696 27072
rect 6748 27010 6776 27639
rect 6840 27441 6868 30359
rect 10692 30048 10744 30054
rect 10692 29990 10744 29996
rect 8852 29844 8904 29850
rect 8852 29786 8904 29792
rect 9864 29844 9916 29850
rect 9864 29786 9916 29792
rect 7196 29776 7248 29782
rect 7196 29718 7248 29724
rect 7012 29640 7064 29646
rect 7012 29582 7064 29588
rect 6918 28792 6974 28801
rect 6918 28727 6974 28736
rect 6932 27878 6960 28727
rect 6920 27872 6972 27878
rect 6920 27814 6972 27820
rect 7024 27577 7052 29582
rect 7208 29170 7236 29718
rect 7470 29608 7526 29617
rect 7470 29543 7526 29552
rect 7484 29170 7512 29543
rect 8864 29170 8892 29786
rect 9404 29776 9456 29782
rect 9404 29718 9456 29724
rect 9678 29744 9734 29753
rect 9128 29572 9180 29578
rect 9128 29514 9180 29520
rect 9140 29306 9168 29514
rect 9128 29300 9180 29306
rect 9128 29242 9180 29248
rect 9036 29232 9088 29238
rect 9140 29209 9168 29242
rect 9036 29174 9088 29180
rect 9126 29200 9182 29209
rect 7196 29164 7248 29170
rect 7196 29106 7248 29112
rect 7472 29164 7524 29170
rect 7472 29106 7524 29112
rect 7564 29164 7616 29170
rect 7564 29106 7616 29112
rect 8024 29164 8076 29170
rect 8024 29106 8076 29112
rect 8852 29164 8904 29170
rect 8852 29106 8904 29112
rect 7104 28960 7156 28966
rect 7104 28902 7156 28908
rect 7116 28558 7144 28902
rect 7104 28552 7156 28558
rect 7196 28552 7248 28558
rect 7104 28494 7156 28500
rect 7194 28520 7196 28529
rect 7248 28520 7250 28529
rect 7116 28014 7144 28494
rect 7194 28455 7250 28464
rect 7196 28416 7248 28422
rect 7194 28384 7196 28393
rect 7472 28416 7524 28422
rect 7248 28384 7250 28393
rect 7472 28358 7524 28364
rect 7194 28319 7250 28328
rect 7208 28218 7236 28319
rect 7196 28212 7248 28218
rect 7196 28154 7248 28160
rect 7484 28082 7512 28358
rect 7576 28150 7604 29106
rect 8036 28762 8064 29106
rect 8668 29096 8720 29102
rect 8668 29038 8720 29044
rect 8392 29028 8444 29034
rect 8392 28970 8444 28976
rect 8208 28960 8260 28966
rect 8208 28902 8260 28908
rect 8024 28756 8076 28762
rect 8024 28698 8076 28704
rect 8220 28558 8248 28902
rect 8208 28552 8260 28558
rect 8208 28494 8260 28500
rect 8300 28552 8352 28558
rect 8300 28494 8352 28500
rect 7748 28416 7800 28422
rect 7748 28358 7800 28364
rect 7564 28144 7616 28150
rect 7564 28086 7616 28092
rect 7760 28082 7788 28358
rect 7196 28076 7248 28082
rect 7196 28018 7248 28024
rect 7472 28076 7524 28082
rect 7472 28018 7524 28024
rect 7748 28076 7800 28082
rect 7748 28018 7800 28024
rect 8024 28076 8076 28082
rect 8024 28018 8076 28024
rect 7104 28008 7156 28014
rect 7104 27950 7156 27956
rect 7010 27568 7066 27577
rect 7010 27503 7066 27512
rect 6920 27464 6972 27470
rect 6826 27432 6882 27441
rect 7208 27441 7236 28018
rect 7484 27849 7512 28018
rect 7564 28008 7616 28014
rect 7760 27985 7788 28018
rect 7564 27950 7616 27956
rect 7746 27976 7802 27985
rect 7470 27840 7526 27849
rect 7470 27775 7526 27784
rect 7288 27668 7340 27674
rect 7288 27610 7340 27616
rect 7380 27668 7432 27674
rect 7380 27610 7432 27616
rect 6920 27406 6972 27412
rect 7194 27432 7250 27441
rect 6826 27367 6882 27376
rect 6826 27160 6882 27169
rect 6826 27095 6882 27104
rect 6552 26988 6604 26994
rect 6552 26930 6604 26936
rect 6656 26982 6776 27010
rect 6366 26888 6422 26897
rect 6366 26823 6422 26832
rect 6368 26512 6420 26518
rect 6368 26454 6420 26460
rect 6380 25906 6408 26454
rect 6460 26376 6512 26382
rect 6460 26318 6512 26324
rect 6368 25900 6420 25906
rect 6368 25842 6420 25848
rect 6472 25362 6500 26318
rect 6564 26042 6592 26930
rect 6656 26246 6684 26982
rect 6840 26926 6868 27095
rect 6828 26920 6880 26926
rect 6828 26862 6880 26868
rect 6828 26784 6880 26790
rect 6828 26726 6880 26732
rect 6736 26580 6788 26586
rect 6736 26522 6788 26528
rect 6748 26246 6776 26522
rect 6840 26296 6868 26726
rect 6932 26466 6960 27406
rect 7194 27367 7250 27376
rect 7196 27328 7248 27334
rect 7010 27296 7066 27305
rect 7196 27270 7248 27276
rect 7010 27231 7066 27240
rect 7024 27130 7052 27231
rect 7012 27124 7064 27130
rect 7012 27066 7064 27072
rect 7104 27056 7156 27062
rect 7104 26998 7156 27004
rect 7012 26988 7064 26994
rect 7012 26930 7064 26936
rect 7024 26586 7052 26930
rect 7012 26580 7064 26586
rect 7012 26522 7064 26528
rect 6932 26438 7052 26466
rect 6920 26308 6972 26314
rect 6840 26268 6920 26296
rect 6920 26250 6972 26256
rect 6644 26240 6696 26246
rect 6642 26208 6644 26217
rect 6736 26240 6788 26246
rect 6696 26208 6698 26217
rect 6736 26182 6788 26188
rect 6642 26143 6698 26152
rect 6552 26036 6604 26042
rect 6552 25978 6604 25984
rect 6644 26036 6696 26042
rect 6644 25978 6696 25984
rect 6564 25906 6592 25978
rect 6552 25900 6604 25906
rect 6552 25842 6604 25848
rect 6552 25492 6604 25498
rect 6552 25434 6604 25440
rect 6460 25356 6512 25362
rect 6460 25298 6512 25304
rect 6564 25294 6592 25434
rect 6656 25294 6684 25978
rect 6748 25498 6776 26182
rect 6920 25900 6972 25906
rect 6920 25842 6972 25848
rect 6828 25764 6880 25770
rect 6828 25706 6880 25712
rect 6736 25492 6788 25498
rect 6736 25434 6788 25440
rect 6840 25294 6868 25706
rect 6932 25498 6960 25842
rect 6920 25492 6972 25498
rect 6920 25434 6972 25440
rect 6552 25288 6604 25294
rect 6552 25230 6604 25236
rect 6644 25288 6696 25294
rect 6644 25230 6696 25236
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 6460 25152 6512 25158
rect 6460 25094 6512 25100
rect 6826 25120 6882 25129
rect 6366 23760 6422 23769
rect 6366 23695 6368 23704
rect 6420 23695 6422 23704
rect 6368 23666 6420 23672
rect 6366 23624 6422 23633
rect 6366 23559 6368 23568
rect 6420 23559 6422 23568
rect 6368 23530 6420 23536
rect 6276 22636 6328 22642
rect 6276 22578 6328 22584
rect 6092 22500 6144 22506
rect 6092 22442 6144 22448
rect 6000 22024 6052 22030
rect 6000 21966 6052 21972
rect 6104 21962 6132 22442
rect 5908 21956 5960 21962
rect 5908 21898 5960 21904
rect 6092 21956 6144 21962
rect 6092 21898 6144 21904
rect 6104 21604 6132 21898
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 6196 21729 6224 21830
rect 6182 21720 6238 21729
rect 6182 21655 6238 21664
rect 6104 21576 6224 21604
rect 6090 21312 6146 21321
rect 6090 21247 6146 21256
rect 5906 21176 5962 21185
rect 6104 21146 6132 21247
rect 5906 21111 5962 21120
rect 6000 21140 6052 21146
rect 5920 20874 5948 21111
rect 6000 21082 6052 21088
rect 6092 21140 6144 21146
rect 6092 21082 6144 21088
rect 6012 20874 6040 21082
rect 6092 20936 6144 20942
rect 6092 20878 6144 20884
rect 5908 20868 5960 20874
rect 5908 20810 5960 20816
rect 6000 20868 6052 20874
rect 6000 20810 6052 20816
rect 5816 16176 5868 16182
rect 5816 16118 5868 16124
rect 5920 16046 5948 20810
rect 5998 20360 6054 20369
rect 5998 20295 6054 20304
rect 6012 19718 6040 20295
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 6000 19304 6052 19310
rect 6000 19246 6052 19252
rect 6012 16726 6040 19246
rect 6104 18766 6132 20878
rect 6196 18834 6224 21576
rect 6472 21554 6500 25094
rect 6826 25055 6882 25064
rect 6644 24948 6696 24954
rect 6644 24890 6696 24896
rect 6552 24608 6604 24614
rect 6552 24550 6604 24556
rect 6564 24206 6592 24550
rect 6552 24200 6604 24206
rect 6552 24142 6604 24148
rect 6550 24032 6606 24041
rect 6550 23967 6606 23976
rect 6564 23118 6592 23967
rect 6552 23112 6604 23118
rect 6552 23054 6604 23060
rect 6550 22808 6606 22817
rect 6656 22778 6684 24890
rect 6736 24336 6788 24342
rect 6736 24278 6788 24284
rect 6748 24138 6776 24278
rect 6736 24132 6788 24138
rect 6736 24074 6788 24080
rect 6736 23520 6788 23526
rect 6736 23462 6788 23468
rect 6748 23322 6776 23462
rect 6736 23316 6788 23322
rect 6736 23258 6788 23264
rect 6840 23118 6868 25055
rect 6920 24676 6972 24682
rect 6920 24618 6972 24624
rect 6932 24410 6960 24618
rect 6920 24404 6972 24410
rect 6920 24346 6972 24352
rect 6932 24206 6960 24346
rect 7024 24206 7052 26438
rect 7116 26296 7144 26998
rect 7208 26994 7236 27270
rect 7300 27130 7328 27610
rect 7392 27470 7420 27610
rect 7472 27600 7524 27606
rect 7472 27542 7524 27548
rect 7380 27464 7432 27470
rect 7380 27406 7432 27412
rect 7288 27124 7340 27130
rect 7288 27066 7340 27072
rect 7196 26988 7248 26994
rect 7196 26930 7248 26936
rect 7300 26450 7328 27066
rect 7288 26444 7340 26450
rect 7288 26386 7340 26392
rect 7288 26308 7340 26314
rect 7116 26268 7288 26296
rect 7288 26250 7340 26256
rect 7196 25900 7248 25906
rect 7196 25842 7248 25848
rect 7104 25832 7156 25838
rect 7102 25800 7104 25809
rect 7156 25800 7158 25809
rect 7102 25735 7158 25744
rect 7208 25702 7236 25842
rect 7104 25696 7156 25702
rect 7104 25638 7156 25644
rect 7196 25696 7248 25702
rect 7196 25638 7248 25644
rect 7116 24562 7144 25638
rect 7196 24880 7248 24886
rect 7300 24868 7328 26250
rect 7248 24840 7328 24868
rect 7196 24822 7248 24828
rect 7116 24534 7328 24562
rect 6920 24200 6972 24206
rect 6920 24142 6972 24148
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 6920 23724 6972 23730
rect 6920 23666 6972 23672
rect 6932 23254 6960 23666
rect 7300 23474 7328 24534
rect 7392 24206 7420 27406
rect 7484 27130 7512 27542
rect 7472 27124 7524 27130
rect 7472 27066 7524 27072
rect 7472 26988 7524 26994
rect 7472 26930 7524 26936
rect 7484 26246 7512 26930
rect 7472 26240 7524 26246
rect 7472 26182 7524 26188
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7484 23594 7512 24006
rect 7576 23730 7604 27950
rect 7746 27911 7802 27920
rect 7840 27872 7892 27878
rect 7840 27814 7892 27820
rect 7852 27674 7880 27814
rect 8036 27713 8064 28018
rect 8022 27704 8078 27713
rect 7840 27668 7892 27674
rect 8022 27639 8078 27648
rect 7840 27610 7892 27616
rect 7852 27146 7880 27610
rect 8024 27600 8076 27606
rect 8024 27542 8076 27548
rect 7932 27464 7984 27470
rect 7932 27406 7984 27412
rect 7944 27334 7972 27406
rect 7932 27328 7984 27334
rect 7930 27296 7932 27305
rect 7984 27296 7986 27305
rect 7930 27231 7986 27240
rect 7852 27118 7972 27146
rect 7656 26988 7708 26994
rect 7656 26930 7708 26936
rect 7840 26988 7892 26994
rect 7840 26930 7892 26936
rect 7668 26790 7696 26930
rect 7748 26920 7800 26926
rect 7748 26862 7800 26868
rect 7656 26784 7708 26790
rect 7656 26726 7708 26732
rect 7760 26382 7788 26862
rect 7852 26586 7880 26930
rect 7840 26580 7892 26586
rect 7840 26522 7892 26528
rect 7748 26376 7800 26382
rect 7748 26318 7800 26324
rect 7746 26072 7802 26081
rect 7746 26007 7802 26016
rect 7656 25968 7708 25974
rect 7656 25910 7708 25916
rect 7668 24342 7696 25910
rect 7760 24698 7788 26007
rect 7852 24818 7880 26522
rect 7944 25158 7972 27118
rect 7932 25152 7984 25158
rect 7932 25094 7984 25100
rect 7840 24812 7892 24818
rect 7840 24754 7892 24760
rect 7760 24670 7880 24698
rect 7748 24608 7800 24614
rect 7748 24550 7800 24556
rect 7656 24336 7708 24342
rect 7656 24278 7708 24284
rect 7564 23724 7616 23730
rect 7564 23666 7616 23672
rect 7472 23588 7524 23594
rect 7472 23530 7524 23536
rect 7564 23520 7616 23526
rect 7300 23446 7512 23474
rect 7564 23462 7616 23468
rect 7378 23352 7434 23361
rect 7378 23287 7434 23296
rect 6920 23248 6972 23254
rect 6920 23190 6972 23196
rect 7196 23248 7248 23254
rect 7196 23190 7248 23196
rect 7286 23216 7342 23225
rect 6736 23112 6788 23118
rect 6736 23054 6788 23060
rect 6828 23112 6880 23118
rect 6920 23112 6972 23118
rect 6828 23054 6880 23060
rect 6918 23080 6920 23089
rect 6972 23080 6974 23089
rect 6748 22982 6776 23054
rect 6974 23038 7052 23066
rect 6918 23015 6974 23024
rect 6736 22976 6788 22982
rect 6736 22918 6788 22924
rect 6748 22778 6776 22918
rect 6918 22808 6974 22817
rect 6550 22743 6606 22752
rect 6644 22772 6696 22778
rect 6564 22710 6592 22743
rect 6644 22714 6696 22720
rect 6736 22772 6788 22778
rect 6918 22743 6974 22752
rect 6736 22714 6788 22720
rect 6552 22704 6604 22710
rect 6552 22646 6604 22652
rect 6550 22264 6606 22273
rect 6550 22199 6606 22208
rect 6460 21548 6512 21554
rect 6460 21490 6512 21496
rect 6368 21344 6420 21350
rect 6368 21286 6420 21292
rect 6380 20942 6408 21286
rect 6460 21072 6512 21078
rect 6460 21014 6512 21020
rect 6368 20936 6420 20942
rect 6274 20904 6330 20913
rect 6368 20878 6420 20884
rect 6274 20839 6330 20848
rect 6288 20806 6316 20839
rect 6276 20800 6328 20806
rect 6276 20742 6328 20748
rect 6368 20800 6420 20806
rect 6368 20742 6420 20748
rect 6380 20534 6408 20742
rect 6368 20528 6420 20534
rect 6368 20470 6420 20476
rect 6276 20324 6328 20330
rect 6276 20266 6328 20272
rect 6288 19990 6316 20266
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6276 19984 6328 19990
rect 6276 19926 6328 19932
rect 6380 19854 6408 20198
rect 6472 19854 6500 21014
rect 6564 19990 6592 22199
rect 6748 21622 6776 22714
rect 6932 22166 6960 22743
rect 6920 22160 6972 22166
rect 6920 22102 6972 22108
rect 6828 22024 6880 22030
rect 6828 21966 6880 21972
rect 6840 21690 6868 21966
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 6736 21616 6788 21622
rect 6736 21558 6788 21564
rect 6736 21480 6788 21486
rect 6736 21422 6788 21428
rect 6932 21434 6960 22102
rect 7024 21554 7052 23038
rect 7208 23032 7236 23190
rect 7286 23151 7288 23160
rect 7340 23151 7342 23160
rect 7288 23122 7340 23128
rect 7208 23004 7328 23032
rect 7194 22944 7250 22953
rect 7194 22879 7250 22888
rect 7208 22642 7236 22879
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 7196 22432 7248 22438
rect 7196 22374 7248 22380
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 6642 20360 6698 20369
rect 6642 20295 6698 20304
rect 6552 19984 6604 19990
rect 6552 19926 6604 19932
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6460 19848 6512 19854
rect 6460 19790 6512 19796
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 6092 18760 6144 18766
rect 6092 18702 6144 18708
rect 6104 18170 6132 18702
rect 6472 18358 6500 19654
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 6564 18873 6592 19110
rect 6550 18864 6606 18873
rect 6550 18799 6606 18808
rect 6460 18352 6512 18358
rect 6460 18294 6512 18300
rect 6564 18222 6592 18799
rect 6276 18216 6328 18222
rect 6104 18142 6224 18170
rect 6276 18158 6328 18164
rect 6552 18216 6604 18222
rect 6552 18158 6604 18164
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 6104 16590 6132 18022
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 5908 16040 5960 16046
rect 5908 15982 5960 15988
rect 6000 15972 6052 15978
rect 6000 15914 6052 15920
rect 5816 15904 5868 15910
rect 6012 15858 6040 15914
rect 5816 15846 5868 15852
rect 5630 15736 5686 15745
rect 5540 15700 5592 15706
rect 5630 15671 5686 15680
rect 5540 15642 5592 15648
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 5540 14952 5592 14958
rect 5446 14920 5502 14929
rect 5540 14894 5592 14900
rect 5446 14855 5502 14864
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5354 13832 5410 13841
rect 5354 13767 5410 13776
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5078 12744 5134 12753
rect 5368 12730 5396 13767
rect 5460 13190 5488 14855
rect 5552 14618 5580 14894
rect 5540 14612 5592 14618
rect 5644 14600 5672 15438
rect 5724 14952 5776 14958
rect 5722 14920 5724 14929
rect 5776 14920 5778 14929
rect 5722 14855 5778 14864
rect 5724 14612 5776 14618
rect 5644 14572 5724 14600
rect 5540 14554 5592 14560
rect 5724 14554 5776 14560
rect 5630 14512 5686 14521
rect 5630 14447 5686 14456
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 14006 5580 14214
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5448 13184 5500 13190
rect 5552 13161 5580 13942
rect 5644 13870 5672 14447
rect 5736 14385 5764 14554
rect 5828 14414 5856 15846
rect 5920 15830 6040 15858
rect 5920 15201 5948 15830
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 5906 15192 5962 15201
rect 5906 15127 5962 15136
rect 5920 14482 5948 15127
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5816 14408 5868 14414
rect 5722 14376 5778 14385
rect 5816 14350 5868 14356
rect 5722 14311 5778 14320
rect 5828 14278 5856 14350
rect 6012 14346 6040 15642
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 5816 14272 5868 14278
rect 6104 14226 6132 16390
rect 6196 16114 6224 18142
rect 6184 16108 6236 16114
rect 6184 16050 6236 16056
rect 6288 15978 6316 18158
rect 6458 17912 6514 17921
rect 6458 17847 6514 17856
rect 6368 17808 6420 17814
rect 6368 17750 6420 17756
rect 6380 17202 6408 17750
rect 6472 17678 6500 17847
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6472 17270 6500 17478
rect 6564 17338 6592 17614
rect 6656 17377 6684 20295
rect 6748 18834 6776 21422
rect 6932 21406 7052 21434
rect 6920 20528 6972 20534
rect 6826 20496 6882 20505
rect 6920 20470 6972 20476
rect 6826 20431 6882 20440
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6736 18692 6788 18698
rect 6736 18634 6788 18640
rect 6642 17368 6698 17377
rect 6552 17332 6604 17338
rect 6642 17303 6698 17312
rect 6552 17274 6604 17280
rect 6460 17264 6512 17270
rect 6460 17206 6512 17212
rect 6642 17232 6698 17241
rect 6368 17196 6420 17202
rect 6642 17167 6644 17176
rect 6368 17138 6420 17144
rect 6696 17167 6698 17176
rect 6644 17138 6696 17144
rect 6276 15972 6328 15978
rect 6276 15914 6328 15920
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6196 15570 6224 15846
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 5816 14214 5868 14220
rect 5920 14198 6132 14226
rect 5722 14104 5778 14113
rect 5722 14039 5724 14048
rect 5776 14039 5778 14048
rect 5724 14010 5776 14016
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5632 13252 5684 13258
rect 5632 13194 5684 13200
rect 5448 13126 5500 13132
rect 5538 13152 5594 13161
rect 5538 13087 5594 13096
rect 5644 12968 5672 13194
rect 5736 13002 5764 13874
rect 5920 13326 5948 14198
rect 6196 14090 6224 14282
rect 6000 14068 6052 14074
rect 6104 14062 6224 14090
rect 6104 14056 6132 14062
rect 6052 14028 6132 14056
rect 6000 14010 6052 14016
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 5828 13172 5856 13262
rect 5828 13144 5948 13172
rect 5736 12974 5856 13002
rect 5078 12679 5080 12688
rect 5132 12679 5134 12688
rect 5184 12702 5396 12730
rect 5460 12940 5672 12968
rect 5080 12650 5132 12656
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 5000 12238 5028 12378
rect 5080 12368 5132 12374
rect 5080 12310 5132 12316
rect 5092 12238 5120 12310
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 5184 12152 5212 12702
rect 5264 12640 5316 12646
rect 5262 12608 5264 12617
rect 5316 12608 5318 12617
rect 5262 12543 5318 12552
rect 5262 12472 5318 12481
rect 5262 12407 5318 12416
rect 5276 12220 5304 12407
rect 5276 12192 5396 12220
rect 5184 12124 5304 12152
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4816 11852 4936 11880
rect 4804 11756 4856 11762
rect 4724 11716 4804 11744
rect 4436 11698 4488 11704
rect 4804 11698 4856 11704
rect 4158 11656 4214 11665
rect 4158 11591 4214 11600
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3988 10742 4016 10950
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 3988 10198 4016 10678
rect 4080 10266 4108 11494
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4908 11336 4936 11852
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5170 11520 5226 11529
rect 4172 11308 4936 11336
rect 4172 11150 4200 11308
rect 5092 11268 5120 11494
rect 5170 11455 5226 11464
rect 4356 11240 5120 11268
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4264 11082 4292 11154
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4356 10674 4384 11240
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4436 11076 4488 11082
rect 4436 11018 4488 11024
rect 4448 10810 4476 11018
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4434 10704 4490 10713
rect 4344 10668 4396 10674
rect 4434 10639 4490 10648
rect 4344 10610 4396 10616
rect 4448 10538 4476 10639
rect 4436 10532 4488 10538
rect 4436 10474 4488 10480
rect 4540 10470 4568 10950
rect 4632 10810 4660 11086
rect 5184 11014 5212 11455
rect 5276 11082 5304 12124
rect 5368 11898 5396 12192
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5368 11393 5396 11698
rect 5354 11384 5410 11393
rect 5354 11319 5410 11328
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 4712 11008 4764 11014
rect 4896 11008 4948 11014
rect 4712 10950 4764 10956
rect 4816 10968 4896 10996
rect 4724 10849 4752 10950
rect 4710 10840 4766 10849
rect 4620 10804 4672 10810
rect 4710 10775 4766 10784
rect 4620 10746 4672 10752
rect 4620 10668 4672 10674
rect 4816 10656 4844 10968
rect 4896 10950 4948 10956
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 4896 10668 4948 10674
rect 4816 10628 4896 10656
rect 4620 10610 4672 10616
rect 4896 10610 4948 10616
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4068 10260 4120 10266
rect 4632 10248 4660 10610
rect 4802 10432 4858 10441
rect 4802 10367 4858 10376
rect 4068 10202 4120 10208
rect 4540 10220 4660 10248
rect 4710 10296 4766 10305
rect 4710 10231 4766 10240
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 4080 10118 4292 10146
rect 3884 10056 3936 10062
rect 3804 10016 3884 10044
rect 3884 9998 3936 10004
rect 3896 9722 3924 9998
rect 3976 9988 4028 9994
rect 4080 9976 4108 10118
rect 4264 10062 4292 10118
rect 4160 10056 4212 10062
rect 4028 9948 4108 9976
rect 4158 10024 4160 10033
rect 4252 10056 4304 10062
rect 4212 10024 4214 10033
rect 4252 9998 4304 10004
rect 4158 9959 4214 9968
rect 3976 9930 4028 9936
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3896 9586 3924 9658
rect 4434 9616 4490 9625
rect 3884 9580 3936 9586
rect 4434 9551 4490 9560
rect 3884 9522 3936 9528
rect 4068 9512 4120 9518
rect 3882 9480 3938 9489
rect 3712 9438 3882 9466
rect 4068 9454 4120 9460
rect 4252 9512 4304 9518
rect 4448 9500 4476 9551
rect 4304 9472 4476 9500
rect 4252 9454 4304 9460
rect 3882 9415 3938 9424
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 3804 7449 3832 9318
rect 3896 8974 3924 9415
rect 4080 9178 4108 9454
rect 4540 9364 4568 10220
rect 4724 9722 4752 10231
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4816 9586 4844 10367
rect 5000 10169 5028 10746
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 4986 10160 5042 10169
rect 4896 10124 4948 10130
rect 4986 10095 5042 10104
rect 4896 10066 4948 10072
rect 4908 9926 4936 10066
rect 5092 9994 5120 10542
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 4896 9920 4948 9926
rect 5184 9908 5212 10406
rect 5276 10062 5304 11018
rect 5354 10976 5410 10985
rect 5354 10911 5410 10920
rect 5368 10674 5396 10911
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5356 10192 5408 10198
rect 5354 10160 5356 10169
rect 5408 10160 5410 10169
rect 5354 10095 5410 10104
rect 5264 10056 5316 10062
rect 5460 10044 5488 12940
rect 5724 12912 5776 12918
rect 5724 12854 5776 12860
rect 5736 12764 5764 12854
rect 5538 12744 5594 12753
rect 5538 12679 5594 12688
rect 5644 12736 5764 12764
rect 5552 10849 5580 12679
rect 5644 12050 5672 12736
rect 5828 12374 5856 12974
rect 5920 12850 5948 13144
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5816 12368 5868 12374
rect 5722 12336 5778 12345
rect 5816 12310 5868 12316
rect 5722 12271 5778 12280
rect 5736 12238 5764 12271
rect 5724 12232 5776 12238
rect 6012 12186 6040 13806
rect 6288 13326 6316 15642
rect 6380 15178 6408 17138
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6564 15638 6592 16934
rect 6748 16232 6776 18634
rect 6840 17184 6868 20431
rect 6932 18034 6960 20470
rect 7024 19009 7052 21406
rect 7010 19000 7066 19009
rect 7010 18935 7066 18944
rect 7010 18864 7066 18873
rect 7010 18799 7066 18808
rect 7024 18766 7052 18799
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 7024 18154 7052 18702
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 6932 18006 7052 18034
rect 6920 17196 6972 17202
rect 6840 17156 6920 17184
rect 6840 16969 6868 17156
rect 6920 17138 6972 17144
rect 6826 16960 6882 16969
rect 6826 16895 6882 16904
rect 7024 16250 7052 18006
rect 7012 16244 7064 16250
rect 6748 16204 6868 16232
rect 6734 16144 6790 16153
rect 6734 16079 6736 16088
rect 6788 16079 6790 16088
rect 6736 16050 6788 16056
rect 6734 15736 6790 15745
rect 6734 15671 6736 15680
rect 6788 15671 6790 15680
rect 6736 15642 6788 15648
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 6642 15600 6698 15609
rect 6642 15535 6698 15544
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6564 15337 6592 15438
rect 6550 15328 6606 15337
rect 6550 15263 6606 15272
rect 6380 15150 6500 15178
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6380 13870 6408 14894
rect 6472 14498 6500 15150
rect 6656 14618 6684 15535
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6748 15162 6776 15438
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6840 14634 6868 16204
rect 7012 16186 7064 16192
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6748 14606 6868 14634
rect 6472 14470 6684 14498
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 6368 13456 6420 13462
rect 6368 13398 6420 13404
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6104 12481 6132 12922
rect 6196 12889 6224 13126
rect 6182 12880 6238 12889
rect 6182 12815 6238 12824
rect 6288 12782 6316 13262
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 6090 12472 6146 12481
rect 6090 12407 6146 12416
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 5724 12174 5776 12180
rect 5828 12158 6040 12186
rect 5722 12064 5778 12073
rect 5644 12022 5722 12050
rect 5722 11999 5778 12008
rect 5630 11928 5686 11937
rect 5630 11863 5632 11872
rect 5684 11863 5686 11872
rect 5724 11892 5776 11898
rect 5632 11834 5684 11840
rect 5724 11834 5776 11840
rect 5630 11792 5686 11801
rect 5630 11727 5632 11736
rect 5684 11727 5686 11736
rect 5632 11698 5684 11704
rect 5632 11144 5684 11150
rect 5630 11112 5632 11121
rect 5684 11112 5686 11121
rect 5630 11047 5686 11056
rect 5736 11014 5764 11834
rect 5828 11082 5856 12158
rect 5908 11620 5960 11626
rect 5908 11562 5960 11568
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5724 11008 5776 11014
rect 5920 10985 5948 11562
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 6012 11393 6040 11494
rect 5998 11384 6054 11393
rect 5998 11319 6054 11328
rect 5724 10950 5776 10956
rect 5906 10976 5962 10985
rect 5906 10911 5962 10920
rect 5538 10840 5594 10849
rect 5538 10775 5594 10784
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5908 10804 5960 10810
rect 6012 10792 6040 11319
rect 5960 10764 6040 10792
rect 5908 10746 5960 10752
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5644 10588 5672 10678
rect 5736 10656 5764 10746
rect 6000 10668 6052 10674
rect 5736 10628 6000 10656
rect 6000 10610 6052 10616
rect 5644 10560 5948 10588
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5264 9998 5316 10004
rect 5386 10016 5488 10044
rect 5386 9976 5414 10016
rect 5368 9948 5414 9976
rect 5184 9880 5304 9908
rect 4896 9862 4948 9868
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5276 9704 5304 9880
rect 5368 9722 5396 9948
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5000 9676 5304 9704
rect 5356 9716 5408 9722
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4540 9336 4660 9364
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4068 9172 4120 9178
rect 3988 9132 4068 9160
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3988 7478 4016 9132
rect 4068 9114 4120 9120
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4172 8566 4200 8910
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4160 8560 4212 8566
rect 4080 8520 4160 8548
rect 3976 7472 4028 7478
rect 3790 7440 3846 7449
rect 4080 7460 4108 8520
rect 4160 8502 4212 8508
rect 4356 8362 4384 8842
rect 4448 8634 4476 8910
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4540 8378 4568 8910
rect 4632 8498 4660 9336
rect 4724 8974 4752 9386
rect 4894 9344 4950 9353
rect 4894 9279 4950 9288
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4816 8634 4844 8910
rect 4908 8838 4936 9279
rect 4896 8832 4948 8838
rect 5000 8820 5028 9676
rect 5356 9658 5408 9664
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5092 8945 5120 9114
rect 5078 8936 5134 8945
rect 5184 8922 5212 9318
rect 5276 9042 5304 9386
rect 5460 9382 5488 9862
rect 5552 9500 5580 10406
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5644 9568 5672 9862
rect 5736 9722 5764 10202
rect 5828 10062 5856 10406
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 5828 9761 5856 9862
rect 5814 9752 5870 9761
rect 5724 9716 5776 9722
rect 5814 9687 5870 9696
rect 5920 9704 5948 10560
rect 6104 10470 6132 12242
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6196 10282 6224 12718
rect 6380 12442 6408 13398
rect 6472 12986 6500 14350
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6458 12880 6514 12889
rect 6564 12850 6592 14350
rect 6656 13734 6684 14470
rect 6748 14414 6776 14606
rect 6828 14544 6880 14550
rect 6826 14512 6828 14521
rect 6880 14512 6882 14521
rect 6826 14447 6882 14456
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6644 13728 6696 13734
rect 6644 13670 6696 13676
rect 6748 13308 6776 14350
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6656 13280 6776 13308
rect 6458 12815 6514 12824
rect 6552 12844 6604 12850
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6472 12322 6500 12815
rect 6552 12786 6604 12792
rect 6552 12708 6604 12714
rect 6552 12650 6604 12656
rect 6380 12294 6500 12322
rect 6564 12306 6592 12650
rect 6656 12617 6684 13280
rect 6736 13184 6788 13190
rect 6734 13152 6736 13161
rect 6788 13152 6790 13161
rect 6734 13087 6790 13096
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6642 12608 6698 12617
rect 6642 12543 6698 12552
rect 6552 12300 6604 12306
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 6288 11354 6316 11698
rect 6380 11354 6408 12294
rect 6552 12242 6604 12248
rect 6656 12238 6684 12543
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6552 12164 6604 12170
rect 6552 12106 6604 12112
rect 6564 11937 6592 12106
rect 6748 11937 6776 12922
rect 6840 12889 6868 14214
rect 6826 12880 6882 12889
rect 6826 12815 6882 12824
rect 6826 12744 6882 12753
rect 6826 12679 6828 12688
rect 6880 12679 6882 12688
rect 6828 12650 6880 12656
rect 6932 12442 6960 16118
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 7024 16017 7052 16050
rect 7010 16008 7066 16017
rect 7010 15943 7066 15952
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7024 15065 7052 15098
rect 7010 15056 7066 15065
rect 7010 14991 7066 15000
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 7024 14414 7052 14894
rect 7012 14408 7064 14414
rect 7012 14350 7064 14356
rect 7012 13796 7064 13802
rect 7012 13738 7064 13744
rect 7024 12850 7052 13738
rect 7116 13002 7144 22374
rect 7208 22030 7236 22374
rect 7196 22024 7248 22030
rect 7196 21966 7248 21972
rect 7300 21434 7328 23004
rect 7392 22642 7420 23287
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 7208 21406 7328 21434
rect 7208 19922 7236 21406
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7300 21078 7328 21286
rect 7288 21072 7340 21078
rect 7288 21014 7340 21020
rect 7392 20806 7420 22578
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7196 19916 7248 19922
rect 7196 19858 7248 19864
rect 7380 19848 7432 19854
rect 7300 19808 7380 19836
rect 7300 17746 7328 19808
rect 7380 19790 7432 19796
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 7392 19514 7420 19654
rect 7380 19508 7432 19514
rect 7380 19450 7432 19456
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7196 17604 7248 17610
rect 7196 17546 7248 17552
rect 7208 17338 7236 17546
rect 7300 17338 7328 17682
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7392 17270 7420 19450
rect 7484 19446 7512 23446
rect 7576 23322 7604 23462
rect 7654 23352 7710 23361
rect 7564 23316 7616 23322
rect 7654 23287 7710 23296
rect 7564 23258 7616 23264
rect 7564 23112 7616 23118
rect 7562 23080 7564 23089
rect 7616 23080 7618 23089
rect 7562 23015 7618 23024
rect 7576 22778 7604 23015
rect 7668 22982 7696 23287
rect 7656 22976 7708 22982
rect 7656 22918 7708 22924
rect 7564 22772 7616 22778
rect 7564 22714 7616 22720
rect 7668 22409 7696 22918
rect 7654 22400 7710 22409
rect 7654 22335 7710 22344
rect 7564 21548 7616 21554
rect 7564 21490 7616 21496
rect 7576 21350 7604 21490
rect 7564 21344 7616 21350
rect 7564 21286 7616 21292
rect 7564 19984 7616 19990
rect 7562 19952 7564 19961
rect 7616 19952 7618 19961
rect 7562 19887 7618 19896
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7576 19496 7604 19654
rect 7656 19508 7708 19514
rect 7576 19468 7656 19496
rect 7472 19440 7524 19446
rect 7576 19417 7604 19468
rect 7656 19450 7708 19456
rect 7472 19382 7524 19388
rect 7562 19408 7618 19417
rect 7562 19343 7618 19352
rect 7564 19304 7616 19310
rect 7564 19246 7616 19252
rect 7472 19236 7524 19242
rect 7472 19178 7524 19184
rect 7484 18970 7512 19178
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7484 18766 7512 18906
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 7472 18624 7524 18630
rect 7470 18592 7472 18601
rect 7524 18592 7526 18601
rect 7470 18527 7526 18536
rect 7472 18148 7524 18154
rect 7472 18090 7524 18096
rect 7484 18057 7512 18090
rect 7470 18048 7526 18057
rect 7470 17983 7526 17992
rect 7576 17354 7604 19246
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7668 18630 7696 18906
rect 7760 18630 7788 24550
rect 7852 23225 7880 24670
rect 7838 23216 7894 23225
rect 7838 23151 7894 23160
rect 7932 23180 7984 23186
rect 7932 23122 7984 23128
rect 7840 23112 7892 23118
rect 7840 23054 7892 23060
rect 7852 22778 7880 23054
rect 7840 22772 7892 22778
rect 7840 22714 7892 22720
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7852 22234 7880 22578
rect 7840 22228 7892 22234
rect 7840 22170 7892 22176
rect 7944 21690 7972 23122
rect 7932 21684 7984 21690
rect 7932 21626 7984 21632
rect 8036 21622 8064 27542
rect 8116 26852 8168 26858
rect 8116 26794 8168 26800
rect 8128 26586 8156 26794
rect 8116 26580 8168 26586
rect 8116 26522 8168 26528
rect 8128 26314 8156 26522
rect 8116 26308 8168 26314
rect 8116 26250 8168 26256
rect 8116 25900 8168 25906
rect 8116 25842 8168 25848
rect 8128 24857 8156 25842
rect 8220 25129 8248 28494
rect 8312 28422 8340 28494
rect 8300 28416 8352 28422
rect 8300 28358 8352 28364
rect 8312 26382 8340 28358
rect 8404 28218 8432 28970
rect 8576 28688 8628 28694
rect 8576 28630 8628 28636
rect 8680 28642 8708 29038
rect 9048 28994 9076 29174
rect 9416 29170 9444 29718
rect 9678 29679 9734 29688
rect 9692 29306 9720 29679
rect 9680 29300 9732 29306
rect 9680 29242 9732 29248
rect 9772 29300 9824 29306
rect 9772 29242 9824 29248
rect 9126 29135 9182 29144
rect 9404 29164 9456 29170
rect 9404 29106 9456 29112
rect 8956 28966 9076 28994
rect 8392 28212 8444 28218
rect 8444 28172 8524 28200
rect 8392 28154 8444 28160
rect 8496 27470 8524 28172
rect 8588 28082 8616 28630
rect 8680 28614 8892 28642
rect 8680 28150 8708 28614
rect 8760 28552 8812 28558
rect 8760 28494 8812 28500
rect 8772 28150 8800 28494
rect 8668 28144 8720 28150
rect 8668 28086 8720 28092
rect 8760 28144 8812 28150
rect 8760 28086 8812 28092
rect 8576 28076 8628 28082
rect 8576 28018 8628 28024
rect 8668 27940 8720 27946
rect 8668 27882 8720 27888
rect 8484 27464 8536 27470
rect 8484 27406 8536 27412
rect 8392 26988 8444 26994
rect 8392 26930 8444 26936
rect 8300 26376 8352 26382
rect 8300 26318 8352 26324
rect 8300 26240 8352 26246
rect 8300 26182 8352 26188
rect 8312 25974 8340 26182
rect 8404 26042 8432 26930
rect 8484 26784 8536 26790
rect 8482 26752 8484 26761
rect 8576 26784 8628 26790
rect 8536 26752 8538 26761
rect 8576 26726 8628 26732
rect 8482 26687 8538 26696
rect 8588 26217 8616 26726
rect 8574 26208 8630 26217
rect 8574 26143 8630 26152
rect 8680 26058 8708 27882
rect 8772 27878 8800 28086
rect 8760 27872 8812 27878
rect 8760 27814 8812 27820
rect 8760 27056 8812 27062
rect 8760 26998 8812 27004
rect 8772 26246 8800 26998
rect 8760 26240 8812 26246
rect 8760 26182 8812 26188
rect 8392 26036 8444 26042
rect 8392 25978 8444 25984
rect 8496 26030 8708 26058
rect 8300 25968 8352 25974
rect 8300 25910 8352 25916
rect 8392 25900 8444 25906
rect 8392 25842 8444 25848
rect 8300 25832 8352 25838
rect 8300 25774 8352 25780
rect 8312 25702 8340 25774
rect 8300 25696 8352 25702
rect 8300 25638 8352 25644
rect 8404 25294 8432 25842
rect 8496 25498 8524 26030
rect 8772 25906 8800 26182
rect 8760 25900 8812 25906
rect 8760 25842 8812 25848
rect 8576 25696 8628 25702
rect 8576 25638 8628 25644
rect 8484 25492 8536 25498
rect 8484 25434 8536 25440
rect 8392 25288 8444 25294
rect 8392 25230 8444 25236
rect 8206 25120 8262 25129
rect 8206 25055 8262 25064
rect 8114 24848 8170 24857
rect 8496 24818 8524 25434
rect 8588 25362 8616 25638
rect 8772 25498 8800 25842
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 8576 25356 8628 25362
rect 8576 25298 8628 25304
rect 8588 24818 8616 25298
rect 8666 25256 8722 25265
rect 8666 25191 8722 25200
rect 8680 24886 8708 25191
rect 8668 24880 8720 24886
rect 8864 24834 8892 28614
rect 8956 26586 8984 28966
rect 9220 28960 9272 28966
rect 9416 28937 9444 29106
rect 9692 29102 9720 29242
rect 9784 29170 9812 29242
rect 9876 29170 9904 29786
rect 10704 29646 10732 29990
rect 11704 29776 11756 29782
rect 11704 29718 11756 29724
rect 10692 29640 10744 29646
rect 10692 29582 10744 29588
rect 10232 29572 10284 29578
rect 10232 29514 10284 29520
rect 10048 29232 10100 29238
rect 10048 29174 10100 29180
rect 9772 29164 9824 29170
rect 9772 29106 9824 29112
rect 9864 29164 9916 29170
rect 9864 29106 9916 29112
rect 9680 29096 9732 29102
rect 9876 29073 9904 29106
rect 9680 29038 9732 29044
rect 9862 29064 9918 29073
rect 9862 28999 9918 29008
rect 9864 28960 9916 28966
rect 9220 28902 9272 28908
rect 9402 28928 9458 28937
rect 9232 28626 9260 28902
rect 9864 28902 9916 28908
rect 9402 28863 9458 28872
rect 9220 28620 9272 28626
rect 9220 28562 9272 28568
rect 9036 28416 9088 28422
rect 9036 28358 9088 28364
rect 9048 28082 9076 28358
rect 9036 28076 9088 28082
rect 9036 28018 9088 28024
rect 9126 27976 9182 27985
rect 9126 27911 9128 27920
rect 9180 27911 9182 27920
rect 9128 27882 9180 27888
rect 9128 27328 9180 27334
rect 9126 27296 9128 27305
rect 9180 27296 9182 27305
rect 9126 27231 9182 27240
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 8944 26580 8996 26586
rect 8944 26522 8996 26528
rect 8956 25838 8984 26522
rect 9048 26042 9076 26930
rect 9140 26194 9168 26930
rect 9232 26382 9260 28562
rect 9772 28552 9824 28558
rect 9772 28494 9824 28500
rect 9588 28484 9640 28490
rect 9588 28426 9640 28432
rect 9404 28416 9456 28422
rect 9600 28393 9628 28426
rect 9404 28358 9456 28364
rect 9586 28384 9642 28393
rect 9416 28150 9444 28358
rect 9586 28319 9642 28328
rect 9784 28218 9812 28494
rect 9876 28218 9904 28902
rect 9956 28416 10008 28422
rect 9956 28358 10008 28364
rect 9772 28212 9824 28218
rect 9772 28154 9824 28160
rect 9864 28212 9916 28218
rect 9864 28154 9916 28160
rect 9404 28144 9456 28150
rect 9404 28086 9456 28092
rect 9588 28144 9640 28150
rect 9588 28086 9640 28092
rect 9312 27872 9364 27878
rect 9312 27814 9364 27820
rect 9324 27538 9352 27814
rect 9312 27532 9364 27538
rect 9312 27474 9364 27480
rect 9324 26994 9352 27474
rect 9416 27334 9444 28086
rect 9496 28076 9548 28082
rect 9496 28018 9548 28024
rect 9404 27328 9456 27334
rect 9404 27270 9456 27276
rect 9312 26988 9364 26994
rect 9312 26930 9364 26936
rect 9324 26450 9352 26930
rect 9416 26926 9444 27270
rect 9508 27130 9536 28018
rect 9600 27878 9628 28086
rect 9680 27940 9732 27946
rect 9680 27882 9732 27888
rect 9588 27872 9640 27878
rect 9588 27814 9640 27820
rect 9600 27606 9628 27814
rect 9588 27600 9640 27606
rect 9588 27542 9640 27548
rect 9600 27470 9628 27542
rect 9692 27470 9720 27882
rect 9588 27464 9640 27470
rect 9588 27406 9640 27412
rect 9680 27464 9732 27470
rect 9680 27406 9732 27412
rect 9784 27418 9812 28154
rect 9876 28082 9904 28154
rect 9864 28076 9916 28082
rect 9864 28018 9916 28024
rect 9968 27538 9996 28358
rect 10060 28082 10088 29174
rect 10244 28994 10272 29514
rect 10508 29504 10560 29510
rect 10508 29446 10560 29452
rect 10152 28966 10272 28994
rect 10152 28490 10180 28966
rect 10416 28756 10468 28762
rect 10416 28698 10468 28704
rect 10140 28484 10192 28490
rect 10140 28426 10192 28432
rect 10152 28393 10180 28426
rect 10138 28384 10194 28393
rect 10138 28319 10194 28328
rect 10048 28076 10100 28082
rect 10048 28018 10100 28024
rect 9956 27532 10008 27538
rect 9956 27474 10008 27480
rect 9496 27124 9548 27130
rect 9496 27066 9548 27072
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 9404 26580 9456 26586
rect 9404 26522 9456 26528
rect 9312 26444 9364 26450
rect 9312 26386 9364 26392
rect 9220 26376 9272 26382
rect 9220 26318 9272 26324
rect 9220 26240 9272 26246
rect 9140 26188 9220 26194
rect 9140 26182 9272 26188
rect 9140 26166 9260 26182
rect 9036 26036 9088 26042
rect 9036 25978 9088 25984
rect 8944 25832 8996 25838
rect 8944 25774 8996 25780
rect 9048 25294 9076 25978
rect 9140 25770 9168 26166
rect 9416 25906 9444 26522
rect 9508 26314 9536 27066
rect 9600 26874 9628 27406
rect 9692 27146 9720 27406
rect 9784 27402 9904 27418
rect 9784 27396 9916 27402
rect 9784 27390 9864 27396
rect 9864 27338 9916 27344
rect 9692 27118 9812 27146
rect 9784 27062 9812 27118
rect 9772 27056 9824 27062
rect 9772 26998 9824 27004
rect 9968 26994 9996 27474
rect 9956 26988 10008 26994
rect 9956 26930 10008 26936
rect 9772 26920 9824 26926
rect 9600 26868 9772 26874
rect 9600 26862 9824 26868
rect 9600 26846 9812 26862
rect 9864 26784 9916 26790
rect 9864 26726 9916 26732
rect 9586 26616 9642 26625
rect 9586 26551 9642 26560
rect 9770 26616 9826 26625
rect 9876 26586 9904 26726
rect 9770 26551 9826 26560
rect 9864 26580 9916 26586
rect 9496 26308 9548 26314
rect 9496 26250 9548 26256
rect 9496 26036 9548 26042
rect 9496 25978 9548 25984
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9508 25838 9536 25978
rect 9496 25832 9548 25838
rect 9496 25774 9548 25780
rect 9128 25764 9180 25770
rect 9128 25706 9180 25712
rect 8944 25288 8996 25294
rect 8944 25230 8996 25236
rect 9036 25288 9088 25294
rect 9036 25230 9088 25236
rect 8668 24822 8720 24828
rect 8114 24783 8170 24792
rect 8484 24812 8536 24818
rect 8484 24754 8536 24760
rect 8576 24812 8628 24818
rect 8576 24754 8628 24760
rect 8772 24806 8892 24834
rect 8484 24676 8536 24682
rect 8484 24618 8536 24624
rect 8496 24070 8524 24618
rect 8484 24064 8536 24070
rect 8484 24006 8536 24012
rect 8496 23730 8524 24006
rect 8484 23724 8536 23730
rect 8484 23666 8536 23672
rect 8300 23520 8352 23526
rect 8300 23462 8352 23468
rect 8312 23202 8340 23462
rect 8128 23174 8340 23202
rect 8128 23118 8156 23174
rect 8116 23112 8168 23118
rect 8116 23054 8168 23060
rect 8208 23112 8260 23118
rect 8208 23054 8260 23060
rect 8114 22944 8170 22953
rect 8114 22879 8170 22888
rect 8024 21616 8076 21622
rect 8024 21558 8076 21564
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 7852 20874 7880 21490
rect 8024 21344 8076 21350
rect 8024 21286 8076 21292
rect 7930 21040 7986 21049
rect 7930 20975 7986 20984
rect 7944 20874 7972 20975
rect 7840 20868 7892 20874
rect 7840 20810 7892 20816
rect 7932 20868 7984 20874
rect 7932 20810 7984 20816
rect 7838 20768 7894 20777
rect 7838 20703 7894 20712
rect 7656 18624 7708 18630
rect 7654 18592 7656 18601
rect 7748 18624 7800 18630
rect 7708 18592 7710 18601
rect 7748 18566 7800 18572
rect 7654 18527 7710 18536
rect 7746 18320 7802 18329
rect 7852 18290 7880 20703
rect 7930 20088 7986 20097
rect 7930 20023 7986 20032
rect 7944 19310 7972 20023
rect 7932 19304 7984 19310
rect 7932 19246 7984 19252
rect 7932 18760 7984 18766
rect 7932 18702 7984 18708
rect 7944 18426 7972 18702
rect 7932 18420 7984 18426
rect 7932 18362 7984 18368
rect 7746 18255 7748 18264
rect 7800 18255 7802 18264
rect 7840 18284 7892 18290
rect 7748 18226 7800 18232
rect 7840 18226 7892 18232
rect 7760 18170 7788 18226
rect 7932 18216 7984 18222
rect 7760 18154 7880 18170
rect 7932 18158 7984 18164
rect 7760 18148 7892 18154
rect 7760 18142 7840 18148
rect 7840 18090 7892 18096
rect 7746 18048 7802 18057
rect 7746 17983 7802 17992
rect 7656 17808 7708 17814
rect 7656 17750 7708 17756
rect 7484 17326 7604 17354
rect 7668 17338 7696 17750
rect 7656 17332 7708 17338
rect 7380 17264 7432 17270
rect 7380 17206 7432 17212
rect 7484 17082 7512 17326
rect 7656 17274 7708 17280
rect 7656 17196 7708 17202
rect 7288 17060 7340 17066
rect 7288 17002 7340 17008
rect 7392 17054 7512 17082
rect 7576 17156 7656 17184
rect 7194 16144 7250 16153
rect 7194 16079 7250 16088
rect 7208 14657 7236 16079
rect 7300 15065 7328 17002
rect 7392 16561 7420 17054
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7484 16794 7512 16934
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7472 16584 7524 16590
rect 7378 16552 7434 16561
rect 7472 16526 7524 16532
rect 7378 16487 7434 16496
rect 7484 15434 7512 16526
rect 7380 15428 7432 15434
rect 7380 15370 7432 15376
rect 7472 15428 7524 15434
rect 7472 15370 7524 15376
rect 7392 15094 7420 15370
rect 7380 15088 7432 15094
rect 7286 15056 7342 15065
rect 7380 15030 7432 15036
rect 7286 14991 7342 15000
rect 7194 14648 7250 14657
rect 7194 14583 7250 14592
rect 7300 14482 7328 14991
rect 7392 14618 7420 15030
rect 7484 15026 7512 15370
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7470 14784 7526 14793
rect 7470 14719 7526 14728
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7288 14476 7340 14482
rect 7288 14418 7340 14424
rect 7288 14340 7340 14346
rect 7288 14282 7340 14288
rect 7300 14074 7328 14282
rect 7484 14278 7512 14719
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7378 14104 7434 14113
rect 7288 14068 7340 14074
rect 7378 14039 7434 14048
rect 7288 14010 7340 14016
rect 7392 13870 7420 14039
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 7208 13161 7236 13806
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7288 13456 7340 13462
rect 7286 13424 7288 13433
rect 7340 13424 7342 13433
rect 7484 13394 7512 13670
rect 7286 13359 7342 13368
rect 7472 13388 7524 13394
rect 7194 13152 7250 13161
rect 7194 13087 7250 13096
rect 7116 12974 7236 13002
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6550 11928 6606 11937
rect 6550 11863 6606 11872
rect 6734 11928 6790 11937
rect 6734 11863 6790 11872
rect 6460 11824 6512 11830
rect 6512 11784 6684 11812
rect 6460 11766 6512 11772
rect 6458 11656 6514 11665
rect 6458 11591 6460 11600
rect 6512 11591 6514 11600
rect 6460 11562 6512 11568
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6288 11234 6316 11290
rect 6564 11286 6592 11494
rect 6552 11280 6604 11286
rect 6288 11206 6500 11234
rect 6656 11257 6684 11784
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6552 11222 6604 11228
rect 6642 11248 6698 11257
rect 6368 11144 6420 11150
rect 6366 11112 6368 11121
rect 6420 11112 6422 11121
rect 6366 11047 6422 11056
rect 6366 10976 6422 10985
rect 6366 10911 6422 10920
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6172 10254 6224 10282
rect 6000 9716 6052 9722
rect 5724 9658 5776 9664
rect 5828 9654 5856 9687
rect 5920 9676 6000 9704
rect 6000 9658 6052 9664
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5644 9540 5764 9568
rect 5552 9472 5672 9500
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5448 9104 5500 9110
rect 5500 9064 5580 9092
rect 5448 9046 5500 9052
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5184 8894 5396 8922
rect 5078 8871 5134 8880
rect 5000 8809 5304 8820
rect 5000 8800 5318 8809
rect 5000 8792 5262 8800
rect 4896 8774 4948 8780
rect 4874 8732 5182 8741
rect 5262 8735 5318 8744
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4802 8528 4858 8537
rect 4620 8492 4672 8498
rect 4802 8463 4858 8472
rect 4986 8528 5042 8537
rect 4986 8463 5042 8472
rect 5264 8492 5316 8498
rect 4620 8434 4672 8440
rect 4344 8356 4396 8362
rect 4540 8350 4660 8378
rect 4344 8298 4396 8304
rect 4632 8265 4660 8350
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4618 8256 4674 8265
rect 4214 8188 4522 8197
rect 4618 8191 4674 8200
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4724 7732 4752 8298
rect 4816 8090 4844 8463
rect 5000 8430 5028 8463
rect 5264 8434 5316 8440
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 5276 8022 5304 8434
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 4724 7704 4844 7732
rect 4160 7472 4212 7478
rect 4080 7432 4160 7460
rect 3976 7414 4028 7420
rect 4160 7414 4212 7420
rect 4250 7440 4306 7449
rect 3790 7375 3846 7384
rect 3988 6934 4016 7414
rect 4816 7410 4844 7704
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4986 7440 5042 7449
rect 4250 7375 4252 7384
rect 4304 7375 4306 7384
rect 4712 7404 4764 7410
rect 4252 7346 4304 7352
rect 4712 7346 4764 7352
rect 4804 7404 4856 7410
rect 4986 7375 4988 7384
rect 4804 7346 4856 7352
rect 5040 7375 5042 7384
rect 4988 7346 5040 7352
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4724 7002 4752 7346
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 5092 7002 5120 7210
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 5368 5778 5396 8894
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5460 8566 5488 8774
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5552 8498 5580 9064
rect 5644 8974 5672 9472
rect 5736 9330 5764 9540
rect 6104 9382 6132 10202
rect 6172 10044 6200 10254
rect 6288 10062 6316 10406
rect 6276 10056 6328 10062
rect 6172 10016 6224 10044
rect 6092 9376 6144 9382
rect 5736 9302 6040 9330
rect 6092 9318 6144 9324
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5446 8392 5502 8401
rect 5446 8327 5502 8336
rect 5460 6934 5488 8327
rect 5552 7750 5580 8434
rect 5644 7954 5672 8910
rect 5736 8498 5764 8910
rect 5828 8906 5856 9114
rect 6012 9110 6040 9302
rect 6090 9208 6146 9217
rect 6090 9143 6146 9152
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 5816 8900 5868 8906
rect 5816 8842 5868 8848
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 5920 8634 5948 8842
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 6012 8498 6040 9046
rect 6104 8974 6132 9143
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 5814 8392 5870 8401
rect 5814 8327 5870 8336
rect 5828 8294 5856 8327
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5552 7410 5580 7686
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5552 5710 5580 7142
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 5828 3126 5856 8230
rect 5920 8022 5948 8230
rect 6012 8022 6040 8434
rect 6104 8265 6132 8774
rect 6090 8256 6146 8265
rect 6090 8191 6146 8200
rect 5908 8016 5960 8022
rect 5908 7958 5960 7964
rect 6000 8016 6052 8022
rect 6000 7958 6052 7964
rect 5920 7410 5948 7958
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5920 7274 5948 7346
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 6092 7200 6144 7206
rect 6196 7188 6224 10016
rect 6276 9998 6328 10004
rect 6274 9752 6330 9761
rect 6274 9687 6330 9696
rect 6288 9654 6316 9687
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6380 8673 6408 10911
rect 6472 9761 6500 11206
rect 6642 11183 6698 11192
rect 6644 11076 6696 11082
rect 6644 11018 6696 11024
rect 6656 10985 6684 11018
rect 6642 10976 6698 10985
rect 6748 10962 6776 11494
rect 6840 11354 6868 12378
rect 6918 12336 6974 12345
rect 6918 12271 6974 12280
rect 6932 12102 6960 12271
rect 7024 12238 7052 12582
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 7010 11928 7066 11937
rect 7010 11863 7012 11872
rect 7064 11863 7066 11872
rect 7012 11834 7064 11840
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7024 11665 7052 11698
rect 7010 11656 7066 11665
rect 7010 11591 7066 11600
rect 7010 11520 7066 11529
rect 7010 11455 7066 11464
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 7024 11150 7052 11455
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 7116 10996 7144 12718
rect 7208 11830 7236 12974
rect 7300 12850 7328 13359
rect 7472 13330 7524 13336
rect 7380 13252 7432 13258
rect 7380 13194 7432 13200
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7392 12730 7420 13194
rect 7300 12702 7420 12730
rect 7300 12238 7328 12702
rect 7484 12238 7512 13330
rect 7576 12288 7604 17156
rect 7656 17138 7708 17144
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7668 15570 7696 16934
rect 7760 16561 7788 17983
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 7852 17678 7880 17818
rect 7840 17672 7892 17678
rect 7840 17614 7892 17620
rect 7944 16810 7972 18158
rect 8036 17814 8064 21286
rect 8128 19922 8156 22879
rect 8220 22438 8248 23054
rect 8300 22976 8352 22982
rect 8352 22936 8432 22964
rect 8300 22918 8352 22924
rect 8298 22536 8354 22545
rect 8298 22471 8354 22480
rect 8208 22432 8260 22438
rect 8208 22374 8260 22380
rect 8208 21344 8260 21350
rect 8208 21286 8260 21292
rect 8220 21078 8248 21286
rect 8208 21072 8260 21078
rect 8208 21014 8260 21020
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 8220 20534 8248 20878
rect 8208 20528 8260 20534
rect 8208 20470 8260 20476
rect 8312 20466 8340 22471
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 8116 19916 8168 19922
rect 8116 19858 8168 19864
rect 8220 19825 8248 19994
rect 8206 19816 8262 19825
rect 8206 19751 8262 19760
rect 8116 19440 8168 19446
rect 8116 19382 8168 19388
rect 8128 18714 8156 19382
rect 8220 18834 8248 19751
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 8128 18686 8248 18714
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 8128 18222 8156 18362
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8024 17808 8076 17814
rect 8024 17750 8076 17756
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 7852 16782 7972 16810
rect 8036 16794 8064 17274
rect 8220 17202 8248 18686
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 8312 17105 8340 20402
rect 8404 19334 8432 22936
rect 8588 21486 8616 24754
rect 8666 24576 8722 24585
rect 8666 24511 8722 24520
rect 8680 24206 8708 24511
rect 8668 24200 8720 24206
rect 8668 24142 8720 24148
rect 8772 23712 8800 24806
rect 8956 24410 8984 25230
rect 9036 24948 9088 24954
rect 9036 24890 9088 24896
rect 9048 24449 9076 24890
rect 9034 24440 9090 24449
rect 8944 24404 8996 24410
rect 9034 24375 9090 24384
rect 8944 24346 8996 24352
rect 8850 24304 8906 24313
rect 8850 24239 8906 24248
rect 8864 24138 8892 24239
rect 8956 24206 8984 24346
rect 8944 24200 8996 24206
rect 8996 24160 9076 24188
rect 8944 24142 8996 24148
rect 8852 24132 8904 24138
rect 8852 24074 8904 24080
rect 9048 23730 9076 24160
rect 9140 24138 9168 25706
rect 9600 25650 9628 26551
rect 9680 25900 9732 25906
rect 9680 25842 9732 25848
rect 9232 25622 9628 25650
rect 9232 24857 9260 25622
rect 9692 25498 9720 25842
rect 9312 25492 9364 25498
rect 9312 25434 9364 25440
rect 9680 25492 9732 25498
rect 9680 25434 9732 25440
rect 9218 24848 9274 24857
rect 9218 24783 9274 24792
rect 9324 24410 9352 25434
rect 9588 25424 9640 25430
rect 9586 25392 9588 25401
rect 9640 25392 9642 25401
rect 9784 25378 9812 26551
rect 9864 26522 9916 26528
rect 9586 25327 9642 25336
rect 9692 25350 9812 25378
rect 9968 25362 9996 26930
rect 10060 26246 10088 28018
rect 10232 28008 10284 28014
rect 10232 27950 10284 27956
rect 10140 27940 10192 27946
rect 10140 27882 10192 27888
rect 10152 27849 10180 27882
rect 10138 27840 10194 27849
rect 10138 27775 10194 27784
rect 10244 27713 10272 27950
rect 10428 27878 10456 28698
rect 10520 28558 10548 29446
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 10968 29164 11020 29170
rect 10968 29106 11020 29112
rect 10508 28552 10560 28558
rect 10508 28494 10560 28500
rect 10416 27872 10468 27878
rect 10336 27832 10416 27860
rect 10230 27704 10286 27713
rect 10230 27639 10286 27648
rect 10140 27464 10192 27470
rect 10140 27406 10192 27412
rect 10232 27464 10284 27470
rect 10232 27406 10284 27412
rect 10152 26450 10180 27406
rect 10244 27305 10272 27406
rect 10230 27296 10286 27305
rect 10230 27231 10286 27240
rect 10244 27130 10272 27231
rect 10232 27124 10284 27130
rect 10232 27066 10284 27072
rect 10232 26784 10284 26790
rect 10232 26726 10284 26732
rect 10140 26444 10192 26450
rect 10140 26386 10192 26392
rect 10048 26240 10100 26246
rect 10048 26182 10100 26188
rect 9956 25356 10008 25362
rect 9496 25288 9548 25294
rect 9692 25276 9720 25350
rect 9956 25298 10008 25304
rect 10152 25294 10180 26386
rect 9496 25230 9548 25236
rect 9600 25248 9720 25276
rect 10140 25288 10192 25294
rect 9770 25256 9826 25265
rect 9402 25120 9458 25129
rect 9402 25055 9458 25064
rect 9312 24404 9364 24410
rect 9312 24346 9364 24352
rect 9324 24206 9352 24346
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 9128 24132 9180 24138
rect 9128 24074 9180 24080
rect 9416 23730 9444 25055
rect 9508 24614 9536 25230
rect 9496 24608 9548 24614
rect 9494 24576 9496 24585
rect 9548 24576 9550 24585
rect 9494 24511 9550 24520
rect 8852 23724 8904 23730
rect 8772 23684 8852 23712
rect 8772 23526 8800 23684
rect 8852 23666 8904 23672
rect 9036 23724 9088 23730
rect 9036 23666 9088 23672
rect 9404 23724 9456 23730
rect 9404 23666 9456 23672
rect 8760 23520 8812 23526
rect 8760 23462 8812 23468
rect 9036 23520 9088 23526
rect 9036 23462 9088 23468
rect 9048 23089 9076 23462
rect 9034 23080 9090 23089
rect 9034 23015 9090 23024
rect 8668 22636 8720 22642
rect 8852 22636 8904 22642
rect 8668 22578 8720 22584
rect 8772 22596 8852 22624
rect 8680 22234 8708 22578
rect 8668 22228 8720 22234
rect 8668 22170 8720 22176
rect 8668 22024 8720 22030
rect 8666 21992 8668 22001
rect 8720 21992 8722 22001
rect 8666 21927 8722 21936
rect 8668 21888 8720 21894
rect 8668 21830 8720 21836
rect 8576 21480 8628 21486
rect 8576 21422 8628 21428
rect 8574 21176 8630 21185
rect 8680 21146 8708 21830
rect 8772 21418 8800 22596
rect 8852 22578 8904 22584
rect 8944 22636 8996 22642
rect 8944 22578 8996 22584
rect 8956 22506 8984 22578
rect 8944 22500 8996 22506
rect 8944 22442 8996 22448
rect 8852 22160 8904 22166
rect 8852 22102 8904 22108
rect 8760 21412 8812 21418
rect 8760 21354 8812 21360
rect 8574 21111 8630 21120
rect 8668 21140 8720 21146
rect 8588 19446 8616 21111
rect 8668 21082 8720 21088
rect 8772 20874 8800 21354
rect 8760 20868 8812 20874
rect 8760 20810 8812 20816
rect 8864 20398 8892 22102
rect 8956 22030 8984 22442
rect 8944 22024 8996 22030
rect 8944 21966 8996 21972
rect 8942 21856 8998 21865
rect 8942 21791 8998 21800
rect 8956 21078 8984 21791
rect 8944 21072 8996 21078
rect 8944 21014 8996 21020
rect 8956 20777 8984 21014
rect 8942 20768 8998 20777
rect 8942 20703 8998 20712
rect 8942 20632 8998 20641
rect 8942 20567 8998 20576
rect 8852 20392 8904 20398
rect 8852 20334 8904 20340
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8576 19440 8628 19446
rect 8576 19382 8628 19388
rect 8404 19306 8616 19334
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8298 17096 8354 17105
rect 8298 17031 8354 17040
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8024 16788 8076 16794
rect 7746 16552 7802 16561
rect 7746 16487 7802 16496
rect 7852 15858 7880 16782
rect 8024 16730 8076 16736
rect 8022 16008 8078 16017
rect 8022 15943 8078 15952
rect 7760 15830 7880 15858
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7760 14906 7788 15830
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7668 14878 7788 14906
rect 7668 14822 7696 14878
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7760 14482 7788 14758
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 7668 14113 7696 14350
rect 7654 14104 7710 14113
rect 7654 14039 7710 14048
rect 7748 14000 7800 14006
rect 7746 13968 7748 13977
rect 7800 13968 7802 13977
rect 7746 13903 7802 13912
rect 7656 13864 7708 13870
rect 7654 13832 7656 13841
rect 7708 13832 7710 13841
rect 7654 13767 7710 13776
rect 7852 13530 7880 15642
rect 8036 14958 8064 15943
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 7930 14648 7986 14657
rect 7930 14583 7986 14592
rect 7944 14482 7972 14583
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 7840 13524 7892 13530
rect 7892 13484 7972 13512
rect 7840 13466 7892 13472
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7668 13258 7696 13330
rect 7656 13252 7708 13258
rect 7656 13194 7708 13200
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7668 12481 7696 12854
rect 7760 12628 7788 13398
rect 7840 13252 7892 13258
rect 7840 13194 7892 13200
rect 7852 12753 7880 13194
rect 7838 12744 7894 12753
rect 7838 12679 7894 12688
rect 7944 12646 7972 13484
rect 7932 12640 7984 12646
rect 7760 12600 7880 12628
rect 7654 12472 7710 12481
rect 7654 12407 7710 12416
rect 7576 12260 7788 12288
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7654 12200 7710 12209
rect 7196 11824 7248 11830
rect 7196 11766 7248 11772
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7208 11354 7236 11562
rect 7300 11558 7328 12174
rect 7654 12135 7710 12144
rect 7562 12064 7618 12073
rect 7562 11999 7618 12008
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7470 11248 7526 11257
rect 7288 11212 7340 11218
rect 7470 11183 7472 11192
rect 7288 11154 7340 11160
rect 7524 11183 7526 11192
rect 7472 11154 7524 11160
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7300 11098 7328 11154
rect 6932 10968 7144 10996
rect 6748 10934 6868 10962
rect 6642 10911 6698 10920
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6736 10668 6788 10674
rect 6840 10656 6868 10934
rect 6932 10810 6960 10968
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6840 10628 6960 10656
rect 6736 10610 6788 10616
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6564 9897 6592 10542
rect 6656 10198 6684 10610
rect 6748 10441 6776 10610
rect 6932 10538 6960 10628
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 7116 10441 7144 10542
rect 6734 10432 6790 10441
rect 6734 10367 6790 10376
rect 7102 10432 7158 10441
rect 7102 10367 7158 10376
rect 6734 10296 6790 10305
rect 6734 10231 6736 10240
rect 6788 10231 6790 10240
rect 6736 10202 6788 10208
rect 6644 10192 6696 10198
rect 6920 10192 6972 10198
rect 6644 10134 6696 10140
rect 6918 10160 6920 10169
rect 6972 10160 6974 10169
rect 6550 9888 6606 9897
rect 6550 9823 6606 9832
rect 6458 9752 6514 9761
rect 6458 9687 6514 9696
rect 6656 9466 6684 10134
rect 6918 10095 6974 10104
rect 6920 10056 6972 10062
rect 6918 10024 6920 10033
rect 6972 10024 6974 10033
rect 6918 9959 6974 9968
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 6736 9716 6788 9722
rect 6788 9676 6960 9704
rect 6736 9658 6788 9664
rect 6656 9438 6868 9466
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6472 9178 6500 9318
rect 6656 9217 6684 9318
rect 6642 9208 6698 9217
rect 6460 9172 6512 9178
rect 6642 9143 6698 9152
rect 6736 9172 6788 9178
rect 6460 9114 6512 9120
rect 6472 8974 6500 9114
rect 6656 8974 6684 9143
rect 6736 9114 6788 9120
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6644 8832 6696 8838
rect 6642 8800 6644 8809
rect 6696 8800 6698 8809
rect 6642 8735 6698 8744
rect 6366 8664 6422 8673
rect 6276 8628 6328 8634
rect 6366 8599 6422 8608
rect 6276 8570 6328 8576
rect 6288 7886 6316 8570
rect 6748 8401 6776 9114
rect 6840 8634 6868 9438
rect 6932 9042 6960 9676
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 7024 8838 7052 9522
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6734 8392 6790 8401
rect 6734 8327 6790 8336
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6380 7546 6408 7754
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6656 7478 6684 7686
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6748 7410 6776 7822
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6932 7546 6960 7754
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 7024 7410 7052 8774
rect 7116 7886 7144 9930
rect 7208 9110 7236 11086
rect 7300 11070 7420 11098
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7300 10674 7328 10950
rect 7392 10713 7420 11070
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7484 10810 7512 11018
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7576 10742 7604 11999
rect 7668 11830 7696 12135
rect 7656 11824 7708 11830
rect 7656 11766 7708 11772
rect 7654 11656 7710 11665
rect 7654 11591 7710 11600
rect 7668 11132 7696 11591
rect 7760 11286 7788 12260
rect 7852 12170 7880 12600
rect 7930 12608 7932 12617
rect 7984 12608 7986 12617
rect 7930 12543 7986 12552
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 7944 12170 7972 12378
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 7932 12164 7984 12170
rect 7932 12106 7984 12112
rect 7852 11898 7880 12106
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7748 11144 7800 11150
rect 7668 11104 7748 11132
rect 7748 11086 7800 11092
rect 7654 10976 7710 10985
rect 7654 10911 7710 10920
rect 7564 10736 7616 10742
rect 7378 10704 7434 10713
rect 7288 10668 7340 10674
rect 7564 10678 7616 10684
rect 7378 10639 7434 10648
rect 7288 10610 7340 10616
rect 7392 10470 7420 10639
rect 7668 10606 7696 10911
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7760 10198 7788 10610
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7470 9616 7526 9625
rect 7288 9580 7340 9586
rect 7470 9551 7526 9560
rect 7288 9522 7340 9528
rect 7300 9450 7328 9522
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7484 9382 7512 9551
rect 7576 9382 7604 9862
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7484 9217 7512 9318
rect 7470 9208 7526 9217
rect 7470 9143 7526 9152
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 7576 9024 7604 9318
rect 7392 8996 7604 9024
rect 7392 8566 7420 8996
rect 7668 8838 7696 9522
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7760 8838 7788 9386
rect 7852 9024 7880 11494
rect 7944 11014 7972 12106
rect 8036 11558 8064 14758
rect 8128 12073 8156 14962
rect 8220 14074 8248 16934
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8312 15978 8340 16594
rect 8404 16590 8432 16934
rect 8496 16794 8524 19110
rect 8588 17678 8616 19306
rect 8680 18222 8708 19790
rect 8760 19780 8812 19786
rect 8760 19722 8812 19728
rect 8772 19446 8800 19722
rect 8760 19440 8812 19446
rect 8760 19382 8812 19388
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 8772 18086 8800 18634
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8496 16182 8524 16730
rect 8484 16176 8536 16182
rect 8484 16118 8536 16124
rect 8300 15972 8352 15978
rect 8300 15914 8352 15920
rect 8312 15502 8340 15914
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8482 15464 8538 15473
rect 8482 15399 8538 15408
rect 8496 15366 8524 15399
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8404 15026 8432 15302
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8312 14618 8340 14962
rect 8496 14906 8524 14962
rect 8404 14878 8524 14906
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8404 14482 8432 14878
rect 8588 14804 8616 17614
rect 8668 17128 8720 17134
rect 8666 17096 8668 17105
rect 8720 17096 8722 17105
rect 8666 17031 8722 17040
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8680 15473 8708 16050
rect 8666 15464 8722 15473
rect 8666 15399 8722 15408
rect 8666 15328 8722 15337
rect 8666 15263 8722 15272
rect 8680 14890 8708 15263
rect 8772 15094 8800 17750
rect 8864 16114 8892 20198
rect 8956 19854 8984 20567
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8944 18760 8996 18766
rect 8944 18702 8996 18708
rect 8956 18426 8984 18702
rect 8944 18420 8996 18426
rect 8944 18362 8996 18368
rect 9048 18329 9076 23015
rect 9416 22778 9444 23666
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 9600 22658 9628 25248
rect 10140 25230 10192 25236
rect 9770 25191 9826 25200
rect 9956 25220 10008 25226
rect 9680 24812 9732 24818
rect 9680 24754 9732 24760
rect 9692 24449 9720 24754
rect 9784 24750 9812 25191
rect 9956 25162 10008 25168
rect 9862 24984 9918 24993
rect 9968 24954 9996 25162
rect 10140 25152 10192 25158
rect 10140 25094 10192 25100
rect 9862 24919 9918 24928
rect 9956 24948 10008 24954
rect 9772 24744 9824 24750
rect 9772 24686 9824 24692
rect 9770 24576 9826 24585
rect 9770 24511 9826 24520
rect 9678 24440 9734 24449
rect 9678 24375 9734 24384
rect 9680 24336 9732 24342
rect 9680 24278 9732 24284
rect 9692 24177 9720 24278
rect 9678 24168 9734 24177
rect 9678 24103 9734 24112
rect 9784 23662 9812 24511
rect 9772 23656 9824 23662
rect 9772 23598 9824 23604
rect 9772 23520 9824 23526
rect 9772 23462 9824 23468
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 9324 22630 9628 22658
rect 9126 22536 9182 22545
rect 9126 22471 9128 22480
rect 9180 22471 9182 22480
rect 9128 22442 9180 22448
rect 9324 22094 9352 22630
rect 9692 22522 9720 23258
rect 9784 22710 9812 23462
rect 9772 22704 9824 22710
rect 9772 22646 9824 22652
rect 9508 22494 9720 22522
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 9140 22066 9352 22094
rect 9034 18320 9090 18329
rect 9034 18255 9090 18264
rect 9140 17542 9168 22066
rect 9220 21956 9272 21962
rect 9220 21898 9272 21904
rect 9232 21185 9260 21898
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9324 21554 9352 21830
rect 9312 21548 9364 21554
rect 9312 21490 9364 21496
rect 9324 21457 9352 21490
rect 9310 21448 9366 21457
rect 9310 21383 9366 21392
rect 9218 21176 9274 21185
rect 9218 21111 9220 21120
rect 9272 21111 9274 21120
rect 9220 21082 9272 21088
rect 9310 21040 9366 21049
rect 9220 21004 9272 21010
rect 9310 20975 9366 20984
rect 9220 20946 9272 20952
rect 9232 20874 9260 20946
rect 9220 20868 9272 20874
rect 9220 20810 9272 20816
rect 9218 20632 9274 20641
rect 9218 20567 9274 20576
rect 9232 20262 9260 20567
rect 9220 20256 9272 20262
rect 9220 20198 9272 20204
rect 9220 18692 9272 18698
rect 9220 18634 9272 18640
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 8942 16824 8998 16833
rect 8942 16759 8998 16768
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8864 15162 8892 15846
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 8760 15088 8812 15094
rect 8760 15030 8812 15036
rect 8852 15020 8904 15026
rect 8852 14962 8904 14968
rect 8864 14906 8892 14962
rect 8668 14884 8720 14890
rect 8668 14826 8720 14832
rect 8772 14878 8892 14906
rect 8496 14776 8616 14804
rect 8666 14784 8722 14793
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 8220 12986 8248 13126
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 8114 12064 8170 12073
rect 8114 11999 8170 12008
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8128 11370 8156 11999
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8036 11342 8156 11370
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 7944 9450 7972 9522
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 7852 8996 7972 9024
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7380 8560 7432 8566
rect 7380 8502 7432 8508
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7484 7478 7512 8570
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 7668 7410 7696 8366
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 6380 7274 6408 7346
rect 6368 7268 6420 7274
rect 6368 7210 6420 7216
rect 6144 7160 6224 7188
rect 6828 7200 6880 7206
rect 6092 7142 6144 7148
rect 7012 7200 7064 7206
rect 6880 7160 6960 7188
rect 6828 7142 6880 7148
rect 6932 6361 6960 7160
rect 7012 7142 7064 7148
rect 7024 6934 7052 7142
rect 7668 7002 7696 7346
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 7760 6798 7788 8774
rect 7852 8498 7880 8774
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7944 8242 7972 8996
rect 8036 8362 8064 11342
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 8128 10266 8156 11018
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8220 10146 8248 11494
rect 8128 10118 8248 10146
rect 8128 8401 8156 10118
rect 8312 9450 8340 14350
rect 8392 14000 8444 14006
rect 8392 13942 8444 13948
rect 8404 11014 8432 13942
rect 8496 13818 8524 14776
rect 8666 14719 8722 14728
rect 8574 14512 8630 14521
rect 8574 14447 8630 14456
rect 8588 13938 8616 14447
rect 8680 13938 8708 14719
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 8496 13790 8616 13818
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8496 13326 8524 13670
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 8404 8945 8432 10542
rect 8496 10130 8524 13262
rect 8588 12850 8616 13790
rect 8668 13796 8720 13802
rect 8668 13738 8720 13744
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8588 11529 8616 12242
rect 8680 11665 8708 13738
rect 8772 13530 8800 14878
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8864 14346 8892 14758
rect 8956 14550 8984 16759
rect 9140 16250 9168 17138
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 8944 14544 8996 14550
rect 8944 14486 8996 14492
rect 9048 14498 9076 16050
rect 9128 15632 9180 15638
rect 9128 15574 9180 15580
rect 9140 14618 9168 15574
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 8852 14340 8904 14346
rect 8852 14282 8904 14288
rect 8852 13728 8904 13734
rect 8956 13716 8984 14486
rect 9048 14470 9168 14498
rect 9036 13728 9088 13734
rect 8956 13688 9036 13716
rect 8852 13670 8904 13676
rect 9036 13670 9088 13676
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8864 13258 8892 13670
rect 9140 13546 9168 14470
rect 9048 13518 9168 13546
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8772 12714 8800 12786
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8666 11656 8722 11665
rect 8666 11591 8722 11600
rect 8668 11552 8720 11558
rect 8574 11520 8630 11529
rect 8668 11494 8720 11500
rect 8574 11455 8630 11464
rect 8680 11393 8708 11494
rect 8666 11384 8722 11393
rect 8666 11319 8722 11328
rect 8772 11268 8800 12038
rect 8574 11248 8630 11257
rect 8574 11183 8630 11192
rect 8680 11240 8800 11268
rect 8588 11150 8616 11183
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8680 10849 8708 11240
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 8666 10840 8722 10849
rect 8666 10775 8722 10784
rect 8574 10296 8630 10305
rect 8574 10231 8630 10240
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8588 9704 8616 10231
rect 8496 9676 8616 9704
rect 8496 9353 8524 9676
rect 8574 9616 8630 9625
rect 8574 9551 8630 9560
rect 8482 9344 8538 9353
rect 8482 9279 8538 9288
rect 8390 8936 8446 8945
rect 8208 8900 8260 8906
rect 8390 8871 8446 8880
rect 8208 8842 8260 8848
rect 8220 8498 8248 8842
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8392 8424 8444 8430
rect 8114 8392 8170 8401
rect 8024 8356 8076 8362
rect 8392 8366 8444 8372
rect 8114 8327 8170 8336
rect 8024 8298 8076 8304
rect 8116 8288 8168 8294
rect 7944 8214 8064 8242
rect 8404 8265 8432 8366
rect 8484 8288 8536 8294
rect 8116 8230 8168 8236
rect 8206 8256 8262 8265
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7840 8016 7892 8022
rect 7840 7958 7892 7964
rect 7852 7410 7880 7958
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7944 7002 7972 8026
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 6918 6352 6974 6361
rect 6918 6287 6974 6296
rect 7378 6352 7434 6361
rect 7378 6287 7434 6296
rect 7102 6080 7158 6089
rect 7102 6015 7158 6024
rect 7116 5642 7144 6015
rect 7392 5710 7420 6287
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7104 5636 7156 5642
rect 7104 5578 7156 5584
rect 8036 5098 8064 8214
rect 8128 7954 8156 8230
rect 8206 8191 8262 8200
rect 8390 8256 8446 8265
rect 8484 8230 8536 8236
rect 8390 8191 8446 8200
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8128 7410 8156 7890
rect 8220 7585 8248 8191
rect 8496 7886 8524 8230
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8206 7576 8262 7585
rect 8206 7511 8262 7520
rect 8220 7410 8248 7511
rect 8496 7410 8524 7822
rect 8588 7410 8616 9551
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 8206 6760 8262 6769
rect 8206 6695 8262 6704
rect 8220 5914 8248 6695
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8220 5302 8248 5850
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 8312 5166 8340 5510
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 8404 5030 8432 5510
rect 8496 5234 8524 5782
rect 8680 5710 8708 10775
rect 8772 9489 8800 11086
rect 8864 9926 8892 13194
rect 8942 13152 8998 13161
rect 8942 13087 8998 13096
rect 8956 12850 8984 13087
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8956 9738 8984 11154
rect 9048 10810 9076 13518
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9140 12238 9168 12582
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9126 11792 9182 11801
rect 9126 11727 9182 11736
rect 9140 11558 9168 11727
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 9036 9988 9088 9994
rect 9036 9930 9088 9936
rect 8864 9710 8984 9738
rect 8758 9480 8814 9489
rect 8758 9415 8814 9424
rect 8864 9353 8892 9710
rect 8944 9648 8996 9654
rect 8942 9616 8944 9625
rect 8996 9616 8998 9625
rect 8942 9551 8998 9560
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8850 9344 8906 9353
rect 8850 9279 8906 9288
rect 8758 9072 8814 9081
rect 8758 9007 8814 9016
rect 8772 8634 8800 9007
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8758 8528 8814 8537
rect 8758 8463 8814 8472
rect 8852 8492 8904 8498
rect 8772 7392 8800 8463
rect 8852 8434 8904 8440
rect 8864 8362 8892 8434
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8864 8090 8892 8298
rect 8956 8090 8984 9454
rect 9048 9178 9076 9930
rect 9140 9625 9168 10950
rect 9232 10266 9260 18634
rect 9324 15638 9352 20975
rect 9416 20058 9444 22170
rect 9508 21865 9536 22494
rect 9680 22432 9732 22438
rect 9680 22374 9732 22380
rect 9692 22114 9720 22374
rect 9600 22086 9720 22114
rect 9600 22030 9628 22086
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9680 22024 9732 22030
rect 9680 21966 9732 21972
rect 9494 21856 9550 21865
rect 9494 21791 9550 21800
rect 9692 21622 9720 21966
rect 9680 21616 9732 21622
rect 9680 21558 9732 21564
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9496 21412 9548 21418
rect 9496 21354 9548 21360
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 9416 19718 9444 19994
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 9416 18290 9444 19654
rect 9508 18766 9536 21354
rect 9600 20233 9628 21490
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 9692 20924 9720 21286
rect 9784 20992 9812 22646
rect 9876 22438 9904 24919
rect 9956 24890 10008 24896
rect 9968 24614 9996 24890
rect 10048 24880 10100 24886
rect 10152 24857 10180 25094
rect 10048 24822 10100 24828
rect 10138 24848 10194 24857
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 9956 24064 10008 24070
rect 9956 24006 10008 24012
rect 9968 23662 9996 24006
rect 9956 23656 10008 23662
rect 9956 23598 10008 23604
rect 9956 22568 10008 22574
rect 9956 22510 10008 22516
rect 9864 22432 9916 22438
rect 9968 22409 9996 22510
rect 9864 22374 9916 22380
rect 9954 22400 10010 22409
rect 9954 22335 10010 22344
rect 9968 22094 9996 22335
rect 9876 22066 9996 22094
rect 9876 22030 9904 22066
rect 9864 22024 9916 22030
rect 9864 21966 9916 21972
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9876 21350 9904 21830
rect 9864 21344 9916 21350
rect 9864 21286 9916 21292
rect 9784 20964 9904 20992
rect 9692 20896 9812 20924
rect 9784 20754 9812 20896
rect 9876 20874 9904 20964
rect 9864 20868 9916 20874
rect 9864 20810 9916 20816
rect 9862 20768 9918 20777
rect 9784 20726 9862 20754
rect 9862 20703 9918 20712
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 9586 20224 9642 20233
rect 9586 20159 9642 20168
rect 9680 19916 9732 19922
rect 9784 19904 9812 20538
rect 9864 20256 9916 20262
rect 9864 20198 9916 20204
rect 9732 19876 9812 19904
rect 9680 19858 9732 19864
rect 9772 19780 9824 19786
rect 9772 19722 9824 19728
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9312 15632 9364 15638
rect 9312 15574 9364 15580
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9324 15026 9352 15302
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9324 14074 9352 14350
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9324 13841 9352 13874
rect 9310 13832 9366 13841
rect 9310 13767 9366 13776
rect 9310 13696 9366 13705
rect 9310 13631 9366 13640
rect 9324 13161 9352 13631
rect 9416 13410 9444 18226
rect 9600 16674 9628 19654
rect 9678 19544 9734 19553
rect 9678 19479 9734 19488
rect 9692 19446 9720 19479
rect 9680 19440 9732 19446
rect 9680 19382 9732 19388
rect 9678 19272 9734 19281
rect 9678 19207 9734 19216
rect 9692 18766 9720 19207
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9692 17241 9720 17682
rect 9678 17232 9734 17241
rect 9678 17167 9734 17176
rect 9784 17116 9812 19722
rect 9876 18601 9904 20198
rect 9968 19718 9996 21966
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 9956 19440 10008 19446
rect 9956 19382 10008 19388
rect 9968 19242 9996 19382
rect 9956 19236 10008 19242
rect 9956 19178 10008 19184
rect 10060 18902 10088 24822
rect 10138 24783 10194 24792
rect 10140 24268 10192 24274
rect 10140 24210 10192 24216
rect 10152 23798 10180 24210
rect 10140 23792 10192 23798
rect 10140 23734 10192 23740
rect 10244 22642 10272 26726
rect 10336 25906 10364 27832
rect 10416 27814 10468 27820
rect 10520 27452 10548 28494
rect 10612 27849 10640 29106
rect 10692 28960 10744 28966
rect 10692 28902 10744 28908
rect 10784 28960 10836 28966
rect 10784 28902 10836 28908
rect 10598 27840 10654 27849
rect 10598 27775 10654 27784
rect 10600 27464 10652 27470
rect 10520 27424 10600 27452
rect 10600 27406 10652 27412
rect 10416 27396 10468 27402
rect 10416 27338 10468 27344
rect 10428 27130 10456 27338
rect 10416 27124 10468 27130
rect 10416 27066 10468 27072
rect 10416 26920 10468 26926
rect 10416 26862 10468 26868
rect 10324 25900 10376 25906
rect 10324 25842 10376 25848
rect 10428 25786 10456 26862
rect 10506 26208 10562 26217
rect 10506 26143 10562 26152
rect 10520 25906 10548 26143
rect 10508 25900 10560 25906
rect 10508 25842 10560 25848
rect 10336 25758 10456 25786
rect 10336 23780 10364 25758
rect 10508 25288 10560 25294
rect 10508 25230 10560 25236
rect 10416 25152 10468 25158
rect 10416 25094 10468 25100
rect 10428 23905 10456 25094
rect 10520 24993 10548 25230
rect 10506 24984 10562 24993
rect 10506 24919 10562 24928
rect 10612 24206 10640 27406
rect 10704 26382 10732 28902
rect 10796 28762 10824 28902
rect 10784 28756 10836 28762
rect 10784 28698 10836 28704
rect 10796 28558 10824 28698
rect 10784 28552 10836 28558
rect 10784 28494 10836 28500
rect 10876 28552 10928 28558
rect 10876 28494 10928 28500
rect 10782 28112 10838 28121
rect 10782 28047 10784 28056
rect 10836 28047 10838 28056
rect 10784 28018 10836 28024
rect 10888 27878 10916 28494
rect 10876 27872 10928 27878
rect 10782 27840 10838 27849
rect 10876 27814 10928 27820
rect 10782 27775 10838 27784
rect 10796 26790 10824 27775
rect 10888 27402 10916 27814
rect 10980 27606 11008 29106
rect 11152 29096 11204 29102
rect 11152 29038 11204 29044
rect 11164 28694 11192 29038
rect 11244 29028 11296 29034
rect 11244 28970 11296 28976
rect 11152 28688 11204 28694
rect 11152 28630 11204 28636
rect 11058 28520 11114 28529
rect 11058 28455 11114 28464
rect 11072 28422 11100 28455
rect 11060 28416 11112 28422
rect 11060 28358 11112 28364
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 11072 27674 11100 28154
rect 11256 28150 11284 28970
rect 11520 28960 11572 28966
rect 11520 28902 11572 28908
rect 11532 28558 11560 28902
rect 11428 28552 11480 28558
rect 11428 28494 11480 28500
rect 11520 28552 11572 28558
rect 11520 28494 11572 28500
rect 11334 28384 11390 28393
rect 11334 28319 11390 28328
rect 11244 28144 11296 28150
rect 11244 28086 11296 28092
rect 11152 28076 11204 28082
rect 11152 28018 11204 28024
rect 11164 27849 11192 28018
rect 11244 28008 11296 28014
rect 11244 27950 11296 27956
rect 11150 27840 11206 27849
rect 11150 27775 11206 27784
rect 11060 27668 11112 27674
rect 11060 27610 11112 27616
rect 10968 27600 11020 27606
rect 10968 27542 11020 27548
rect 11058 27568 11114 27577
rect 10876 27396 10928 27402
rect 10876 27338 10928 27344
rect 10784 26784 10836 26790
rect 10784 26726 10836 26732
rect 10796 26625 10824 26726
rect 10782 26616 10838 26625
rect 10782 26551 10838 26560
rect 10692 26376 10744 26382
rect 10692 26318 10744 26324
rect 10784 26376 10836 26382
rect 10784 26318 10836 26324
rect 10704 25129 10732 26318
rect 10796 25702 10824 26318
rect 10784 25696 10836 25702
rect 10784 25638 10836 25644
rect 10690 25120 10746 25129
rect 10690 25055 10746 25064
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 10704 24206 10732 24550
rect 10508 24200 10560 24206
rect 10508 24142 10560 24148
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10692 24200 10744 24206
rect 10692 24142 10744 24148
rect 10414 23896 10470 23905
rect 10414 23831 10470 23840
rect 10336 23752 10456 23780
rect 10324 23656 10376 23662
rect 10324 23598 10376 23604
rect 10428 23610 10456 23752
rect 10520 23730 10548 24142
rect 10612 23848 10640 24142
rect 10784 24132 10836 24138
rect 10888 24120 10916 27338
rect 10980 26994 11008 27542
rect 11058 27503 11114 27512
rect 11072 27334 11100 27503
rect 11060 27328 11112 27334
rect 11060 27270 11112 27276
rect 11152 27328 11204 27334
rect 11152 27270 11204 27276
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 11060 26988 11112 26994
rect 11060 26930 11112 26936
rect 11072 26897 11100 26930
rect 11058 26888 11114 26897
rect 11058 26823 11114 26832
rect 11060 26512 11112 26518
rect 11060 26454 11112 26460
rect 10966 25800 11022 25809
rect 10966 25735 11022 25744
rect 10980 25702 11008 25735
rect 10968 25696 11020 25702
rect 10968 25638 11020 25644
rect 10836 24092 10916 24120
rect 10784 24074 10836 24080
rect 10980 24018 11008 25638
rect 10796 23990 11008 24018
rect 10692 23860 10744 23866
rect 10612 23820 10692 23848
rect 10692 23802 10744 23808
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10232 22636 10284 22642
rect 10232 22578 10284 22584
rect 10140 22160 10192 22166
rect 10140 22102 10192 22108
rect 10048 18896 10100 18902
rect 10048 18838 10100 18844
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 9862 18592 9918 18601
rect 9862 18527 9918 18536
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 9876 17270 9904 18362
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 9864 17128 9916 17134
rect 9784 17088 9864 17116
rect 9864 17070 9916 17076
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9784 16726 9812 16934
rect 9772 16720 9824 16726
rect 9600 16646 9720 16674
rect 9772 16662 9824 16668
rect 9876 16658 9904 17070
rect 9968 16969 9996 18634
rect 10152 17354 10180 22102
rect 10232 21344 10284 21350
rect 10232 21286 10284 21292
rect 10244 20806 10272 21286
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 10230 19952 10286 19961
rect 10230 19887 10232 19896
rect 10284 19887 10286 19896
rect 10232 19858 10284 19864
rect 10232 19372 10284 19378
rect 10232 19314 10284 19320
rect 10244 18970 10272 19314
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 10336 18766 10364 23598
rect 10428 23582 10640 23610
rect 10414 23216 10470 23225
rect 10414 23151 10470 23160
rect 10428 21729 10456 23151
rect 10506 22808 10562 22817
rect 10506 22743 10562 22752
rect 10520 22710 10548 22743
rect 10508 22704 10560 22710
rect 10508 22646 10560 22652
rect 10520 21894 10548 22646
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 10414 21720 10470 21729
rect 10414 21655 10470 21664
rect 10508 21616 10560 21622
rect 10414 21584 10470 21593
rect 10508 21558 10560 21564
rect 10414 21519 10470 21528
rect 10428 21486 10456 21519
rect 10416 21480 10468 21486
rect 10416 21422 10468 21428
rect 10428 21010 10456 21422
rect 10520 21146 10548 21558
rect 10508 21140 10560 21146
rect 10508 21082 10560 21088
rect 10416 21004 10468 21010
rect 10416 20946 10468 20952
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10520 20602 10548 20946
rect 10508 20596 10560 20602
rect 10508 20538 10560 20544
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10428 17678 10456 20402
rect 10506 20360 10562 20369
rect 10506 20295 10508 20304
rect 10560 20295 10562 20304
rect 10508 20266 10560 20272
rect 10508 19848 10560 19854
rect 10508 19790 10560 19796
rect 10520 19514 10548 19790
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10506 19000 10562 19009
rect 10506 18935 10508 18944
rect 10560 18935 10562 18944
rect 10508 18906 10560 18912
rect 10612 18902 10640 23582
rect 10796 23118 10824 23990
rect 10968 23724 11020 23730
rect 10968 23666 11020 23672
rect 10980 23497 11008 23666
rect 10966 23488 11022 23497
rect 10966 23423 11022 23432
rect 11072 23118 11100 26454
rect 11164 25514 11192 27270
rect 11256 27062 11284 27950
rect 11348 27606 11376 28319
rect 11440 28218 11468 28494
rect 11612 28484 11664 28490
rect 11612 28426 11664 28432
rect 11428 28212 11480 28218
rect 11428 28154 11480 28160
rect 11520 28076 11572 28082
rect 11520 28018 11572 28024
rect 11428 27940 11480 27946
rect 11428 27882 11480 27888
rect 11440 27713 11468 27882
rect 11426 27704 11482 27713
rect 11426 27639 11482 27648
rect 11336 27600 11388 27606
rect 11336 27542 11388 27548
rect 11532 27470 11560 28018
rect 11336 27464 11388 27470
rect 11336 27406 11388 27412
rect 11520 27464 11572 27470
rect 11520 27406 11572 27412
rect 11348 27169 11376 27406
rect 11428 27328 11480 27334
rect 11428 27270 11480 27276
rect 11334 27160 11390 27169
rect 11334 27095 11390 27104
rect 11244 27056 11296 27062
rect 11244 26998 11296 27004
rect 11242 26888 11298 26897
rect 11242 26823 11298 26832
rect 11256 26382 11284 26823
rect 11244 26376 11296 26382
rect 11244 26318 11296 26324
rect 11440 26314 11468 27270
rect 11428 26308 11480 26314
rect 11428 26250 11480 26256
rect 11520 26308 11572 26314
rect 11520 26250 11572 26256
rect 11336 26240 11388 26246
rect 11336 26182 11388 26188
rect 11348 25906 11376 26182
rect 11440 26042 11468 26250
rect 11428 26036 11480 26042
rect 11428 25978 11480 25984
rect 11532 25974 11560 26250
rect 11520 25968 11572 25974
rect 11520 25910 11572 25916
rect 11336 25900 11388 25906
rect 11336 25842 11388 25848
rect 11428 25900 11480 25906
rect 11428 25842 11480 25848
rect 11164 25486 11376 25514
rect 11440 25498 11468 25842
rect 11520 25832 11572 25838
rect 11520 25774 11572 25780
rect 11244 25424 11296 25430
rect 11244 25366 11296 25372
rect 11152 25356 11204 25362
rect 11152 25298 11204 25304
rect 11164 24410 11192 25298
rect 11256 25294 11284 25366
rect 11244 25288 11296 25294
rect 11244 25230 11296 25236
rect 11152 24404 11204 24410
rect 11152 24346 11204 24352
rect 11256 24206 11284 25230
rect 11348 24614 11376 25486
rect 11428 25492 11480 25498
rect 11428 25434 11480 25440
rect 11532 25294 11560 25774
rect 11428 25288 11480 25294
rect 11428 25230 11480 25236
rect 11520 25288 11572 25294
rect 11520 25230 11572 25236
rect 11336 24608 11388 24614
rect 11336 24550 11388 24556
rect 11244 24200 11296 24206
rect 11244 24142 11296 24148
rect 11150 23896 11206 23905
rect 11150 23831 11206 23840
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 11060 22976 11112 22982
rect 11060 22918 11112 22924
rect 10692 22772 10744 22778
rect 10692 22714 10744 22720
rect 10704 21962 10732 22714
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10692 21956 10744 21962
rect 10692 21898 10744 21904
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10704 21078 10732 21490
rect 10692 21072 10744 21078
rect 10692 21014 10744 21020
rect 10704 19961 10732 21014
rect 10690 19952 10746 19961
rect 10690 19887 10746 19896
rect 10692 19712 10744 19718
rect 10692 19654 10744 19660
rect 10600 18896 10652 18902
rect 10600 18838 10652 18844
rect 10508 18148 10560 18154
rect 10508 18090 10560 18096
rect 10520 18057 10548 18090
rect 10600 18080 10652 18086
rect 10506 18048 10562 18057
rect 10600 18022 10652 18028
rect 10506 17983 10562 17992
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10520 17678 10548 17750
rect 10416 17672 10468 17678
rect 10508 17672 10560 17678
rect 10416 17614 10468 17620
rect 10506 17640 10508 17649
rect 10560 17640 10562 17649
rect 10506 17575 10562 17584
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 10060 17326 10180 17354
rect 9954 16960 10010 16969
rect 9954 16895 10010 16904
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9508 16182 9536 16390
rect 9496 16176 9548 16182
rect 9496 16118 9548 16124
rect 9494 15328 9550 15337
rect 9494 15263 9550 15272
rect 9508 14793 9536 15263
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9600 14822 9628 14962
rect 9588 14816 9640 14822
rect 9494 14784 9550 14793
rect 9588 14758 9640 14764
rect 9494 14719 9550 14728
rect 9494 14648 9550 14657
rect 9494 14583 9550 14592
rect 9508 14550 9536 14583
rect 9692 14550 9720 16646
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9876 16250 9904 16390
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9770 15736 9826 15745
rect 9770 15671 9826 15680
rect 9784 15502 9812 15671
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9496 14544 9548 14550
rect 9496 14486 9548 14492
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9508 13954 9536 14486
rect 9784 14414 9812 15302
rect 9876 15201 9904 16186
rect 9968 15337 9996 16458
rect 10060 15502 10088 17326
rect 10140 17264 10192 17270
rect 10140 17206 10192 17212
rect 10152 16250 10180 17206
rect 10244 17134 10272 17478
rect 10336 17338 10364 17478
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10230 16960 10286 16969
rect 10230 16895 10286 16904
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10244 15638 10272 16895
rect 10428 16794 10456 17138
rect 10520 16833 10548 17138
rect 10506 16824 10562 16833
rect 10416 16788 10468 16794
rect 10506 16759 10562 16768
rect 10416 16730 10468 16736
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 9954 15328 10010 15337
rect 10138 15328 10194 15337
rect 9954 15263 10010 15272
rect 10060 15286 10138 15314
rect 9862 15192 9918 15201
rect 9862 15127 9918 15136
rect 10060 15094 10088 15286
rect 10138 15263 10194 15272
rect 10048 15088 10100 15094
rect 9968 15048 10048 15076
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9876 14657 9904 14758
rect 9862 14648 9918 14657
rect 9862 14583 9918 14592
rect 9968 14482 9996 15048
rect 10048 15030 10100 15036
rect 10244 15008 10272 15574
rect 10336 15366 10364 15846
rect 10416 15632 10468 15638
rect 10416 15574 10468 15580
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10428 15178 10456 15574
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10336 15150 10456 15178
rect 10336 15026 10364 15150
rect 10198 14980 10272 15008
rect 10324 15020 10376 15026
rect 10198 14940 10226 14980
rect 10324 14962 10376 14968
rect 10060 14912 10226 14940
rect 10060 14822 10088 14912
rect 10329 14906 10357 14962
rect 10329 14878 10364 14906
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9772 14408 9824 14414
rect 10232 14408 10284 14414
rect 9772 14350 9824 14356
rect 10138 14376 10194 14385
rect 9508 13938 9628 13954
rect 9508 13932 9640 13938
rect 9508 13926 9588 13932
rect 9588 13874 9640 13880
rect 9496 13864 9548 13870
rect 9494 13832 9496 13841
rect 9548 13832 9550 13841
rect 9494 13767 9550 13776
rect 9586 13696 9642 13705
rect 9586 13631 9642 13640
rect 9600 13530 9628 13631
rect 9784 13530 9812 14350
rect 9956 14340 10008 14346
rect 10232 14350 10284 14356
rect 10138 14311 10194 14320
rect 9956 14282 10008 14288
rect 9862 14240 9918 14249
rect 9862 14175 9918 14184
rect 9876 13938 9904 14175
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9862 13832 9918 13841
rect 9862 13767 9918 13776
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9416 13382 9628 13410
rect 9310 13152 9366 13161
rect 9310 13087 9366 13096
rect 9494 13152 9550 13161
rect 9494 13087 9550 13096
rect 9508 12850 9536 13087
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9312 12776 9364 12782
rect 9310 12744 9312 12753
rect 9364 12744 9366 12753
rect 9310 12679 9366 12688
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9496 12640 9548 12646
rect 9600 12628 9628 13382
rect 9876 13326 9904 13767
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9876 12850 9904 13262
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9678 12744 9734 12753
rect 9862 12744 9918 12753
rect 9734 12714 9812 12730
rect 9734 12708 9824 12714
rect 9734 12702 9772 12708
rect 9678 12679 9734 12688
rect 9862 12679 9918 12688
rect 9772 12650 9824 12656
rect 9600 12600 9720 12628
rect 9496 12582 9548 12588
rect 9324 12442 9352 12582
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9508 12356 9536 12582
rect 9463 12328 9536 12356
rect 9463 12322 9491 12328
rect 9324 12294 9491 12322
rect 9324 12238 9352 12294
rect 9692 12238 9720 12600
rect 9770 12608 9826 12617
rect 9770 12543 9826 12552
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9324 11150 9352 12174
rect 9404 12096 9456 12102
rect 9680 12096 9732 12102
rect 9404 12038 9456 12044
rect 9586 12064 9642 12073
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9312 10736 9364 10742
rect 9416 10713 9444 12038
rect 9680 12038 9732 12044
rect 9586 11999 9642 12008
rect 9600 11762 9628 11999
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9692 11694 9720 12038
rect 9680 11688 9732 11694
rect 9494 11656 9550 11665
rect 9680 11630 9732 11636
rect 9494 11591 9550 11600
rect 9312 10678 9364 10684
rect 9402 10704 9458 10713
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9324 9722 9352 10678
rect 9402 10639 9458 10648
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9126 9616 9182 9625
rect 9126 9551 9182 9560
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 9140 8974 9168 9386
rect 9232 9178 9260 9658
rect 9416 9353 9444 10406
rect 9508 10130 9536 11591
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9692 11354 9720 11494
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9600 10266 9628 10542
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9692 10062 9720 10406
rect 9680 10056 9732 10062
rect 9494 10024 9550 10033
rect 9680 9998 9732 10004
rect 9494 9959 9550 9968
rect 9508 9518 9536 9959
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9402 9344 9458 9353
rect 9402 9279 9458 9288
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9508 9058 9536 9454
rect 9232 9030 9536 9058
rect 9232 8974 9260 9030
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9220 8968 9272 8974
rect 9496 8968 9548 8974
rect 9220 8910 9272 8916
rect 9402 8936 9458 8945
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 9048 8498 9076 8842
rect 9232 8786 9260 8910
rect 9496 8910 9548 8916
rect 9402 8871 9404 8880
rect 9456 8871 9458 8880
rect 9404 8842 9456 8848
rect 9140 8758 9260 8786
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9034 8392 9090 8401
rect 9034 8327 9090 8336
rect 9048 8090 9076 8327
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8956 7410 8984 7822
rect 8852 7404 8904 7410
rect 8772 7364 8852 7392
rect 8852 7346 8904 7352
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 8956 7274 8984 7346
rect 8944 7268 8996 7274
rect 8944 7210 8996 7216
rect 9048 7206 9076 7346
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9140 5710 9168 8758
rect 9220 8628 9272 8634
rect 9508 8616 9536 8910
rect 9220 8570 9272 8576
rect 9416 8588 9536 8616
rect 9232 8265 9260 8570
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9218 8256 9274 8265
rect 9218 8191 9274 8200
rect 9232 7886 9260 8191
rect 9324 8022 9352 8502
rect 9416 8362 9444 8588
rect 9600 8537 9628 9454
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9692 8906 9720 9318
rect 9784 9042 9812 12543
rect 9876 10062 9904 12679
rect 9968 11898 9996 14282
rect 10152 13938 10180 14311
rect 10244 14074 10272 14350
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10060 13274 10088 13670
rect 10152 13394 10180 13670
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10060 13258 10180 13274
rect 10060 13252 10192 13258
rect 10060 13246 10140 13252
rect 10140 13194 10192 13200
rect 10046 12880 10102 12889
rect 10046 12815 10048 12824
rect 10100 12815 10102 12824
rect 10048 12786 10100 12792
rect 10048 12640 10100 12646
rect 10152 12617 10180 13194
rect 10048 12582 10100 12588
rect 10138 12608 10194 12617
rect 10060 12458 10088 12582
rect 10138 12543 10194 12552
rect 10244 12458 10272 13466
rect 10060 12430 10272 12458
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9956 11688 10008 11694
rect 10060 11665 10088 11698
rect 9956 11630 10008 11636
rect 10046 11656 10102 11665
rect 9968 11558 9996 11630
rect 10046 11591 10102 11600
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 10152 10674 10180 12430
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 10244 11898 10272 12242
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10232 11144 10284 11150
rect 10230 11112 10232 11121
rect 10284 11112 10286 11121
rect 10230 11047 10286 11056
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9692 8566 9720 8842
rect 9876 8838 9904 9522
rect 9968 8974 9996 10610
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 10060 9722 10088 9930
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9864 8832 9916 8838
rect 10060 8809 10088 9522
rect 10152 9110 10180 10202
rect 10230 10024 10286 10033
rect 10336 9994 10364 14878
rect 10414 14376 10470 14385
rect 10414 14311 10470 14320
rect 10428 14278 10456 14311
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10428 12918 10456 14010
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10520 12753 10548 15506
rect 10612 15502 10640 18022
rect 10704 16794 10732 19654
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10796 16114 10824 22374
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10888 21321 10916 21966
rect 10980 21962 11008 22510
rect 10968 21956 11020 21962
rect 10968 21898 11020 21904
rect 11072 21842 11100 22918
rect 11164 22098 11192 23831
rect 11244 22976 11296 22982
rect 11244 22918 11296 22924
rect 11256 22642 11284 22918
rect 11244 22636 11296 22642
rect 11244 22578 11296 22584
rect 11152 22092 11204 22098
rect 11152 22034 11204 22040
rect 11244 21888 11296 21894
rect 11072 21814 11192 21842
rect 11244 21830 11296 21836
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 10966 21584 11022 21593
rect 10966 21519 10968 21528
rect 11020 21519 11022 21528
rect 10968 21490 11020 21496
rect 11072 21434 11100 21626
rect 10980 21406 11100 21434
rect 10874 21312 10930 21321
rect 10874 21247 10930 21256
rect 10876 20392 10928 20398
rect 10876 20334 10928 20340
rect 10888 19446 10916 20334
rect 10876 19440 10928 19446
rect 10876 19382 10928 19388
rect 10874 19272 10930 19281
rect 10874 19207 10930 19216
rect 10888 18358 10916 19207
rect 10980 19174 11008 21406
rect 11058 20768 11114 20777
rect 11058 20703 11114 20712
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 11072 18850 11100 20703
rect 11164 20330 11192 21814
rect 11256 21146 11284 21830
rect 11244 21140 11296 21146
rect 11244 21082 11296 21088
rect 11152 20324 11204 20330
rect 11152 20266 11204 20272
rect 11256 20262 11284 21082
rect 11244 20256 11296 20262
rect 11244 20198 11296 20204
rect 11348 20074 11376 24550
rect 11440 24410 11468 25230
rect 11624 25106 11652 28426
rect 11716 27130 11744 29718
rect 12716 29164 12768 29170
rect 12716 29106 12768 29112
rect 13268 29164 13320 29170
rect 13268 29106 13320 29112
rect 12072 29028 12124 29034
rect 12072 28970 12124 28976
rect 11980 28960 12032 28966
rect 11980 28902 12032 28908
rect 11888 28688 11940 28694
rect 11888 28630 11940 28636
rect 11900 27849 11928 28630
rect 11992 28558 12020 28902
rect 12084 28694 12112 28970
rect 12452 28966 12664 28994
rect 12452 28762 12480 28966
rect 12530 28928 12586 28937
rect 12530 28863 12586 28872
rect 12544 28762 12572 28863
rect 12440 28756 12492 28762
rect 12440 28698 12492 28704
rect 12532 28756 12584 28762
rect 12532 28698 12584 28704
rect 12072 28688 12124 28694
rect 12072 28630 12124 28636
rect 12346 28656 12402 28665
rect 12530 28656 12586 28665
rect 12402 28614 12480 28642
rect 12346 28591 12402 28600
rect 11980 28552 12032 28558
rect 11980 28494 12032 28500
rect 12348 28552 12400 28558
rect 12348 28494 12400 28500
rect 11980 28416 12032 28422
rect 11980 28358 12032 28364
rect 11886 27840 11942 27849
rect 11886 27775 11942 27784
rect 11794 27704 11850 27713
rect 11794 27639 11850 27648
rect 11808 27384 11836 27639
rect 11992 27470 12020 28358
rect 12164 27872 12216 27878
rect 12164 27814 12216 27820
rect 12256 27872 12308 27878
rect 12256 27814 12308 27820
rect 11980 27464 12032 27470
rect 11980 27406 12032 27412
rect 11888 27396 11940 27402
rect 11808 27356 11888 27384
rect 11808 27130 11836 27356
rect 11888 27338 11940 27344
rect 11704 27124 11756 27130
rect 11704 27066 11756 27072
rect 11796 27124 11848 27130
rect 11796 27066 11848 27072
rect 11704 26376 11756 26382
rect 11808 26364 11836 27066
rect 11756 26336 11836 26364
rect 11888 26376 11940 26382
rect 11704 26318 11756 26324
rect 11888 26318 11940 26324
rect 11716 25838 11744 26318
rect 11900 26246 11928 26318
rect 11888 26240 11940 26246
rect 11888 26182 11940 26188
rect 11796 26036 11848 26042
rect 11796 25978 11848 25984
rect 11704 25832 11756 25838
rect 11704 25774 11756 25780
rect 11704 25424 11756 25430
rect 11704 25366 11756 25372
rect 11532 25078 11652 25106
rect 11532 24954 11560 25078
rect 11520 24948 11572 24954
rect 11520 24890 11572 24896
rect 11532 24818 11560 24890
rect 11716 24818 11744 25366
rect 11808 25294 11836 25978
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11796 25152 11848 25158
rect 11796 25094 11848 25100
rect 11808 24818 11836 25094
rect 11520 24812 11572 24818
rect 11520 24754 11572 24760
rect 11704 24812 11756 24818
rect 11704 24754 11756 24760
rect 11796 24812 11848 24818
rect 11796 24754 11848 24760
rect 11520 24676 11572 24682
rect 11520 24618 11572 24624
rect 11428 24404 11480 24410
rect 11428 24346 11480 24352
rect 11440 24070 11468 24346
rect 11532 24342 11560 24618
rect 11520 24336 11572 24342
rect 11520 24278 11572 24284
rect 11428 24064 11480 24070
rect 11428 24006 11480 24012
rect 11440 23798 11468 24006
rect 11428 23792 11480 23798
rect 11428 23734 11480 23740
rect 11532 23202 11560 24278
rect 11716 23866 11744 24754
rect 11888 24132 11940 24138
rect 11940 24092 12020 24120
rect 11888 24074 11940 24080
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11704 23860 11756 23866
rect 11624 23820 11704 23848
rect 11624 23730 11652 23820
rect 11704 23802 11756 23808
rect 11612 23724 11664 23730
rect 11612 23666 11664 23672
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 11716 23526 11744 23666
rect 11808 23633 11836 24006
rect 11992 23730 12020 24092
rect 12072 23860 12124 23866
rect 12072 23802 12124 23808
rect 12084 23769 12112 23802
rect 12070 23760 12126 23769
rect 11888 23724 11940 23730
rect 11888 23666 11940 23672
rect 11980 23724 12032 23730
rect 12070 23695 12126 23704
rect 11980 23666 12032 23672
rect 11794 23624 11850 23633
rect 11794 23559 11850 23568
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 11612 23316 11664 23322
rect 11612 23258 11664 23264
rect 11440 23174 11560 23202
rect 11440 22574 11468 23174
rect 11518 23080 11574 23089
rect 11518 23015 11520 23024
rect 11572 23015 11574 23024
rect 11520 22986 11572 22992
rect 11624 22778 11652 23258
rect 11796 23248 11848 23254
rect 11900 23225 11928 23666
rect 11796 23190 11848 23196
rect 11886 23216 11942 23225
rect 11704 22976 11756 22982
rect 11704 22918 11756 22924
rect 11612 22772 11664 22778
rect 11612 22714 11664 22720
rect 11428 22568 11480 22574
rect 11428 22510 11480 22516
rect 11716 22273 11744 22918
rect 11808 22438 11836 23190
rect 11886 23151 11942 23160
rect 11980 23112 12032 23118
rect 11980 23054 12032 23060
rect 11888 22976 11940 22982
rect 11992 22953 12020 23054
rect 12072 23044 12124 23050
rect 12072 22986 12124 22992
rect 11888 22918 11940 22924
rect 11978 22944 12034 22953
rect 11900 22642 11928 22918
rect 11978 22879 12034 22888
rect 12084 22642 12112 22986
rect 11888 22636 11940 22642
rect 11888 22578 11940 22584
rect 12072 22636 12124 22642
rect 12072 22578 12124 22584
rect 12072 22500 12124 22506
rect 12072 22442 12124 22448
rect 11796 22432 11848 22438
rect 11796 22374 11848 22380
rect 11980 22432 12032 22438
rect 11980 22374 12032 22380
rect 11702 22264 11758 22273
rect 11702 22199 11758 22208
rect 11992 22098 12020 22374
rect 11980 22092 12032 22098
rect 11980 22034 12032 22040
rect 11612 22024 11664 22030
rect 11610 21992 11612 22001
rect 11888 22024 11940 22030
rect 11664 21992 11666 22001
rect 12084 22012 12112 22442
rect 12176 22438 12204 27814
rect 12268 27713 12296 27814
rect 12254 27704 12310 27713
rect 12254 27639 12310 27648
rect 12256 27600 12308 27606
rect 12256 27542 12308 27548
rect 12268 27305 12296 27542
rect 12360 27470 12388 28494
rect 12452 28422 12480 28614
rect 12530 28591 12586 28600
rect 12544 28490 12572 28591
rect 12532 28484 12584 28490
rect 12532 28426 12584 28432
rect 12440 28416 12492 28422
rect 12440 28358 12492 28364
rect 12544 28218 12572 28426
rect 12532 28212 12584 28218
rect 12452 28172 12532 28200
rect 12348 27464 12400 27470
rect 12346 27432 12348 27441
rect 12400 27432 12402 27441
rect 12346 27367 12402 27376
rect 12254 27296 12310 27305
rect 12254 27231 12310 27240
rect 12452 27112 12480 28172
rect 12532 28154 12584 28160
rect 12532 28076 12584 28082
rect 12532 28018 12584 28024
rect 12544 27674 12572 28018
rect 12532 27668 12584 27674
rect 12532 27610 12584 27616
rect 12636 27606 12664 28966
rect 12728 28762 12756 29106
rect 12900 29028 12952 29034
rect 12900 28970 12952 28976
rect 12808 28960 12860 28966
rect 12808 28902 12860 28908
rect 12716 28756 12768 28762
rect 12716 28698 12768 28704
rect 12716 28620 12768 28626
rect 12820 28608 12848 28902
rect 12768 28580 12848 28608
rect 12716 28562 12768 28568
rect 12820 28404 12848 28580
rect 12912 28642 12940 28970
rect 13176 28688 13228 28694
rect 13174 28656 13176 28665
rect 13228 28656 13230 28665
rect 12912 28614 13124 28642
rect 12912 28558 12940 28614
rect 12900 28552 12952 28558
rect 12900 28494 12952 28500
rect 12992 28552 13044 28558
rect 12992 28494 13044 28500
rect 12820 28376 12940 28404
rect 12716 28076 12768 28082
rect 12716 28018 12768 28024
rect 12624 27600 12676 27606
rect 12624 27542 12676 27548
rect 12532 27464 12584 27470
rect 12532 27406 12584 27412
rect 12544 27130 12572 27406
rect 12728 27169 12756 28018
rect 12808 28008 12860 28014
rect 12808 27950 12860 27956
rect 12820 27878 12848 27950
rect 12808 27872 12860 27878
rect 12808 27814 12860 27820
rect 12808 27464 12860 27470
rect 12806 27432 12808 27441
rect 12860 27432 12862 27441
rect 12806 27367 12862 27376
rect 12714 27160 12770 27169
rect 12360 27084 12480 27112
rect 12532 27124 12584 27130
rect 12256 26512 12308 26518
rect 12256 26454 12308 26460
rect 12268 25945 12296 26454
rect 12254 25936 12310 25945
rect 12254 25871 12310 25880
rect 12360 25294 12388 27084
rect 12714 27095 12770 27104
rect 12532 27066 12584 27072
rect 12440 26988 12492 26994
rect 12440 26930 12492 26936
rect 12452 25401 12480 26930
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 12532 26036 12584 26042
rect 12532 25978 12584 25984
rect 12438 25392 12494 25401
rect 12438 25327 12494 25336
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12256 25220 12308 25226
rect 12256 25162 12308 25168
rect 12268 24954 12296 25162
rect 12256 24948 12308 24954
rect 12256 24890 12308 24896
rect 12360 24818 12388 25230
rect 12544 25158 12572 25978
rect 12624 25832 12676 25838
rect 12624 25774 12676 25780
rect 12636 25430 12664 25774
rect 12624 25424 12676 25430
rect 12624 25366 12676 25372
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 12532 25152 12584 25158
rect 12532 25094 12584 25100
rect 12636 24970 12664 25230
rect 12544 24942 12664 24970
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 12256 24744 12308 24750
rect 12256 24686 12308 24692
rect 12346 24712 12402 24721
rect 12268 24614 12296 24686
rect 12544 24698 12572 24942
rect 12544 24670 12664 24698
rect 12346 24647 12402 24656
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 12360 23225 12388 24647
rect 12440 24608 12492 24614
rect 12440 24550 12492 24556
rect 12452 23798 12480 24550
rect 12636 24138 12664 24670
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12440 23792 12492 23798
rect 12440 23734 12492 23740
rect 12346 23216 12402 23225
rect 12268 23160 12346 23168
rect 12268 23151 12402 23160
rect 12268 23140 12388 23151
rect 12268 22642 12296 23140
rect 12348 22772 12400 22778
rect 12348 22714 12400 22720
rect 12256 22636 12308 22642
rect 12256 22578 12308 22584
rect 12256 22500 12308 22506
rect 12256 22442 12308 22448
rect 12164 22432 12216 22438
rect 12164 22374 12216 22380
rect 12164 22024 12216 22030
rect 12084 21984 12164 22012
rect 11888 21966 11940 21972
rect 12164 21966 12216 21972
rect 11610 21927 11666 21936
rect 11520 21888 11572 21894
rect 11900 21865 11928 21966
rect 12164 21888 12216 21894
rect 11520 21830 11572 21836
rect 11886 21856 11942 21865
rect 11428 21412 11480 21418
rect 11428 21354 11480 21360
rect 11440 20534 11468 21354
rect 11428 20528 11480 20534
rect 11428 20470 11480 20476
rect 11428 20392 11480 20398
rect 11428 20334 11480 20340
rect 11256 20046 11376 20074
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 11164 19446 11192 19858
rect 11152 19440 11204 19446
rect 11152 19382 11204 19388
rect 11152 19304 11204 19310
rect 11150 19272 11152 19281
rect 11204 19272 11206 19281
rect 11150 19207 11206 19216
rect 11164 18970 11192 19207
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 10980 18822 11100 18850
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 10888 16998 10916 17750
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10980 16810 11008 18822
rect 11256 18766 11284 20046
rect 11440 19258 11468 20334
rect 11532 19846 11560 21830
rect 12164 21830 12216 21836
rect 11886 21791 11942 21800
rect 11704 21684 11756 21690
rect 11704 21626 11756 21632
rect 11612 21548 11664 21554
rect 11612 21490 11664 21496
rect 11624 20330 11652 21490
rect 11716 21010 11744 21626
rect 11794 21584 11850 21593
rect 11794 21519 11796 21528
rect 11848 21519 11850 21528
rect 12072 21548 12124 21554
rect 11796 21490 11848 21496
rect 12072 21490 12124 21496
rect 11980 21412 12032 21418
rect 11980 21354 12032 21360
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11808 21185 11836 21286
rect 11794 21176 11850 21185
rect 11794 21111 11850 21120
rect 11704 21004 11756 21010
rect 11704 20946 11756 20952
rect 11704 20800 11756 20806
rect 11704 20742 11756 20748
rect 11716 20466 11744 20742
rect 11808 20466 11836 21111
rect 11992 20942 12020 21354
rect 11980 20936 12032 20942
rect 11886 20904 11942 20913
rect 11980 20878 12032 20884
rect 11886 20839 11942 20848
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11612 20324 11664 20330
rect 11612 20266 11664 20272
rect 11704 20324 11756 20330
rect 11704 20266 11756 20272
rect 11716 20210 11744 20266
rect 11624 20182 11744 20210
rect 11794 20224 11850 20233
rect 11624 19961 11652 20182
rect 11794 20159 11850 20168
rect 11610 19952 11666 19961
rect 11610 19887 11666 19896
rect 11532 19818 11744 19846
rect 11348 19230 11468 19258
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 11072 18193 11100 18634
rect 11244 18216 11296 18222
rect 11058 18184 11114 18193
rect 11244 18158 11296 18164
rect 11058 18119 11114 18128
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11058 17504 11114 17513
rect 11058 17439 11114 17448
rect 11072 17338 11100 17439
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 11058 17232 11114 17241
rect 11058 17167 11060 17176
rect 11112 17167 11114 17176
rect 11060 17138 11112 17144
rect 10888 16782 11008 16810
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10598 15328 10654 15337
rect 10598 15263 10654 15272
rect 10612 14550 10640 15263
rect 10704 14822 10732 15846
rect 10784 15496 10836 15502
rect 10888 15484 10916 16782
rect 11058 16552 11114 16561
rect 11058 16487 11114 16496
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10836 15456 10916 15484
rect 10784 15438 10836 15444
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10796 15026 10824 15302
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10888 14822 10916 15302
rect 10980 15162 11008 16050
rect 11072 15552 11100 16487
rect 11164 16454 11192 17818
rect 11256 17377 11284 18158
rect 11242 17368 11298 17377
rect 11242 17303 11298 17312
rect 11256 17202 11284 17303
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11348 16574 11376 19230
rect 11532 18290 11560 19246
rect 11716 19224 11744 19818
rect 11808 19786 11836 20159
rect 11900 19961 11928 20839
rect 12084 20806 12112 21490
rect 12176 21010 12204 21830
rect 12164 21004 12216 21010
rect 12164 20946 12216 20952
rect 12072 20800 12124 20806
rect 12072 20742 12124 20748
rect 12084 20346 12112 20742
rect 12268 20466 12296 22442
rect 12360 21962 12388 22714
rect 12348 21956 12400 21962
rect 12348 21898 12400 21904
rect 12346 21584 12402 21593
rect 12346 21519 12402 21528
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 12084 20318 12204 20346
rect 11886 19952 11942 19961
rect 11886 19887 11942 19896
rect 12072 19916 12124 19922
rect 11900 19854 11928 19887
rect 12176 19904 12204 20318
rect 12360 19922 12388 21519
rect 12452 21457 12480 23734
rect 12624 23724 12676 23730
rect 12728 23712 12756 26318
rect 12808 26308 12860 26314
rect 12912 26296 12940 28376
rect 13004 28218 13032 28494
rect 12992 28212 13044 28218
rect 12992 28154 13044 28160
rect 12992 27872 13044 27878
rect 12992 27814 13044 27820
rect 13004 27606 13032 27814
rect 12992 27600 13044 27606
rect 12992 27542 13044 27548
rect 12992 26920 13044 26926
rect 12992 26862 13044 26868
rect 13004 26790 13032 26862
rect 12992 26784 13044 26790
rect 12992 26726 13044 26732
rect 13004 26625 13032 26726
rect 12990 26616 13046 26625
rect 12990 26551 13046 26560
rect 13096 26518 13124 28614
rect 13174 28591 13230 28600
rect 13174 27024 13230 27033
rect 13174 26959 13176 26968
rect 13228 26959 13230 26968
rect 13176 26930 13228 26936
rect 13084 26512 13136 26518
rect 13084 26454 13136 26460
rect 12860 26268 12940 26296
rect 12808 26250 12860 26256
rect 13176 26240 13228 26246
rect 13176 26182 13228 26188
rect 12992 25696 13044 25702
rect 12992 25638 13044 25644
rect 13084 25696 13136 25702
rect 13084 25638 13136 25644
rect 12808 25492 12860 25498
rect 12808 25434 12860 25440
rect 12820 24070 12848 25434
rect 13004 25294 13032 25638
rect 13096 25498 13124 25638
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 12992 25288 13044 25294
rect 12992 25230 13044 25236
rect 13084 25288 13136 25294
rect 13084 25230 13136 25236
rect 12992 25152 13044 25158
rect 12992 25094 13044 25100
rect 13004 24614 13032 25094
rect 13096 24682 13124 25230
rect 13084 24676 13136 24682
rect 13084 24618 13136 24624
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 12898 24440 12954 24449
rect 13004 24410 13032 24550
rect 12898 24375 12954 24384
rect 12992 24404 13044 24410
rect 12808 24064 12860 24070
rect 12808 24006 12860 24012
rect 12676 23684 12756 23712
rect 12624 23666 12676 23672
rect 12530 23624 12586 23633
rect 12530 23559 12586 23568
rect 12544 22506 12572 23559
rect 12636 22982 12664 23666
rect 12806 23488 12862 23497
rect 12806 23423 12862 23432
rect 12820 23118 12848 23423
rect 12808 23112 12860 23118
rect 12808 23054 12860 23060
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12624 22568 12676 22574
rect 12624 22510 12676 22516
rect 12532 22500 12584 22506
rect 12532 22442 12584 22448
rect 12530 22400 12586 22409
rect 12530 22335 12586 22344
rect 12544 22012 12572 22335
rect 12636 22137 12664 22510
rect 12716 22432 12768 22438
rect 12820 22409 12848 23054
rect 12912 22778 12940 24375
rect 12992 24346 13044 24352
rect 13188 24274 13216 26182
rect 13280 24993 13308 29106
rect 13358 28248 13414 28257
rect 13358 28183 13360 28192
rect 13412 28183 13414 28192
rect 13360 28154 13412 28160
rect 13360 27328 13412 27334
rect 13360 27270 13412 27276
rect 13372 27062 13400 27270
rect 13360 27056 13412 27062
rect 13360 26998 13412 27004
rect 13360 26920 13412 26926
rect 13360 26862 13412 26868
rect 13372 26382 13400 26862
rect 13360 26376 13412 26382
rect 13464 26353 13492 30738
rect 13740 28994 13768 30767
rect 14832 30660 14884 30666
rect 14832 30602 14884 30608
rect 14096 30592 14148 30598
rect 14096 30534 14148 30540
rect 14108 30394 14136 30534
rect 14096 30388 14148 30394
rect 14096 30330 14148 30336
rect 14002 29200 14058 29209
rect 14002 29135 14058 29144
rect 13740 28966 13860 28994
rect 13544 28620 13596 28626
rect 13544 28562 13596 28568
rect 13556 27878 13584 28562
rect 13728 28008 13780 28014
rect 13728 27950 13780 27956
rect 13544 27872 13596 27878
rect 13544 27814 13596 27820
rect 13740 27441 13768 27950
rect 13726 27432 13782 27441
rect 13726 27367 13782 27376
rect 13728 27124 13780 27130
rect 13728 27066 13780 27072
rect 13636 27056 13688 27062
rect 13636 26998 13688 27004
rect 13544 26784 13596 26790
rect 13544 26726 13596 26732
rect 13360 26318 13412 26324
rect 13450 26344 13506 26353
rect 13372 26081 13400 26318
rect 13450 26279 13506 26288
rect 13358 26072 13414 26081
rect 13358 26007 13414 26016
rect 13360 25220 13412 25226
rect 13360 25162 13412 25168
rect 13266 24984 13322 24993
rect 13266 24919 13322 24928
rect 13268 24812 13320 24818
rect 13268 24754 13320 24760
rect 13280 24721 13308 24754
rect 13266 24712 13322 24721
rect 13266 24647 13322 24656
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 13084 24132 13136 24138
rect 13084 24074 13136 24080
rect 12992 23860 13044 23866
rect 12992 23802 13044 23808
rect 13004 23730 13032 23802
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 13096 23497 13124 24074
rect 13188 23730 13216 24210
rect 13176 23724 13228 23730
rect 13176 23666 13228 23672
rect 13082 23488 13138 23497
rect 13082 23423 13138 23432
rect 13082 22808 13138 22817
rect 12900 22772 12952 22778
rect 12952 22732 13032 22760
rect 13138 22766 13216 22794
rect 13372 22778 13400 25162
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13464 24585 13492 24754
rect 13450 24576 13506 24585
rect 13450 24511 13506 24520
rect 13450 23352 13506 23361
rect 13450 23287 13506 23296
rect 13464 23118 13492 23287
rect 13452 23112 13504 23118
rect 13452 23054 13504 23060
rect 13082 22743 13138 22752
rect 12900 22714 12952 22720
rect 12900 22500 12952 22506
rect 12900 22442 12952 22448
rect 12716 22374 12768 22380
rect 12806 22400 12862 22409
rect 12728 22234 12756 22374
rect 12806 22335 12862 22344
rect 12716 22228 12768 22234
rect 12716 22170 12768 22176
rect 12808 22228 12860 22234
rect 12808 22170 12860 22176
rect 12622 22128 12678 22137
rect 12622 22063 12678 22072
rect 12624 22024 12676 22030
rect 12544 21984 12624 22012
rect 12624 21966 12676 21972
rect 12820 21842 12848 22170
rect 12728 21814 12848 21842
rect 12624 21480 12676 21486
rect 12438 21448 12494 21457
rect 12438 21383 12494 21392
rect 12622 21448 12624 21457
rect 12676 21448 12678 21457
rect 12622 21383 12678 21392
rect 12636 21010 12664 21383
rect 12728 21350 12756 21814
rect 12806 21720 12862 21729
rect 12806 21655 12862 21664
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12820 21146 12848 21655
rect 12912 21554 12940 22442
rect 13004 22438 13032 22732
rect 13084 22704 13136 22710
rect 13084 22646 13136 22652
rect 12992 22432 13044 22438
rect 12992 22374 13044 22380
rect 12992 22160 13044 22166
rect 12992 22102 13044 22108
rect 13004 21554 13032 22102
rect 13096 22001 13124 22646
rect 13188 22137 13216 22766
rect 13360 22772 13412 22778
rect 13360 22714 13412 22720
rect 13452 22772 13504 22778
rect 13452 22714 13504 22720
rect 13268 22568 13320 22574
rect 13268 22510 13320 22516
rect 13174 22128 13230 22137
rect 13174 22063 13230 22072
rect 13082 21992 13138 22001
rect 13082 21927 13138 21936
rect 13176 21956 13228 21962
rect 13176 21898 13228 21904
rect 12900 21548 12952 21554
rect 12900 21490 12952 21496
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 12898 21448 12954 21457
rect 13188 21434 13216 21898
rect 13280 21690 13308 22510
rect 13360 22432 13412 22438
rect 13360 22374 13412 22380
rect 13268 21684 13320 21690
rect 13268 21626 13320 21632
rect 13372 21554 13400 22374
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13360 21548 13412 21554
rect 13360 21490 13412 21496
rect 12898 21383 12954 21392
rect 13004 21406 13216 21434
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 12808 21140 12860 21146
rect 12808 21082 12860 21088
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 12440 20596 12492 20602
rect 12492 20556 12572 20584
rect 12440 20538 12492 20544
rect 12544 20330 12572 20556
rect 12728 20472 12756 21082
rect 12808 21004 12860 21010
rect 12808 20946 12860 20952
rect 12820 20777 12848 20946
rect 12912 20942 12940 21383
rect 13004 21298 13032 21406
rect 13176 21344 13228 21350
rect 13004 21270 13124 21298
rect 13176 21286 13228 21292
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12806 20768 12862 20777
rect 12806 20703 12862 20712
rect 12898 20632 12954 20641
rect 12898 20567 12954 20576
rect 12636 20444 12756 20472
rect 12440 20324 12492 20330
rect 12440 20266 12492 20272
rect 12532 20324 12584 20330
rect 12532 20266 12584 20272
rect 12348 19916 12400 19922
rect 12176 19876 12296 19904
rect 12072 19858 12124 19864
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11796 19780 11848 19786
rect 11796 19722 11848 19728
rect 11980 19712 12032 19718
rect 11980 19654 12032 19660
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11624 19196 11744 19224
rect 11624 19156 11652 19196
rect 11613 19128 11652 19156
rect 11613 18986 11641 19128
rect 11900 19122 11928 19314
rect 11992 19310 12020 19654
rect 12084 19378 12112 19858
rect 12072 19372 12124 19378
rect 12268 19334 12296 19876
rect 12348 19858 12400 19864
rect 12072 19314 12124 19320
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 12176 19306 12296 19334
rect 12360 19360 12388 19858
rect 12452 19553 12480 20266
rect 12532 19780 12584 19786
rect 12532 19722 12584 19728
rect 12544 19689 12572 19722
rect 12530 19680 12586 19689
rect 12530 19615 12586 19624
rect 12438 19544 12494 19553
rect 12438 19479 12494 19488
rect 12532 19372 12584 19378
rect 12360 19332 12480 19360
rect 12072 19236 12124 19242
rect 12072 19178 12124 19184
rect 11808 19094 11928 19122
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 11613 18958 11652 18986
rect 11520 18284 11572 18290
rect 11520 18226 11572 18232
rect 11520 18148 11572 18154
rect 11520 18090 11572 18096
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11440 17377 11468 17818
rect 11426 17368 11482 17377
rect 11426 17303 11482 17312
rect 11348 16546 11468 16574
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11164 15910 11192 15982
rect 11152 15904 11204 15910
rect 11150 15872 11152 15881
rect 11204 15872 11206 15881
rect 11150 15807 11206 15816
rect 11072 15524 11376 15552
rect 11242 15192 11298 15201
rect 10968 15156 11020 15162
rect 11242 15127 11298 15136
rect 10968 15098 11020 15104
rect 11256 15094 11284 15127
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 10692 14816 10744 14822
rect 10876 14816 10928 14822
rect 10692 14758 10744 14764
rect 10796 14776 10876 14804
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10600 14340 10652 14346
rect 10600 14282 10652 14288
rect 10612 14113 10640 14282
rect 10598 14104 10654 14113
rect 10598 14039 10654 14048
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10506 12744 10562 12753
rect 10612 12714 10640 13670
rect 10506 12679 10562 12688
rect 10600 12708 10652 12714
rect 10600 12650 10652 12656
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10520 11830 10548 12106
rect 10508 11824 10560 11830
rect 10508 11766 10560 11772
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10428 11665 10456 11698
rect 10414 11656 10470 11665
rect 10414 11591 10470 11600
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10428 11354 10456 11494
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10520 11150 10548 11494
rect 10612 11150 10640 12650
rect 10704 12050 10732 14758
rect 10796 12170 10824 14776
rect 10876 14758 10928 14764
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10888 14113 10916 14418
rect 10980 14346 11008 14962
rect 11060 14884 11112 14890
rect 11060 14826 11112 14832
rect 11072 14793 11100 14826
rect 11058 14784 11114 14793
rect 11058 14719 11114 14728
rect 11164 14634 11192 14962
rect 11072 14606 11192 14634
rect 11244 14612 11296 14618
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 10874 14104 10930 14113
rect 10874 14039 10930 14048
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10888 13841 10916 13874
rect 11072 13870 11100 14606
rect 11244 14554 11296 14560
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 11060 13864 11112 13870
rect 10874 13832 10930 13841
rect 11060 13806 11112 13812
rect 10874 13767 10930 13776
rect 11164 13716 11192 14486
rect 11256 14074 11284 14554
rect 11348 14550 11376 15524
rect 11336 14544 11388 14550
rect 11336 14486 11388 14492
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11348 14074 11376 14214
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11256 13841 11284 14010
rect 11242 13832 11298 13841
rect 11440 13802 11468 16546
rect 11532 16017 11560 18090
rect 11624 17882 11652 18958
rect 11808 18601 11836 19094
rect 11886 19000 11942 19009
rect 11886 18935 11888 18944
rect 11940 18935 11942 18944
rect 11888 18906 11940 18912
rect 11992 18816 12020 19110
rect 12084 18970 12112 19178
rect 12176 19009 12204 19306
rect 12162 19000 12218 19009
rect 12072 18964 12124 18970
rect 12162 18935 12218 18944
rect 12072 18906 12124 18912
rect 12072 18828 12124 18834
rect 11992 18788 12072 18816
rect 12072 18770 12124 18776
rect 12176 18714 12204 18935
rect 11992 18686 12204 18714
rect 12256 18760 12308 18766
rect 12452 18748 12480 19332
rect 12532 19314 12584 19320
rect 12544 19281 12572 19314
rect 12530 19272 12586 19281
rect 12530 19207 12586 19216
rect 12636 19174 12664 20444
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12728 19718 12756 20334
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12820 19514 12848 19994
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12806 19272 12862 19281
rect 12806 19207 12862 19216
rect 12624 19168 12676 19174
rect 12530 19136 12586 19145
rect 12624 19110 12676 19116
rect 12530 19071 12586 19080
rect 12544 18902 12572 19071
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 12636 18766 12664 18906
rect 12820 18766 12848 19207
rect 12308 18720 12480 18748
rect 12624 18760 12676 18766
rect 12256 18702 12308 18708
rect 12624 18702 12676 18708
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 11888 18624 11940 18630
rect 11794 18592 11850 18601
rect 11888 18566 11940 18572
rect 11794 18527 11850 18536
rect 11900 18426 11928 18566
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11612 17876 11664 17882
rect 11612 17818 11664 17824
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 11624 17105 11652 17682
rect 11716 17241 11744 18362
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11808 17678 11836 18226
rect 11796 17672 11848 17678
rect 11796 17614 11848 17620
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11702 17232 11758 17241
rect 11702 17167 11704 17176
rect 11756 17167 11758 17176
rect 11704 17138 11756 17144
rect 11610 17096 11666 17105
rect 11808 17082 11836 17274
rect 11610 17031 11666 17040
rect 11716 17054 11836 17082
rect 11716 16522 11744 17054
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11808 16561 11836 16730
rect 11794 16552 11850 16561
rect 11704 16516 11756 16522
rect 11794 16487 11850 16496
rect 11704 16458 11756 16464
rect 11610 16280 11666 16289
rect 11610 16215 11666 16224
rect 11624 16046 11652 16215
rect 11612 16040 11664 16046
rect 11518 16008 11574 16017
rect 11612 15982 11664 15988
rect 11518 15943 11574 15952
rect 11808 15910 11836 16487
rect 11900 16289 11928 18226
rect 11992 17814 12020 18686
rect 12624 18624 12676 18630
rect 12268 18550 12572 18578
rect 12912 18578 12940 20567
rect 12624 18566 12676 18572
rect 12162 18456 12218 18465
rect 12162 18391 12164 18400
rect 12216 18391 12218 18400
rect 12164 18362 12216 18368
rect 12176 18290 12204 18362
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12268 18222 12296 18550
rect 12346 18456 12402 18465
rect 12346 18391 12402 18400
rect 12440 18420 12492 18426
rect 12256 18216 12308 18222
rect 12162 18184 12218 18193
rect 12256 18158 12308 18164
rect 12360 18154 12388 18391
rect 12440 18362 12492 18368
rect 12162 18119 12218 18128
rect 12348 18148 12400 18154
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 11980 17808 12032 17814
rect 11980 17750 12032 17756
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 11992 16726 12020 17138
rect 11980 16720 12032 16726
rect 11980 16662 12032 16668
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11886 16280 11942 16289
rect 11886 16215 11942 16224
rect 11992 16164 12020 16526
rect 11900 16136 12020 16164
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11900 15722 11928 16136
rect 11978 16008 12034 16017
rect 11978 15943 12034 15952
rect 11808 15694 11928 15722
rect 11518 15328 11574 15337
rect 11518 15263 11574 15272
rect 11532 14346 11560 15263
rect 11808 15026 11836 15694
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11704 14612 11756 14618
rect 11900 14600 11928 14962
rect 11992 14634 12020 15943
rect 12084 14822 12112 17818
rect 12176 17270 12204 18119
rect 12348 18090 12400 18096
rect 12452 17882 12480 18362
rect 12544 18222 12572 18550
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 12348 17740 12400 17746
rect 12400 17700 12480 17728
rect 12348 17682 12400 17688
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12360 17270 12388 17478
rect 12164 17264 12216 17270
rect 12164 17206 12216 17212
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12164 17128 12216 17134
rect 12162 17096 12164 17105
rect 12452 17116 12480 17700
rect 12216 17096 12218 17105
rect 12162 17031 12218 17040
rect 12360 17088 12480 17116
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12176 16794 12204 16934
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 12164 16108 12216 16114
rect 12164 16050 12216 16056
rect 12176 15502 12204 16050
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12268 15337 12296 16934
rect 12360 15570 12388 17088
rect 12544 16561 12572 17750
rect 12636 17338 12664 18566
rect 12820 18550 12940 18578
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12728 18329 12756 18362
rect 12714 18320 12770 18329
rect 12714 18255 12770 18264
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12728 17678 12756 17818
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12820 17610 12848 18550
rect 12900 18420 12952 18426
rect 12900 18362 12952 18368
rect 12808 17604 12860 17610
rect 12808 17546 12860 17552
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12728 17218 12756 17274
rect 12636 17190 12756 17218
rect 12530 16552 12586 16561
rect 12530 16487 12586 16496
rect 12440 16448 12492 16454
rect 12438 16416 12440 16425
rect 12492 16416 12494 16425
rect 12438 16351 12494 16360
rect 12532 16176 12584 16182
rect 12532 16118 12584 16124
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 12254 15328 12310 15337
rect 12254 15263 12310 15272
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11992 14606 12112 14634
rect 11756 14572 11928 14600
rect 11704 14554 11756 14560
rect 11520 14340 11572 14346
rect 11520 14282 11572 14288
rect 11518 14104 11574 14113
rect 11518 14039 11520 14048
rect 11572 14039 11574 14048
rect 11520 14010 11572 14016
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11242 13767 11298 13776
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 11428 13796 11480 13802
rect 11428 13738 11480 13744
rect 10888 13688 11192 13716
rect 10888 13190 10916 13688
rect 11348 13682 11376 13738
rect 11348 13654 11468 13682
rect 11440 13530 11468 13654
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11256 13376 11284 13466
rect 11164 13348 11284 13376
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10888 12782 10916 13126
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10888 12170 10916 12582
rect 10784 12164 10836 12170
rect 10784 12106 10836 12112
rect 10876 12164 10928 12170
rect 10876 12106 10928 12112
rect 10874 12064 10930 12073
rect 10704 12022 10824 12050
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 10704 11218 10732 11562
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10506 10432 10562 10441
rect 10506 10367 10562 10376
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10230 9959 10286 9968
rect 10324 9988 10376 9994
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 9864 8774 9916 8780
rect 10046 8800 10102 8809
rect 9680 8560 9732 8566
rect 9586 8528 9642 8537
rect 9496 8492 9548 8498
rect 9680 8502 9732 8508
rect 9876 8498 9904 8774
rect 10046 8735 10102 8744
rect 9954 8528 10010 8537
rect 9586 8463 9642 8472
rect 9864 8492 9916 8498
rect 9496 8434 9548 8440
rect 9954 8463 10010 8472
rect 9864 8434 9916 8440
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9312 8016 9364 8022
rect 9312 7958 9364 7964
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9508 7585 9536 8434
rect 9968 8430 9996 8463
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9600 7886 9628 8366
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9956 7812 10008 7818
rect 9956 7754 10008 7760
rect 9494 7576 9550 7585
rect 9494 7511 9550 7520
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9508 7002 9536 7346
rect 9968 7342 9996 7754
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9876 7002 9904 7210
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9310 6896 9366 6905
rect 9310 6831 9366 6840
rect 9494 6896 9550 6905
rect 9494 6831 9550 6840
rect 9588 6860 9640 6866
rect 9324 6798 9352 6831
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9310 6080 9366 6089
rect 9310 6015 9366 6024
rect 9324 5778 9352 6015
rect 9416 5914 9444 6734
rect 9508 6662 9536 6831
rect 9588 6802 9640 6808
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 9600 5166 9628 6802
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 9600 4690 9628 5102
rect 10060 5098 10088 8735
rect 10152 6458 10180 9046
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10048 5092 10100 5098
rect 10048 5034 10100 5040
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9956 4616 10008 4622
rect 9954 4584 9956 4593
rect 10008 4584 10010 4593
rect 9954 4519 10010 4528
rect 10244 3738 10272 9959
rect 10324 9930 10376 9936
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10336 8498 10364 9522
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10428 7886 10456 10202
rect 10520 9704 10548 10367
rect 10612 10130 10640 11086
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10520 9676 10640 9704
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10520 9450 10548 9522
rect 10508 9444 10560 9450
rect 10508 9386 10560 9392
rect 10520 8362 10548 9386
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10428 7410 10456 7822
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10520 7206 10548 7414
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10612 6798 10640 9676
rect 10704 7206 10732 11154
rect 10796 8022 10824 12022
rect 10874 11999 10930 12008
rect 10888 11665 10916 11999
rect 10980 11898 11008 13194
rect 11164 12889 11192 13348
rect 11440 13308 11468 13466
rect 11256 13280 11468 13308
rect 11150 12880 11206 12889
rect 11150 12815 11206 12824
rect 11256 12782 11284 13280
rect 11426 12880 11482 12889
rect 11426 12815 11428 12824
rect 11480 12815 11482 12824
rect 11428 12786 11480 12792
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11152 12640 11204 12646
rect 11334 12608 11390 12617
rect 11204 12588 11334 12594
rect 11152 12582 11334 12588
rect 11164 12566 11334 12582
rect 11334 12543 11390 12552
rect 11440 12442 11468 12786
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11428 12232 11480 12238
rect 11426 12200 11428 12209
rect 11480 12200 11482 12209
rect 11426 12135 11482 12144
rect 11058 12064 11114 12073
rect 11058 11999 11114 12008
rect 11242 12064 11298 12073
rect 11242 11999 11298 12008
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 10874 11656 10930 11665
rect 10874 11591 10930 11600
rect 10888 11150 10916 11591
rect 10876 11144 10928 11150
rect 10874 11112 10876 11121
rect 10928 11112 10930 11121
rect 10874 11047 10930 11056
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10980 10130 11008 10610
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10888 9518 10916 9862
rect 10968 9716 11020 9722
rect 11072 9704 11100 11999
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 11164 11558 11192 11834
rect 11256 11558 11284 11999
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11440 11354 11468 11698
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11440 10470 11468 10610
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11242 10024 11298 10033
rect 11242 9959 11298 9968
rect 11256 9926 11284 9959
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11020 9676 11100 9704
rect 11242 9752 11298 9761
rect 11242 9687 11298 9696
rect 10968 9658 11020 9664
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10980 9042 11008 9522
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10980 8566 11008 8842
rect 11072 8809 11100 9676
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 11164 9217 11192 9386
rect 11150 9208 11206 9217
rect 11150 9143 11206 9152
rect 11152 8832 11204 8838
rect 11058 8800 11114 8809
rect 11152 8774 11204 8780
rect 11058 8735 11114 8744
rect 10968 8560 11020 8566
rect 11060 8560 11112 8566
rect 10968 8502 11020 8508
rect 11058 8528 11060 8537
rect 11112 8528 11114 8537
rect 11164 8498 11192 8774
rect 11058 8463 11114 8472
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10888 8294 10916 8366
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10784 8016 10836 8022
rect 10784 7958 10836 7964
rect 10888 7206 10916 8026
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10704 7002 10732 7142
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10612 6186 10640 6734
rect 10704 6322 10732 6938
rect 10980 6882 11008 7686
rect 11256 7002 11284 9687
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11348 8634 11376 8910
rect 11440 8906 11468 10406
rect 11428 8900 11480 8906
rect 11428 8842 11480 8848
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11426 8392 11482 8401
rect 11426 8327 11428 8336
rect 11480 8327 11482 8336
rect 11428 8298 11480 8304
rect 11532 8294 11560 13806
rect 11624 11778 11652 14554
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11716 14346 11744 14418
rect 11900 14414 11928 14572
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11704 14340 11756 14346
rect 11704 14282 11756 14288
rect 11702 14104 11758 14113
rect 11702 14039 11758 14048
rect 11716 13938 11744 14039
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11716 13326 11744 13738
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11702 13016 11758 13025
rect 11702 12951 11758 12960
rect 11808 12968 11836 14350
rect 11992 14090 12020 14486
rect 12084 14414 12112 14606
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 11900 14062 12020 14090
rect 11900 13326 11928 14062
rect 11980 14000 12032 14006
rect 11978 13968 11980 13977
rect 12032 13968 12034 13977
rect 12176 13954 12204 15098
rect 12256 14952 12308 14958
rect 12254 14920 12256 14929
rect 12308 14920 12310 14929
rect 12254 14855 12310 14864
rect 12254 14648 12310 14657
rect 12254 14583 12310 14592
rect 12268 14482 12296 14583
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 12268 14074 12296 14282
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 11978 13903 12034 13912
rect 12084 13926 12204 13954
rect 11978 13832 12034 13841
rect 11978 13767 12034 13776
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11716 12306 11744 12951
rect 11808 12940 11928 12968
rect 11900 12850 11928 12940
rect 11992 12850 12020 13767
rect 12084 13530 12112 13926
rect 12164 13864 12216 13870
rect 12162 13832 12164 13841
rect 12216 13832 12218 13841
rect 12162 13767 12218 13776
rect 12360 13716 12388 15506
rect 12452 15502 12480 15914
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 14618 12480 14894
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12544 14074 12572 16118
rect 12636 16046 12664 17190
rect 12820 16998 12848 17546
rect 12912 17105 12940 18362
rect 13004 17921 13032 21082
rect 13096 20618 13124 21270
rect 13188 20777 13216 21286
rect 13174 20768 13230 20777
rect 13174 20703 13230 20712
rect 13096 20590 13216 20618
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 13096 19242 13124 20198
rect 13084 19236 13136 19242
rect 13084 19178 13136 19184
rect 13082 18456 13138 18465
rect 13082 18391 13138 18400
rect 12990 17912 13046 17921
rect 13096 17882 13124 18391
rect 12990 17847 13046 17856
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 12992 17808 13044 17814
rect 12992 17750 13044 17756
rect 13004 17377 13032 17750
rect 12990 17368 13046 17377
rect 12990 17303 13046 17312
rect 12898 17096 12954 17105
rect 12898 17031 12954 17040
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12728 14793 12756 16934
rect 13004 16590 13032 17303
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 12820 16250 12848 16526
rect 12900 16448 12952 16454
rect 13096 16402 13124 17818
rect 13188 16794 13216 20590
rect 13280 19718 13308 21490
rect 13358 21176 13414 21185
rect 13358 21111 13414 21120
rect 13372 21078 13400 21111
rect 13360 21072 13412 21078
rect 13360 21014 13412 21020
rect 13360 20936 13412 20942
rect 13358 20904 13360 20913
rect 13412 20904 13414 20913
rect 13358 20839 13414 20848
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13372 19854 13400 20538
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13268 19712 13320 19718
rect 13268 19654 13320 19660
rect 13358 19680 13414 19689
rect 13358 19615 13414 19624
rect 13372 19514 13400 19615
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 13280 19310 13308 19450
rect 13268 19304 13320 19310
rect 13268 19246 13320 19252
rect 13280 18970 13308 19246
rect 13268 18964 13320 18970
rect 13268 18906 13320 18912
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 13280 17921 13308 18770
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13266 17912 13322 17921
rect 13266 17847 13322 17856
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13280 16833 13308 17614
rect 13372 17542 13400 18022
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 13266 16824 13322 16833
rect 13176 16788 13228 16794
rect 13266 16759 13322 16768
rect 13176 16730 13228 16736
rect 12900 16390 12952 16396
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12820 15706 12848 16050
rect 12912 15978 12940 16390
rect 13004 16374 13124 16402
rect 12900 15972 12952 15978
rect 12900 15914 12952 15920
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 13004 15620 13032 16374
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 12912 15592 13032 15620
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12820 15337 12848 15370
rect 12806 15328 12862 15337
rect 12806 15263 12862 15272
rect 12714 14784 12770 14793
rect 12714 14719 12770 14728
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12636 14346 12664 14486
rect 12624 14340 12676 14346
rect 12912 14328 12940 15592
rect 13096 15552 13124 16186
rect 13188 16046 13216 16730
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 12624 14282 12676 14288
rect 12728 14300 12940 14328
rect 13004 15524 13124 15552
rect 13266 15600 13322 15609
rect 13266 15535 13322 15544
rect 12622 14240 12678 14249
rect 12622 14175 12678 14184
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12438 13968 12494 13977
rect 12438 13903 12440 13912
rect 12492 13903 12494 13912
rect 12532 13932 12584 13938
rect 12440 13874 12492 13880
rect 12532 13874 12584 13880
rect 12544 13818 12572 13874
rect 12176 13688 12388 13716
rect 12452 13790 12572 13818
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11808 12753 11836 12786
rect 11794 12744 11850 12753
rect 12070 12744 12126 12753
rect 11794 12679 11850 12688
rect 11900 12702 12070 12730
rect 11808 12374 11836 12679
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11716 12209 11744 12242
rect 11702 12200 11758 12209
rect 11702 12135 11758 12144
rect 11900 12102 11928 12702
rect 12070 12679 12126 12688
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 12084 12306 12112 12582
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12176 12186 12204 13688
rect 12452 13530 12480 13790
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12084 12158 12204 12186
rect 12268 12186 12296 13262
rect 12544 12918 12572 13398
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12360 12345 12388 12786
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12346 12336 12402 12345
rect 12346 12271 12402 12280
rect 12268 12158 12388 12186
rect 11888 12096 11940 12102
rect 11794 12064 11850 12073
rect 11888 12038 11940 12044
rect 11794 11999 11850 12008
rect 11624 11750 11744 11778
rect 11808 11762 11836 11999
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11716 11642 11744 11750
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 12084 11694 12112 12158
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12072 11688 12124 11694
rect 11624 10742 11652 11630
rect 11716 11614 11836 11642
rect 12072 11630 12124 11636
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 11702 10704 11758 10713
rect 11702 10639 11704 10648
rect 11756 10639 11758 10648
rect 11704 10610 11756 10616
rect 11716 10470 11744 10610
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11702 9208 11758 9217
rect 11808 9178 11836 11614
rect 12176 11558 12204 12038
rect 12360 11762 12388 12158
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12268 11626 12296 11698
rect 12256 11620 12308 11626
rect 12256 11562 12308 11568
rect 11888 11552 11940 11558
rect 12164 11552 12216 11558
rect 11888 11494 11940 11500
rect 12070 11520 12126 11529
rect 11900 11354 11928 11494
rect 12164 11494 12216 11500
rect 12070 11455 12126 11464
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 12084 11014 12112 11455
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 11992 10674 12020 10950
rect 12176 10826 12204 11018
rect 12084 10798 12204 10826
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 12084 10305 12112 10798
rect 12256 10736 12308 10742
rect 12256 10678 12308 10684
rect 12268 10470 12296 10678
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12070 10296 12126 10305
rect 12070 10231 12126 10240
rect 11978 9480 12034 9489
rect 11978 9415 12034 9424
rect 11702 9143 11758 9152
rect 11796 9172 11848 9178
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11532 8090 11560 8230
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11624 7954 11652 8978
rect 11716 8673 11744 9143
rect 11796 9114 11848 9120
rect 11702 8664 11758 8673
rect 11702 8599 11704 8608
rect 11756 8599 11758 8608
rect 11704 8570 11756 8576
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11716 8090 11744 8434
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11808 7886 11836 9114
rect 11992 8673 12020 9415
rect 11978 8664 12034 8673
rect 11888 8628 11940 8634
rect 11978 8599 12034 8608
rect 11888 8570 11940 8576
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11518 7168 11574 7177
rect 11518 7103 11574 7112
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 10980 6854 11284 6882
rect 11256 6798 11284 6854
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 10796 6633 10824 6734
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10876 6656 10928 6662
rect 10782 6624 10838 6633
rect 10876 6598 10928 6604
rect 10782 6559 10838 6568
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10600 6180 10652 6186
rect 10600 6122 10652 6128
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 10888 2689 10916 6598
rect 10980 5302 11008 6666
rect 11150 6624 11206 6633
rect 11150 6559 11206 6568
rect 11058 6216 11114 6225
rect 11058 6151 11114 6160
rect 11072 5846 11100 6151
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11164 5681 11192 6559
rect 11256 6186 11284 6734
rect 11440 6254 11468 6938
rect 11532 6934 11560 7103
rect 11520 6928 11572 6934
rect 11900 6882 11928 8570
rect 11978 8120 12034 8129
rect 12084 8106 12112 10231
rect 12176 9110 12204 10406
rect 12254 9480 12310 9489
rect 12254 9415 12310 9424
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12176 8294 12204 9046
rect 12268 9042 12296 9415
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12360 8906 12388 11698
rect 12452 10062 12480 12718
rect 12544 12646 12572 12718
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12544 11676 12572 12310
rect 12636 11830 12664 14175
rect 12624 11824 12676 11830
rect 12624 11766 12676 11772
rect 12544 11648 12664 11676
rect 12530 10432 12586 10441
rect 12530 10367 12586 10376
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12544 9722 12572 10367
rect 12636 9761 12664 11648
rect 12728 10810 12756 14300
rect 12806 13968 12862 13977
rect 12806 13903 12808 13912
rect 12860 13903 12862 13912
rect 12808 13874 12860 13880
rect 12808 13796 12860 13802
rect 13004 13784 13032 15524
rect 13084 15428 13136 15434
rect 13084 15370 13136 15376
rect 13096 14618 13124 15370
rect 13280 14958 13308 15535
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 13096 14414 13124 14554
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 12808 13738 12860 13744
rect 12912 13756 13032 13784
rect 12820 13394 12848 13738
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 12820 11898 12848 12242
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12912 11558 12940 13756
rect 13096 13394 13124 14350
rect 13188 14074 13216 14826
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13280 14414 13308 14758
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13266 13968 13322 13977
rect 13176 13932 13228 13938
rect 13266 13903 13322 13912
rect 13176 13874 13228 13880
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 13004 13297 13032 13330
rect 12990 13288 13046 13297
rect 12990 13223 13046 13232
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 13096 13025 13124 13194
rect 13082 13016 13138 13025
rect 13082 12951 13138 12960
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 13082 12744 13138 12753
rect 13004 11694 13032 12718
rect 13082 12679 13138 12688
rect 13096 12374 13124 12679
rect 13084 12368 13136 12374
rect 13084 12310 13136 12316
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 13096 11762 13124 12174
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 12900 11552 12952 11558
rect 12952 11512 13032 11540
rect 12900 11494 12952 11500
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12728 10305 12756 10542
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12714 10296 12770 10305
rect 12714 10231 12770 10240
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12622 9752 12678 9761
rect 12532 9716 12584 9722
rect 12622 9687 12678 9696
rect 12532 9658 12584 9664
rect 12440 9444 12492 9450
rect 12440 9386 12492 9392
rect 12452 9110 12480 9386
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 12452 8820 12480 9046
rect 12544 8974 12572 9658
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12452 8792 12572 8820
rect 12254 8528 12310 8537
rect 12254 8463 12256 8472
rect 12308 8463 12310 8472
rect 12438 8528 12494 8537
rect 12544 8498 12572 8792
rect 12438 8463 12494 8472
rect 12532 8492 12584 8498
rect 12256 8434 12308 8440
rect 12452 8378 12480 8463
rect 12532 8434 12584 8440
rect 12348 8356 12400 8362
rect 12452 8350 12572 8378
rect 12636 8362 12664 9687
rect 12348 8298 12400 8304
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12084 8078 12204 8106
rect 11978 8055 12034 8064
rect 11992 7970 12020 8055
rect 11992 7942 12112 7970
rect 11520 6870 11572 6876
rect 11532 6798 11560 6870
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11808 6854 11928 6882
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11532 6322 11560 6598
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11244 6180 11296 6186
rect 11244 6122 11296 6128
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11242 5944 11298 5953
rect 11242 5879 11298 5888
rect 11256 5710 11284 5879
rect 11348 5817 11376 6054
rect 11334 5808 11390 5817
rect 11334 5743 11390 5752
rect 11244 5704 11296 5710
rect 11150 5672 11206 5681
rect 11244 5646 11296 5652
rect 11150 5607 11206 5616
rect 10968 5296 11020 5302
rect 10968 5238 11020 5244
rect 10980 4622 11008 5238
rect 11348 5166 11376 5743
rect 11440 5642 11468 6190
rect 11532 5846 11560 6258
rect 11716 6118 11744 6802
rect 11808 6633 11836 6854
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11794 6624 11850 6633
rect 11794 6559 11850 6568
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11520 5840 11572 5846
rect 11520 5782 11572 5788
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11624 5642 11652 5714
rect 11428 5636 11480 5642
rect 11428 5578 11480 5584
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11900 5574 11928 6666
rect 12084 6338 12112 7942
rect 11992 6310 12112 6338
rect 11992 6118 12020 6310
rect 11980 6112 12032 6118
rect 11978 6080 11980 6089
rect 12032 6080 12034 6089
rect 11978 6015 12034 6024
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11900 5234 11928 5510
rect 12084 5370 12112 5646
rect 12176 5545 12204 8078
rect 12268 8022 12296 8230
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 12360 6662 12388 8298
rect 12544 7410 12572 8350
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12636 7886 12664 8026
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12622 7440 12678 7449
rect 12532 7404 12584 7410
rect 12622 7375 12678 7384
rect 12532 7346 12584 7352
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12544 5778 12572 7346
rect 12636 7342 12664 7375
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12624 7200 12676 7206
rect 12622 7168 12624 7177
rect 12676 7168 12678 7177
rect 12622 7103 12678 7112
rect 12728 6905 12756 9998
rect 12820 9586 12848 10474
rect 12912 10266 12940 11290
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 13004 10198 13032 11512
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 13096 10470 13124 10610
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12912 9654 12940 9998
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12820 8265 12848 9522
rect 12912 8974 12940 9590
rect 13004 9382 13032 9590
rect 13096 9586 13124 10406
rect 13188 9674 13216 13874
rect 13280 13326 13308 13903
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13372 12434 13400 17478
rect 13464 16590 13492 22714
rect 13556 21457 13584 26726
rect 13648 26586 13676 26998
rect 13740 26994 13768 27066
rect 13832 27033 13860 28966
rect 13912 28688 13964 28694
rect 13912 28630 13964 28636
rect 13924 27878 13952 28630
rect 13912 27872 13964 27878
rect 13912 27814 13964 27820
rect 13924 27713 13952 27814
rect 13910 27704 13966 27713
rect 13910 27639 13966 27648
rect 13818 27024 13874 27033
rect 13728 26988 13780 26994
rect 14016 27010 14044 29135
rect 14280 28552 14332 28558
rect 14280 28494 14332 28500
rect 14556 28552 14608 28558
rect 14556 28494 14608 28500
rect 14096 28416 14148 28422
rect 14096 28358 14148 28364
rect 14108 28082 14136 28358
rect 14292 28150 14320 28494
rect 14464 28416 14516 28422
rect 14568 28393 14596 28494
rect 14464 28358 14516 28364
rect 14554 28384 14610 28393
rect 14280 28144 14332 28150
rect 14280 28086 14332 28092
rect 14096 28076 14148 28082
rect 14096 28018 14148 28024
rect 14476 27962 14504 28358
rect 14554 28319 14610 28328
rect 14556 28212 14608 28218
rect 14556 28154 14608 28160
rect 13818 26959 13874 26968
rect 13924 26994 14044 27010
rect 14292 27934 14504 27962
rect 13924 26988 14056 26994
rect 13924 26982 14004 26988
rect 13728 26930 13780 26936
rect 13636 26580 13688 26586
rect 13636 26522 13688 26528
rect 13740 26466 13768 26930
rect 13924 26858 13952 26982
rect 14004 26930 14056 26936
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 13912 26852 13964 26858
rect 13912 26794 13964 26800
rect 14004 26852 14056 26858
rect 14004 26794 14056 26800
rect 13820 26784 13872 26790
rect 13820 26726 13872 26732
rect 13648 26438 13768 26466
rect 13648 22030 13676 26438
rect 13728 26376 13780 26382
rect 13728 26318 13780 26324
rect 13740 26042 13768 26318
rect 13728 26036 13780 26042
rect 13728 25978 13780 25984
rect 13728 25492 13780 25498
rect 13728 25434 13780 25440
rect 13740 25401 13768 25434
rect 13726 25392 13782 25401
rect 13726 25327 13728 25336
rect 13780 25327 13782 25336
rect 13728 25298 13780 25304
rect 13832 24818 13860 26726
rect 13912 25696 13964 25702
rect 13912 25638 13964 25644
rect 13924 24886 13952 25638
rect 13912 24880 13964 24886
rect 13912 24822 13964 24828
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13924 24750 13952 24822
rect 13912 24744 13964 24750
rect 13912 24686 13964 24692
rect 14016 24426 14044 26794
rect 14200 26518 14228 26930
rect 14292 26761 14320 27934
rect 14372 27872 14424 27878
rect 14372 27814 14424 27820
rect 14464 27872 14516 27878
rect 14464 27814 14516 27820
rect 14384 27033 14412 27814
rect 14476 27062 14504 27814
rect 14568 27674 14596 28154
rect 14844 28082 14872 30602
rect 15014 30560 15070 30569
rect 15014 30495 15070 30504
rect 15028 28422 15056 30495
rect 15934 30152 15990 30161
rect 15934 30087 15990 30096
rect 15948 29306 15976 30087
rect 17144 29850 17172 31282
rect 18512 30728 18564 30734
rect 18512 30670 18564 30676
rect 17316 30252 17368 30258
rect 17316 30194 17368 30200
rect 17132 29844 17184 29850
rect 17132 29786 17184 29792
rect 17328 29714 17356 30194
rect 17316 29708 17368 29714
rect 17316 29650 17368 29656
rect 16580 29640 16632 29646
rect 16580 29582 16632 29588
rect 17500 29640 17552 29646
rect 17500 29582 17552 29588
rect 15936 29300 15988 29306
rect 15936 29242 15988 29248
rect 16396 29300 16448 29306
rect 16396 29242 16448 29248
rect 16304 29164 16356 29170
rect 16304 29106 16356 29112
rect 15844 28960 15896 28966
rect 15844 28902 15896 28908
rect 15292 28552 15344 28558
rect 15292 28494 15344 28500
rect 15016 28416 15068 28422
rect 15016 28358 15068 28364
rect 15028 28082 15056 28358
rect 14832 28076 14884 28082
rect 14832 28018 14884 28024
rect 15016 28076 15068 28082
rect 15016 28018 15068 28024
rect 15108 28076 15160 28082
rect 15108 28018 15160 28024
rect 14648 27872 14700 27878
rect 14646 27840 14648 27849
rect 14700 27840 14702 27849
rect 14646 27775 14702 27784
rect 14556 27668 14608 27674
rect 14556 27610 14608 27616
rect 14844 27418 14872 28018
rect 15014 27976 15070 27985
rect 15014 27911 15070 27920
rect 15028 27674 15056 27911
rect 15016 27668 15068 27674
rect 15016 27610 15068 27616
rect 14924 27532 14976 27538
rect 14976 27492 15056 27520
rect 14924 27474 14976 27480
rect 14568 27390 14872 27418
rect 14924 27396 14976 27402
rect 14568 27334 14596 27390
rect 14924 27338 14976 27344
rect 14556 27328 14608 27334
rect 14556 27270 14608 27276
rect 14648 27328 14700 27334
rect 14648 27270 14700 27276
rect 14464 27056 14516 27062
rect 14370 27024 14426 27033
rect 14464 26998 14516 27004
rect 14370 26959 14426 26968
rect 14278 26752 14334 26761
rect 14278 26687 14334 26696
rect 14188 26512 14240 26518
rect 14188 26454 14240 26460
rect 14280 25900 14332 25906
rect 14280 25842 14332 25848
rect 14188 25152 14240 25158
rect 14186 25120 14188 25129
rect 14240 25120 14242 25129
rect 14186 25055 14242 25064
rect 14188 24880 14240 24886
rect 14188 24822 14240 24828
rect 13924 24398 14044 24426
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13740 23730 13768 24006
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 13728 23520 13780 23526
rect 13728 23462 13780 23468
rect 13740 22234 13768 23462
rect 13820 23316 13872 23322
rect 13820 23258 13872 23264
rect 13832 22778 13860 23258
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 13728 22228 13780 22234
rect 13728 22170 13780 22176
rect 13636 22024 13688 22030
rect 13636 21966 13688 21972
rect 13818 21992 13874 22001
rect 13818 21927 13874 21936
rect 13832 21894 13860 21927
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13634 21720 13690 21729
rect 13634 21655 13690 21664
rect 13818 21720 13874 21729
rect 13818 21655 13820 21664
rect 13542 21448 13598 21457
rect 13542 21383 13598 21392
rect 13648 21350 13676 21655
rect 13872 21655 13874 21664
rect 13820 21626 13872 21632
rect 13728 21480 13780 21486
rect 13728 21422 13780 21428
rect 13636 21344 13688 21350
rect 13636 21286 13688 21292
rect 13542 20904 13598 20913
rect 13542 20839 13598 20848
rect 13636 20868 13688 20874
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13556 15552 13584 20839
rect 13636 20810 13688 20816
rect 13648 20777 13676 20810
rect 13634 20768 13690 20777
rect 13634 20703 13690 20712
rect 13636 20324 13688 20330
rect 13740 20312 13768 21422
rect 13924 21146 13952 24398
rect 14200 24290 14228 24822
rect 14292 24449 14320 25842
rect 14384 25294 14412 26959
rect 14462 26752 14518 26761
rect 14462 26687 14518 26696
rect 14476 26518 14504 26687
rect 14464 26512 14516 26518
rect 14464 26454 14516 26460
rect 14660 26081 14688 27270
rect 14936 27130 14964 27338
rect 15028 27130 15056 27492
rect 15120 27169 15148 28018
rect 15304 28014 15332 28494
rect 15856 28490 15884 28902
rect 16028 28756 16080 28762
rect 16028 28698 16080 28704
rect 16040 28490 16068 28698
rect 15844 28484 15896 28490
rect 15844 28426 15896 28432
rect 16028 28484 16080 28490
rect 16028 28426 16080 28432
rect 15292 28008 15344 28014
rect 15292 27950 15344 27956
rect 15198 27704 15254 27713
rect 15198 27639 15200 27648
rect 15252 27639 15254 27648
rect 15200 27610 15252 27616
rect 15200 27464 15252 27470
rect 15384 27464 15436 27470
rect 15200 27406 15252 27412
rect 15290 27432 15346 27441
rect 15106 27160 15162 27169
rect 14924 27124 14976 27130
rect 14924 27066 14976 27072
rect 15016 27124 15068 27130
rect 15106 27095 15162 27104
rect 15016 27066 15068 27072
rect 14832 27056 14884 27062
rect 14832 26998 14884 27004
rect 14740 26852 14792 26858
rect 14740 26794 14792 26800
rect 14646 26072 14702 26081
rect 14646 26007 14702 26016
rect 14462 25528 14518 25537
rect 14462 25463 14518 25472
rect 14372 25288 14424 25294
rect 14372 25230 14424 25236
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 14384 24614 14412 25094
rect 14372 24608 14424 24614
rect 14372 24550 14424 24556
rect 14278 24440 14334 24449
rect 14278 24375 14334 24384
rect 14476 24342 14504 25463
rect 14556 25288 14608 25294
rect 14556 25230 14608 25236
rect 14568 24857 14596 25230
rect 14554 24848 14610 24857
rect 14554 24783 14610 24792
rect 14648 24812 14700 24818
rect 14648 24754 14700 24760
rect 14660 24614 14688 24754
rect 14556 24608 14608 24614
rect 14556 24550 14608 24556
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14464 24336 14516 24342
rect 14200 24262 14412 24290
rect 14464 24278 14516 24284
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14188 24200 14240 24206
rect 14188 24142 14240 24148
rect 14002 24032 14058 24041
rect 14002 23967 14058 23976
rect 14016 23254 14044 23967
rect 14004 23248 14056 23254
rect 14004 23190 14056 23196
rect 14004 23044 14056 23050
rect 14004 22986 14056 22992
rect 13912 21140 13964 21146
rect 13912 21082 13964 21088
rect 13912 20936 13964 20942
rect 14016 20913 14044 22986
rect 13912 20878 13964 20884
rect 14002 20904 14058 20913
rect 13820 20868 13872 20874
rect 13820 20810 13872 20816
rect 13688 20284 13768 20312
rect 13636 20266 13688 20272
rect 13636 20052 13688 20058
rect 13832 20040 13860 20810
rect 13924 20244 13952 20878
rect 14002 20839 14058 20848
rect 14016 20398 14044 20839
rect 14108 20472 14136 24142
rect 14200 23730 14228 24142
rect 14280 24132 14332 24138
rect 14280 24074 14332 24080
rect 14292 23730 14320 24074
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 14280 23724 14332 23730
rect 14280 23666 14332 23672
rect 14200 23526 14228 23666
rect 14188 23520 14240 23526
rect 14188 23462 14240 23468
rect 14384 23338 14412 24262
rect 14464 23588 14516 23594
rect 14464 23530 14516 23536
rect 14200 23310 14412 23338
rect 14200 20806 14228 23310
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 14292 22506 14320 22646
rect 14384 22574 14412 23054
rect 14372 22568 14424 22574
rect 14372 22510 14424 22516
rect 14280 22500 14332 22506
rect 14280 22442 14332 22448
rect 14372 22432 14424 22438
rect 14372 22374 14424 22380
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 14292 21729 14320 21966
rect 14278 21720 14334 21729
rect 14278 21655 14334 21664
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14188 20800 14240 20806
rect 14188 20742 14240 20748
rect 14108 20444 14228 20472
rect 14004 20392 14056 20398
rect 14004 20334 14056 20340
rect 14094 20360 14150 20369
rect 14094 20295 14150 20304
rect 14004 20256 14056 20262
rect 13924 20216 14004 20244
rect 14004 20198 14056 20204
rect 13688 20012 13860 20040
rect 14004 20052 14056 20058
rect 13636 19994 13688 20000
rect 14108 20040 14136 20295
rect 14056 20012 14136 20040
rect 14004 19994 14056 20000
rect 14200 19854 14228 20444
rect 14292 20233 14320 21286
rect 14278 20224 14334 20233
rect 14278 20159 14334 20168
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13740 18714 13768 19654
rect 13832 19514 13860 19790
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13910 19408 13966 19417
rect 13910 19343 13966 19352
rect 13924 19310 13952 19343
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13464 15524 13584 15552
rect 13648 18686 13768 18714
rect 13464 14890 13492 15524
rect 13544 15428 13596 15434
rect 13544 15370 13596 15376
rect 13556 15094 13584 15370
rect 13544 15088 13596 15094
rect 13648 15065 13676 18686
rect 13728 18624 13780 18630
rect 13726 18592 13728 18601
rect 13780 18592 13782 18601
rect 13726 18527 13782 18536
rect 13832 18442 13860 19110
rect 13740 18414 13860 18442
rect 13544 15030 13596 15036
rect 13634 15056 13690 15065
rect 13740 15026 13768 18414
rect 14016 18068 14044 19654
rect 14108 18970 14136 19654
rect 14200 19378 14228 19654
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14188 19236 14240 19242
rect 14384 19224 14412 22374
rect 14476 20942 14504 23530
rect 14568 23497 14596 24550
rect 14554 23488 14610 23497
rect 14554 23423 14610 23432
rect 14556 23044 14608 23050
rect 14556 22986 14608 22992
rect 14568 22574 14596 22986
rect 14556 22568 14608 22574
rect 14556 22510 14608 22516
rect 14568 21162 14596 22510
rect 14660 21468 14688 24550
rect 14752 21593 14780 26794
rect 14844 26586 14872 26998
rect 15014 26616 15070 26625
rect 14832 26580 14884 26586
rect 15212 26586 15240 27406
rect 15384 27406 15436 27412
rect 15290 27367 15346 27376
rect 15014 26551 15016 26560
rect 14832 26522 14884 26528
rect 15068 26551 15070 26560
rect 15200 26580 15252 26586
rect 15016 26522 15068 26528
rect 15200 26522 15252 26528
rect 14844 26450 14964 26466
rect 14832 26444 14964 26450
rect 14884 26438 14964 26444
rect 14832 26386 14884 26392
rect 14832 26308 14884 26314
rect 14832 26250 14884 26256
rect 14844 26217 14872 26250
rect 14830 26208 14886 26217
rect 14830 26143 14886 26152
rect 14844 25265 14872 26143
rect 14936 25401 14964 26438
rect 15304 26382 15332 27367
rect 15016 26376 15068 26382
rect 15016 26318 15068 26324
rect 15292 26376 15344 26382
rect 15292 26318 15344 26324
rect 14922 25392 14978 25401
rect 14922 25327 14978 25336
rect 14830 25256 14886 25265
rect 14830 25191 14886 25200
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14844 23866 14872 24754
rect 14924 24744 14976 24750
rect 14924 24686 14976 24692
rect 14832 23860 14884 23866
rect 14832 23802 14884 23808
rect 14738 21584 14794 21593
rect 14738 21519 14794 21528
rect 14660 21440 14872 21468
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14646 21176 14702 21185
rect 14568 21134 14646 21162
rect 14752 21146 14780 21286
rect 14646 21111 14702 21120
rect 14740 21140 14792 21146
rect 14556 21004 14608 21010
rect 14556 20946 14608 20952
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14464 20800 14516 20806
rect 14568 20788 14596 20946
rect 14660 20942 14688 21111
rect 14740 21082 14792 21088
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14568 20760 14688 20788
rect 14464 20742 14516 20748
rect 14476 20534 14504 20742
rect 14464 20528 14516 20534
rect 14464 20470 14516 20476
rect 14660 20466 14688 20760
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14752 20398 14780 21082
rect 14464 20392 14516 20398
rect 14462 20360 14464 20369
rect 14740 20392 14792 20398
rect 14516 20360 14518 20369
rect 14740 20334 14792 20340
rect 14462 20295 14518 20304
rect 14844 20244 14872 21440
rect 14936 21418 14964 24686
rect 15028 23118 15056 26318
rect 15292 25424 15344 25430
rect 15292 25366 15344 25372
rect 15200 25288 15252 25294
rect 15198 25256 15200 25265
rect 15252 25256 15254 25265
rect 15198 25191 15254 25200
rect 15108 24812 15160 24818
rect 15108 24754 15160 24760
rect 15120 24342 15148 24754
rect 15108 24336 15160 24342
rect 15108 24278 15160 24284
rect 15120 24041 15148 24278
rect 15106 24032 15162 24041
rect 15106 23967 15162 23976
rect 15108 23724 15160 23730
rect 15108 23666 15160 23672
rect 15120 23594 15148 23666
rect 15304 23633 15332 25366
rect 15396 24993 15424 27406
rect 15568 26920 15620 26926
rect 15568 26862 15620 26868
rect 15382 24984 15438 24993
rect 15382 24919 15438 24928
rect 15474 24848 15530 24857
rect 15474 24783 15530 24792
rect 15290 23624 15346 23633
rect 15108 23588 15160 23594
rect 15290 23559 15346 23568
rect 15108 23530 15160 23536
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 15016 21956 15068 21962
rect 15016 21898 15068 21904
rect 14924 21412 14976 21418
rect 14924 21354 14976 21360
rect 15028 21049 15056 21898
rect 15014 21040 15070 21049
rect 15014 20975 15070 20984
rect 15120 20754 15148 23530
rect 15292 23520 15344 23526
rect 15292 23462 15344 23468
rect 15200 23044 15252 23050
rect 15200 22986 15252 22992
rect 15212 21486 15240 22986
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 15198 21040 15254 21049
rect 15198 20975 15254 20984
rect 15028 20726 15148 20754
rect 15028 20641 15056 20726
rect 15014 20632 15070 20641
rect 15212 20618 15240 20975
rect 15120 20602 15240 20618
rect 15014 20567 15070 20576
rect 15108 20596 15240 20602
rect 15160 20590 15240 20596
rect 15108 20538 15160 20544
rect 15200 20528 15252 20534
rect 15200 20470 15252 20476
rect 14924 20392 14976 20398
rect 14924 20334 14976 20340
rect 14752 20216 14872 20244
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14660 19961 14688 19994
rect 14646 19952 14702 19961
rect 14464 19916 14516 19922
rect 14646 19887 14702 19896
rect 14464 19858 14516 19864
rect 14240 19196 14412 19224
rect 14188 19178 14240 19184
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14200 18766 14228 19178
rect 14476 19174 14504 19858
rect 14554 19816 14610 19825
rect 14554 19751 14610 19760
rect 14568 19718 14596 19751
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14660 19446 14688 19654
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14464 18964 14516 18970
rect 14516 18924 14596 18952
rect 14464 18906 14516 18912
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14292 18426 14320 18770
rect 14370 18592 14426 18601
rect 14370 18527 14426 18536
rect 14280 18420 14332 18426
rect 14280 18362 14332 18368
rect 14016 18040 14228 18068
rect 14094 17912 14150 17921
rect 14094 17847 14150 17856
rect 13912 17604 13964 17610
rect 13912 17546 13964 17552
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13634 14991 13690 15000
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13452 14884 13504 14890
rect 13452 14826 13504 14832
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13464 13870 13492 14010
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13556 13394 13584 14758
rect 13648 14074 13676 14826
rect 13740 14249 13768 14962
rect 13832 14657 13860 17138
rect 13924 17066 13952 17546
rect 13912 17060 13964 17066
rect 13912 17002 13964 17008
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 14016 16794 14044 16934
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 14004 15972 14056 15978
rect 14004 15914 14056 15920
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13924 15570 13952 15846
rect 14016 15745 14044 15914
rect 14002 15736 14058 15745
rect 14002 15671 14058 15680
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 13910 15464 13966 15473
rect 13910 15399 13966 15408
rect 13818 14648 13874 14657
rect 13818 14583 13874 14592
rect 13726 14240 13782 14249
rect 13726 14175 13782 14184
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 13648 13530 13676 14010
rect 13728 13932 13780 13938
rect 13832 13920 13860 14583
rect 13780 13892 13860 13920
rect 13728 13874 13780 13880
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13924 13274 13952 15399
rect 13556 13246 13952 13274
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13280 12406 13400 12434
rect 13280 10062 13308 12406
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13372 11558 13400 11698
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13188 9646 13308 9674
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12912 8673 12940 8774
rect 12898 8664 12954 8673
rect 12898 8599 12954 8608
rect 13004 8498 13032 9318
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12806 8256 12862 8265
rect 12806 8191 12862 8200
rect 12714 6896 12770 6905
rect 12714 6831 12770 6840
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12162 5536 12218 5545
rect 12162 5471 12218 5480
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 12624 4752 12676 4758
rect 12622 4720 12624 4729
rect 12676 4720 12678 4729
rect 12622 4655 12678 4664
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12820 4282 12848 4558
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 12912 3777 12940 8434
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13004 7546 13032 7822
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 13096 7410 13124 9522
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13188 8945 13216 9454
rect 13174 8936 13230 8945
rect 13174 8871 13230 8880
rect 13188 8838 13216 8871
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13188 7562 13216 8434
rect 13280 8430 13308 9646
rect 13372 9586 13400 11494
rect 13464 11336 13492 13126
rect 13556 12434 13584 13246
rect 13912 13184 13964 13190
rect 13818 13152 13874 13161
rect 13912 13126 13964 13132
rect 13818 13087 13874 13096
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13556 12406 13676 12434
rect 13544 11348 13596 11354
rect 13464 11308 13544 11336
rect 13544 11290 13596 11296
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13280 7834 13308 8366
rect 13372 7954 13400 8910
rect 13556 8498 13584 11290
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13648 8090 13676 12406
rect 13740 11898 13768 12582
rect 13832 12238 13860 13087
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13818 11928 13874 11937
rect 13728 11892 13780 11898
rect 13818 11863 13874 11872
rect 13728 11834 13780 11840
rect 13832 11529 13860 11863
rect 13818 11520 13874 11529
rect 13818 11455 13874 11464
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13740 9178 13768 9454
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13740 8430 13768 8570
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13280 7806 13492 7834
rect 13358 7576 13414 7585
rect 13188 7546 13308 7562
rect 13188 7540 13320 7546
rect 13188 7534 13268 7540
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 13004 6798 13032 7142
rect 13096 7002 13124 7346
rect 13188 7274 13216 7534
rect 13358 7511 13414 7520
rect 13268 7482 13320 7488
rect 13372 7478 13400 7511
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 13176 7268 13228 7274
rect 13176 7210 13228 7216
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 13372 6866 13400 7414
rect 13464 7342 13492 7806
rect 13648 7585 13676 7890
rect 13634 7576 13690 7585
rect 13634 7511 13690 7520
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13452 6928 13504 6934
rect 13452 6870 13504 6876
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 13268 5840 13320 5846
rect 13268 5782 13320 5788
rect 13280 5574 13308 5782
rect 13464 5642 13492 6870
rect 13452 5636 13504 5642
rect 13452 5578 13504 5584
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 12898 3768 12954 3777
rect 12898 3703 12954 3712
rect 13556 3369 13584 7346
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13648 6769 13676 6938
rect 13634 6760 13690 6769
rect 13634 6695 13690 6704
rect 13740 5409 13768 8366
rect 13832 7750 13860 9930
rect 13924 9330 13952 13126
rect 14016 10742 14044 15506
rect 14108 15094 14136 17847
rect 14200 17610 14228 18040
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14188 17604 14240 17610
rect 14188 17546 14240 17552
rect 14292 17105 14320 17614
rect 14278 17096 14334 17105
rect 14278 17031 14334 17040
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14200 15366 14228 16934
rect 14278 16688 14334 16697
rect 14278 16623 14334 16632
rect 14292 16182 14320 16623
rect 14384 16590 14412 18527
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14476 17746 14504 18022
rect 14464 17740 14516 17746
rect 14464 17682 14516 17688
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14280 16176 14332 16182
rect 14280 16118 14332 16124
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14096 15088 14148 15094
rect 14372 15088 14424 15094
rect 14096 15030 14148 15036
rect 14186 15056 14242 15065
rect 14372 15030 14424 15036
rect 14186 14991 14242 15000
rect 14280 15020 14332 15026
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14108 13258 14136 14350
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 14108 12986 14136 13194
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 14108 11218 14136 11766
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 14004 10736 14056 10742
rect 14004 10678 14056 10684
rect 14096 9376 14148 9382
rect 13924 9302 14044 9330
rect 14096 9318 14148 9324
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13832 7410 13860 7686
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13924 7274 13952 8434
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13924 6322 13952 6734
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 14016 6118 14044 9302
rect 14108 8974 14136 9318
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 14094 8664 14150 8673
rect 14094 8599 14150 8608
rect 14108 8498 14136 8599
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14096 7812 14148 7818
rect 14096 7754 14148 7760
rect 14108 7177 14136 7754
rect 14094 7168 14150 7177
rect 14094 7103 14150 7112
rect 14200 6458 14228 14991
rect 14280 14962 14332 14968
rect 14292 14793 14320 14962
rect 14278 14784 14334 14793
rect 14278 14719 14334 14728
rect 14278 14648 14334 14657
rect 14278 14583 14334 14592
rect 14292 13802 14320 14583
rect 14280 13796 14332 13802
rect 14280 13738 14332 13744
rect 14384 13190 14412 15030
rect 14372 13184 14424 13190
rect 14278 13152 14334 13161
rect 14372 13126 14424 13132
rect 14278 13087 14334 13096
rect 14292 11642 14320 13087
rect 14370 13016 14426 13025
rect 14370 12951 14426 12960
rect 14384 12481 14412 12951
rect 14370 12472 14426 12481
rect 14370 12407 14426 12416
rect 14476 12434 14504 17138
rect 14568 13938 14596 18924
rect 14648 18692 14700 18698
rect 14648 18634 14700 18640
rect 14660 18601 14688 18634
rect 14646 18592 14702 18601
rect 14646 18527 14702 18536
rect 14752 18290 14780 20216
rect 14936 20074 14964 20334
rect 14844 20046 14964 20074
rect 14844 19242 14872 20046
rect 14924 19848 14976 19854
rect 14924 19790 14976 19796
rect 14936 19514 14964 19790
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 15016 19440 15068 19446
rect 14922 19408 14978 19417
rect 15212 19402 15240 20470
rect 15016 19382 15068 19388
rect 15200 19396 15252 19402
rect 14922 19343 14978 19352
rect 14832 19236 14884 19242
rect 14832 19178 14884 19184
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14648 18216 14700 18222
rect 14648 18158 14700 18164
rect 14660 18034 14688 18158
rect 14738 18048 14794 18057
rect 14660 18006 14738 18034
rect 14738 17983 14794 17992
rect 14844 17898 14872 18226
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14752 17870 14872 17898
rect 14660 14822 14688 17818
rect 14752 17814 14780 17870
rect 14740 17808 14792 17814
rect 14740 17750 14792 17756
rect 14832 17808 14884 17814
rect 14832 17750 14884 17756
rect 14844 17649 14872 17750
rect 14830 17640 14886 17649
rect 14740 17604 14792 17610
rect 14830 17575 14886 17584
rect 14740 17546 14792 17552
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14648 14544 14700 14550
rect 14648 14486 14700 14492
rect 14660 14346 14688 14486
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14646 13968 14702 13977
rect 14556 13932 14608 13938
rect 14752 13954 14780 17546
rect 14936 17134 14964 19343
rect 15028 18970 15056 19382
rect 15304 19378 15332 23462
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 15396 20806 15424 23054
rect 15488 22438 15516 24783
rect 15580 23594 15608 26862
rect 15752 25764 15804 25770
rect 15752 25706 15804 25712
rect 15658 23760 15714 23769
rect 15658 23695 15660 23704
rect 15712 23695 15714 23704
rect 15660 23666 15712 23672
rect 15568 23588 15620 23594
rect 15568 23530 15620 23536
rect 15764 23526 15792 25706
rect 15856 24857 15884 28426
rect 16212 28416 16264 28422
rect 16212 28358 16264 28364
rect 16026 27704 16082 27713
rect 16026 27639 16028 27648
rect 16080 27639 16082 27648
rect 16028 27610 16080 27616
rect 16118 27160 16174 27169
rect 16118 27095 16174 27104
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 15948 25945 15976 26930
rect 16028 26784 16080 26790
rect 16028 26726 16080 26732
rect 16040 26586 16068 26726
rect 16028 26580 16080 26586
rect 16028 26522 16080 26528
rect 16040 26489 16068 26522
rect 16026 26480 16082 26489
rect 16026 26415 16082 26424
rect 15934 25936 15990 25945
rect 15934 25871 15990 25880
rect 15948 25140 15976 25871
rect 16040 25294 16068 26415
rect 16132 26314 16160 27095
rect 16120 26308 16172 26314
rect 16120 26250 16172 26256
rect 16132 25430 16160 26250
rect 16120 25424 16172 25430
rect 16120 25366 16172 25372
rect 16028 25288 16080 25294
rect 16028 25230 16080 25236
rect 16120 25220 16172 25226
rect 16120 25162 16172 25168
rect 15948 25112 16068 25140
rect 15842 24848 15898 24857
rect 15842 24783 15898 24792
rect 15936 24676 15988 24682
rect 15936 24618 15988 24624
rect 15752 23520 15804 23526
rect 15752 23462 15804 23468
rect 15660 22976 15712 22982
rect 15660 22918 15712 22924
rect 15476 22432 15528 22438
rect 15476 22374 15528 22380
rect 15672 22030 15700 22918
rect 15752 22092 15804 22098
rect 15752 22034 15804 22040
rect 15660 22024 15712 22030
rect 15660 21966 15712 21972
rect 15476 21548 15528 21554
rect 15476 21490 15528 21496
rect 15488 21078 15516 21490
rect 15476 21072 15528 21078
rect 15476 21014 15528 21020
rect 15384 20800 15436 20806
rect 15672 20754 15700 21966
rect 15384 20742 15436 20748
rect 15488 20726 15700 20754
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15200 19338 15252 19344
rect 15292 19372 15344 19378
rect 15292 19314 15344 19320
rect 15108 19168 15160 19174
rect 15106 19136 15108 19145
rect 15200 19168 15252 19174
rect 15160 19136 15162 19145
rect 15200 19110 15252 19116
rect 15106 19071 15162 19080
rect 15212 18986 15240 19110
rect 15016 18964 15068 18970
rect 15016 18906 15068 18912
rect 15120 18958 15240 18986
rect 15290 19000 15346 19009
rect 15028 18086 15056 18906
rect 15016 18080 15068 18086
rect 15016 18022 15068 18028
rect 15120 17898 15148 18958
rect 15290 18935 15346 18944
rect 15304 18426 15332 18935
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15028 17870 15148 17898
rect 15212 17882 15240 18022
rect 15200 17876 15252 17882
rect 15028 17338 15056 17870
rect 15200 17818 15252 17824
rect 15106 17776 15162 17785
rect 15106 17711 15162 17720
rect 15016 17332 15068 17338
rect 15016 17274 15068 17280
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14844 16726 14872 17070
rect 14832 16720 14884 16726
rect 14832 16662 14884 16668
rect 14936 15706 14964 17070
rect 15016 16720 15068 16726
rect 15016 16662 15068 16668
rect 15120 16674 15148 17711
rect 15212 17678 15240 17818
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15304 17338 15332 17750
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15396 16726 15424 20198
rect 15488 18290 15516 20726
rect 15764 20602 15792 22034
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15752 20596 15804 20602
rect 15752 20538 15804 20544
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15488 17377 15516 17478
rect 15474 17368 15530 17377
rect 15474 17303 15530 17312
rect 15580 16833 15608 20402
rect 15660 20256 15712 20262
rect 15660 20198 15712 20204
rect 15672 19922 15700 20198
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15752 19440 15804 19446
rect 15752 19382 15804 19388
rect 15658 18456 15714 18465
rect 15658 18391 15714 18400
rect 15672 18290 15700 18391
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15566 16824 15622 16833
rect 15672 16794 15700 17274
rect 15566 16759 15622 16768
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15384 16720 15436 16726
rect 15028 16522 15056 16662
rect 15120 16646 15332 16674
rect 15384 16662 15436 16668
rect 15108 16584 15160 16590
rect 15200 16584 15252 16590
rect 15108 16526 15160 16532
rect 15198 16552 15200 16561
rect 15304 16572 15332 16646
rect 15252 16552 15254 16561
rect 15304 16544 15424 16572
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 15028 16425 15056 16458
rect 15014 16416 15070 16425
rect 15014 16351 15070 16360
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 15028 15858 15056 16050
rect 15120 15960 15148 16526
rect 15198 16487 15254 16496
rect 15396 16114 15424 16544
rect 15476 16516 15528 16522
rect 15476 16458 15528 16464
rect 15384 16108 15436 16114
rect 15384 16050 15436 16056
rect 15120 15932 15332 15960
rect 15028 15830 15240 15858
rect 15212 15706 15240 15830
rect 15304 15706 15332 15932
rect 15396 15722 15424 16050
rect 15488 16028 15516 16458
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15488 16000 15608 16028
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15292 15700 15344 15706
rect 15396 15694 15516 15722
rect 15292 15642 15344 15648
rect 15016 15496 15068 15502
rect 15014 15464 15016 15473
rect 15068 15464 15070 15473
rect 15014 15399 15070 15408
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 14936 14074 14964 14826
rect 15028 14618 15056 15399
rect 15016 14612 15068 14618
rect 15016 14554 15068 14560
rect 15120 14521 15148 15642
rect 15384 15632 15436 15638
rect 15384 15574 15436 15580
rect 15396 15502 15424 15574
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15488 15348 15516 15694
rect 15396 15320 15516 15348
rect 15198 15056 15254 15065
rect 15198 14991 15254 15000
rect 15106 14512 15162 14521
rect 15106 14447 15162 14456
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 14702 13926 14780 13954
rect 14830 13968 14886 13977
rect 14646 13903 14702 13912
rect 14830 13903 14886 13912
rect 14556 13874 14608 13880
rect 14568 13530 14596 13874
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14752 13326 14780 13670
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14554 12472 14610 12481
rect 14476 12416 14554 12434
rect 14752 12434 14780 13262
rect 14844 13025 14872 13903
rect 14936 13734 14964 14010
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14830 13016 14886 13025
rect 14830 12951 14886 12960
rect 14936 12782 14964 13126
rect 15028 12832 15056 13806
rect 15120 13002 15148 14447
rect 15212 14278 15240 14991
rect 15292 14816 15344 14822
rect 15290 14784 15292 14793
rect 15344 14784 15346 14793
rect 15290 14719 15346 14728
rect 15396 14346 15424 15320
rect 15580 14600 15608 16000
rect 15672 15688 15700 16390
rect 15764 15978 15792 19382
rect 15752 15972 15804 15978
rect 15752 15914 15804 15920
rect 15672 15660 15792 15688
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15488 14572 15608 14600
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 15304 13326 15332 13738
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15382 13152 15438 13161
rect 15382 13087 15438 13096
rect 15290 13016 15346 13025
rect 15120 12974 15240 13002
rect 15108 12844 15160 12850
rect 15028 12804 15108 12832
rect 15108 12786 15160 12792
rect 14924 12776 14976 12782
rect 15212 12730 15240 12974
rect 15290 12951 15346 12960
rect 15304 12850 15332 12951
rect 15396 12850 15424 13087
rect 15488 12986 15516 14572
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 14924 12718 14976 12724
rect 14832 12708 14884 12714
rect 14832 12650 14884 12656
rect 15028 12702 15240 12730
rect 14476 12407 14610 12416
rect 14476 12406 14596 12407
rect 14660 12406 14780 12434
rect 14476 11937 14504 12406
rect 14554 12336 14610 12345
rect 14554 12271 14610 12280
rect 14462 11928 14518 11937
rect 14462 11863 14518 11872
rect 14568 11830 14596 12271
rect 14556 11824 14608 11830
rect 14462 11792 14518 11801
rect 14556 11766 14608 11772
rect 14462 11727 14518 11736
rect 14292 11614 14412 11642
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14292 11218 14320 11494
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 14384 10690 14412 11614
rect 14476 11150 14504 11727
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14292 10662 14412 10690
rect 14556 10668 14608 10674
rect 14292 9489 14320 10662
rect 14556 10610 14608 10616
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14384 9654 14412 10542
rect 14462 10296 14518 10305
rect 14462 10231 14518 10240
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14278 9480 14334 9489
rect 14278 9415 14334 9424
rect 14278 9208 14334 9217
rect 14278 9143 14334 9152
rect 14292 8945 14320 9143
rect 14476 9058 14504 10231
rect 14568 10130 14596 10610
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14554 9208 14610 9217
rect 14554 9143 14556 9152
rect 14608 9143 14610 9152
rect 14556 9114 14608 9120
rect 14476 9030 14596 9058
rect 14372 8968 14424 8974
rect 14278 8936 14334 8945
rect 14372 8910 14424 8916
rect 14278 8871 14334 8880
rect 14384 8634 14412 8910
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14568 8401 14596 9030
rect 14554 8392 14610 8401
rect 14554 8327 14610 8336
rect 14464 8016 14516 8022
rect 14464 7958 14516 7964
rect 14554 7984 14610 7993
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 14384 7546 14412 7822
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14476 7478 14504 7958
rect 14554 7919 14556 7928
rect 14608 7919 14610 7928
rect 14556 7890 14608 7896
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14464 7472 14516 7478
rect 14464 7414 14516 7420
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14108 5574 14136 6394
rect 14200 5914 14228 6394
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 13726 5400 13782 5409
rect 13726 5335 13782 5344
rect 14292 5234 14320 7210
rect 14464 6724 14516 6730
rect 14464 6666 14516 6672
rect 14476 5914 14504 6666
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14372 5296 14424 5302
rect 14370 5264 14372 5273
rect 14424 5264 14426 5273
rect 14280 5228 14332 5234
rect 14476 5234 14504 5510
rect 14370 5199 14426 5208
rect 14464 5228 14516 5234
rect 14280 5170 14332 5176
rect 14464 5170 14516 5176
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14384 4758 14412 4966
rect 14568 4842 14596 7754
rect 14660 5098 14688 12406
rect 14738 11792 14794 11801
rect 14844 11762 14872 12650
rect 15028 11880 15056 12702
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 14936 11852 15056 11880
rect 15108 11892 15160 11898
rect 14738 11727 14794 11736
rect 14832 11756 14884 11762
rect 14752 11558 14780 11727
rect 14832 11698 14884 11704
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14844 11286 14872 11698
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14844 9500 14872 11086
rect 14752 9472 14872 9500
rect 14648 5092 14700 5098
rect 14648 5034 14700 5040
rect 14476 4826 14596 4842
rect 14660 4826 14688 5034
rect 14752 4826 14780 9472
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14844 8838 14872 9318
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14936 8378 14964 11852
rect 15108 11834 15160 11840
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 15028 11665 15056 11698
rect 15014 11656 15070 11665
rect 15014 11591 15070 11600
rect 15016 11008 15068 11014
rect 15120 10985 15148 11834
rect 15016 10950 15068 10956
rect 15106 10976 15162 10985
rect 15028 8673 15056 10950
rect 15106 10911 15162 10920
rect 15212 10674 15240 12582
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15106 9616 15162 9625
rect 15106 9551 15162 9560
rect 15120 9110 15148 9551
rect 15108 9104 15160 9110
rect 15108 9046 15160 9052
rect 15014 8664 15070 8673
rect 15014 8599 15070 8608
rect 15014 8528 15070 8537
rect 15198 8528 15254 8537
rect 15108 8492 15160 8498
rect 15070 8472 15108 8480
rect 15014 8463 15108 8472
rect 15028 8452 15108 8463
rect 15198 8463 15200 8472
rect 15108 8434 15160 8440
rect 15252 8463 15254 8472
rect 15200 8434 15252 8440
rect 14844 8350 14964 8378
rect 15014 8392 15070 8401
rect 14844 7002 14872 8350
rect 15014 8327 15070 8336
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 14936 6458 14964 8230
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 15028 5234 15056 8327
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 15120 6798 15148 8230
rect 15212 7732 15240 8434
rect 15304 8294 15332 12786
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15488 12434 15516 12582
rect 15396 12406 15516 12434
rect 15396 9364 15424 12406
rect 15474 11928 15530 11937
rect 15474 11863 15530 11872
rect 15488 11830 15516 11863
rect 15476 11824 15528 11830
rect 15476 11766 15528 11772
rect 15476 11688 15528 11694
rect 15476 11630 15528 11636
rect 15488 11558 15516 11630
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15488 11286 15516 11494
rect 15580 11354 15608 14282
rect 15672 12918 15700 15506
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15672 12646 15700 12854
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15488 10470 15516 10950
rect 15580 10470 15608 11290
rect 15764 11150 15792 15660
rect 15856 15366 15884 21490
rect 15948 21146 15976 24618
rect 16040 22982 16068 25112
rect 16132 24886 16160 25162
rect 16120 24880 16172 24886
rect 16120 24822 16172 24828
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 16028 22976 16080 22982
rect 16028 22918 16080 22924
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 15948 21010 15976 21082
rect 15936 21004 15988 21010
rect 15936 20946 15988 20952
rect 16132 20890 16160 23666
rect 16224 22438 16252 28358
rect 16316 27606 16344 29106
rect 16408 28558 16436 29242
rect 16396 28552 16448 28558
rect 16396 28494 16448 28500
rect 16592 28082 16620 29582
rect 17224 29572 17276 29578
rect 17224 29514 17276 29520
rect 16856 29504 16908 29510
rect 16856 29446 16908 29452
rect 16868 29238 16896 29446
rect 16856 29232 16908 29238
rect 16856 29174 16908 29180
rect 17236 29034 17264 29514
rect 17408 29504 17460 29510
rect 17408 29446 17460 29452
rect 17420 29170 17448 29446
rect 17408 29164 17460 29170
rect 17408 29106 17460 29112
rect 17224 29028 17276 29034
rect 17224 28970 17276 28976
rect 17316 28756 17368 28762
rect 17316 28698 17368 28704
rect 17328 28490 17356 28698
rect 17316 28484 17368 28490
rect 17316 28426 17368 28432
rect 16580 28076 16632 28082
rect 16580 28018 16632 28024
rect 16672 28008 16724 28014
rect 16672 27950 16724 27956
rect 16396 27668 16448 27674
rect 16396 27610 16448 27616
rect 16304 27600 16356 27606
rect 16304 27542 16356 27548
rect 16304 27328 16356 27334
rect 16304 27270 16356 27276
rect 16316 26489 16344 27270
rect 16302 26480 16358 26489
rect 16302 26415 16358 26424
rect 16304 26376 16356 26382
rect 16408 26330 16436 27610
rect 16488 27464 16540 27470
rect 16488 27406 16540 27412
rect 16500 26858 16528 27406
rect 16488 26852 16540 26858
rect 16488 26794 16540 26800
rect 16356 26324 16436 26330
rect 16304 26318 16436 26324
rect 16316 26302 16436 26318
rect 16488 26308 16540 26314
rect 16316 24818 16344 26302
rect 16488 26250 16540 26256
rect 16396 25288 16448 25294
rect 16396 25230 16448 25236
rect 16408 25158 16436 25230
rect 16396 25152 16448 25158
rect 16396 25094 16448 25100
rect 16408 24954 16436 25094
rect 16396 24948 16448 24954
rect 16396 24890 16448 24896
rect 16304 24812 16356 24818
rect 16304 24754 16356 24760
rect 16316 24410 16344 24754
rect 16304 24404 16356 24410
rect 16304 24346 16356 24352
rect 16396 24404 16448 24410
rect 16396 24346 16448 24352
rect 16304 23316 16356 23322
rect 16304 23258 16356 23264
rect 16212 22432 16264 22438
rect 16212 22374 16264 22380
rect 15948 20862 16160 20890
rect 15948 19553 15976 20862
rect 16120 20800 16172 20806
rect 16120 20742 16172 20748
rect 16028 20528 16080 20534
rect 16028 20470 16080 20476
rect 16040 20058 16068 20470
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 15934 19544 15990 19553
rect 15934 19479 15990 19488
rect 15948 17270 15976 19479
rect 16132 19394 16160 20742
rect 16210 20632 16266 20641
rect 16210 20567 16266 20576
rect 16224 19514 16252 20567
rect 16316 20398 16344 23258
rect 16408 23118 16436 24346
rect 16500 23798 16528 26250
rect 16684 25974 16712 27950
rect 16856 27872 16908 27878
rect 16856 27814 16908 27820
rect 16868 26994 16896 27814
rect 17224 27464 17276 27470
rect 16946 27432 17002 27441
rect 17224 27406 17276 27412
rect 16946 27367 16948 27376
rect 17000 27367 17002 27376
rect 16948 27338 17000 27344
rect 16856 26988 16908 26994
rect 16856 26930 16908 26936
rect 16762 26072 16818 26081
rect 16762 26007 16818 26016
rect 16672 25968 16724 25974
rect 16672 25910 16724 25916
rect 16776 25906 16804 26007
rect 16764 25900 16816 25906
rect 16764 25842 16816 25848
rect 16672 25288 16724 25294
rect 16672 25230 16724 25236
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16488 23792 16540 23798
rect 16488 23734 16540 23740
rect 16592 23474 16620 25094
rect 16684 24954 16712 25230
rect 16776 25129 16804 25842
rect 16868 25673 16896 26930
rect 17132 26920 17184 26926
rect 17132 26862 17184 26868
rect 16946 25936 17002 25945
rect 16946 25871 16948 25880
rect 17000 25871 17002 25880
rect 16948 25842 17000 25848
rect 16854 25664 16910 25673
rect 16854 25599 16910 25608
rect 16856 25152 16908 25158
rect 16762 25120 16818 25129
rect 16856 25094 16908 25100
rect 16762 25055 16818 25064
rect 16672 24948 16724 24954
rect 16672 24890 16724 24896
rect 16868 24818 16896 25094
rect 16960 24818 16988 25842
rect 17038 25664 17094 25673
rect 17038 25599 17094 25608
rect 17052 25362 17080 25599
rect 17040 25356 17092 25362
rect 17040 25298 17092 25304
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 16948 24812 17000 24818
rect 16948 24754 17000 24760
rect 16500 23446 16620 23474
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16396 22976 16448 22982
rect 16396 22918 16448 22924
rect 16408 22574 16436 22918
rect 16500 22642 16528 23446
rect 16578 23352 16634 23361
rect 16578 23287 16580 23296
rect 16632 23287 16634 23296
rect 16580 23258 16632 23264
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 16488 22636 16540 22642
rect 16488 22578 16540 22584
rect 16396 22568 16448 22574
rect 16396 22510 16448 22516
rect 16396 22432 16448 22438
rect 16396 22374 16448 22380
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16028 19372 16080 19378
rect 16132 19366 16252 19394
rect 16028 19314 16080 19320
rect 16040 19009 16068 19314
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16026 19000 16082 19009
rect 16026 18935 16082 18944
rect 16026 18728 16082 18737
rect 16026 18663 16082 18672
rect 16040 18465 16068 18663
rect 16026 18456 16082 18465
rect 16026 18391 16082 18400
rect 16132 18358 16160 19110
rect 16120 18352 16172 18358
rect 16120 18294 16172 18300
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 15936 17264 15988 17270
rect 15936 17206 15988 17212
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 16040 16794 16068 16934
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 15948 16640 15976 16730
rect 16028 16652 16080 16658
rect 15948 16612 16028 16640
rect 16028 16594 16080 16600
rect 15934 16552 15990 16561
rect 15934 16487 15990 16496
rect 15948 16454 15976 16487
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15936 15972 15988 15978
rect 15936 15914 15988 15920
rect 15948 15745 15976 15914
rect 15934 15736 15990 15745
rect 15934 15671 15990 15680
rect 15934 15600 15990 15609
rect 15934 15535 15990 15544
rect 15844 15360 15896 15366
rect 15844 15302 15896 15308
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 15856 13802 15884 15098
rect 15948 13938 15976 15535
rect 16040 14278 16068 16594
rect 16132 16017 16160 17478
rect 16118 16008 16174 16017
rect 16118 15943 16174 15952
rect 16224 15638 16252 19366
rect 16316 18834 16344 20334
rect 16408 19145 16436 22374
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16500 20602 16528 20946
rect 16488 20596 16540 20602
rect 16488 20538 16540 20544
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 16500 20058 16528 20402
rect 16592 20097 16620 23122
rect 16578 20088 16634 20097
rect 16488 20052 16540 20058
rect 16578 20023 16634 20032
rect 16488 19994 16540 20000
rect 16684 19854 16712 24754
rect 16946 24712 17002 24721
rect 16946 24647 17002 24656
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16868 23186 16896 23666
rect 16856 23180 16908 23186
rect 16856 23122 16908 23128
rect 16960 22982 16988 24647
rect 17038 23760 17094 23769
rect 17038 23695 17094 23704
rect 16948 22976 17000 22982
rect 16762 22944 16818 22953
rect 16948 22918 17000 22924
rect 16762 22879 16818 22888
rect 16776 21185 16804 22879
rect 16946 22808 17002 22817
rect 16946 22743 17002 22752
rect 16854 22128 16910 22137
rect 16854 22063 16910 22072
rect 16868 21350 16896 22063
rect 16856 21344 16908 21350
rect 16960 21321 16988 22743
rect 16856 21286 16908 21292
rect 16946 21312 17002 21321
rect 16762 21176 16818 21185
rect 16762 21111 16818 21120
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16776 20330 16804 20402
rect 16764 20324 16816 20330
rect 16764 20266 16816 20272
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 16500 19514 16528 19790
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16394 19136 16450 19145
rect 16394 19071 16450 19080
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 16302 17776 16358 17785
rect 16302 17711 16304 17720
rect 16356 17711 16358 17720
rect 16304 17682 16356 17688
rect 16396 17264 16448 17270
rect 16396 17206 16448 17212
rect 16408 16674 16436 17206
rect 16500 16794 16528 18906
rect 16592 18902 16620 19246
rect 16580 18896 16632 18902
rect 16580 18838 16632 18844
rect 16684 17542 16712 19654
rect 16776 18970 16804 19790
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16776 18222 16804 18566
rect 16868 18358 16896 21286
rect 16946 21247 17002 21256
rect 17052 20602 17080 23695
rect 17144 22166 17172 26862
rect 17236 26314 17264 27406
rect 17316 27328 17368 27334
rect 17316 27270 17368 27276
rect 17328 27062 17356 27270
rect 17316 27056 17368 27062
rect 17316 26998 17368 27004
rect 17408 26784 17460 26790
rect 17408 26726 17460 26732
rect 17420 26602 17448 26726
rect 17328 26574 17448 26602
rect 17224 26308 17276 26314
rect 17224 26250 17276 26256
rect 17224 25764 17276 25770
rect 17224 25706 17276 25712
rect 17236 25430 17264 25706
rect 17224 25424 17276 25430
rect 17224 25366 17276 25372
rect 17224 25288 17276 25294
rect 17224 25230 17276 25236
rect 17236 23361 17264 25230
rect 17222 23352 17278 23361
rect 17222 23287 17278 23296
rect 17224 22636 17276 22642
rect 17224 22578 17276 22584
rect 17132 22160 17184 22166
rect 17132 22102 17184 22108
rect 17144 21486 17172 22102
rect 17132 21480 17184 21486
rect 17132 21422 17184 21428
rect 17040 20596 17092 20602
rect 17040 20538 17092 20544
rect 17236 20466 17264 22578
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 16856 18352 16908 18358
rect 16856 18294 16908 18300
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16592 16794 16620 17138
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16408 16646 16528 16674
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 16396 16516 16448 16522
rect 16396 16458 16448 16464
rect 16316 16046 16344 16458
rect 16408 16182 16436 16458
rect 16396 16176 16448 16182
rect 16396 16118 16448 16124
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16132 14550 16160 15438
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15844 13796 15896 13802
rect 15844 13738 15896 13744
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15856 12442 15884 13262
rect 15948 13258 15976 13874
rect 16040 13870 16068 14214
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 15936 13252 15988 13258
rect 15936 13194 15988 13200
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15842 12336 15898 12345
rect 15842 12271 15898 12280
rect 15856 12073 15884 12271
rect 15842 12064 15898 12073
rect 15842 11999 15898 12008
rect 15948 11286 15976 12786
rect 16040 12306 16068 12786
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 15488 9489 15516 10202
rect 15566 9616 15622 9625
rect 15566 9551 15568 9560
rect 15620 9551 15622 9560
rect 15568 9522 15620 9528
rect 15474 9480 15530 9489
rect 15474 9415 15530 9424
rect 15396 9336 15516 9364
rect 15382 8392 15438 8401
rect 15382 8327 15384 8336
rect 15436 8327 15438 8336
rect 15384 8298 15436 8304
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15382 8256 15438 8265
rect 15382 8191 15438 8200
rect 15212 7704 15332 7732
rect 15198 6896 15254 6905
rect 15198 6831 15254 6840
rect 15212 6798 15240 6831
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15120 5846 15148 6258
rect 15108 5840 15160 5846
rect 15108 5782 15160 5788
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 14464 4820 14596 4826
rect 14516 4814 14596 4820
rect 14464 4762 14516 4768
rect 14372 4752 14424 4758
rect 14372 4694 14424 4700
rect 14568 4622 14596 4814
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14660 4622 14688 4762
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 15120 3641 15148 5782
rect 15304 5710 15332 7704
rect 15396 7324 15424 8191
rect 15488 7478 15516 9336
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15580 8294 15608 8434
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15672 7993 15700 10950
rect 15856 10577 15884 11086
rect 15948 10742 15976 11222
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 16040 10690 16068 12242
rect 16132 11830 16160 14486
rect 16224 14414 16252 14758
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16316 14006 16344 15982
rect 16408 15162 16436 16118
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16500 14618 16528 16646
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16396 14408 16448 14414
rect 16396 14350 16448 14356
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 16224 12646 16252 13874
rect 16304 13796 16356 13802
rect 16304 13738 16356 13744
rect 16316 12646 16344 13738
rect 16408 12782 16436 14350
rect 16500 12850 16528 14350
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16396 12776 16448 12782
rect 16396 12718 16448 12724
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16408 12442 16436 12718
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16592 12102 16620 16594
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16684 16250 16712 16526
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16776 15858 16804 18158
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16868 17066 16896 17614
rect 16856 17060 16908 17066
rect 16856 17002 16908 17008
rect 16684 15830 16804 15858
rect 16684 14822 16712 15830
rect 16762 15736 16818 15745
rect 16762 15671 16764 15680
rect 16816 15671 16818 15680
rect 16764 15642 16816 15648
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16776 14929 16804 15098
rect 16762 14920 16818 14929
rect 16762 14855 16818 14864
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16762 14784 16818 14793
rect 16762 14719 16818 14728
rect 16776 14618 16804 14719
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16684 13938 16712 14554
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16684 12442 16712 13194
rect 16764 12912 16816 12918
rect 16868 12900 16896 17002
rect 16960 16998 16988 20402
rect 17130 20360 17186 20369
rect 17130 20295 17132 20304
rect 17184 20295 17186 20304
rect 17132 20266 17184 20272
rect 17236 20058 17264 20402
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17040 19984 17092 19990
rect 17040 19926 17092 19932
rect 17052 19174 17080 19926
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 17328 18714 17356 26574
rect 17408 26512 17460 26518
rect 17408 26454 17460 26460
rect 17420 25974 17448 26454
rect 17408 25968 17460 25974
rect 17408 25910 17460 25916
rect 17420 25294 17448 25910
rect 17512 25770 17540 29582
rect 18420 29572 18472 29578
rect 18420 29514 18472 29520
rect 18432 29238 18460 29514
rect 18420 29232 18472 29238
rect 18420 29174 18472 29180
rect 18142 29064 18198 29073
rect 18142 28999 18144 29008
rect 18196 28999 18198 29008
rect 18144 28970 18196 28976
rect 18420 28960 18472 28966
rect 18420 28902 18472 28908
rect 18432 28778 18460 28902
rect 18064 28750 18460 28778
rect 17960 28688 18012 28694
rect 17960 28630 18012 28636
rect 17684 28416 17736 28422
rect 17684 28358 17736 28364
rect 17592 27668 17644 27674
rect 17592 27610 17644 27616
rect 17604 27334 17632 27610
rect 17592 27328 17644 27334
rect 17592 27270 17644 27276
rect 17592 26308 17644 26314
rect 17592 26250 17644 26256
rect 17500 25764 17552 25770
rect 17500 25706 17552 25712
rect 17498 25664 17554 25673
rect 17498 25599 17554 25608
rect 17512 25498 17540 25599
rect 17500 25492 17552 25498
rect 17500 25434 17552 25440
rect 17408 25288 17460 25294
rect 17408 25230 17460 25236
rect 17500 25288 17552 25294
rect 17500 25230 17552 25236
rect 17512 24857 17540 25230
rect 17498 24848 17554 24857
rect 17604 24818 17632 26250
rect 17498 24783 17554 24792
rect 17592 24812 17644 24818
rect 17408 24608 17460 24614
rect 17406 24576 17408 24585
rect 17460 24576 17462 24585
rect 17406 24511 17462 24520
rect 17512 24041 17540 24783
rect 17592 24754 17644 24760
rect 17498 24032 17554 24041
rect 17498 23967 17554 23976
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17512 22760 17540 23462
rect 17604 23186 17632 24754
rect 17696 23798 17724 28358
rect 17776 27940 17828 27946
rect 17776 27882 17828 27888
rect 17788 27470 17816 27882
rect 17972 27878 18000 28630
rect 18064 28558 18092 28750
rect 18432 28694 18460 28750
rect 18420 28688 18472 28694
rect 18248 28626 18368 28642
rect 18420 28630 18472 28636
rect 18236 28620 18368 28626
rect 18288 28614 18368 28620
rect 18236 28562 18288 28568
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 18236 28484 18288 28490
rect 18236 28426 18288 28432
rect 18142 28112 18198 28121
rect 18142 28047 18198 28056
rect 18156 28014 18184 28047
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 17960 27872 18012 27878
rect 18012 27832 18092 27860
rect 17960 27814 18012 27820
rect 17960 27668 18012 27674
rect 17960 27610 18012 27616
rect 17776 27464 17828 27470
rect 17972 27441 18000 27610
rect 17776 27406 17828 27412
rect 17958 27432 18014 27441
rect 17868 27396 17920 27402
rect 17958 27367 18014 27376
rect 17868 27338 17920 27344
rect 17776 26784 17828 26790
rect 17776 26726 17828 26732
rect 17788 26353 17816 26726
rect 17774 26344 17830 26353
rect 17774 26279 17830 26288
rect 17776 25288 17828 25294
rect 17776 25230 17828 25236
rect 17684 23792 17736 23798
rect 17684 23734 17736 23740
rect 17592 23180 17644 23186
rect 17592 23122 17644 23128
rect 17590 23080 17646 23089
rect 17696 23050 17724 23734
rect 17788 23474 17816 25230
rect 17880 24954 17908 27338
rect 18064 25242 18092 27832
rect 18248 26994 18276 28426
rect 18340 28150 18368 28614
rect 18420 28552 18472 28558
rect 18420 28494 18472 28500
rect 18432 28257 18460 28494
rect 18418 28248 18474 28257
rect 18418 28183 18474 28192
rect 18328 28144 18380 28150
rect 18328 28086 18380 28092
rect 18420 27532 18472 27538
rect 18420 27474 18472 27480
rect 18236 26988 18288 26994
rect 18236 26930 18288 26936
rect 18248 26382 18276 26930
rect 18432 26908 18460 27474
rect 18524 27441 18552 30670
rect 19352 30258 19380 31282
rect 21928 30394 21956 31282
rect 23110 31240 23166 31249
rect 23110 31175 23166 31184
rect 21916 30388 21968 30394
rect 21916 30330 21968 30336
rect 23018 30288 23074 30297
rect 18696 30252 18748 30258
rect 18696 30194 18748 30200
rect 19340 30252 19392 30258
rect 19340 30194 19392 30200
rect 20536 30252 20588 30258
rect 23018 30223 23074 30232
rect 20536 30194 20588 30200
rect 18708 29850 18736 30194
rect 18880 30048 18932 30054
rect 18880 29990 18932 29996
rect 18696 29844 18748 29850
rect 18696 29786 18748 29792
rect 18892 29646 18920 29990
rect 20548 29850 20576 30194
rect 20628 30048 20680 30054
rect 20628 29990 20680 29996
rect 20904 30048 20956 30054
rect 20904 29990 20956 29996
rect 22192 30048 22244 30054
rect 22192 29990 22244 29996
rect 20536 29844 20588 29850
rect 20536 29786 20588 29792
rect 20640 29714 20668 29990
rect 20628 29708 20680 29714
rect 20628 29650 20680 29656
rect 18880 29640 18932 29646
rect 18880 29582 18932 29588
rect 20166 29336 20222 29345
rect 20166 29271 20222 29280
rect 20180 29170 20208 29271
rect 20168 29164 20220 29170
rect 20168 29106 20220 29112
rect 19616 28960 19668 28966
rect 19616 28902 19668 28908
rect 19892 28960 19944 28966
rect 20180 28937 20208 29106
rect 19892 28902 19944 28908
rect 20166 28928 20222 28937
rect 19522 28792 19578 28801
rect 19432 28756 19484 28762
rect 19522 28727 19578 28736
rect 19432 28698 19484 28704
rect 19340 28688 19392 28694
rect 19340 28630 19392 28636
rect 18972 28416 19024 28422
rect 19352 28393 19380 28630
rect 19444 28422 19472 28698
rect 19432 28416 19484 28422
rect 18972 28358 19024 28364
rect 19338 28384 19394 28393
rect 18604 27872 18656 27878
rect 18604 27814 18656 27820
rect 18616 27713 18644 27814
rect 18602 27704 18658 27713
rect 18602 27639 18658 27648
rect 18880 27668 18932 27674
rect 18880 27614 18932 27616
rect 18800 27610 18932 27614
rect 18800 27586 18920 27610
rect 18800 27520 18828 27586
rect 18984 27520 19012 28358
rect 19432 28358 19484 28364
rect 19338 28319 19394 28328
rect 19156 28076 19208 28082
rect 19156 28018 19208 28024
rect 19168 27577 19196 28018
rect 19248 28008 19300 28014
rect 19248 27950 19300 27956
rect 18792 27492 18828 27520
rect 18892 27492 19012 27520
rect 19154 27568 19210 27577
rect 19260 27538 19288 27950
rect 19340 27668 19392 27674
rect 19340 27610 19392 27616
rect 19444 27614 19472 28358
rect 19536 28064 19564 28727
rect 19628 28665 19656 28902
rect 19904 28762 19932 28902
rect 20166 28863 20222 28872
rect 19892 28756 19944 28762
rect 19892 28698 19944 28704
rect 19984 28756 20036 28762
rect 19984 28698 20036 28704
rect 19614 28656 19670 28665
rect 19614 28591 19670 28600
rect 19616 28076 19668 28082
rect 19536 28036 19616 28064
rect 19616 28018 19668 28024
rect 19904 27878 19932 28698
rect 19996 28422 20024 28698
rect 20352 28688 20404 28694
rect 20352 28630 20404 28636
rect 20168 28620 20220 28626
rect 20220 28580 20300 28608
rect 20168 28562 20220 28568
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 20168 28416 20220 28422
rect 20168 28358 20220 28364
rect 19892 27872 19944 27878
rect 19944 27832 20116 27860
rect 19892 27814 19944 27820
rect 19352 27554 19380 27610
rect 19444 27586 19748 27614
rect 19720 27554 19748 27586
rect 19982 27568 20038 27577
rect 19154 27503 19210 27512
rect 19248 27532 19300 27538
rect 18696 27464 18748 27470
rect 18510 27432 18566 27441
rect 18696 27406 18748 27412
rect 18510 27367 18566 27376
rect 18524 27062 18552 27367
rect 18602 27296 18658 27305
rect 18602 27231 18658 27240
rect 18616 27062 18644 27231
rect 18512 27056 18564 27062
rect 18512 26998 18564 27004
rect 18604 27056 18656 27062
rect 18604 26998 18656 27004
rect 18432 26880 18644 26908
rect 18510 26752 18566 26761
rect 18510 26687 18566 26696
rect 18420 26580 18472 26586
rect 18420 26522 18472 26528
rect 18236 26376 18288 26382
rect 18236 26318 18288 26324
rect 18328 26240 18380 26246
rect 18328 26182 18380 26188
rect 17972 25214 18092 25242
rect 17868 24948 17920 24954
rect 17868 24890 17920 24896
rect 17972 24721 18000 25214
rect 18052 25152 18104 25158
rect 18052 25094 18104 25100
rect 18236 25152 18288 25158
rect 18236 25094 18288 25100
rect 18064 24818 18092 25094
rect 18248 24886 18276 25094
rect 18236 24880 18288 24886
rect 18236 24822 18288 24828
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 17958 24712 18014 24721
rect 18064 24682 18092 24754
rect 17958 24647 18014 24656
rect 18052 24676 18104 24682
rect 18052 24618 18104 24624
rect 18156 24410 18184 24754
rect 18248 24614 18276 24822
rect 18236 24608 18288 24614
rect 18236 24550 18288 24556
rect 18144 24404 18196 24410
rect 18144 24346 18196 24352
rect 18144 23860 18196 23866
rect 18144 23802 18196 23808
rect 18052 23588 18104 23594
rect 18052 23530 18104 23536
rect 17958 23488 18014 23497
rect 17788 23446 17908 23474
rect 17776 23316 17828 23322
rect 17776 23258 17828 23264
rect 17590 23015 17592 23024
rect 17644 23015 17646 23024
rect 17684 23044 17736 23050
rect 17592 22986 17644 22992
rect 17684 22986 17736 22992
rect 17512 22732 17724 22760
rect 17498 22672 17554 22681
rect 17696 22642 17724 22732
rect 17498 22607 17500 22616
rect 17552 22607 17554 22616
rect 17684 22636 17736 22642
rect 17500 22578 17552 22584
rect 17684 22578 17736 22584
rect 17406 21720 17462 21729
rect 17406 21655 17462 21664
rect 17420 21554 17448 21655
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17408 21344 17460 21350
rect 17408 21286 17460 21292
rect 17052 18686 17356 18714
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 16960 16266 16988 16662
rect 17052 16425 17080 18686
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 17144 16833 17172 18566
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17236 18290 17264 18362
rect 17328 18329 17356 18362
rect 17314 18320 17370 18329
rect 17224 18284 17276 18290
rect 17314 18255 17370 18264
rect 17224 18226 17276 18232
rect 17236 17746 17264 18226
rect 17316 17876 17368 17882
rect 17316 17818 17368 17824
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 17130 16824 17186 16833
rect 17130 16759 17186 16768
rect 17328 16658 17356 17818
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17132 16516 17184 16522
rect 17132 16458 17184 16464
rect 17038 16416 17094 16425
rect 17038 16351 17094 16360
rect 16960 16238 17080 16266
rect 16948 16176 17000 16182
rect 16948 16118 17000 16124
rect 16960 15473 16988 16118
rect 17052 15910 17080 16238
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 16946 15464 17002 15473
rect 16946 15399 17002 15408
rect 17144 14958 17172 16458
rect 17224 15428 17276 15434
rect 17224 15370 17276 15376
rect 17132 14952 17184 14958
rect 17132 14894 17184 14900
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 16960 14414 16988 14758
rect 17052 14482 17080 14758
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 16948 14408 17000 14414
rect 17144 14362 17172 14758
rect 16948 14350 17000 14356
rect 17052 14334 17172 14362
rect 17052 13025 17080 14334
rect 17236 14113 17264 15370
rect 17222 14104 17278 14113
rect 17222 14039 17278 14048
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17038 13016 17094 13025
rect 17038 12951 17094 12960
rect 16868 12872 17080 12900
rect 16764 12854 16816 12860
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16120 11824 16172 11830
rect 16120 11766 16172 11772
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 16316 11393 16344 11630
rect 16302 11384 16358 11393
rect 16408 11354 16436 11698
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16578 11520 16634 11529
rect 16500 11393 16528 11494
rect 16578 11455 16634 11464
rect 16486 11384 16542 11393
rect 16302 11319 16358 11328
rect 16396 11348 16448 11354
rect 16316 11234 16344 11319
rect 16486 11319 16542 11328
rect 16396 11290 16448 11296
rect 16486 11248 16542 11257
rect 16316 11206 16436 11234
rect 16040 10662 16160 10690
rect 15842 10568 15898 10577
rect 15842 10503 15898 10512
rect 16026 10568 16082 10577
rect 16132 10538 16160 10662
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16026 10503 16082 10512
rect 16120 10532 16172 10538
rect 16040 10266 16068 10503
rect 16120 10474 16172 10480
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15856 9722 15884 9998
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 15948 9178 15976 10202
rect 16040 9994 16068 10202
rect 16028 9988 16080 9994
rect 16028 9930 16080 9936
rect 16040 9674 16068 9930
rect 16040 9646 16160 9674
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15948 8956 15976 9114
rect 16040 9081 16068 9522
rect 16132 9382 16160 9646
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16026 9072 16082 9081
rect 16026 9007 16082 9016
rect 15948 8928 16068 8956
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15658 7984 15714 7993
rect 15764 7954 15792 8434
rect 15856 8090 15884 8434
rect 16040 8294 16068 8928
rect 15936 8288 15988 8294
rect 15934 8256 15936 8265
rect 16028 8288 16080 8294
rect 15988 8256 15990 8265
rect 16028 8230 16080 8236
rect 15934 8191 15990 8200
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15658 7919 15714 7928
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15476 7472 15528 7478
rect 15476 7414 15528 7420
rect 15396 7296 15516 7324
rect 15488 7002 15516 7296
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 15488 6254 15516 6666
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15672 6322 15700 6598
rect 15764 6458 15792 7890
rect 16224 7886 16252 10610
rect 16304 10464 16356 10470
rect 16302 10432 16304 10441
rect 16356 10432 16358 10441
rect 16302 10367 16358 10376
rect 16408 10282 16436 11206
rect 16486 11183 16542 11192
rect 16500 11150 16528 11183
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16316 10254 16436 10282
rect 16316 9602 16344 10254
rect 16592 10062 16620 11455
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16684 10010 16712 12378
rect 16776 12306 16804 12854
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16776 10849 16804 11494
rect 16762 10840 16818 10849
rect 16762 10775 16818 10784
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16776 10470 16804 10610
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16776 10169 16804 10406
rect 16762 10160 16818 10169
rect 16762 10095 16818 10104
rect 16408 9897 16436 9998
rect 16488 9988 16540 9994
rect 16684 9982 16804 10010
rect 16488 9930 16540 9936
rect 16394 9888 16450 9897
rect 16394 9823 16450 9832
rect 16500 9722 16528 9930
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 16316 9574 16528 9602
rect 16592 9586 16620 9862
rect 16684 9722 16712 9862
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16670 9616 16726 9625
rect 16302 9480 16358 9489
rect 16302 9415 16358 9424
rect 16316 9081 16344 9415
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16302 9072 16358 9081
rect 16302 9007 16358 9016
rect 16408 8838 16436 9114
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15856 6730 15884 7686
rect 16224 7546 16252 7822
rect 16304 7812 16356 7818
rect 16304 7754 16356 7760
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16224 6798 16252 7482
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 15844 6724 15896 6730
rect 15844 6666 15896 6672
rect 16028 6724 16080 6730
rect 16028 6666 16080 6672
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15488 6118 15516 6190
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15764 4690 15792 5102
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15856 4049 15884 6666
rect 16040 5166 16068 6666
rect 16120 5296 16172 5302
rect 16120 5238 16172 5244
rect 16028 5160 16080 5166
rect 16028 5102 16080 5108
rect 16132 4826 16160 5238
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16224 4622 16252 4966
rect 16316 4826 16344 7754
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16408 7342 16436 7686
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 15842 4040 15898 4049
rect 15842 3975 15898 3984
rect 15106 3632 15162 3641
rect 16500 3602 16528 9574
rect 16580 9580 16632 9586
rect 16670 9551 16726 9560
rect 16580 9522 16632 9528
rect 16684 9518 16712 9551
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16592 8430 16620 9318
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16684 8498 16712 8910
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16684 7585 16712 8026
rect 16670 7576 16726 7585
rect 16670 7511 16726 7520
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16592 6866 16620 7346
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16684 5574 16712 5850
rect 16776 5574 16804 9982
rect 16868 9178 16896 11494
rect 16960 11268 16988 12718
rect 17052 11762 17080 12872
rect 17236 12628 17264 13262
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17328 12753 17356 12786
rect 17314 12744 17370 12753
rect 17314 12679 17370 12688
rect 17316 12640 17368 12646
rect 17236 12600 17316 12628
rect 17316 12582 17368 12588
rect 17224 12368 17276 12374
rect 17224 12310 17276 12316
rect 17132 12164 17184 12170
rect 17132 12106 17184 12112
rect 17144 11898 17172 12106
rect 17236 12073 17264 12310
rect 17222 12064 17278 12073
rect 17222 11999 17278 12008
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17224 11688 17276 11694
rect 17130 11656 17186 11665
rect 17224 11630 17276 11636
rect 17130 11591 17186 11600
rect 16960 11240 17080 11268
rect 16948 11144 17000 11150
rect 16946 11112 16948 11121
rect 17000 11112 17002 11121
rect 16946 11047 17002 11056
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16868 8838 16896 8910
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16868 7313 16896 8774
rect 16960 8634 16988 10202
rect 17052 9178 17080 11240
rect 17144 9994 17172 11591
rect 17132 9988 17184 9994
rect 17132 9930 17184 9936
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 16960 8022 16988 8570
rect 16948 8016 17000 8022
rect 16948 7958 17000 7964
rect 17052 7886 17080 9114
rect 17130 8936 17186 8945
rect 17236 8906 17264 11630
rect 17420 11626 17448 21286
rect 17512 18902 17540 22578
rect 17788 22438 17816 23258
rect 17880 22817 17908 23446
rect 17958 23423 18014 23432
rect 17866 22808 17922 22817
rect 17866 22743 17922 22752
rect 17776 22432 17828 22438
rect 17776 22374 17828 22380
rect 17788 22094 17816 22374
rect 17696 22066 17816 22094
rect 17696 22030 17724 22066
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17592 21956 17644 21962
rect 17592 21898 17644 21904
rect 17868 21956 17920 21962
rect 17868 21898 17920 21904
rect 17604 19514 17632 21898
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17776 21888 17828 21894
rect 17776 21830 17828 21836
rect 17696 21457 17724 21830
rect 17788 21622 17816 21830
rect 17776 21616 17828 21622
rect 17776 21558 17828 21564
rect 17776 21480 17828 21486
rect 17682 21448 17738 21457
rect 17776 21422 17828 21428
rect 17682 21383 17738 21392
rect 17788 21350 17816 21422
rect 17684 21344 17736 21350
rect 17682 21312 17684 21321
rect 17776 21344 17828 21350
rect 17736 21312 17738 21321
rect 17776 21286 17828 21292
rect 17682 21247 17738 21256
rect 17682 21040 17738 21049
rect 17682 20975 17738 20984
rect 17592 19508 17644 19514
rect 17696 19496 17724 20975
rect 17880 20777 17908 21898
rect 17866 20768 17922 20777
rect 17866 20703 17922 20712
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17788 19718 17816 20198
rect 17776 19712 17828 19718
rect 17776 19654 17828 19660
rect 17696 19468 17816 19496
rect 17592 19450 17644 19456
rect 17500 18896 17552 18902
rect 17500 18838 17552 18844
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17512 18630 17540 18702
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17500 18148 17552 18154
rect 17500 18090 17552 18096
rect 17512 16590 17540 18090
rect 17604 17202 17632 19450
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17592 17196 17644 17202
rect 17592 17138 17644 17144
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17512 11898 17540 16390
rect 17696 16114 17724 19314
rect 17788 19242 17816 19468
rect 17776 19236 17828 19242
rect 17776 19178 17828 19184
rect 17774 19136 17830 19145
rect 17774 19071 17830 19080
rect 17788 18970 17816 19071
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17788 18222 17816 18702
rect 17776 18216 17828 18222
rect 17776 18158 17828 18164
rect 17880 17338 17908 20703
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 17788 16998 17816 17274
rect 17972 17270 18000 23423
rect 18064 23322 18092 23530
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 18156 22778 18184 23802
rect 18236 22976 18288 22982
rect 18236 22918 18288 22924
rect 18144 22772 18196 22778
rect 18144 22714 18196 22720
rect 18248 22681 18276 22918
rect 18234 22672 18290 22681
rect 18234 22607 18290 22616
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 18236 21548 18288 21554
rect 18236 21490 18288 21496
rect 18064 19378 18092 21490
rect 18144 21344 18196 21350
rect 18144 21286 18196 21292
rect 18156 20806 18184 21286
rect 18248 20913 18276 21490
rect 18234 20904 18290 20913
rect 18234 20839 18290 20848
rect 18144 20800 18196 20806
rect 18144 20742 18196 20748
rect 18340 20398 18368 26182
rect 18432 25906 18460 26522
rect 18524 26246 18552 26687
rect 18616 26364 18644 26880
rect 18708 26518 18736 27406
rect 18792 27282 18820 27492
rect 18892 27316 18920 27492
rect 19168 27452 19196 27503
rect 19352 27526 19472 27554
rect 19248 27474 19300 27480
rect 19076 27424 19196 27452
rect 18892 27288 19012 27316
rect 18792 27254 18828 27282
rect 18800 26976 18828 27254
rect 18800 26948 18920 26976
rect 18788 26852 18840 26858
rect 18788 26794 18840 26800
rect 18800 26761 18828 26794
rect 18786 26752 18842 26761
rect 18786 26687 18842 26696
rect 18696 26512 18748 26518
rect 18696 26454 18748 26460
rect 18800 26382 18828 26687
rect 18892 26382 18920 26948
rect 18696 26376 18748 26382
rect 18616 26336 18696 26364
rect 18696 26318 18748 26324
rect 18788 26376 18840 26382
rect 18788 26318 18840 26324
rect 18880 26376 18932 26382
rect 18880 26318 18932 26324
rect 18512 26240 18564 26246
rect 18512 26182 18564 26188
rect 18420 25900 18472 25906
rect 18420 25842 18472 25848
rect 18420 25356 18472 25362
rect 18420 25298 18472 25304
rect 18432 25158 18460 25298
rect 18524 25294 18552 26182
rect 18696 25832 18748 25838
rect 18696 25774 18748 25780
rect 18512 25288 18564 25294
rect 18512 25230 18564 25236
rect 18420 25152 18472 25158
rect 18420 25094 18472 25100
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18432 23225 18460 24754
rect 18708 23662 18736 25774
rect 18880 24064 18932 24070
rect 18880 24006 18932 24012
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18696 23656 18748 23662
rect 18696 23598 18748 23604
rect 18512 23520 18564 23526
rect 18512 23462 18564 23468
rect 18418 23216 18474 23225
rect 18524 23186 18552 23462
rect 18418 23151 18474 23160
rect 18512 23180 18564 23186
rect 18512 23122 18564 23128
rect 18512 21548 18564 21554
rect 18512 21490 18564 21496
rect 18420 21480 18472 21486
rect 18420 21422 18472 21428
rect 18432 21350 18460 21422
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18432 21010 18460 21286
rect 18420 21004 18472 21010
rect 18420 20946 18472 20952
rect 18524 20942 18552 21490
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18328 20392 18380 20398
rect 18328 20334 18380 20340
rect 18326 20088 18382 20097
rect 18326 20023 18382 20032
rect 18142 19952 18198 19961
rect 18142 19887 18198 19896
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 18064 18086 18092 18566
rect 18156 18329 18184 19887
rect 18142 18320 18198 18329
rect 18142 18255 18198 18264
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 18142 18048 18198 18057
rect 18064 17882 18092 18022
rect 18142 17983 18198 17992
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 18064 17270 18092 17478
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 17868 17128 17920 17134
rect 18064 17116 18092 17206
rect 17868 17070 17920 17076
rect 17972 17088 18092 17116
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 17880 16794 17908 17070
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 17972 16590 18000 17088
rect 18156 17066 18184 17983
rect 18234 17368 18290 17377
rect 18234 17303 18290 17312
rect 18248 17134 18276 17303
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 18144 17060 18196 17066
rect 18144 17002 18196 17008
rect 18340 16946 18368 20023
rect 18524 19334 18552 20878
rect 18156 16918 18368 16946
rect 18432 19306 18552 19334
rect 17960 16584 18012 16590
rect 17960 16526 18012 16532
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 17590 15056 17646 15065
rect 17696 15026 17724 16050
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17788 15026 17816 15098
rect 17866 15056 17922 15065
rect 17590 14991 17646 15000
rect 17684 15020 17736 15026
rect 17604 14618 17632 14991
rect 17684 14962 17736 14968
rect 17776 15020 17828 15026
rect 17866 14991 17922 15000
rect 17776 14962 17828 14968
rect 17684 14884 17736 14890
rect 17684 14826 17736 14832
rect 17776 14884 17828 14890
rect 17776 14826 17828 14832
rect 17696 14657 17724 14826
rect 17682 14648 17738 14657
rect 17592 14612 17644 14618
rect 17682 14583 17738 14592
rect 17592 14554 17644 14560
rect 17788 14482 17816 14826
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17590 13424 17646 13433
rect 17590 13359 17646 13368
rect 17604 13258 17632 13359
rect 17592 13252 17644 13258
rect 17592 13194 17644 13200
rect 17592 12708 17644 12714
rect 17592 12650 17644 12656
rect 17604 12238 17632 12650
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17316 11620 17368 11626
rect 17316 11562 17368 11568
rect 17408 11620 17460 11626
rect 17408 11562 17460 11568
rect 17328 11286 17356 11562
rect 17316 11280 17368 11286
rect 17316 11222 17368 11228
rect 17512 11150 17540 11834
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17590 11112 17646 11121
rect 17316 11076 17368 11082
rect 17590 11047 17646 11056
rect 17316 11018 17368 11024
rect 17130 8871 17186 8880
rect 17224 8900 17276 8906
rect 17144 8786 17172 8871
rect 17224 8842 17276 8848
rect 17144 8758 17264 8786
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17144 8090 17172 8434
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 16854 7304 16910 7313
rect 16854 7239 16910 7248
rect 17144 6322 17172 7890
rect 17236 7886 17264 8758
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17222 7304 17278 7313
rect 17222 7239 17278 7248
rect 17236 6633 17264 7239
rect 17222 6624 17278 6633
rect 17222 6559 17278 6568
rect 17328 6322 17356 11018
rect 17498 10840 17554 10849
rect 17498 10775 17554 10784
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17420 10452 17448 10610
rect 17512 10554 17540 10775
rect 17604 10674 17632 11047
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 17512 10526 17632 10554
rect 17500 10464 17552 10470
rect 17420 10424 17500 10452
rect 17500 10406 17552 10412
rect 17512 10266 17540 10406
rect 17408 10260 17460 10266
rect 17408 10202 17460 10208
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17420 10169 17448 10202
rect 17406 10160 17462 10169
rect 17406 10095 17462 10104
rect 17604 8945 17632 10526
rect 17590 8936 17646 8945
rect 17590 8871 17646 8880
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17236 5778 17264 6190
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 17038 5672 17094 5681
rect 17144 5658 17172 5714
rect 17144 5630 17264 5658
rect 17038 5607 17040 5616
rect 17092 5607 17094 5616
rect 17040 5578 17092 5584
rect 17236 5574 17264 5630
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 15106 3567 15162 3576
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 13542 3360 13598 3369
rect 13542 3295 13598 3304
rect 16592 3194 16620 4082
rect 16776 3670 16804 4082
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 17420 3233 17448 8570
rect 17696 8498 17724 14214
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17788 12714 17816 13466
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17774 12472 17830 12481
rect 17774 12407 17830 12416
rect 17880 12434 17908 14991
rect 17972 13977 18000 15506
rect 17958 13968 18014 13977
rect 17958 13903 18014 13912
rect 17958 13696 18014 13705
rect 17958 13631 18014 13640
rect 17972 12782 18000 13631
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 17788 10470 17816 12407
rect 17880 12406 18000 12434
rect 17866 11928 17922 11937
rect 17972 11898 18000 12406
rect 17866 11863 17922 11872
rect 17960 11892 18012 11898
rect 17880 11830 17908 11863
rect 17960 11834 18012 11840
rect 17868 11824 17920 11830
rect 17868 11766 17920 11772
rect 17972 11694 18000 11834
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17880 9586 17908 11630
rect 18064 10538 18092 16526
rect 18156 15910 18184 16918
rect 18432 16810 18460 19306
rect 18616 18442 18644 23598
rect 18892 23594 18920 24006
rect 18984 23730 19012 27288
rect 19076 23730 19104 27424
rect 19444 27402 19472 27526
rect 19524 27532 19576 27538
rect 19720 27526 19840 27554
rect 19576 27492 19656 27520
rect 19524 27474 19576 27480
rect 19628 27441 19656 27492
rect 19614 27432 19670 27441
rect 19432 27396 19484 27402
rect 19614 27367 19670 27376
rect 19432 27338 19484 27344
rect 19248 27328 19300 27334
rect 19248 27270 19300 27276
rect 19154 27024 19210 27033
rect 19260 26994 19288 27270
rect 19154 26959 19210 26968
rect 19248 26988 19300 26994
rect 19168 26790 19196 26959
rect 19248 26930 19300 26936
rect 19248 26852 19300 26858
rect 19248 26794 19300 26800
rect 19156 26784 19208 26790
rect 19156 26726 19208 26732
rect 19154 26344 19210 26353
rect 19154 26279 19210 26288
rect 19168 25537 19196 26279
rect 19154 25528 19210 25537
rect 19154 25463 19210 25472
rect 19156 25356 19208 25362
rect 19156 25298 19208 25304
rect 19168 24818 19196 25298
rect 19156 24812 19208 24818
rect 19156 24754 19208 24760
rect 19260 24721 19288 26794
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 19352 25702 19380 25842
rect 19340 25696 19392 25702
rect 19340 25638 19392 25644
rect 19352 25537 19380 25638
rect 19338 25528 19394 25537
rect 19338 25463 19394 25472
rect 19444 25294 19472 27338
rect 19616 27328 19668 27334
rect 19708 27328 19760 27334
rect 19616 27270 19668 27276
rect 19706 27296 19708 27305
rect 19760 27296 19762 27305
rect 19524 27056 19576 27062
rect 19524 26998 19576 27004
rect 19628 27000 19656 27270
rect 19706 27231 19762 27240
rect 19536 26908 19564 26998
rect 19616 26994 19668 27000
rect 19812 26976 19840 27526
rect 19982 27503 20038 27512
rect 19996 27470 20024 27503
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 19984 27328 20036 27334
rect 19890 27296 19946 27305
rect 19984 27270 20036 27276
rect 19890 27231 19946 27240
rect 19616 26936 19668 26942
rect 19720 26948 19840 26976
rect 19536 26880 19656 26908
rect 19628 26790 19656 26880
rect 19524 26784 19576 26790
rect 19524 26726 19576 26732
rect 19616 26784 19668 26790
rect 19616 26726 19668 26732
rect 19536 26586 19564 26726
rect 19524 26580 19576 26586
rect 19524 26522 19576 26528
rect 19522 26072 19578 26081
rect 19522 26007 19578 26016
rect 19536 25770 19564 26007
rect 19614 25936 19670 25945
rect 19614 25871 19616 25880
rect 19668 25871 19670 25880
rect 19616 25842 19668 25848
rect 19524 25764 19576 25770
rect 19524 25706 19576 25712
rect 19720 25498 19748 26948
rect 19904 26926 19932 27231
rect 19996 26994 20024 27270
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 19892 26920 19944 26926
rect 19892 26862 19944 26868
rect 19800 26784 19852 26790
rect 19800 26726 19852 26732
rect 19892 26784 19944 26790
rect 19892 26726 19944 26732
rect 19812 26330 19840 26726
rect 19904 26450 19932 26726
rect 19892 26444 19944 26450
rect 19892 26386 19944 26392
rect 19984 26444 20036 26450
rect 19984 26386 20036 26392
rect 19996 26330 20024 26386
rect 19812 26302 20024 26330
rect 19800 26036 19852 26042
rect 19800 25978 19852 25984
rect 19708 25492 19760 25498
rect 19708 25434 19760 25440
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19708 25288 19760 25294
rect 19708 25230 19760 25236
rect 19720 24993 19748 25230
rect 19706 24984 19762 24993
rect 19706 24919 19762 24928
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19616 24812 19668 24818
rect 19616 24754 19668 24760
rect 19246 24712 19302 24721
rect 19246 24647 19302 24656
rect 19248 24608 19300 24614
rect 19248 24550 19300 24556
rect 18972 23724 19024 23730
rect 18972 23666 19024 23672
rect 19064 23724 19116 23730
rect 19064 23666 19116 23672
rect 18788 23588 18840 23594
rect 18788 23530 18840 23536
rect 18880 23588 18932 23594
rect 18880 23530 18932 23536
rect 18694 23488 18750 23497
rect 18694 23423 18750 23432
rect 18708 22642 18736 23423
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18800 22506 18828 23530
rect 18984 23225 19012 23666
rect 18970 23216 19026 23225
rect 18970 23151 19026 23160
rect 19064 23112 19116 23118
rect 19064 23054 19116 23060
rect 19156 23112 19208 23118
rect 19156 23054 19208 23060
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18972 22976 19024 22982
rect 18972 22918 19024 22924
rect 18892 22681 18920 22918
rect 18878 22672 18934 22681
rect 18878 22607 18934 22616
rect 18788 22500 18840 22506
rect 18788 22442 18840 22448
rect 18800 22098 18828 22442
rect 18878 22400 18934 22409
rect 18878 22335 18934 22344
rect 18788 22092 18840 22098
rect 18788 22034 18840 22040
rect 18788 21616 18840 21622
rect 18788 21558 18840 21564
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18248 16782 18460 16810
rect 18524 18414 18644 18442
rect 18248 15994 18276 16782
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18432 16522 18460 16594
rect 18420 16516 18472 16522
rect 18420 16458 18472 16464
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 18418 16416 18474 16425
rect 18340 16114 18368 16390
rect 18418 16351 18474 16360
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18248 15966 18368 15994
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 18156 12481 18184 15642
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 18248 14346 18276 14962
rect 18236 14340 18288 14346
rect 18236 14282 18288 14288
rect 18340 14226 18368 15966
rect 18432 15026 18460 16351
rect 18524 15706 18552 18414
rect 18604 18352 18656 18358
rect 18604 18294 18656 18300
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18248 14198 18368 14226
rect 18248 13802 18276 14198
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 18328 13728 18380 13734
rect 18328 13670 18380 13676
rect 18142 12472 18198 12481
rect 18142 12407 18198 12416
rect 18340 11830 18368 13670
rect 18328 11824 18380 11830
rect 18328 11766 18380 11772
rect 18432 10742 18460 14758
rect 18524 14618 18552 14758
rect 18616 14657 18644 18294
rect 18708 18086 18736 18906
rect 18800 18290 18828 21558
rect 18892 19242 18920 22335
rect 18984 22234 19012 22918
rect 18972 22228 19024 22234
rect 18972 22170 19024 22176
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18880 19236 18932 19242
rect 18880 19178 18932 19184
rect 18984 18290 19012 19450
rect 18788 18284 18840 18290
rect 18788 18226 18840 18232
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18694 16688 18750 16697
rect 18694 16623 18750 16632
rect 18708 16590 18736 16623
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18800 16046 18828 16730
rect 18970 16552 19026 16561
rect 18970 16487 19026 16496
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18602 14648 18658 14657
rect 18512 14612 18564 14618
rect 18602 14583 18658 14592
rect 18512 14554 18564 14560
rect 18708 14498 18736 15846
rect 18800 15502 18828 15982
rect 18892 15638 18920 16390
rect 18880 15632 18932 15638
rect 18880 15574 18932 15580
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 18878 15192 18934 15201
rect 18878 15127 18934 15136
rect 18892 15026 18920 15127
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18786 14920 18842 14929
rect 18786 14855 18788 14864
rect 18840 14855 18842 14864
rect 18880 14884 18932 14890
rect 18788 14826 18840 14832
rect 18880 14826 18932 14832
rect 18786 14648 18842 14657
rect 18892 14618 18920 14826
rect 18786 14583 18842 14592
rect 18880 14612 18932 14618
rect 18524 14470 18736 14498
rect 18524 12850 18552 14470
rect 18800 14414 18828 14583
rect 18880 14554 18932 14560
rect 18878 14512 18934 14521
rect 18878 14447 18934 14456
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18786 13968 18842 13977
rect 18696 13932 18748 13938
rect 18786 13903 18788 13912
rect 18696 13874 18748 13880
rect 18840 13903 18842 13912
rect 18788 13874 18840 13880
rect 18708 13530 18736 13874
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 18604 13456 18656 13462
rect 18604 13398 18656 13404
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18616 12434 18644 13398
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18708 12850 18736 13126
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 18788 12776 18840 12782
rect 18786 12744 18788 12753
rect 18840 12744 18842 12753
rect 18786 12679 18842 12688
rect 18892 12646 18920 14447
rect 18984 13938 19012 16487
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 18984 13326 19012 13874
rect 18972 13320 19024 13326
rect 18972 13262 19024 13268
rect 18970 13016 19026 13025
rect 18970 12951 19026 12960
rect 18984 12753 19012 12951
rect 18970 12744 19026 12753
rect 18970 12679 19026 12688
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18616 12406 18736 12434
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18524 11762 18552 12038
rect 18512 11756 18564 11762
rect 18708 11744 18736 12406
rect 18800 12374 18828 12582
rect 18788 12368 18840 12374
rect 18788 12310 18840 12316
rect 19076 12102 19104 23054
rect 19168 22778 19196 23054
rect 19156 22772 19208 22778
rect 19156 22714 19208 22720
rect 19168 22137 19196 22714
rect 19154 22128 19210 22137
rect 19154 22063 19210 22072
rect 19156 22024 19208 22030
rect 19156 21966 19208 21972
rect 19168 21554 19196 21966
rect 19260 21865 19288 24550
rect 19352 24410 19380 24754
rect 19430 24712 19486 24721
rect 19430 24647 19486 24656
rect 19444 24614 19472 24647
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19340 24404 19392 24410
rect 19340 24346 19392 24352
rect 19628 24342 19656 24754
rect 19812 24721 19840 25978
rect 19890 25936 19946 25945
rect 19890 25871 19892 25880
rect 19944 25871 19946 25880
rect 19892 25842 19944 25848
rect 19984 25696 20036 25702
rect 19984 25638 20036 25644
rect 19892 25424 19944 25430
rect 19892 25366 19944 25372
rect 19904 24954 19932 25366
rect 19996 25294 20024 25638
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 19892 24948 19944 24954
rect 19892 24890 19944 24896
rect 19904 24818 19932 24890
rect 19892 24812 19944 24818
rect 19892 24754 19944 24760
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 19798 24712 19854 24721
rect 19798 24647 19854 24656
rect 19892 24608 19944 24614
rect 19996 24596 20024 24754
rect 19944 24568 20024 24596
rect 19892 24550 19944 24556
rect 19616 24336 19668 24342
rect 19616 24278 19668 24284
rect 19524 24064 19576 24070
rect 19524 24006 19576 24012
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19352 22953 19380 23462
rect 19536 23186 19564 24006
rect 19524 23180 19576 23186
rect 19524 23122 19576 23128
rect 19430 23080 19486 23089
rect 19628 23066 19656 24278
rect 19708 23316 19760 23322
rect 19708 23258 19760 23264
rect 19430 23015 19486 23024
rect 19536 23038 19656 23066
rect 19338 22944 19394 22953
rect 19338 22879 19394 22888
rect 19444 22778 19472 23015
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19536 22642 19564 23038
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19524 22636 19576 22642
rect 19524 22578 19576 22584
rect 19352 22409 19380 22578
rect 19338 22400 19394 22409
rect 19338 22335 19394 22344
rect 19444 22273 19472 22578
rect 19628 22574 19656 22714
rect 19616 22568 19668 22574
rect 19616 22510 19668 22516
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19430 22264 19486 22273
rect 19430 22199 19486 22208
rect 19338 22128 19394 22137
rect 19338 22063 19394 22072
rect 19352 21944 19380 22063
rect 19352 21916 19472 21944
rect 19246 21856 19302 21865
rect 19246 21791 19302 21800
rect 19338 21720 19394 21729
rect 19338 21655 19340 21664
rect 19392 21655 19394 21664
rect 19340 21626 19392 21632
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19340 21548 19392 21554
rect 19340 21490 19392 21496
rect 19260 21049 19288 21490
rect 19246 21040 19302 21049
rect 19246 20975 19302 20984
rect 19352 20913 19380 21490
rect 19444 21486 19472 21916
rect 19536 21554 19564 22374
rect 19614 22128 19670 22137
rect 19614 22063 19616 22072
rect 19668 22063 19670 22072
rect 19616 22034 19668 22040
rect 19720 21672 19748 23258
rect 19904 22794 19932 24550
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 19996 22982 20024 23462
rect 19984 22976 20036 22982
rect 19984 22918 20036 22924
rect 19904 22766 20024 22794
rect 19800 22636 19852 22642
rect 19800 22578 19852 22584
rect 19812 21690 19840 22578
rect 19996 22574 20024 22766
rect 19892 22568 19944 22574
rect 19892 22510 19944 22516
rect 19984 22568 20036 22574
rect 19984 22510 20036 22516
rect 19904 22030 19932 22510
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 19628 21644 19748 21672
rect 19800 21684 19852 21690
rect 19524 21548 19576 21554
rect 19524 21490 19576 21496
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19536 21049 19564 21286
rect 19522 21040 19578 21049
rect 19522 20975 19578 20984
rect 19338 20904 19394 20913
rect 19338 20839 19394 20848
rect 19522 20904 19578 20913
rect 19522 20839 19578 20848
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 19156 20256 19208 20262
rect 19156 20198 19208 20204
rect 19168 16182 19196 20198
rect 19352 18698 19380 20402
rect 19444 19922 19472 20742
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19430 19680 19486 19689
rect 19430 19615 19486 19624
rect 19248 18692 19300 18698
rect 19248 18634 19300 18640
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19260 18057 19288 18634
rect 19246 18048 19302 18057
rect 19246 17983 19302 17992
rect 19352 17898 19380 18634
rect 19444 18057 19472 19615
rect 19536 18290 19564 20839
rect 19628 20058 19656 21644
rect 19800 21626 19852 21632
rect 19890 21584 19946 21593
rect 19890 21519 19892 21528
rect 19944 21519 19946 21528
rect 19892 21490 19944 21496
rect 19996 21457 20024 22102
rect 19706 21448 19762 21457
rect 19982 21448 20038 21457
rect 19706 21383 19762 21392
rect 19892 21412 19944 21418
rect 19720 21049 19748 21383
rect 19982 21383 20038 21392
rect 19892 21354 19944 21360
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 19812 21146 19840 21286
rect 19800 21140 19852 21146
rect 19800 21082 19852 21088
rect 19706 21040 19762 21049
rect 19904 20992 19932 21354
rect 19706 20975 19762 20984
rect 19812 20964 19932 20992
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 19720 20777 19748 20878
rect 19706 20768 19762 20777
rect 19706 20703 19762 20712
rect 19812 20398 19840 20964
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 19800 20392 19852 20398
rect 19800 20334 19852 20340
rect 19706 20088 19762 20097
rect 19616 20052 19668 20058
rect 19706 20023 19762 20032
rect 19616 19994 19668 20000
rect 19616 19236 19668 19242
rect 19616 19178 19668 19184
rect 19524 18284 19576 18290
rect 19524 18226 19576 18232
rect 19524 18080 19576 18086
rect 19430 18048 19486 18057
rect 19524 18022 19576 18028
rect 19430 17983 19486 17992
rect 19260 17870 19380 17898
rect 19156 16176 19208 16182
rect 19156 16118 19208 16124
rect 19156 14884 19208 14890
rect 19156 14826 19208 14832
rect 19168 14657 19196 14826
rect 19154 14648 19210 14657
rect 19154 14583 19210 14592
rect 19260 14362 19288 17870
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19338 16824 19394 16833
rect 19338 16759 19394 16768
rect 19352 16250 19380 16759
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19168 14334 19288 14362
rect 19352 14346 19380 15370
rect 19444 14396 19472 17614
rect 19536 15201 19564 18022
rect 19628 17202 19656 19178
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19720 16266 19748 20023
rect 19628 16238 19748 16266
rect 19628 15434 19656 16238
rect 19708 16176 19760 16182
rect 19706 16144 19708 16153
rect 19760 16144 19762 16153
rect 19706 16079 19762 16088
rect 19720 16046 19748 16079
rect 19708 16040 19760 16046
rect 19708 15982 19760 15988
rect 19706 15736 19762 15745
rect 19706 15671 19762 15680
rect 19616 15428 19668 15434
rect 19616 15370 19668 15376
rect 19720 15366 19748 15671
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19522 15192 19578 15201
rect 19522 15127 19578 15136
rect 19614 15056 19670 15065
rect 19614 14991 19616 15000
rect 19668 14991 19670 15000
rect 19616 14962 19668 14968
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19536 14521 19564 14554
rect 19522 14512 19578 14521
rect 19628 14498 19656 14758
rect 19812 14532 19840 20334
rect 19892 20324 19944 20330
rect 19892 20266 19944 20272
rect 19904 20097 19932 20266
rect 19890 20088 19946 20097
rect 19890 20023 19946 20032
rect 19892 19916 19944 19922
rect 19892 19858 19944 19864
rect 19904 19718 19932 19858
rect 19996 19854 20024 20402
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19892 19168 19944 19174
rect 19892 19110 19944 19116
rect 19904 18766 19932 19110
rect 19892 18760 19944 18766
rect 19892 18702 19944 18708
rect 19892 18352 19944 18358
rect 19892 18294 19944 18300
rect 19904 17678 19932 18294
rect 19996 18086 20024 19314
rect 20088 19242 20116 27832
rect 20180 27441 20208 28358
rect 20272 28150 20300 28580
rect 20364 28393 20392 28630
rect 20536 28552 20588 28558
rect 20536 28494 20588 28500
rect 20548 28393 20576 28494
rect 20350 28384 20406 28393
rect 20350 28319 20406 28328
rect 20534 28384 20590 28393
rect 20534 28319 20590 28328
rect 20260 28144 20312 28150
rect 20260 28086 20312 28092
rect 20442 28112 20498 28121
rect 20272 27674 20300 28086
rect 20442 28047 20498 28056
rect 20536 28076 20588 28082
rect 20352 28008 20404 28014
rect 20352 27950 20404 27956
rect 20260 27668 20312 27674
rect 20260 27610 20312 27616
rect 20260 27532 20312 27538
rect 20260 27474 20312 27480
rect 20166 27432 20222 27441
rect 20166 27367 20222 27376
rect 20166 26888 20222 26897
rect 20166 26823 20222 26832
rect 20180 26790 20208 26823
rect 20168 26784 20220 26790
rect 20168 26726 20220 26732
rect 20168 26512 20220 26518
rect 20272 26500 20300 27474
rect 20220 26472 20300 26500
rect 20168 26454 20220 26460
rect 20258 26208 20314 26217
rect 20258 26143 20314 26152
rect 20272 25906 20300 26143
rect 20260 25900 20312 25906
rect 20260 25842 20312 25848
rect 20260 25696 20312 25702
rect 20260 25638 20312 25644
rect 20168 25492 20220 25498
rect 20168 25434 20220 25440
rect 20180 24954 20208 25434
rect 20272 25401 20300 25638
rect 20258 25392 20314 25401
rect 20258 25327 20314 25336
rect 20258 24984 20314 24993
rect 20168 24948 20220 24954
rect 20258 24919 20314 24928
rect 20168 24890 20220 24896
rect 20272 24886 20300 24919
rect 20260 24880 20312 24886
rect 20260 24822 20312 24828
rect 20168 24608 20220 24614
rect 20168 24550 20220 24556
rect 20180 24274 20208 24550
rect 20168 24268 20220 24274
rect 20168 24210 20220 24216
rect 20364 24154 20392 27950
rect 20456 27878 20484 28047
rect 20536 28018 20588 28024
rect 20444 27872 20496 27878
rect 20444 27814 20496 27820
rect 20456 27674 20484 27814
rect 20444 27668 20496 27674
rect 20444 27610 20496 27616
rect 20444 26988 20496 26994
rect 20444 26930 20496 26936
rect 20456 26382 20484 26930
rect 20444 26376 20496 26382
rect 20444 26318 20496 26324
rect 20442 26072 20498 26081
rect 20442 26007 20498 26016
rect 20456 25906 20484 26007
rect 20444 25900 20496 25906
rect 20444 25842 20496 25848
rect 20444 25696 20496 25702
rect 20444 25638 20496 25644
rect 20456 25498 20484 25638
rect 20444 25492 20496 25498
rect 20548 25480 20576 28018
rect 20640 26897 20668 29650
rect 20916 29646 20944 29990
rect 20904 29640 20956 29646
rect 20904 29582 20956 29588
rect 21272 29640 21324 29646
rect 21272 29582 21324 29588
rect 20720 27056 20772 27062
rect 20720 26998 20772 27004
rect 20626 26888 20682 26897
rect 20626 26823 20682 26832
rect 20732 25838 20760 26998
rect 20812 26920 20864 26926
rect 20812 26862 20864 26868
rect 20824 26042 20852 26862
rect 21178 26344 21234 26353
rect 21178 26279 21180 26288
rect 21232 26279 21234 26288
rect 21180 26250 21232 26256
rect 20812 26036 20864 26042
rect 20812 25978 20864 25984
rect 20996 25900 21048 25906
rect 20996 25842 21048 25848
rect 21180 25900 21232 25906
rect 21180 25842 21232 25848
rect 20720 25832 20772 25838
rect 20720 25774 20772 25780
rect 20812 25832 20864 25838
rect 21008 25809 21036 25842
rect 20812 25774 20864 25780
rect 20994 25800 21050 25809
rect 20824 25498 20852 25774
rect 20994 25735 21050 25744
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 20812 25492 20864 25498
rect 20548 25452 20668 25480
rect 20444 25434 20496 25440
rect 20534 25392 20590 25401
rect 20534 25327 20590 25336
rect 20548 25294 20576 25327
rect 20536 25288 20588 25294
rect 20536 25230 20588 25236
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 20548 24410 20576 24550
rect 20536 24404 20588 24410
rect 20536 24346 20588 24352
rect 20548 24177 20576 24346
rect 20180 24126 20392 24154
rect 20534 24168 20590 24177
rect 20180 22953 20208 24126
rect 20534 24103 20590 24112
rect 20352 23316 20404 23322
rect 20352 23258 20404 23264
rect 20260 23112 20312 23118
rect 20260 23054 20312 23060
rect 20166 22944 20222 22953
rect 20166 22879 20222 22888
rect 20272 22778 20300 23054
rect 20260 22772 20312 22778
rect 20260 22714 20312 22720
rect 20168 22636 20220 22642
rect 20168 22578 20220 22584
rect 20180 22234 20208 22578
rect 20260 22432 20312 22438
rect 20260 22374 20312 22380
rect 20168 22228 20220 22234
rect 20168 22170 20220 22176
rect 20166 22128 20222 22137
rect 20272 22098 20300 22374
rect 20166 22063 20168 22072
rect 20220 22063 20222 22072
rect 20260 22092 20312 22098
rect 20168 22034 20220 22040
rect 20260 22034 20312 22040
rect 20364 21842 20392 23258
rect 20640 22930 20668 25452
rect 20812 25434 20864 25440
rect 20720 25424 20772 25430
rect 20720 25366 20772 25372
rect 20732 24614 20760 25366
rect 20720 24608 20772 24614
rect 20720 24550 20772 24556
rect 20824 24410 20852 25434
rect 20812 24404 20864 24410
rect 20812 24346 20864 24352
rect 21008 24256 21036 25638
rect 21192 25430 21220 25842
rect 21088 25424 21140 25430
rect 21088 25366 21140 25372
rect 21180 25424 21232 25430
rect 21180 25366 21232 25372
rect 21100 24324 21128 25366
rect 21180 25288 21232 25294
rect 21180 25230 21232 25236
rect 21192 24562 21220 25230
rect 21284 24682 21312 29582
rect 22204 29510 22232 29990
rect 22468 29572 22520 29578
rect 22468 29514 22520 29520
rect 22100 29504 22152 29510
rect 22100 29446 22152 29452
rect 22192 29504 22244 29510
rect 22192 29446 22244 29452
rect 22376 29504 22428 29510
rect 22376 29446 22428 29452
rect 22112 29238 22140 29446
rect 22100 29232 22152 29238
rect 22100 29174 22152 29180
rect 22204 29170 22232 29446
rect 22388 29170 22416 29446
rect 22480 29306 22508 29514
rect 22468 29300 22520 29306
rect 22468 29242 22520 29248
rect 21916 29164 21968 29170
rect 21916 29106 21968 29112
rect 22192 29164 22244 29170
rect 22192 29106 22244 29112
rect 22376 29164 22428 29170
rect 22376 29106 22428 29112
rect 21928 29073 21956 29106
rect 21914 29064 21970 29073
rect 21914 28999 21970 29008
rect 22190 29064 22246 29073
rect 22190 28999 22246 29008
rect 21732 28620 21784 28626
rect 21732 28562 21784 28568
rect 21744 27946 21772 28562
rect 22100 28008 22152 28014
rect 21822 27976 21878 27985
rect 21732 27940 21784 27946
rect 22100 27950 22152 27956
rect 21822 27911 21824 27920
rect 21732 27882 21784 27888
rect 21876 27911 21878 27920
rect 21824 27882 21876 27888
rect 22112 27849 22140 27950
rect 22098 27840 22154 27849
rect 22098 27775 22154 27784
rect 22098 27704 22154 27713
rect 22098 27639 22154 27648
rect 22006 27432 22062 27441
rect 22006 27367 22062 27376
rect 22020 27334 22048 27367
rect 22008 27328 22060 27334
rect 22008 27270 22060 27276
rect 22112 27169 22140 27639
rect 22204 27577 22232 28999
rect 22558 28520 22614 28529
rect 22558 28455 22614 28464
rect 22376 28212 22428 28218
rect 22376 28154 22428 28160
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22190 27568 22246 27577
rect 22190 27503 22246 27512
rect 22296 27402 22324 28018
rect 22388 27538 22416 28154
rect 22572 28082 22600 28455
rect 22560 28076 22612 28082
rect 22560 28018 22612 28024
rect 22468 27668 22520 27674
rect 22468 27610 22520 27616
rect 22376 27532 22428 27538
rect 22376 27474 22428 27480
rect 22284 27396 22336 27402
rect 22284 27338 22336 27344
rect 22098 27160 22154 27169
rect 22296 27130 22324 27338
rect 22098 27095 22154 27104
rect 22284 27124 22336 27130
rect 22284 27066 22336 27072
rect 21822 27024 21878 27033
rect 21456 26988 21508 26994
rect 21822 26959 21878 26968
rect 21456 26930 21508 26936
rect 21364 26512 21416 26518
rect 21364 26454 21416 26460
rect 21376 25809 21404 26454
rect 21362 25800 21418 25809
rect 21362 25735 21418 25744
rect 21468 25702 21496 26930
rect 21732 26512 21784 26518
rect 21732 26454 21784 26460
rect 21744 26382 21772 26454
rect 21836 26382 21864 26959
rect 22008 26852 22060 26858
rect 22008 26794 22060 26800
rect 21916 26444 21968 26450
rect 21916 26386 21968 26392
rect 21732 26376 21784 26382
rect 21732 26318 21784 26324
rect 21824 26376 21876 26382
rect 21824 26318 21876 26324
rect 21548 26308 21600 26314
rect 21548 26250 21600 26256
rect 21560 25702 21588 26250
rect 21364 25696 21416 25702
rect 21364 25638 21416 25644
rect 21456 25696 21508 25702
rect 21456 25638 21508 25644
rect 21548 25696 21600 25702
rect 21548 25638 21600 25644
rect 21376 25498 21404 25638
rect 21364 25492 21416 25498
rect 21364 25434 21416 25440
rect 21468 25362 21496 25638
rect 21456 25356 21508 25362
rect 21456 25298 21508 25304
rect 21548 25288 21600 25294
rect 21548 25230 21600 25236
rect 21454 24984 21510 24993
rect 21454 24919 21510 24928
rect 21468 24842 21496 24919
rect 21456 24836 21508 24842
rect 21364 24812 21416 24818
rect 21560 24834 21588 25230
rect 21560 24806 21772 24834
rect 21456 24778 21508 24784
rect 21364 24754 21416 24760
rect 21272 24676 21324 24682
rect 21272 24618 21324 24624
rect 21376 24585 21404 24754
rect 21456 24744 21508 24750
rect 21456 24686 21508 24692
rect 21362 24576 21418 24585
rect 21192 24534 21312 24562
rect 21180 24336 21232 24342
rect 21100 24296 21180 24324
rect 21180 24278 21232 24284
rect 21008 24228 21128 24256
rect 20812 24200 20864 24206
rect 20812 24142 20864 24148
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 20732 23526 20760 23802
rect 20824 23769 20852 24142
rect 20996 24064 21048 24070
rect 20996 24006 21048 24012
rect 20810 23760 20866 23769
rect 20810 23695 20866 23704
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 20824 23338 20852 23695
rect 20902 23488 20958 23497
rect 20902 23423 20958 23432
rect 20732 23322 20852 23338
rect 20720 23316 20852 23322
rect 20772 23310 20852 23316
rect 20720 23258 20772 23264
rect 20916 23254 20944 23423
rect 20812 23248 20864 23254
rect 20812 23190 20864 23196
rect 20904 23248 20956 23254
rect 20904 23190 20956 23196
rect 20720 23044 20772 23050
rect 20720 22986 20772 22992
rect 20732 22953 20760 22986
rect 20180 21814 20392 21842
rect 20456 22902 20668 22930
rect 20718 22944 20774 22953
rect 20180 19446 20208 21814
rect 20258 21720 20314 21729
rect 20258 21655 20314 21664
rect 20352 21684 20404 21690
rect 20272 21622 20300 21655
rect 20352 21626 20404 21632
rect 20260 21616 20312 21622
rect 20260 21558 20312 21564
rect 20258 21448 20314 21457
rect 20258 21383 20314 21392
rect 20272 21350 20300 21383
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 20260 21140 20312 21146
rect 20260 21082 20312 21088
rect 20272 20466 20300 21082
rect 20364 20777 20392 21626
rect 20456 20806 20484 22902
rect 20718 22879 20774 22888
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20628 22704 20680 22710
rect 20628 22646 20680 22652
rect 20640 22094 20668 22646
rect 20732 22409 20760 22714
rect 20718 22400 20774 22409
rect 20718 22335 20774 22344
rect 20548 22066 20668 22094
rect 20720 22092 20772 22098
rect 20444 20800 20496 20806
rect 20350 20768 20406 20777
rect 20444 20742 20496 20748
rect 20350 20703 20406 20712
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20352 20256 20404 20262
rect 20456 20244 20484 20742
rect 20404 20216 20484 20244
rect 20352 20198 20404 20204
rect 20260 20052 20312 20058
rect 20260 19994 20312 20000
rect 20168 19440 20220 19446
rect 20168 19382 20220 19388
rect 20168 19304 20220 19310
rect 20166 19272 20168 19281
rect 20220 19272 20222 19281
rect 20076 19236 20128 19242
rect 20166 19207 20222 19216
rect 20076 19178 20128 19184
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 20076 18284 20128 18290
rect 20076 18226 20128 18232
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19892 17536 19944 17542
rect 19892 17478 19944 17484
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19904 15910 19932 17478
rect 19996 16697 20024 17478
rect 19982 16688 20038 16697
rect 19982 16623 20038 16632
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19996 16182 20024 16390
rect 19984 16176 20036 16182
rect 19984 16118 20036 16124
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 20088 15065 20116 18226
rect 20074 15056 20130 15065
rect 20074 14991 20130 15000
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 19984 14544 20036 14550
rect 19812 14504 19984 14532
rect 19628 14470 19748 14498
rect 19984 14486 20036 14492
rect 19522 14447 19578 14456
rect 19720 14414 19748 14470
rect 20088 14414 20116 14758
rect 19708 14408 19760 14414
rect 19444 14368 19564 14396
rect 19340 14340 19392 14346
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19076 11898 19104 12038
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 18708 11716 19012 11744
rect 18512 11698 18564 11704
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18616 11150 18644 11494
rect 18604 11144 18656 11150
rect 18510 11112 18566 11121
rect 18604 11086 18656 11092
rect 18708 11082 18736 11494
rect 18510 11047 18566 11056
rect 18696 11076 18748 11082
rect 18420 10736 18472 10742
rect 18420 10678 18472 10684
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 18052 10532 18104 10538
rect 18052 10474 18104 10480
rect 18064 10130 18092 10474
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 18156 9586 18184 10542
rect 18420 10532 18472 10538
rect 18420 10474 18472 10480
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18248 9586 18276 9862
rect 17868 9580 17920 9586
rect 18144 9580 18196 9586
rect 17868 9522 17920 9528
rect 18064 9540 18144 9568
rect 17776 9444 17828 9450
rect 17776 9386 17828 9392
rect 17788 8945 17816 9386
rect 17774 8936 17830 8945
rect 17774 8871 17776 8880
rect 17828 8871 17830 8880
rect 17776 8842 17828 8848
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17500 8288 17552 8294
rect 17500 8230 17552 8236
rect 17512 6118 17540 8230
rect 17880 8090 17908 9522
rect 18064 8650 18092 9540
rect 18144 9522 18196 9528
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18156 9110 18184 9318
rect 18144 9104 18196 9110
rect 18144 9046 18196 9052
rect 18248 8922 18276 9522
rect 17972 8622 18092 8650
rect 18156 8894 18276 8922
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17972 7954 18000 8622
rect 18050 8528 18106 8537
rect 18050 8463 18106 8472
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17592 7812 17644 7818
rect 17592 7754 17644 7760
rect 17604 7478 17632 7754
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 17774 6896 17830 6905
rect 17774 6831 17830 6840
rect 17788 6798 17816 6831
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17592 6724 17644 6730
rect 17592 6666 17644 6672
rect 17604 6497 17632 6666
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17590 6488 17646 6497
rect 17590 6423 17646 6432
rect 17696 6254 17724 6598
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17788 6118 17816 6258
rect 17500 6112 17552 6118
rect 17776 6112 17828 6118
rect 17500 6054 17552 6060
rect 17774 6080 17776 6089
rect 17868 6112 17920 6118
rect 17828 6080 17830 6089
rect 17868 6054 17920 6060
rect 17774 6015 17830 6024
rect 17880 5642 17908 6054
rect 17972 5817 18000 6734
rect 18064 6662 18092 8463
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 17958 5808 18014 5817
rect 17958 5743 18014 5752
rect 17868 5636 17920 5642
rect 17868 5578 17920 5584
rect 18064 5030 18092 5850
rect 18156 5166 18184 8894
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 18156 4622 18184 5102
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17696 3602 17724 3878
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17406 3224 17462 3233
rect 16580 3188 16632 3194
rect 17406 3159 17462 3168
rect 16580 3130 16632 3136
rect 10874 2680 10930 2689
rect 10874 2615 10930 2624
rect 17696 2446 17724 3538
rect 18248 3534 18276 8774
rect 18340 6882 18368 9522
rect 18432 9178 18460 10474
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 18524 9042 18552 11047
rect 18696 11018 18748 11024
rect 18800 10985 18828 11494
rect 18786 10976 18842 10985
rect 18786 10911 18842 10920
rect 18880 10736 18932 10742
rect 18880 10678 18932 10684
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18800 10577 18828 10610
rect 18786 10568 18842 10577
rect 18786 10503 18842 10512
rect 18602 9480 18658 9489
rect 18602 9415 18658 9424
rect 18616 9178 18644 9415
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18512 9036 18564 9042
rect 18564 8996 18644 9024
rect 18512 8978 18564 8984
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18524 7002 18552 7754
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18340 6854 18552 6882
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18432 6361 18460 6598
rect 18418 6352 18474 6361
rect 18418 6287 18474 6296
rect 18432 5953 18460 6287
rect 18418 5944 18474 5953
rect 18418 5879 18474 5888
rect 18524 5710 18552 6854
rect 18616 6458 18644 8996
rect 18708 8945 18736 9114
rect 18694 8936 18750 8945
rect 18694 8871 18750 8880
rect 18786 7848 18842 7857
rect 18786 7783 18842 7792
rect 18800 7546 18828 7783
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18892 6934 18920 10678
rect 18984 9518 19012 11716
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18880 6928 18932 6934
rect 18880 6870 18932 6876
rect 18708 6730 18920 6746
rect 18696 6724 18932 6730
rect 18748 6718 18880 6724
rect 18696 6666 18748 6672
rect 18880 6666 18932 6672
rect 18984 6662 19012 9454
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18788 6248 18840 6254
rect 18788 6190 18840 6196
rect 18800 5710 18828 6190
rect 18984 6118 19012 6598
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 18984 5778 19012 6054
rect 19076 5914 19104 10542
rect 19168 10062 19196 14334
rect 19340 14282 19392 14288
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19260 10985 19288 14214
rect 19352 13705 19380 14282
rect 19338 13696 19394 13705
rect 19338 13631 19394 13640
rect 19536 13326 19564 14368
rect 19708 14350 19760 14356
rect 19800 14408 19852 14414
rect 19800 14350 19852 14356
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19614 12336 19670 12345
rect 19614 12271 19670 12280
rect 19430 12200 19486 12209
rect 19340 12164 19392 12170
rect 19628 12170 19656 12271
rect 19430 12135 19432 12144
rect 19340 12106 19392 12112
rect 19484 12135 19486 12144
rect 19616 12164 19668 12170
rect 19432 12106 19484 12112
rect 19616 12106 19668 12112
rect 19352 11694 19380 12106
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19430 11928 19486 11937
rect 19430 11863 19486 11872
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 19352 11393 19380 11630
rect 19338 11384 19394 11393
rect 19338 11319 19394 11328
rect 19246 10976 19302 10985
rect 19246 10911 19302 10920
rect 19444 10810 19472 11863
rect 19536 11354 19564 12038
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19614 11248 19670 11257
rect 19614 11183 19670 11192
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19352 10470 19380 10610
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 19168 9722 19196 9998
rect 19260 9897 19288 10406
rect 19628 10130 19656 11183
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 19246 9888 19302 9897
rect 19246 9823 19302 9832
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 19352 9625 19380 9930
rect 19444 9761 19472 9930
rect 19430 9752 19486 9761
rect 19430 9687 19486 9696
rect 19614 9752 19670 9761
rect 19614 9687 19670 9696
rect 19338 9616 19394 9625
rect 19338 9551 19394 9560
rect 19352 9382 19380 9551
rect 19522 9480 19578 9489
rect 19522 9415 19578 9424
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19432 8560 19484 8566
rect 19430 8528 19432 8537
rect 19484 8528 19486 8537
rect 19430 8463 19486 8472
rect 19340 7812 19392 7818
rect 19340 7754 19392 7760
rect 19352 7478 19380 7754
rect 19340 7472 19392 7478
rect 19338 7440 19340 7449
rect 19392 7440 19394 7449
rect 19338 7375 19394 7384
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 19260 6934 19288 7142
rect 19248 6928 19300 6934
rect 19248 6870 19300 6876
rect 19260 6322 19288 6870
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19536 6254 19564 9415
rect 19628 6322 19656 9687
rect 19720 6390 19748 14350
rect 19812 13433 19840 14350
rect 19892 14000 19944 14006
rect 19890 13968 19892 13977
rect 19944 13968 19946 13977
rect 19890 13903 19946 13912
rect 20076 13728 20128 13734
rect 20076 13670 20128 13676
rect 20088 13530 20116 13670
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 19798 13424 19854 13433
rect 19798 13359 19854 13368
rect 19800 13320 19852 13326
rect 19800 13262 19852 13268
rect 19812 10792 19840 13262
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 20088 12442 20116 12786
rect 20076 12436 20128 12442
rect 20076 12378 20128 12384
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19890 11112 19946 11121
rect 19890 11047 19892 11056
rect 19944 11047 19946 11056
rect 19892 11018 19944 11024
rect 19812 10764 19932 10792
rect 19798 10568 19854 10577
rect 19798 10503 19854 10512
rect 19812 10266 19840 10503
rect 19904 10470 19932 10764
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19800 10260 19852 10266
rect 19800 10202 19852 10208
rect 19996 9586 20024 11290
rect 20076 10192 20128 10198
rect 20076 10134 20128 10140
rect 20088 9994 20116 10134
rect 20076 9988 20128 9994
rect 20076 9930 20128 9936
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 19812 8634 19840 9522
rect 19984 9444 20036 9450
rect 19984 9386 20036 9392
rect 19890 8664 19946 8673
rect 19800 8628 19852 8634
rect 19890 8599 19892 8608
rect 19800 8570 19852 8576
rect 19944 8599 19946 8608
rect 19892 8570 19944 8576
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19812 7936 19840 8434
rect 19904 8294 19932 8570
rect 19892 8288 19944 8294
rect 19892 8230 19944 8236
rect 19996 8090 20024 9386
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19984 7948 20036 7954
rect 19812 7908 19984 7936
rect 19984 7890 20036 7896
rect 20088 6798 20116 9930
rect 20180 8430 20208 19110
rect 20272 18426 20300 19994
rect 20352 19440 20404 19446
rect 20352 19382 20404 19388
rect 20442 19408 20498 19417
rect 20364 18698 20392 19382
rect 20442 19343 20444 19352
rect 20496 19343 20498 19352
rect 20444 19314 20496 19320
rect 20444 19236 20496 19242
rect 20444 19178 20496 19184
rect 20352 18692 20404 18698
rect 20352 18634 20404 18640
rect 20260 18420 20312 18426
rect 20260 18362 20312 18368
rect 20272 18290 20300 18362
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20272 17134 20300 17818
rect 20260 17128 20312 17134
rect 20260 17070 20312 17076
rect 20260 16720 20312 16726
rect 20258 16688 20260 16697
rect 20312 16688 20314 16697
rect 20258 16623 20314 16632
rect 20456 16574 20484 19178
rect 20548 18698 20576 22066
rect 20824 22094 20852 23190
rect 21008 22710 21036 24006
rect 20996 22704 21048 22710
rect 20916 22664 20996 22692
rect 20916 22574 20944 22664
rect 20996 22646 21048 22652
rect 20904 22568 20956 22574
rect 21100 22556 21128 24228
rect 21192 24206 21220 24278
rect 21180 24200 21232 24206
rect 21284 24177 21312 24534
rect 21362 24511 21418 24520
rect 21180 24142 21232 24148
rect 21270 24168 21326 24177
rect 21270 24103 21326 24112
rect 21272 24064 21324 24070
rect 21272 24006 21324 24012
rect 21180 23112 21232 23118
rect 21180 23054 21232 23060
rect 21192 22642 21220 23054
rect 21180 22636 21232 22642
rect 21180 22578 21232 22584
rect 20904 22510 20956 22516
rect 21008 22528 21128 22556
rect 20904 22432 20956 22438
rect 21008 22420 21036 22528
rect 21284 22438 21312 24006
rect 20956 22392 21036 22420
rect 21272 22432 21324 22438
rect 20904 22374 20956 22380
rect 21272 22374 21324 22380
rect 21180 22228 21232 22234
rect 21180 22170 21232 22176
rect 21192 22098 21220 22170
rect 20824 22066 21036 22094
rect 20720 22034 20772 22040
rect 20628 22024 20680 22030
rect 20628 21966 20680 21972
rect 20640 19553 20668 21966
rect 20732 21486 20760 22034
rect 20812 21616 20864 21622
rect 20810 21584 20812 21593
rect 20864 21584 20866 21593
rect 20810 21519 20866 21528
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20824 21010 20852 21286
rect 20812 21004 20864 21010
rect 20812 20946 20864 20952
rect 20904 20528 20956 20534
rect 20732 20476 20904 20482
rect 20732 20470 20956 20476
rect 20732 20466 20944 20470
rect 20720 20460 20944 20466
rect 20772 20454 20944 20460
rect 20720 20402 20772 20408
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20732 20058 20760 20198
rect 20720 20052 20772 20058
rect 20720 19994 20772 20000
rect 20904 20052 20956 20058
rect 20904 19994 20956 20000
rect 20810 19680 20866 19689
rect 20810 19615 20866 19624
rect 20626 19544 20682 19553
rect 20626 19479 20682 19488
rect 20718 19408 20774 19417
rect 20718 19343 20774 19352
rect 20536 18692 20588 18698
rect 20536 18634 20588 18640
rect 20548 17610 20576 18634
rect 20732 18630 20760 19343
rect 20824 19310 20852 19615
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20640 17746 20668 18022
rect 20628 17740 20680 17746
rect 20628 17682 20680 17688
rect 20536 17604 20588 17610
rect 20536 17546 20588 17552
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20640 17134 20668 17546
rect 20628 17128 20680 17134
rect 20628 17070 20680 17076
rect 20272 16546 20484 16574
rect 20272 15745 20300 16546
rect 20536 16516 20588 16522
rect 20536 16458 20588 16464
rect 20548 16402 20576 16458
rect 20364 16374 20576 16402
rect 20258 15736 20314 15745
rect 20258 15671 20314 15680
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20272 9654 20300 15302
rect 20364 14521 20392 16374
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20456 15706 20484 15846
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20444 15496 20496 15502
rect 20444 15438 20496 15444
rect 20456 15178 20484 15438
rect 20548 15366 20576 16050
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20456 15150 20576 15178
rect 20640 15162 20668 17070
rect 20810 16416 20866 16425
rect 20810 16351 20866 16360
rect 20718 16144 20774 16153
rect 20718 16079 20720 16088
rect 20772 16079 20774 16088
rect 20720 16050 20772 16056
rect 20718 16008 20774 16017
rect 20718 15943 20774 15952
rect 20732 15337 20760 15943
rect 20824 15366 20852 16351
rect 20916 16266 20944 19994
rect 21008 19854 21036 22066
rect 21180 22092 21232 22098
rect 21180 22034 21232 22040
rect 21376 22030 21404 24511
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 21364 21888 21416 21894
rect 21364 21830 21416 21836
rect 21180 21548 21232 21554
rect 21180 21490 21232 21496
rect 21192 21146 21220 21490
rect 21180 21140 21232 21146
rect 21180 21082 21232 21088
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 21180 21004 21232 21010
rect 21180 20946 21232 20952
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 21100 20097 21128 20402
rect 21086 20088 21142 20097
rect 21086 20023 21142 20032
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 21088 19848 21140 19854
rect 21088 19790 21140 19796
rect 20996 19236 21048 19242
rect 20996 19178 21048 19184
rect 21008 18766 21036 19178
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 20996 18080 21048 18086
rect 20996 18022 21048 18028
rect 21008 16590 21036 18022
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 20916 16238 21036 16266
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20812 15360 20864 15366
rect 20718 15328 20774 15337
rect 20812 15302 20864 15308
rect 20718 15263 20774 15272
rect 20444 15088 20496 15094
rect 20444 15030 20496 15036
rect 20350 14512 20406 14521
rect 20350 14447 20406 14456
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20364 13977 20392 14350
rect 20456 14249 20484 15030
rect 20548 14278 20576 15150
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20626 15056 20682 15065
rect 20626 14991 20682 15000
rect 20536 14272 20588 14278
rect 20442 14240 20498 14249
rect 20536 14214 20588 14220
rect 20442 14175 20498 14184
rect 20536 14000 20588 14006
rect 20350 13968 20406 13977
rect 20536 13942 20588 13948
rect 20350 13903 20406 13912
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20352 13796 20404 13802
rect 20352 13738 20404 13744
rect 20364 13394 20392 13738
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20364 11665 20392 11698
rect 20350 11656 20406 11665
rect 20350 11591 20406 11600
rect 20456 11354 20484 13874
rect 20548 13734 20576 13942
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 20548 12986 20576 13194
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 20548 11762 20576 12378
rect 20640 11762 20668 14991
rect 20812 14612 20864 14618
rect 20812 14554 20864 14560
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20732 13870 20760 14486
rect 20824 14074 20852 14554
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20810 13696 20866 13705
rect 20732 11898 20760 13670
rect 20810 13631 20866 13640
rect 20824 13326 20852 13631
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 20536 11552 20588 11558
rect 20536 11494 20588 11500
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20548 11218 20576 11494
rect 20444 11212 20496 11218
rect 20444 11154 20496 11160
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 20350 11112 20406 11121
rect 20456 11098 20484 11154
rect 20732 11150 20760 11834
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20720 11144 20772 11150
rect 20456 11070 20576 11098
rect 20720 11086 20772 11092
rect 20350 11047 20406 11056
rect 20364 10996 20392 11047
rect 20364 10968 20484 10996
rect 20350 10840 20406 10849
rect 20350 10775 20352 10784
rect 20404 10775 20406 10784
rect 20352 10746 20404 10752
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20364 10198 20392 10406
rect 20352 10192 20404 10198
rect 20352 10134 20404 10140
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20260 9648 20312 9654
rect 20364 9625 20392 9998
rect 20456 9926 20484 10968
rect 20548 10962 20576 11070
rect 20548 10934 20760 10962
rect 20534 10840 20590 10849
rect 20732 10810 20760 10934
rect 20720 10804 20772 10810
rect 20590 10784 20668 10792
rect 20534 10775 20536 10784
rect 20588 10764 20668 10784
rect 20536 10746 20588 10752
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 20548 9722 20576 10610
rect 20640 10470 20668 10764
rect 20720 10746 20772 10752
rect 20720 10532 20772 10538
rect 20720 10474 20772 10480
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20626 10296 20682 10305
rect 20732 10266 20760 10474
rect 20626 10231 20682 10240
rect 20720 10260 20772 10266
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20260 9590 20312 9596
rect 20350 9616 20406 9625
rect 20350 9551 20406 9560
rect 20444 9580 20496 9586
rect 20444 9522 20496 9528
rect 20350 9208 20406 9217
rect 20350 9143 20406 9152
rect 20364 8673 20392 9143
rect 20350 8664 20406 8673
rect 20350 8599 20406 8608
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20180 8090 20208 8366
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20180 7342 20208 7822
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 20258 6896 20314 6905
rect 20258 6831 20260 6840
rect 20312 6831 20314 6840
rect 20260 6802 20312 6808
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 19996 6390 20024 6734
rect 19708 6384 19760 6390
rect 19708 6326 19760 6332
rect 19984 6384 20036 6390
rect 19984 6326 20036 6332
rect 19616 6316 19668 6322
rect 19616 6258 19668 6264
rect 19524 6248 19576 6254
rect 19524 6190 19576 6196
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 18972 5772 19024 5778
rect 18972 5714 19024 5720
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18788 5704 18840 5710
rect 19536 5681 19564 6190
rect 18788 5646 18840 5652
rect 19522 5672 19578 5681
rect 18524 5234 18552 5646
rect 19628 5642 19656 6258
rect 20088 6118 20116 6734
rect 20076 6112 20128 6118
rect 20076 6054 20128 6060
rect 20352 6112 20404 6118
rect 20352 6054 20404 6060
rect 20364 5846 20392 6054
rect 20352 5840 20404 5846
rect 20352 5782 20404 5788
rect 20456 5710 20484 9522
rect 20640 7886 20668 10231
rect 20720 10202 20772 10208
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 20534 6760 20590 6769
rect 20534 6695 20590 6704
rect 20548 6662 20576 6695
rect 20640 6662 20668 6938
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20534 6488 20590 6497
rect 20534 6423 20590 6432
rect 20548 6322 20576 6423
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20640 6186 20668 6598
rect 20732 6390 20760 10202
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20628 6180 20680 6186
rect 20628 6122 20680 6128
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20718 5672 20774 5681
rect 19522 5607 19578 5616
rect 19616 5636 19668 5642
rect 20718 5607 20774 5616
rect 19616 5578 19668 5584
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 19708 4616 19760 4622
rect 20732 4593 20760 5607
rect 20824 4622 20852 11290
rect 20916 11121 20944 16050
rect 21008 12434 21036 16238
rect 21100 14074 21128 19790
rect 21192 19786 21220 20946
rect 21180 19780 21232 19786
rect 21180 19722 21232 19728
rect 21284 19666 21312 21082
rect 21192 19638 21312 19666
rect 21192 18442 21220 19638
rect 21272 18964 21324 18970
rect 21272 18906 21324 18912
rect 21284 18873 21312 18906
rect 21270 18864 21326 18873
rect 21270 18799 21326 18808
rect 21192 18414 21312 18442
rect 21180 18352 21232 18358
rect 21180 18294 21232 18300
rect 21192 15910 21220 18294
rect 21284 15910 21312 18414
rect 21180 15904 21232 15910
rect 21180 15846 21232 15852
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21376 15722 21404 21830
rect 21468 20330 21496 24686
rect 21640 24608 21692 24614
rect 21640 24550 21692 24556
rect 21548 24404 21600 24410
rect 21548 24346 21600 24352
rect 21560 21146 21588 24346
rect 21652 24274 21680 24550
rect 21640 24268 21692 24274
rect 21640 24210 21692 24216
rect 21638 24168 21694 24177
rect 21638 24103 21694 24112
rect 21652 23202 21680 24103
rect 21744 23798 21772 24806
rect 21836 24800 21864 26318
rect 21928 26217 21956 26386
rect 21914 26208 21970 26217
rect 21914 26143 21970 26152
rect 21916 26036 21968 26042
rect 21916 25978 21968 25984
rect 21928 25906 21956 25978
rect 21916 25900 21968 25906
rect 21916 25842 21968 25848
rect 21916 25288 21968 25294
rect 21914 25256 21916 25265
rect 21968 25256 21970 25265
rect 21914 25191 21970 25200
rect 21836 24772 21956 24800
rect 21824 24676 21876 24682
rect 21824 24618 21876 24624
rect 21732 23792 21784 23798
rect 21732 23734 21784 23740
rect 21744 23322 21772 23734
rect 21836 23497 21864 24618
rect 21928 24313 21956 24772
rect 21914 24304 21970 24313
rect 21914 24239 21970 24248
rect 21914 24168 21970 24177
rect 21914 24103 21970 24112
rect 21928 24070 21956 24103
rect 21916 24064 21968 24070
rect 21916 24006 21968 24012
rect 21822 23488 21878 23497
rect 21822 23423 21878 23432
rect 21732 23316 21784 23322
rect 21732 23258 21784 23264
rect 21652 23174 21772 23202
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 21548 21140 21600 21146
rect 21548 21082 21600 21088
rect 21652 21049 21680 22510
rect 21638 21040 21694 21049
rect 21638 20975 21694 20984
rect 21548 20868 21600 20874
rect 21548 20810 21600 20816
rect 21640 20868 21692 20874
rect 21640 20810 21692 20816
rect 21456 20324 21508 20330
rect 21456 20266 21508 20272
rect 21560 20040 21588 20810
rect 21652 20466 21680 20810
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 21640 20324 21692 20330
rect 21640 20266 21692 20272
rect 21468 20012 21588 20040
rect 21468 19145 21496 20012
rect 21652 19972 21680 20266
rect 21560 19944 21680 19972
rect 21454 19136 21510 19145
rect 21454 19071 21510 19080
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21468 18426 21496 18702
rect 21456 18420 21508 18426
rect 21456 18362 21508 18368
rect 21456 18148 21508 18154
rect 21456 18090 21508 18096
rect 21192 15694 21404 15722
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 21100 12918 21128 13874
rect 21088 12912 21140 12918
rect 21088 12854 21140 12860
rect 21008 12406 21128 12434
rect 20996 12164 21048 12170
rect 20996 12106 21048 12112
rect 20902 11112 20958 11121
rect 20902 11047 20958 11056
rect 20902 10976 20958 10985
rect 20902 10911 20958 10920
rect 20916 10606 20944 10911
rect 20904 10600 20956 10606
rect 20904 10542 20956 10548
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 21008 10418 21036 12106
rect 21100 10985 21128 12406
rect 21192 11218 21220 15694
rect 21468 15586 21496 18090
rect 21560 17678 21588 19944
rect 21744 19904 21772 23174
rect 21824 23112 21876 23118
rect 22020 23066 22048 26794
rect 22480 26790 22508 27610
rect 22572 27130 22600 28018
rect 22928 27328 22980 27334
rect 22928 27270 22980 27276
rect 22560 27124 22612 27130
rect 22560 27066 22612 27072
rect 22560 26988 22612 26994
rect 22560 26930 22612 26936
rect 22468 26784 22520 26790
rect 22468 26726 22520 26732
rect 22480 25922 22508 26726
rect 22388 25894 22508 25922
rect 22100 25152 22152 25158
rect 22100 25094 22152 25100
rect 22112 24886 22140 25094
rect 22100 24880 22152 24886
rect 22100 24822 22152 24828
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 22100 24676 22152 24682
rect 22100 24618 22152 24624
rect 22112 24585 22140 24618
rect 22098 24576 22154 24585
rect 22098 24511 22154 24520
rect 22204 24410 22232 24754
rect 22282 24712 22338 24721
rect 22282 24647 22338 24656
rect 22192 24404 22244 24410
rect 22192 24346 22244 24352
rect 22296 23730 22324 24647
rect 22284 23724 22336 23730
rect 22284 23666 22336 23672
rect 22192 23520 22244 23526
rect 22192 23462 22244 23468
rect 22204 23118 22232 23462
rect 22282 23216 22338 23225
rect 22388 23186 22416 25894
rect 22572 24954 22600 26930
rect 22836 26784 22888 26790
rect 22742 26752 22798 26761
rect 22836 26726 22888 26732
rect 22742 26687 22798 26696
rect 22756 26450 22784 26687
rect 22848 26586 22876 26726
rect 22836 26580 22888 26586
rect 22836 26522 22888 26528
rect 22744 26444 22796 26450
rect 22744 26386 22796 26392
rect 22742 26344 22798 26353
rect 22742 26279 22798 26288
rect 22652 25900 22704 25906
rect 22652 25842 22704 25848
rect 22664 25430 22692 25842
rect 22756 25498 22784 26279
rect 22836 26240 22888 26246
rect 22836 26182 22888 26188
rect 22848 26042 22876 26182
rect 22836 26036 22888 26042
rect 22836 25978 22888 25984
rect 22940 25786 22968 27270
rect 22848 25758 22968 25786
rect 22744 25492 22796 25498
rect 22744 25434 22796 25440
rect 22652 25424 22704 25430
rect 22652 25366 22704 25372
rect 22756 25294 22784 25434
rect 22652 25288 22704 25294
rect 22650 25256 22652 25265
rect 22744 25288 22796 25294
rect 22704 25256 22706 25265
rect 22744 25230 22796 25236
rect 22650 25191 22706 25200
rect 22560 24948 22612 24954
rect 22560 24890 22612 24896
rect 22744 24948 22796 24954
rect 22744 24890 22796 24896
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 22560 24812 22612 24818
rect 22756 24800 22784 24890
rect 22560 24754 22612 24760
rect 22664 24772 22784 24800
rect 22282 23151 22338 23160
rect 22376 23180 22428 23186
rect 21824 23054 21876 23060
rect 21836 22098 21864 23054
rect 21928 23038 22048 23066
rect 22192 23112 22244 23118
rect 22192 23054 22244 23060
rect 21928 22982 21956 23038
rect 21916 22976 21968 22982
rect 21916 22918 21968 22924
rect 22008 22976 22060 22982
rect 22008 22918 22060 22924
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22020 22234 22048 22918
rect 22008 22228 22060 22234
rect 22008 22170 22060 22176
rect 21824 22092 21876 22098
rect 21824 22034 21876 22040
rect 22006 21040 22062 21049
rect 22006 20975 22062 20984
rect 21652 19876 21772 19904
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 21652 16810 21680 19876
rect 21730 19272 21786 19281
rect 21730 19207 21786 19216
rect 21744 18834 21772 19207
rect 21916 18964 21968 18970
rect 21916 18906 21968 18912
rect 21732 18828 21784 18834
rect 21732 18770 21784 18776
rect 21824 18760 21876 18766
rect 21824 18702 21876 18708
rect 21836 18426 21864 18702
rect 21824 18420 21876 18426
rect 21824 18362 21876 18368
rect 21928 17746 21956 18906
rect 22020 18737 22048 20975
rect 22006 18728 22062 18737
rect 22006 18663 22062 18672
rect 22006 18048 22062 18057
rect 22006 17983 22062 17992
rect 21916 17740 21968 17746
rect 21916 17682 21968 17688
rect 21824 17604 21876 17610
rect 21824 17546 21876 17552
rect 21652 16782 21772 16810
rect 21640 16720 21692 16726
rect 21640 16662 21692 16668
rect 21546 16008 21602 16017
rect 21546 15943 21602 15952
rect 21376 15558 21496 15586
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21284 13938 21312 14758
rect 21376 13938 21404 15558
rect 21456 14340 21508 14346
rect 21456 14282 21508 14288
rect 21468 14249 21496 14282
rect 21454 14240 21510 14249
rect 21454 14175 21510 14184
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21364 13932 21416 13938
rect 21364 13874 21416 13880
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21468 13841 21496 13874
rect 21454 13832 21510 13841
rect 21454 13767 21510 13776
rect 21560 13705 21588 15943
rect 21652 15638 21680 16662
rect 21640 15632 21692 15638
rect 21640 15574 21692 15580
rect 21640 15088 21692 15094
rect 21640 15030 21692 15036
rect 21652 14346 21680 15030
rect 21640 14340 21692 14346
rect 21640 14282 21692 14288
rect 21652 13802 21680 14282
rect 21744 13938 21772 16782
rect 21836 15706 21864 17546
rect 22020 17270 22048 17983
rect 22008 17264 22060 17270
rect 22008 17206 22060 17212
rect 22112 15994 22140 22918
rect 22296 22624 22324 23151
rect 22376 23122 22428 23128
rect 22480 22778 22508 24754
rect 22572 23322 22600 24754
rect 22664 24410 22692 24772
rect 22848 24698 22876 25758
rect 22928 25696 22980 25702
rect 22928 25638 22980 25644
rect 22940 24886 22968 25638
rect 22928 24880 22980 24886
rect 22928 24822 22980 24828
rect 22756 24682 22876 24698
rect 22744 24676 22876 24682
rect 22796 24670 22876 24676
rect 22744 24618 22796 24624
rect 22652 24404 22704 24410
rect 22652 24346 22704 24352
rect 22560 23316 22612 23322
rect 22560 23258 22612 23264
rect 22756 23225 22784 24618
rect 22836 24608 22888 24614
rect 22836 24550 22888 24556
rect 22848 23322 22876 24550
rect 22836 23316 22888 23322
rect 22836 23258 22888 23264
rect 22742 23216 22798 23225
rect 22742 23151 22798 23160
rect 22560 23044 22612 23050
rect 22560 22986 22612 22992
rect 22652 23044 22704 23050
rect 22652 22986 22704 22992
rect 22468 22772 22520 22778
rect 22468 22714 22520 22720
rect 22376 22636 22428 22642
rect 22296 22596 22376 22624
rect 22376 22578 22428 22584
rect 22284 22432 22336 22438
rect 22284 22374 22336 22380
rect 22296 22030 22324 22374
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22204 21146 22232 21966
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 22388 21078 22416 22578
rect 22572 22506 22600 22986
rect 22664 22545 22692 22986
rect 22744 22976 22796 22982
rect 22742 22944 22744 22953
rect 22836 22976 22888 22982
rect 22796 22944 22798 22953
rect 22836 22918 22888 22924
rect 22742 22879 22798 22888
rect 22744 22636 22796 22642
rect 22744 22578 22796 22584
rect 22650 22536 22706 22545
rect 22560 22500 22612 22506
rect 22650 22471 22706 22480
rect 22560 22442 22612 22448
rect 22572 22030 22600 22442
rect 22756 22273 22784 22578
rect 22742 22264 22798 22273
rect 22652 22228 22704 22234
rect 22742 22199 22798 22208
rect 22652 22170 22704 22176
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 22376 21072 22428 21078
rect 22376 21014 22428 21020
rect 22572 21010 22600 21830
rect 22560 21004 22612 21010
rect 22560 20946 22612 20952
rect 22558 20496 22614 20505
rect 22558 20431 22560 20440
rect 22612 20431 22614 20440
rect 22560 20402 22612 20408
rect 22284 20392 22336 20398
rect 22284 20334 22336 20340
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 22204 18154 22232 19858
rect 22192 18148 22244 18154
rect 22192 18090 22244 18096
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 22204 17542 22232 17818
rect 22296 17746 22324 20334
rect 22558 19952 22614 19961
rect 22558 19887 22614 19896
rect 22572 19378 22600 19887
rect 22560 19372 22612 19378
rect 22560 19314 22612 19320
rect 22376 19168 22428 19174
rect 22664 19122 22692 22170
rect 22742 21720 22798 21729
rect 22742 21655 22798 21664
rect 22756 20913 22784 21655
rect 22742 20904 22798 20913
rect 22742 20839 22798 20848
rect 22756 19174 22784 20839
rect 22376 19110 22428 19116
rect 22388 18086 22416 19110
rect 22572 19094 22692 19122
rect 22744 19168 22796 19174
rect 22744 19110 22796 19116
rect 22466 19000 22522 19009
rect 22466 18935 22468 18944
rect 22520 18935 22522 18944
rect 22468 18906 22520 18912
rect 22468 18760 22520 18766
rect 22466 18728 22468 18737
rect 22520 18728 22522 18737
rect 22466 18663 22522 18672
rect 22572 18306 22600 19094
rect 22652 18964 22704 18970
rect 22652 18906 22704 18912
rect 22480 18278 22600 18306
rect 22376 18080 22428 18086
rect 22376 18022 22428 18028
rect 22284 17740 22336 17746
rect 22284 17682 22336 17688
rect 22480 17678 22508 18278
rect 22558 18184 22614 18193
rect 22558 18119 22614 18128
rect 22468 17672 22520 17678
rect 22468 17614 22520 17620
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22284 17060 22336 17066
rect 22284 17002 22336 17008
rect 22296 16794 22324 17002
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22480 16658 22508 17614
rect 22572 17270 22600 18119
rect 22664 17882 22692 18906
rect 22744 18896 22796 18902
rect 22744 18838 22796 18844
rect 22756 18358 22784 18838
rect 22744 18352 22796 18358
rect 22744 18294 22796 18300
rect 22652 17876 22704 17882
rect 22652 17818 22704 17824
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 22560 17264 22612 17270
rect 22560 17206 22612 17212
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22112 15966 22232 15994
rect 21916 15904 21968 15910
rect 21916 15846 21968 15852
rect 21824 15700 21876 15706
rect 21824 15642 21876 15648
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 21732 13932 21784 13938
rect 21732 13874 21784 13880
rect 21836 13818 21864 15370
rect 21640 13796 21692 13802
rect 21640 13738 21692 13744
rect 21744 13790 21864 13818
rect 21546 13696 21602 13705
rect 21546 13631 21602 13640
rect 21744 13546 21772 13790
rect 21824 13728 21876 13734
rect 21824 13670 21876 13676
rect 21468 13518 21772 13546
rect 21272 13456 21324 13462
rect 21272 13398 21324 13404
rect 21284 13258 21312 13398
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21272 13252 21324 13258
rect 21272 13194 21324 13200
rect 21376 13138 21404 13262
rect 21284 13110 21404 13138
rect 21284 12306 21312 13110
rect 21468 12442 21496 13518
rect 21640 13456 21692 13462
rect 21640 13398 21692 13404
rect 21548 13184 21600 13190
rect 21548 13126 21600 13132
rect 21456 12436 21508 12442
rect 21456 12378 21508 12384
rect 21454 12336 21510 12345
rect 21272 12300 21324 12306
rect 21454 12271 21510 12280
rect 21272 12242 21324 12248
rect 21180 11212 21232 11218
rect 21180 11154 21232 11160
rect 21086 10976 21142 10985
rect 21086 10911 21142 10920
rect 21100 10742 21128 10911
rect 21088 10736 21140 10742
rect 21088 10678 21140 10684
rect 21178 10568 21234 10577
rect 21178 10503 21234 10512
rect 21192 10470 21220 10503
rect 21180 10464 21232 10470
rect 20916 9674 20944 10406
rect 21008 10390 21128 10418
rect 21180 10406 21232 10412
rect 20916 9646 21036 9674
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20916 8566 20944 9522
rect 21008 9382 21036 9646
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 20904 8560 20956 8566
rect 20904 8502 20956 8508
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 20904 8424 20956 8430
rect 20904 8366 20956 8372
rect 20916 5914 20944 8366
rect 21008 8090 21036 8434
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 21008 7721 21036 8026
rect 20994 7712 21050 7721
rect 20994 7647 21050 7656
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 21008 5710 21036 5850
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 21100 5370 21128 10390
rect 21180 9580 21232 9586
rect 21284 9568 21312 12242
rect 21468 12238 21496 12271
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 21560 11898 21588 13126
rect 21652 12782 21680 13398
rect 21732 13388 21784 13394
rect 21732 13330 21784 13336
rect 21744 13297 21772 13330
rect 21730 13288 21786 13297
rect 21730 13223 21786 13232
rect 21836 13025 21864 13670
rect 21822 13016 21878 13025
rect 21822 12951 21878 12960
rect 21928 12782 21956 15846
rect 22006 15736 22062 15745
rect 22006 15671 22062 15680
rect 22020 15502 22048 15671
rect 22204 15570 22232 15966
rect 22296 15638 22324 16458
rect 22468 15904 22520 15910
rect 22468 15846 22520 15852
rect 22480 15706 22508 15846
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 22192 15564 22244 15570
rect 22664 15552 22692 17682
rect 22742 17640 22798 17649
rect 22742 17575 22798 17584
rect 22192 15506 22244 15512
rect 22572 15524 22692 15552
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 21640 12776 21692 12782
rect 21640 12718 21692 12724
rect 21916 12776 21968 12782
rect 21916 12718 21968 12724
rect 21640 12640 21692 12646
rect 22020 12594 22048 15438
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 22112 13870 22140 14962
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22098 13288 22154 13297
rect 22098 13223 22154 13232
rect 22112 12850 22140 13223
rect 22204 12850 22232 15506
rect 22468 15428 22520 15434
rect 22468 15370 22520 15376
rect 22480 15162 22508 15370
rect 22572 15178 22600 15524
rect 22652 15428 22704 15434
rect 22652 15370 22704 15376
rect 22664 15337 22692 15370
rect 22650 15328 22706 15337
rect 22756 15314 22784 17575
rect 22848 16182 22876 22918
rect 22940 18970 22968 24822
rect 23032 24721 23060 30223
rect 23124 25906 23152 31175
rect 23570 30968 23626 30977
rect 23570 30903 23626 30912
rect 23202 29472 23258 29481
rect 23202 29407 23258 29416
rect 23216 28558 23244 29407
rect 23294 28656 23350 28665
rect 23294 28591 23350 28600
rect 23204 28552 23256 28558
rect 23204 28494 23256 28500
rect 23308 28150 23336 28591
rect 23388 28552 23440 28558
rect 23388 28494 23440 28500
rect 23584 28506 23612 30903
rect 23676 29850 23704 31282
rect 23664 29844 23716 29850
rect 23664 29786 23716 29792
rect 24492 29572 24544 29578
rect 24492 29514 24544 29520
rect 24504 29306 24532 29514
rect 25332 29510 25360 31282
rect 26976 30796 27028 30802
rect 26976 30738 27028 30744
rect 26148 30252 26200 30258
rect 26148 30194 26200 30200
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 25320 29504 25372 29510
rect 25320 29446 25372 29452
rect 24492 29300 24544 29306
rect 24492 29242 24544 29248
rect 25332 29170 25360 29446
rect 25320 29164 25372 29170
rect 25320 29106 25372 29112
rect 23756 29096 23808 29102
rect 24400 29096 24452 29102
rect 23808 29056 24072 29084
rect 23756 29038 23808 29044
rect 23756 28960 23808 28966
rect 23756 28902 23808 28908
rect 23768 28558 23796 28902
rect 23756 28552 23808 28558
rect 23296 28144 23348 28150
rect 23296 28086 23348 28092
rect 23400 27878 23428 28494
rect 23480 28484 23532 28490
rect 23584 28478 23704 28506
rect 23756 28494 23808 28500
rect 23480 28426 23532 28432
rect 23388 27872 23440 27878
rect 23492 27849 23520 28426
rect 23572 28416 23624 28422
rect 23572 28358 23624 28364
rect 23388 27814 23440 27820
rect 23478 27840 23534 27849
rect 23478 27775 23534 27784
rect 23584 27713 23612 28358
rect 23570 27704 23626 27713
rect 23570 27639 23626 27648
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 23296 26988 23348 26994
rect 23296 26930 23348 26936
rect 23204 26784 23256 26790
rect 23204 26726 23256 26732
rect 23216 26450 23244 26726
rect 23204 26444 23256 26450
rect 23204 26386 23256 26392
rect 23308 26314 23336 26930
rect 23480 26512 23532 26518
rect 23480 26454 23532 26460
rect 23296 26308 23348 26314
rect 23296 26250 23348 26256
rect 23492 25906 23520 26454
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 23124 25294 23152 25842
rect 23478 25800 23534 25809
rect 23478 25735 23534 25744
rect 23492 25430 23520 25735
rect 23480 25424 23532 25430
rect 23480 25366 23532 25372
rect 23584 25378 23612 27406
rect 23676 25702 23704 28478
rect 23768 28082 23796 28494
rect 23940 28416 23992 28422
rect 23940 28358 23992 28364
rect 23756 28076 23808 28082
rect 23756 28018 23808 28024
rect 23952 27470 23980 28358
rect 23940 27464 23992 27470
rect 23846 27432 23902 27441
rect 23940 27406 23992 27412
rect 23846 27367 23848 27376
rect 23900 27367 23902 27376
rect 23848 27338 23900 27344
rect 23952 27334 23980 27406
rect 23940 27328 23992 27334
rect 23940 27270 23992 27276
rect 23756 27056 23808 27062
rect 23756 26998 23808 27004
rect 23768 26790 23796 26998
rect 23756 26784 23808 26790
rect 23756 26726 23808 26732
rect 23768 26450 23796 26726
rect 23756 26444 23808 26450
rect 23756 26386 23808 26392
rect 23848 25764 23900 25770
rect 23848 25706 23900 25712
rect 23664 25696 23716 25702
rect 23664 25638 23716 25644
rect 23676 25498 23704 25638
rect 23664 25492 23716 25498
rect 23664 25434 23716 25440
rect 23754 25392 23810 25401
rect 23112 25288 23164 25294
rect 23492 25276 23520 25366
rect 23584 25350 23704 25378
rect 23492 25248 23612 25276
rect 23112 25230 23164 25236
rect 23204 25152 23256 25158
rect 23204 25094 23256 25100
rect 23388 25152 23440 25158
rect 23388 25094 23440 25100
rect 23112 24812 23164 24818
rect 23112 24754 23164 24760
rect 23018 24712 23074 24721
rect 23018 24647 23074 24656
rect 23032 24206 23060 24647
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 23124 24070 23152 24754
rect 23216 24750 23244 25094
rect 23400 24800 23428 25094
rect 23480 24812 23532 24818
rect 23308 24772 23480 24800
rect 23204 24744 23256 24750
rect 23204 24686 23256 24692
rect 23112 24064 23164 24070
rect 23112 24006 23164 24012
rect 23020 22432 23072 22438
rect 23020 22374 23072 22380
rect 23032 22234 23060 22374
rect 23020 22228 23072 22234
rect 23020 22170 23072 22176
rect 23124 22094 23152 24006
rect 23032 22066 23152 22094
rect 23032 20398 23060 22066
rect 23216 22030 23244 24686
rect 23308 24614 23336 24772
rect 23480 24754 23532 24760
rect 23386 24712 23442 24721
rect 23584 24698 23612 25248
rect 23386 24647 23442 24656
rect 23492 24670 23612 24698
rect 23400 24614 23428 24647
rect 23296 24608 23348 24614
rect 23296 24550 23348 24556
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23386 23896 23442 23905
rect 23386 23831 23442 23840
rect 23296 23656 23348 23662
rect 23296 23598 23348 23604
rect 23308 23118 23336 23598
rect 23400 23594 23428 23831
rect 23388 23588 23440 23594
rect 23388 23530 23440 23536
rect 23296 23112 23348 23118
rect 23296 23054 23348 23060
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 23112 21888 23164 21894
rect 23112 21830 23164 21836
rect 23124 21622 23152 21830
rect 23112 21616 23164 21622
rect 23112 21558 23164 21564
rect 23112 20936 23164 20942
rect 23112 20878 23164 20884
rect 23020 20392 23072 20398
rect 23020 20334 23072 20340
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 23032 19378 23060 20198
rect 23124 19922 23152 20878
rect 23112 19916 23164 19922
rect 23112 19858 23164 19864
rect 23020 19372 23072 19378
rect 23020 19314 23072 19320
rect 22928 18964 22980 18970
rect 22928 18906 22980 18912
rect 22928 18692 22980 18698
rect 22928 18634 22980 18640
rect 22836 16176 22888 16182
rect 22836 16118 22888 16124
rect 22848 15450 22876 16118
rect 22940 16046 22968 18634
rect 22928 16040 22980 16046
rect 22928 15982 22980 15988
rect 22926 15736 22982 15745
rect 23032 15706 23060 19314
rect 23112 18760 23164 18766
rect 23112 18702 23164 18708
rect 23124 17082 23152 18702
rect 23216 17678 23244 21966
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23308 19417 23336 20402
rect 23294 19408 23350 19417
rect 23294 19343 23350 19352
rect 23400 18970 23428 22714
rect 23492 21486 23520 24670
rect 23676 24562 23704 25350
rect 23754 25327 23810 25336
rect 23768 24954 23796 25327
rect 23756 24948 23808 24954
rect 23756 24890 23808 24896
rect 23860 24682 23888 25706
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 23848 24676 23900 24682
rect 23848 24618 23900 24624
rect 23676 24534 23888 24562
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23572 24132 23624 24138
rect 23572 24074 23624 24080
rect 23584 23497 23612 24074
rect 23676 24041 23704 24142
rect 23756 24132 23808 24138
rect 23756 24074 23808 24080
rect 23662 24032 23718 24041
rect 23662 23967 23718 23976
rect 23768 23633 23796 24074
rect 23754 23624 23810 23633
rect 23860 23610 23888 24534
rect 23952 23730 23980 24754
rect 24044 23882 24072 29056
rect 24400 29038 24452 29044
rect 24216 27668 24268 27674
rect 24216 27610 24268 27616
rect 24228 27577 24256 27610
rect 24214 27568 24270 27577
rect 24214 27503 24270 27512
rect 24124 27396 24176 27402
rect 24124 27338 24176 27344
rect 24136 25158 24164 27338
rect 24308 26376 24360 26382
rect 24308 26318 24360 26324
rect 24216 25696 24268 25702
rect 24216 25638 24268 25644
rect 24228 25498 24256 25638
rect 24216 25492 24268 25498
rect 24216 25434 24268 25440
rect 24216 25220 24268 25226
rect 24216 25162 24268 25168
rect 24124 25152 24176 25158
rect 24124 25094 24176 25100
rect 24228 24886 24256 25162
rect 24320 24993 24348 26318
rect 24306 24984 24362 24993
rect 24306 24919 24362 24928
rect 24216 24880 24268 24886
rect 24216 24822 24268 24828
rect 24320 24750 24348 24919
rect 24308 24744 24360 24750
rect 24308 24686 24360 24692
rect 24308 24608 24360 24614
rect 24308 24550 24360 24556
rect 24216 24268 24268 24274
rect 24216 24210 24268 24216
rect 24044 23854 24164 23882
rect 23940 23724 23992 23730
rect 23940 23666 23992 23672
rect 24030 23624 24086 23633
rect 23860 23582 23980 23610
rect 23754 23559 23810 23568
rect 23848 23520 23900 23526
rect 23570 23488 23626 23497
rect 23570 23423 23626 23432
rect 23846 23488 23848 23497
rect 23900 23488 23902 23497
rect 23846 23423 23902 23432
rect 23952 23338 23980 23582
rect 24030 23559 24086 23568
rect 24044 23526 24072 23559
rect 24032 23520 24084 23526
rect 24032 23462 24084 23468
rect 23572 23316 23624 23322
rect 23572 23258 23624 23264
rect 23860 23310 23980 23338
rect 23480 21480 23532 21486
rect 23480 21422 23532 21428
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 23492 21146 23520 21286
rect 23480 21140 23532 21146
rect 23480 21082 23532 21088
rect 23584 19334 23612 23258
rect 23756 21956 23808 21962
rect 23756 21898 23808 21904
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 23492 19306 23612 19334
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 23492 18834 23520 19306
rect 23572 19168 23624 19174
rect 23572 19110 23624 19116
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23492 18698 23520 18770
rect 23584 18698 23612 19110
rect 23480 18692 23532 18698
rect 23480 18634 23532 18640
rect 23572 18692 23624 18698
rect 23572 18634 23624 18640
rect 23480 18284 23532 18290
rect 23480 18226 23532 18232
rect 23492 17882 23520 18226
rect 23480 17876 23532 17882
rect 23480 17818 23532 17824
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23202 17232 23258 17241
rect 23202 17167 23204 17176
rect 23256 17167 23258 17176
rect 23204 17138 23256 17144
rect 23492 17134 23520 17818
rect 23480 17128 23532 17134
rect 23124 17054 23244 17082
rect 23480 17070 23532 17076
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 22926 15671 22982 15680
rect 23020 15700 23072 15706
rect 22940 15570 22968 15671
rect 23020 15642 23072 15648
rect 22928 15564 22980 15570
rect 22928 15506 22980 15512
rect 22848 15434 22968 15450
rect 22848 15428 22980 15434
rect 22848 15422 22928 15428
rect 22928 15370 22980 15376
rect 22756 15286 23060 15314
rect 22650 15263 22706 15272
rect 22468 15156 22520 15162
rect 22572 15150 22784 15178
rect 22468 15098 22520 15104
rect 22374 14648 22430 14657
rect 22374 14583 22430 14592
rect 22282 14240 22338 14249
rect 22282 14175 22338 14184
rect 22296 13734 22324 14175
rect 22388 14006 22416 14583
rect 22376 14000 22428 14006
rect 22376 13942 22428 13948
rect 22480 13938 22508 15098
rect 22560 14340 22612 14346
rect 22560 14282 22612 14288
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22572 13734 22600 14282
rect 22652 13864 22704 13870
rect 22652 13806 22704 13812
rect 22284 13728 22336 13734
rect 22468 13728 22520 13734
rect 22284 13670 22336 13676
rect 22374 13696 22430 13705
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 21640 12582 21692 12588
rect 21652 12306 21680 12582
rect 21744 12566 22048 12594
rect 22098 12608 22154 12617
rect 21640 12300 21692 12306
rect 21640 12242 21692 12248
rect 21652 12170 21680 12242
rect 21640 12164 21692 12170
rect 21640 12106 21692 12112
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21376 11558 21404 11834
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21376 10577 21404 10610
rect 21362 10568 21418 10577
rect 21560 10538 21588 11834
rect 21640 11688 21692 11694
rect 21640 11630 21692 11636
rect 21362 10503 21418 10512
rect 21548 10532 21600 10538
rect 21232 9540 21312 9568
rect 21180 9522 21232 9528
rect 21192 6390 21220 9522
rect 21180 6384 21232 6390
rect 21180 6326 21232 6332
rect 21376 5681 21404 10503
rect 21548 10474 21600 10480
rect 21456 9580 21508 9586
rect 21456 9522 21508 9528
rect 21468 8809 21496 9522
rect 21548 9512 21600 9518
rect 21546 9480 21548 9489
rect 21600 9480 21602 9489
rect 21546 9415 21602 9424
rect 21454 8800 21510 8809
rect 21454 8735 21510 8744
rect 21652 7954 21680 11630
rect 21744 9450 21772 12566
rect 22098 12543 22154 12552
rect 22112 12442 22140 12543
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 21824 12164 21876 12170
rect 21824 12106 21876 12112
rect 21836 11529 21864 12106
rect 21822 11520 21878 11529
rect 21822 11455 21878 11464
rect 21824 10668 21876 10674
rect 21928 10656 21956 12378
rect 22100 12232 22152 12238
rect 22100 12174 22152 12180
rect 22008 11620 22060 11626
rect 22008 11562 22060 11568
rect 22020 11286 22048 11562
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 22112 10810 22140 12174
rect 22192 12096 22244 12102
rect 22190 12064 22192 12073
rect 22244 12064 22246 12073
rect 22190 11999 22246 12008
rect 22296 11540 22324 13670
rect 22468 13670 22520 13676
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22374 13631 22430 13640
rect 22388 13462 22416 13631
rect 22376 13456 22428 13462
rect 22376 13398 22428 13404
rect 22376 13252 22428 13258
rect 22376 13194 22428 13200
rect 22388 12730 22416 13194
rect 22480 12850 22508 13670
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22388 12714 22508 12730
rect 22388 12708 22520 12714
rect 22388 12702 22468 12708
rect 22468 12650 22520 12656
rect 22376 12164 22428 12170
rect 22376 12106 22428 12112
rect 22388 11694 22416 12106
rect 22376 11688 22428 11694
rect 22376 11630 22428 11636
rect 22296 11512 22416 11540
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22204 10810 22232 11086
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 21876 10628 21956 10656
rect 22006 10704 22062 10713
rect 22006 10639 22008 10648
rect 21824 10610 21876 10616
rect 22060 10639 22062 10648
rect 22100 10668 22152 10674
rect 22008 10610 22060 10616
rect 22100 10610 22152 10616
rect 21836 10470 21864 10610
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 22112 9674 22140 10610
rect 22204 10606 22232 10746
rect 22296 10606 22324 11018
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 22284 10600 22336 10606
rect 22284 10542 22336 10548
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22192 10192 22244 10198
rect 22192 10134 22244 10140
rect 21836 9646 22140 9674
rect 21732 9444 21784 9450
rect 21732 9386 21784 9392
rect 21836 8378 21864 9646
rect 22204 9586 22232 10134
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 21928 9178 21956 9522
rect 22296 9489 22324 10202
rect 22282 9480 22338 9489
rect 22282 9415 22338 9424
rect 22008 9376 22060 9382
rect 22284 9376 22336 9382
rect 22008 9318 22060 9324
rect 22204 9336 22284 9364
rect 22020 9178 22048 9318
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 22008 9172 22060 9178
rect 22008 9114 22060 9120
rect 22008 8968 22060 8974
rect 22006 8936 22008 8945
rect 22060 8936 22062 8945
rect 22006 8871 22062 8880
rect 21836 8350 21956 8378
rect 21824 8288 21876 8294
rect 21824 8230 21876 8236
rect 21732 8084 21784 8090
rect 21732 8026 21784 8032
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21652 6866 21680 7890
rect 21744 7834 21772 8026
rect 21836 7954 21864 8230
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 21744 7818 21864 7834
rect 21744 7812 21876 7818
rect 21744 7806 21824 7812
rect 21824 7754 21876 7760
rect 21928 7750 21956 8350
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 21640 6860 21692 6866
rect 21640 6802 21692 6808
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 22112 6118 22140 6802
rect 22100 6112 22152 6118
rect 22100 6054 22152 6060
rect 21362 5672 21418 5681
rect 21362 5607 21418 5616
rect 21088 5364 21140 5370
rect 21088 5306 21140 5312
rect 22204 4622 22232 9336
rect 22284 9318 22336 9324
rect 22282 9208 22338 9217
rect 22388 9178 22416 11512
rect 22468 11280 22520 11286
rect 22468 11222 22520 11228
rect 22572 11234 22600 13466
rect 22664 13297 22692 13806
rect 22650 13288 22706 13297
rect 22650 13223 22706 13232
rect 22756 12986 22784 15150
rect 22928 14952 22980 14958
rect 22928 14894 22980 14900
rect 22940 14346 22968 14894
rect 22928 14340 22980 14346
rect 22928 14282 22980 14288
rect 22926 13968 22982 13977
rect 22926 13903 22982 13912
rect 22940 13802 22968 13903
rect 22928 13796 22980 13802
rect 22928 13738 22980 13744
rect 22940 13530 22968 13738
rect 22928 13524 22980 13530
rect 22928 13466 22980 13472
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22664 12617 22692 12718
rect 22650 12608 22706 12617
rect 22650 12543 22706 12552
rect 22756 12238 22784 12922
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22744 12096 22796 12102
rect 22744 12038 22796 12044
rect 22756 11694 22784 12038
rect 22744 11688 22796 11694
rect 22744 11630 22796 11636
rect 22282 9143 22338 9152
rect 22376 9172 22428 9178
rect 22296 8974 22324 9143
rect 22376 9114 22428 9120
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22376 7200 22428 7206
rect 22376 7142 22428 7148
rect 22388 6798 22416 7142
rect 22480 6798 22508 11222
rect 22572 11206 22784 11234
rect 22652 11144 22704 11150
rect 22650 11112 22652 11121
rect 22704 11112 22706 11121
rect 22650 11047 22706 11056
rect 22560 11008 22612 11014
rect 22756 10996 22784 11206
rect 22560 10950 22612 10956
rect 22664 10968 22784 10996
rect 22572 10742 22600 10950
rect 22560 10736 22612 10742
rect 22560 10678 22612 10684
rect 22664 10674 22692 10968
rect 22742 10840 22798 10849
rect 22742 10775 22798 10784
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22560 10532 22612 10538
rect 22560 10474 22612 10480
rect 22572 10062 22600 10474
rect 22650 10296 22706 10305
rect 22650 10231 22706 10240
rect 22664 10130 22692 10231
rect 22652 10124 22704 10130
rect 22652 10066 22704 10072
rect 22560 10056 22612 10062
rect 22560 9998 22612 10004
rect 22756 9602 22784 10775
rect 22848 10062 22876 12582
rect 23032 12306 23060 15286
rect 23124 13870 23152 16934
rect 23216 15502 23244 17054
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23400 16046 23428 16594
rect 23584 16590 23612 18634
rect 23676 17513 23704 19994
rect 23662 17504 23718 17513
rect 23662 17439 23718 17448
rect 23664 16652 23716 16658
rect 23664 16594 23716 16600
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 23478 16280 23534 16289
rect 23478 16215 23480 16224
rect 23532 16215 23534 16224
rect 23480 16186 23532 16192
rect 23388 16040 23440 16046
rect 23388 15982 23440 15988
rect 23492 15910 23520 16186
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 23204 15496 23256 15502
rect 23204 15438 23256 15444
rect 23216 14822 23244 15438
rect 23308 14958 23336 15846
rect 23676 15609 23704 16594
rect 23662 15600 23718 15609
rect 23572 15564 23624 15570
rect 23662 15535 23718 15544
rect 23572 15506 23624 15512
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23388 15088 23440 15094
rect 23388 15030 23440 15036
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 23204 14816 23256 14822
rect 23204 14758 23256 14764
rect 23296 14408 23348 14414
rect 23296 14350 23348 14356
rect 23204 14340 23256 14346
rect 23204 14282 23256 14288
rect 23216 14006 23244 14282
rect 23204 14000 23256 14006
rect 23204 13942 23256 13948
rect 23112 13864 23164 13870
rect 23112 13806 23164 13812
rect 23308 13376 23336 14350
rect 23400 13841 23428 15030
rect 23386 13832 23442 13841
rect 23386 13767 23442 13776
rect 23308 13348 23428 13376
rect 23294 13288 23350 13297
rect 23294 13223 23350 13232
rect 23112 13184 23164 13190
rect 23112 13126 23164 13132
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 22928 11348 22980 11354
rect 22928 11290 22980 11296
rect 22940 10674 22968 11290
rect 23018 11248 23074 11257
rect 23018 11183 23074 11192
rect 22928 10668 22980 10674
rect 22928 10610 22980 10616
rect 23032 10554 23060 11183
rect 23124 11150 23152 13126
rect 23204 12776 23256 12782
rect 23204 12718 23256 12724
rect 23216 12481 23244 12718
rect 23202 12472 23258 12481
rect 23308 12442 23336 13223
rect 23202 12407 23258 12416
rect 23296 12436 23348 12442
rect 23296 12378 23348 12384
rect 23204 12300 23256 12306
rect 23204 12242 23256 12248
rect 23112 11144 23164 11150
rect 23112 11086 23164 11092
rect 22940 10526 23060 10554
rect 22940 10470 22968 10526
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 23020 10464 23072 10470
rect 23020 10406 23072 10412
rect 22940 10130 22968 10406
rect 23032 10305 23060 10406
rect 23018 10296 23074 10305
rect 23018 10231 23074 10240
rect 22928 10124 22980 10130
rect 22928 10066 22980 10072
rect 22836 10056 22888 10062
rect 22836 9998 22888 10004
rect 22664 9574 22784 9602
rect 23020 9580 23072 9586
rect 22560 9376 22612 9382
rect 22558 9344 22560 9353
rect 22612 9344 22614 9353
rect 22558 9279 22614 9288
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22572 8022 22600 8910
rect 22664 8294 22692 9574
rect 23020 9522 23072 9528
rect 22744 9512 22796 9518
rect 22744 9454 22796 9460
rect 22652 8288 22704 8294
rect 22652 8230 22704 8236
rect 22560 8016 22612 8022
rect 22560 7958 22612 7964
rect 22756 7970 22784 9454
rect 22834 8120 22890 8129
rect 22834 8055 22836 8064
rect 22888 8055 22890 8064
rect 22836 8026 22888 8032
rect 22756 7942 22876 7970
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22376 6792 22428 6798
rect 22376 6734 22428 6740
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22572 6458 22600 6734
rect 22652 6656 22704 6662
rect 22652 6598 22704 6604
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22664 6390 22692 6598
rect 22652 6384 22704 6390
rect 22652 6326 22704 6332
rect 22376 6316 22428 6322
rect 22376 6258 22428 6264
rect 22388 5914 22416 6258
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 22756 5409 22784 7822
rect 22742 5400 22798 5409
rect 22742 5335 22798 5344
rect 22468 4752 22520 4758
rect 22468 4694 22520 4700
rect 20812 4616 20864 4622
rect 19708 4558 19760 4564
rect 20718 4584 20774 4593
rect 18512 4480 18564 4486
rect 18512 4422 18564 4428
rect 18524 3534 18552 4422
rect 19720 4282 19748 4558
rect 20812 4558 20864 4564
rect 21180 4616 21232 4622
rect 21180 4558 21232 4564
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 20718 4519 20774 4528
rect 20996 4548 21048 4554
rect 20996 4490 21048 4496
rect 21088 4548 21140 4554
rect 21088 4490 21140 4496
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18800 3670 18828 4082
rect 18788 3664 18840 3670
rect 18788 3606 18840 3612
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 19720 2446 19748 4218
rect 20904 4072 20956 4078
rect 20904 4014 20956 4020
rect 20916 3398 20944 4014
rect 21008 3466 21036 4490
rect 21100 3534 21128 4490
rect 21192 4282 21220 4558
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21180 4276 21232 4282
rect 21180 4218 21232 4224
rect 21376 3534 21404 4422
rect 22480 4146 22508 4694
rect 21916 4140 21968 4146
rect 21916 4082 21968 4088
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 21928 3602 21956 4082
rect 22848 3913 22876 7942
rect 22928 7812 22980 7818
rect 22928 7754 22980 7760
rect 22940 6769 22968 7754
rect 22926 6760 22982 6769
rect 22926 6695 22982 6704
rect 23032 6458 23060 9522
rect 23110 8120 23166 8129
rect 23110 8055 23166 8064
rect 23124 7750 23152 8055
rect 23112 7744 23164 7750
rect 23112 7686 23164 7692
rect 23216 7002 23244 12242
rect 23296 11620 23348 11626
rect 23296 11562 23348 11568
rect 23308 11082 23336 11562
rect 23296 11076 23348 11082
rect 23296 11018 23348 11024
rect 23204 6996 23256 7002
rect 23204 6938 23256 6944
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 23204 6316 23256 6322
rect 23204 6258 23256 6264
rect 23020 6248 23072 6254
rect 23216 6225 23244 6258
rect 23020 6190 23072 6196
rect 23202 6216 23258 6225
rect 23032 5914 23060 6190
rect 23202 6151 23258 6160
rect 23020 5908 23072 5914
rect 23020 5850 23072 5856
rect 23308 5846 23336 11018
rect 23400 10538 23428 13348
rect 23492 12170 23520 15302
rect 23584 15026 23612 15506
rect 23768 15162 23796 21898
rect 23860 21690 23888 23310
rect 24136 22094 24164 23854
rect 24044 22066 24164 22094
rect 23940 22024 23992 22030
rect 23940 21966 23992 21972
rect 23848 21684 23900 21690
rect 23848 21626 23900 21632
rect 23952 21570 23980 21966
rect 23860 21542 23980 21570
rect 23860 21350 23888 21542
rect 24044 21486 24072 22066
rect 24032 21480 24084 21486
rect 24032 21422 24084 21428
rect 23848 21344 23900 21350
rect 23846 21312 23848 21321
rect 23900 21312 23902 21321
rect 23846 21247 23902 21256
rect 24228 20806 24256 24210
rect 24320 21350 24348 24550
rect 24412 21894 24440 29038
rect 24492 28552 24544 28558
rect 24492 28494 24544 28500
rect 24504 24614 24532 28494
rect 25594 28248 25650 28257
rect 25594 28183 25650 28192
rect 25608 28150 25636 28183
rect 25596 28144 25648 28150
rect 25596 28086 25648 28092
rect 24860 28076 24912 28082
rect 24860 28018 24912 28024
rect 25504 28076 25556 28082
rect 25504 28018 25556 28024
rect 24768 28008 24820 28014
rect 24768 27950 24820 27956
rect 24780 27878 24808 27950
rect 24768 27872 24820 27878
rect 24768 27814 24820 27820
rect 24584 25900 24636 25906
rect 24584 25842 24636 25848
rect 24492 24608 24544 24614
rect 24492 24550 24544 24556
rect 24490 24440 24546 24449
rect 24490 24375 24546 24384
rect 24504 23118 24532 24375
rect 24492 23112 24544 23118
rect 24492 23054 24544 23060
rect 24596 22273 24624 25842
rect 24780 25158 24808 27814
rect 24872 26586 24900 28018
rect 25516 27878 25544 28018
rect 25596 27940 25648 27946
rect 25596 27882 25648 27888
rect 25136 27872 25188 27878
rect 25136 27814 25188 27820
rect 25320 27872 25372 27878
rect 25504 27872 25556 27878
rect 25320 27814 25372 27820
rect 25502 27840 25504 27849
rect 25556 27840 25558 27849
rect 24860 26580 24912 26586
rect 24860 26522 24912 26528
rect 25148 25809 25176 27814
rect 25332 27606 25360 27814
rect 25502 27775 25558 27784
rect 25608 27674 25636 27882
rect 25596 27668 25648 27674
rect 25648 27628 25728 27656
rect 25596 27610 25648 27616
rect 25320 27600 25372 27606
rect 25320 27542 25372 27548
rect 25412 26988 25464 26994
rect 25412 26930 25464 26936
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 25228 26784 25280 26790
rect 25228 26726 25280 26732
rect 25134 25800 25190 25809
rect 25134 25735 25190 25744
rect 24952 25696 25004 25702
rect 24952 25638 25004 25644
rect 24860 25492 24912 25498
rect 24860 25434 24912 25440
rect 24768 25152 24820 25158
rect 24768 25094 24820 25100
rect 24676 24132 24728 24138
rect 24676 24074 24728 24080
rect 24688 23769 24716 24074
rect 24674 23760 24730 23769
rect 24674 23695 24730 23704
rect 24676 23316 24728 23322
rect 24676 23258 24728 23264
rect 24582 22264 24638 22273
rect 24582 22199 24638 22208
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24584 21412 24636 21418
rect 24584 21354 24636 21360
rect 24308 21344 24360 21350
rect 24308 21286 24360 21292
rect 24400 21344 24452 21350
rect 24400 21286 24452 21292
rect 24492 21344 24544 21350
rect 24492 21286 24544 21292
rect 24308 21072 24360 21078
rect 24308 21014 24360 21020
rect 24216 20800 24268 20806
rect 24216 20742 24268 20748
rect 23940 20528 23992 20534
rect 23846 20496 23902 20505
rect 23940 20470 23992 20476
rect 23846 20431 23902 20440
rect 23860 19825 23888 20431
rect 23846 19816 23902 19825
rect 23846 19751 23902 19760
rect 23952 19514 23980 20470
rect 24032 20392 24084 20398
rect 24032 20334 24084 20340
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 23940 19168 23992 19174
rect 23940 19110 23992 19116
rect 23848 18760 23900 18766
rect 23848 18702 23900 18708
rect 23860 18426 23888 18702
rect 23848 18420 23900 18426
rect 23848 18362 23900 18368
rect 23848 17264 23900 17270
rect 23848 17206 23900 17212
rect 23860 16998 23888 17206
rect 23848 16992 23900 16998
rect 23952 16969 23980 19110
rect 23848 16934 23900 16940
rect 23938 16960 23994 16969
rect 23860 16794 23888 16934
rect 23938 16895 23994 16904
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 23848 15904 23900 15910
rect 23848 15846 23900 15852
rect 23938 15872 23994 15881
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 23572 15020 23624 15026
rect 23572 14962 23624 14968
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23676 14385 23704 14962
rect 23662 14376 23718 14385
rect 23662 14311 23718 14320
rect 23572 14000 23624 14006
rect 23572 13942 23624 13948
rect 23480 12164 23532 12170
rect 23480 12106 23532 12112
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 23388 10532 23440 10538
rect 23388 10474 23440 10480
rect 23492 10470 23520 11494
rect 23584 10742 23612 13942
rect 23768 12986 23796 14962
rect 23860 14822 23888 15846
rect 23938 15807 23994 15816
rect 23848 14816 23900 14822
rect 23848 14758 23900 14764
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 23676 12442 23704 12718
rect 23756 12640 23808 12646
rect 23756 12582 23808 12588
rect 23664 12436 23716 12442
rect 23664 12378 23716 12384
rect 23768 12306 23796 12582
rect 23756 12300 23808 12306
rect 23756 12242 23808 12248
rect 23664 11348 23716 11354
rect 23664 11290 23716 11296
rect 23572 10736 23624 10742
rect 23572 10678 23624 10684
rect 23572 10600 23624 10606
rect 23572 10542 23624 10548
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 23584 10305 23612 10542
rect 23570 10296 23626 10305
rect 23388 10260 23440 10266
rect 23570 10231 23626 10240
rect 23388 10202 23440 10208
rect 23400 9042 23428 10202
rect 23388 9036 23440 9042
rect 23388 8978 23440 8984
rect 23478 8664 23534 8673
rect 23478 8599 23534 8608
rect 23492 8566 23520 8599
rect 23584 8566 23612 10231
rect 23480 8560 23532 8566
rect 23480 8502 23532 8508
rect 23572 8560 23624 8566
rect 23572 8502 23624 8508
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23400 7449 23428 7482
rect 23386 7440 23442 7449
rect 23676 7410 23704 11290
rect 23756 8288 23808 8294
rect 23754 8256 23756 8265
rect 23808 8256 23810 8265
rect 23754 8191 23810 8200
rect 23386 7375 23442 7384
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 23860 7342 23888 14758
rect 23952 14006 23980 15807
rect 23940 14000 23992 14006
rect 23940 13942 23992 13948
rect 23940 13864 23992 13870
rect 23938 13832 23940 13841
rect 23992 13832 23994 13841
rect 23938 13767 23994 13776
rect 23938 13696 23994 13705
rect 23938 13631 23994 13640
rect 23952 12986 23980 13631
rect 23940 12980 23992 12986
rect 23940 12922 23992 12928
rect 23940 12844 23992 12850
rect 23940 12786 23992 12792
rect 23952 12374 23980 12786
rect 23940 12368 23992 12374
rect 23938 12336 23940 12345
rect 23992 12336 23994 12345
rect 23938 12271 23994 12280
rect 23938 11792 23994 11801
rect 23938 11727 23994 11736
rect 23952 11354 23980 11727
rect 24044 11558 24072 20334
rect 24124 19848 24176 19854
rect 24124 19790 24176 19796
rect 24136 18970 24164 19790
rect 24320 18970 24348 21014
rect 24412 19174 24440 21286
rect 24504 20777 24532 21286
rect 24490 20768 24546 20777
rect 24490 20703 24546 20712
rect 24596 20330 24624 21354
rect 24584 20324 24636 20330
rect 24584 20266 24636 20272
rect 24492 20256 24544 20262
rect 24492 20198 24544 20204
rect 24504 19922 24532 20198
rect 24492 19916 24544 19922
rect 24492 19858 24544 19864
rect 24584 19916 24636 19922
rect 24584 19858 24636 19864
rect 24492 19372 24544 19378
rect 24492 19314 24544 19320
rect 24400 19168 24452 19174
rect 24400 19110 24452 19116
rect 24124 18964 24176 18970
rect 24124 18906 24176 18912
rect 24308 18964 24360 18970
rect 24308 18906 24360 18912
rect 24308 17808 24360 17814
rect 24308 17750 24360 17756
rect 24214 17232 24270 17241
rect 24320 17202 24348 17750
rect 24400 17604 24452 17610
rect 24400 17546 24452 17552
rect 24412 17338 24440 17546
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 24214 17167 24216 17176
rect 24268 17167 24270 17176
rect 24308 17196 24360 17202
rect 24216 17138 24268 17144
rect 24308 17138 24360 17144
rect 24124 17060 24176 17066
rect 24124 17002 24176 17008
rect 24136 13818 24164 17002
rect 24216 16992 24268 16998
rect 24216 16934 24268 16940
rect 24228 13938 24256 16934
rect 24306 16416 24362 16425
rect 24306 16351 24362 16360
rect 24320 16114 24348 16351
rect 24308 16108 24360 16114
rect 24308 16050 24360 16056
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 24320 14521 24348 14554
rect 24306 14512 24362 14521
rect 24306 14447 24362 14456
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24136 13790 24256 13818
rect 24124 13728 24176 13734
rect 24122 13696 24124 13705
rect 24176 13696 24178 13705
rect 24122 13631 24178 13640
rect 24124 13320 24176 13326
rect 24122 13288 24124 13297
rect 24176 13288 24178 13297
rect 24122 13223 24178 13232
rect 24124 12640 24176 12646
rect 24124 12582 24176 12588
rect 24136 11830 24164 12582
rect 24124 11824 24176 11830
rect 24124 11766 24176 11772
rect 24032 11552 24084 11558
rect 24032 11494 24084 11500
rect 23940 11348 23992 11354
rect 23940 11290 23992 11296
rect 24228 11150 24256 13790
rect 24412 13326 24440 17274
rect 24504 16726 24532 19314
rect 24596 18057 24624 19858
rect 24582 18048 24638 18057
rect 24582 17983 24638 17992
rect 24688 16998 24716 23258
rect 24780 22778 24808 25094
rect 24872 24954 24900 25434
rect 24964 25362 24992 25638
rect 24952 25356 25004 25362
rect 24952 25298 25004 25304
rect 24860 24948 24912 24954
rect 24860 24890 24912 24896
rect 24860 24404 24912 24410
rect 24860 24346 24912 24352
rect 24872 23798 24900 24346
rect 24860 23792 24912 23798
rect 24860 23734 24912 23740
rect 24860 23112 24912 23118
rect 24964 23089 24992 25298
rect 25044 25220 25096 25226
rect 25044 25162 25096 25168
rect 25056 23322 25084 25162
rect 25134 25120 25190 25129
rect 25134 25055 25190 25064
rect 25148 24614 25176 25055
rect 25136 24608 25188 24614
rect 25136 24550 25188 24556
rect 25240 24410 25268 26726
rect 25320 26308 25372 26314
rect 25320 26250 25372 26256
rect 25228 24404 25280 24410
rect 25228 24346 25280 24352
rect 25136 24064 25188 24070
rect 25136 24006 25188 24012
rect 25044 23316 25096 23322
rect 25044 23258 25096 23264
rect 25044 23180 25096 23186
rect 25044 23122 25096 23128
rect 24860 23054 24912 23060
rect 24950 23080 25006 23089
rect 24768 22772 24820 22778
rect 24768 22714 24820 22720
rect 24768 21548 24820 21554
rect 24768 21490 24820 21496
rect 24780 20942 24808 21490
rect 24872 21146 24900 23054
rect 24950 23015 25006 23024
rect 25056 22642 25084 23122
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 24952 22228 25004 22234
rect 24952 22170 25004 22176
rect 24860 21140 24912 21146
rect 24860 21082 24912 21088
rect 24768 20936 24820 20942
rect 24768 20878 24820 20884
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24766 20088 24822 20097
rect 24766 20023 24768 20032
rect 24820 20023 24822 20032
rect 24768 19994 24820 20000
rect 24768 19372 24820 19378
rect 24768 19314 24820 19320
rect 24676 16992 24728 16998
rect 24676 16934 24728 16940
rect 24492 16720 24544 16726
rect 24492 16662 24544 16668
rect 24676 15020 24728 15026
rect 24676 14962 24728 14968
rect 24688 14890 24716 14962
rect 24676 14884 24728 14890
rect 24676 14826 24728 14832
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24504 14482 24532 14758
rect 24492 14476 24544 14482
rect 24492 14418 24544 14424
rect 24688 14396 24716 14826
rect 24780 14618 24808 19314
rect 24872 16522 24900 20878
rect 24964 19922 24992 22170
rect 24952 19916 25004 19922
rect 24952 19858 25004 19864
rect 24964 19689 24992 19858
rect 24950 19680 25006 19689
rect 24950 19615 25006 19624
rect 25056 19446 25084 22578
rect 25148 22030 25176 24006
rect 25240 23866 25268 24346
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 25240 22409 25268 22578
rect 25226 22400 25282 22409
rect 25226 22335 25282 22344
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 25134 21448 25190 21457
rect 25134 21383 25190 21392
rect 25044 19440 25096 19446
rect 25044 19382 25096 19388
rect 25044 19304 25096 19310
rect 25044 19246 25096 19252
rect 24950 19136 25006 19145
rect 24950 19071 25006 19080
rect 24860 16516 24912 16522
rect 24860 16458 24912 16464
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 24872 14822 24900 16050
rect 24964 15502 24992 19071
rect 25056 15858 25084 19246
rect 25148 18766 25176 21383
rect 25332 21146 25360 26250
rect 25424 26042 25452 26930
rect 25608 26586 25636 26930
rect 25700 26790 25728 27628
rect 25688 26784 25740 26790
rect 25688 26726 25740 26732
rect 25596 26580 25648 26586
rect 25596 26522 25648 26528
rect 25688 26512 25740 26518
rect 25594 26480 25650 26489
rect 25688 26454 25740 26460
rect 25594 26415 25650 26424
rect 25412 26036 25464 26042
rect 25412 25978 25464 25984
rect 25424 24206 25452 25978
rect 25504 25832 25556 25838
rect 25504 25774 25556 25780
rect 25516 25294 25544 25774
rect 25608 25362 25636 26415
rect 25596 25356 25648 25362
rect 25596 25298 25648 25304
rect 25504 25288 25556 25294
rect 25504 25230 25556 25236
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 25700 24070 25728 26454
rect 25792 25838 25820 29582
rect 25962 28112 26018 28121
rect 25962 28047 26018 28056
rect 25976 27470 26004 28047
rect 26160 27674 26188 30194
rect 26148 27668 26200 27674
rect 26148 27610 26200 27616
rect 26516 27532 26568 27538
rect 26516 27474 26568 27480
rect 25964 27464 26016 27470
rect 25964 27406 26016 27412
rect 25976 26994 26004 27406
rect 25964 26988 26016 26994
rect 25964 26930 26016 26936
rect 25976 26518 26004 26930
rect 26056 26784 26108 26790
rect 26056 26726 26108 26732
rect 25964 26512 26016 26518
rect 25964 26454 26016 26460
rect 25780 25832 25832 25838
rect 25780 25774 25832 25780
rect 25964 25696 26016 25702
rect 25964 25638 26016 25644
rect 25976 25498 26004 25638
rect 25780 25492 25832 25498
rect 25780 25434 25832 25440
rect 25964 25492 26016 25498
rect 25964 25434 26016 25440
rect 25688 24064 25740 24070
rect 25688 24006 25740 24012
rect 25792 23610 25820 25434
rect 25964 24676 26016 24682
rect 25964 24618 26016 24624
rect 25976 23662 26004 24618
rect 26068 23730 26096 26726
rect 26330 26072 26386 26081
rect 26330 26007 26386 26016
rect 26238 25256 26294 25265
rect 26238 25191 26240 25200
rect 26292 25191 26294 25200
rect 26240 25162 26292 25168
rect 26148 25152 26200 25158
rect 26148 25094 26200 25100
rect 26056 23724 26108 23730
rect 26056 23666 26108 23672
rect 25700 23582 25820 23610
rect 25964 23656 26016 23662
rect 25964 23598 26016 23604
rect 25504 23044 25556 23050
rect 25504 22986 25556 22992
rect 25596 23044 25648 23050
rect 25596 22986 25648 22992
rect 25412 22092 25464 22098
rect 25412 22034 25464 22040
rect 25320 21140 25372 21146
rect 25320 21082 25372 21088
rect 25228 19916 25280 19922
rect 25228 19858 25280 19864
rect 25240 19718 25268 19858
rect 25228 19712 25280 19718
rect 25228 19654 25280 19660
rect 25320 19712 25372 19718
rect 25320 19654 25372 19660
rect 25228 19440 25280 19446
rect 25228 19382 25280 19388
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 25148 17678 25176 18702
rect 25136 17672 25188 17678
rect 25136 17614 25188 17620
rect 25134 16824 25190 16833
rect 25134 16759 25190 16768
rect 25148 16522 25176 16759
rect 25136 16516 25188 16522
rect 25136 16458 25188 16464
rect 25240 15881 25268 19382
rect 25226 15872 25282 15881
rect 25056 15830 25176 15858
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24952 14952 25004 14958
rect 24950 14920 24952 14929
rect 25004 14920 25006 14929
rect 24950 14855 25006 14864
rect 24860 14816 24912 14822
rect 24860 14758 24912 14764
rect 24768 14612 24820 14618
rect 24768 14554 24820 14560
rect 24768 14408 24820 14414
rect 24490 14376 24546 14385
rect 24688 14368 24768 14396
rect 24768 14350 24820 14356
rect 24490 14311 24546 14320
rect 24504 14278 24532 14311
rect 24492 14272 24544 14278
rect 24492 14214 24544 14220
rect 24584 13796 24636 13802
rect 24584 13738 24636 13744
rect 24490 13424 24546 13433
rect 24490 13359 24546 13368
rect 24400 13320 24452 13326
rect 24400 13262 24452 13268
rect 24400 12980 24452 12986
rect 24400 12922 24452 12928
rect 24412 12646 24440 12922
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 24400 12436 24452 12442
rect 24400 12378 24452 12384
rect 24216 11144 24268 11150
rect 24214 11112 24216 11121
rect 24268 11112 24270 11121
rect 24214 11047 24270 11056
rect 24032 11008 24084 11014
rect 24032 10950 24084 10956
rect 24306 10976 24362 10985
rect 23938 10840 23994 10849
rect 23938 10775 23994 10784
rect 23952 10742 23980 10775
rect 23940 10736 23992 10742
rect 23940 10678 23992 10684
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23952 8106 23980 8434
rect 24044 8294 24072 10950
rect 24306 10911 24362 10920
rect 24122 10704 24178 10713
rect 24320 10674 24348 10911
rect 24122 10639 24124 10648
rect 24176 10639 24178 10648
rect 24308 10668 24360 10674
rect 24124 10610 24176 10616
rect 24308 10610 24360 10616
rect 24122 10296 24178 10305
rect 24122 10231 24178 10240
rect 24136 9897 24164 10231
rect 24216 10056 24268 10062
rect 24216 9998 24268 10004
rect 24122 9888 24178 9897
rect 24122 9823 24178 9832
rect 24032 8288 24084 8294
rect 24032 8230 24084 8236
rect 23952 8078 24072 8106
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 23572 6656 23624 6662
rect 23572 6598 23624 6604
rect 23388 6112 23440 6118
rect 23388 6054 23440 6060
rect 23296 5840 23348 5846
rect 23296 5782 23348 5788
rect 23400 5710 23428 6054
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 23478 5672 23534 5681
rect 23204 5636 23256 5642
rect 23478 5607 23480 5616
rect 23204 5578 23256 5584
rect 23532 5607 23534 5616
rect 23480 5578 23532 5584
rect 23216 5370 23244 5578
rect 23204 5364 23256 5370
rect 23204 5306 23256 5312
rect 23216 5273 23244 5306
rect 23202 5264 23258 5273
rect 23584 5234 23612 6598
rect 23202 5199 23258 5208
rect 23572 5228 23624 5234
rect 23572 5170 23624 5176
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23940 5228 23992 5234
rect 23940 5170 23992 5176
rect 23768 4622 23796 5170
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23756 4616 23808 4622
rect 23756 4558 23808 4564
rect 23584 3942 23612 4558
rect 23952 4282 23980 5170
rect 23940 4276 23992 4282
rect 23940 4218 23992 4224
rect 23572 3936 23624 3942
rect 22834 3904 22890 3913
rect 23572 3878 23624 3884
rect 22834 3839 22890 3848
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 20996 3460 21048 3466
rect 20996 3402 21048 3408
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 21364 3392 21416 3398
rect 21364 3334 21416 3340
rect 21376 2446 21404 3334
rect 23584 2446 23612 3878
rect 24044 3505 24072 8078
rect 24122 7440 24178 7449
rect 24122 7375 24178 7384
rect 24136 7206 24164 7375
rect 24228 7342 24256 9998
rect 24306 9752 24362 9761
rect 24306 9687 24362 9696
rect 24320 9518 24348 9687
rect 24308 9512 24360 9518
rect 24308 9454 24360 9460
rect 24308 8288 24360 8294
rect 24308 8230 24360 8236
rect 24216 7336 24268 7342
rect 24216 7278 24268 7284
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 24320 6118 24348 8230
rect 24308 6112 24360 6118
rect 24308 6054 24360 6060
rect 24412 5914 24440 12378
rect 24504 12084 24532 13359
rect 24596 13190 24624 13738
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24584 13184 24636 13190
rect 24584 13126 24636 13132
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24688 12714 24716 12922
rect 24766 12880 24822 12889
rect 24872 12850 24900 13330
rect 24766 12815 24768 12824
rect 24820 12815 24822 12824
rect 24860 12844 24912 12850
rect 24768 12786 24820 12792
rect 24860 12786 24912 12792
rect 24676 12708 24728 12714
rect 24676 12650 24728 12656
rect 24688 12434 24716 12650
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 24596 12406 24716 12434
rect 24950 12472 25006 12481
rect 24950 12407 24952 12416
rect 24596 12238 24624 12406
rect 25004 12407 25006 12416
rect 24952 12378 25004 12384
rect 24768 12368 24820 12374
rect 24768 12310 24820 12316
rect 24950 12336 25006 12345
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24504 12056 24624 12084
rect 24492 11552 24544 11558
rect 24492 11494 24544 11500
rect 24504 10130 24532 11494
rect 24596 10674 24624 12056
rect 24780 11558 24808 12310
rect 24950 12271 25006 12280
rect 24860 12232 24912 12238
rect 24860 12174 24912 12180
rect 24872 11898 24900 12174
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24964 11642 24992 12271
rect 25056 11762 25084 12582
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 24964 11614 25084 11642
rect 24768 11552 24820 11558
rect 24768 11494 24820 11500
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24952 10668 25004 10674
rect 24952 10610 25004 10616
rect 24768 10600 24820 10606
rect 24768 10542 24820 10548
rect 24860 10600 24912 10606
rect 24860 10542 24912 10548
rect 24492 10124 24544 10130
rect 24492 10066 24544 10072
rect 24780 9994 24808 10542
rect 24768 9988 24820 9994
rect 24768 9930 24820 9936
rect 24676 9920 24728 9926
rect 24872 9874 24900 10542
rect 24728 9868 24900 9874
rect 24676 9862 24900 9868
rect 24688 9846 24900 9862
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24492 9444 24544 9450
rect 24492 9386 24544 9392
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 24504 5234 24532 9386
rect 24584 8900 24636 8906
rect 24584 8842 24636 8848
rect 24596 8401 24624 8842
rect 24688 8634 24716 9454
rect 24964 8838 24992 10610
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 24766 8664 24822 8673
rect 24676 8628 24728 8634
rect 25056 8650 25084 11614
rect 25148 9450 25176 15830
rect 25226 15807 25282 15816
rect 25228 14476 25280 14482
rect 25228 14418 25280 14424
rect 25240 14346 25268 14418
rect 25228 14340 25280 14346
rect 25228 14282 25280 14288
rect 25240 14074 25268 14282
rect 25228 14068 25280 14074
rect 25228 14010 25280 14016
rect 25332 12434 25360 19654
rect 25424 18086 25452 22034
rect 25516 22001 25544 22986
rect 25502 21992 25558 22001
rect 25502 21927 25558 21936
rect 25504 21344 25556 21350
rect 25504 21286 25556 21292
rect 25412 18080 25464 18086
rect 25412 18022 25464 18028
rect 25424 16794 25452 18022
rect 25412 16788 25464 16794
rect 25412 16730 25464 16736
rect 25412 16516 25464 16522
rect 25412 16458 25464 16464
rect 25424 12481 25452 16458
rect 25516 16130 25544 21286
rect 25608 18057 25636 22986
rect 25700 22098 25728 23582
rect 25780 23520 25832 23526
rect 25780 23462 25832 23468
rect 25792 23322 25820 23462
rect 25780 23316 25832 23322
rect 25780 23258 25832 23264
rect 25792 22778 25820 23258
rect 25976 23118 26004 23598
rect 26056 23180 26108 23186
rect 26056 23122 26108 23128
rect 25964 23112 26016 23118
rect 25964 23054 26016 23060
rect 25780 22772 25832 22778
rect 25780 22714 25832 22720
rect 25688 22092 25740 22098
rect 25688 22034 25740 22040
rect 25872 22092 25924 22098
rect 25872 22034 25924 22040
rect 25686 21992 25742 22001
rect 25686 21927 25688 21936
rect 25740 21927 25742 21936
rect 25688 21898 25740 21904
rect 25594 18048 25650 18057
rect 25594 17983 25650 17992
rect 25516 16102 25636 16130
rect 25502 16008 25558 16017
rect 25502 15943 25558 15952
rect 25516 15910 25544 15943
rect 25504 15904 25556 15910
rect 25504 15846 25556 15852
rect 25504 15496 25556 15502
rect 25504 15438 25556 15444
rect 25240 12406 25360 12434
rect 25410 12472 25466 12481
rect 25410 12407 25466 12416
rect 25136 9444 25188 9450
rect 25136 9386 25188 9392
rect 24766 8599 24768 8608
rect 24676 8570 24728 8576
rect 24820 8599 24822 8608
rect 24964 8622 25084 8650
rect 24768 8570 24820 8576
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 24582 8392 24638 8401
rect 24582 8327 24638 8336
rect 24780 6866 24808 8434
rect 24768 6860 24820 6866
rect 24768 6802 24820 6808
rect 24584 6724 24636 6730
rect 24584 6666 24636 6672
rect 24596 5574 24624 6666
rect 24584 5568 24636 5574
rect 24584 5510 24636 5516
rect 24582 5400 24638 5409
rect 24582 5335 24638 5344
rect 24216 5228 24268 5234
rect 24216 5170 24268 5176
rect 24492 5228 24544 5234
rect 24492 5170 24544 5176
rect 24228 5030 24256 5170
rect 24124 5024 24176 5030
rect 24124 4966 24176 4972
rect 24216 5024 24268 5030
rect 24216 4966 24268 4972
rect 24136 4146 24164 4966
rect 24228 4622 24256 4966
rect 24596 4622 24624 5335
rect 24964 5114 24992 8622
rect 25240 7936 25268 12406
rect 25516 12374 25544 15438
rect 25608 14822 25636 16102
rect 25596 14816 25648 14822
rect 25594 14784 25596 14793
rect 25648 14784 25650 14793
rect 25594 14719 25650 14728
rect 25596 14340 25648 14346
rect 25596 14282 25648 14288
rect 25608 12442 25636 14282
rect 25596 12436 25648 12442
rect 25596 12378 25648 12384
rect 25320 12368 25372 12374
rect 25320 12310 25372 12316
rect 25504 12368 25556 12374
rect 25504 12310 25556 12316
rect 25332 12220 25360 12310
rect 25332 12192 25544 12220
rect 25320 11756 25372 11762
rect 25320 11698 25372 11704
rect 25332 10470 25360 11698
rect 25516 11354 25544 12192
rect 25608 12073 25636 12378
rect 25594 12064 25650 12073
rect 25594 11999 25650 12008
rect 25596 11824 25648 11830
rect 25596 11766 25648 11772
rect 25504 11348 25556 11354
rect 25504 11290 25556 11296
rect 25412 11076 25464 11082
rect 25412 11018 25464 11024
rect 25320 10464 25372 10470
rect 25424 10441 25452 11018
rect 25320 10406 25372 10412
rect 25410 10432 25466 10441
rect 25410 10367 25466 10376
rect 25424 8242 25452 10367
rect 25516 9217 25544 11290
rect 25608 10470 25636 11766
rect 25700 11150 25728 21898
rect 25884 21350 25912 22034
rect 25872 21344 25924 21350
rect 25872 21286 25924 21292
rect 25780 21140 25832 21146
rect 25780 21082 25832 21088
rect 25792 21026 25820 21082
rect 25792 20998 26004 21026
rect 25976 20942 26004 20998
rect 25872 20936 25924 20942
rect 25872 20878 25924 20884
rect 25964 20936 26016 20942
rect 25964 20878 26016 20884
rect 25884 20777 25912 20878
rect 25870 20768 25926 20777
rect 25870 20703 25926 20712
rect 26068 20210 26096 23122
rect 26160 23118 26188 25094
rect 26240 23792 26292 23798
rect 26240 23734 26292 23740
rect 26252 23322 26280 23734
rect 26240 23316 26292 23322
rect 26240 23258 26292 23264
rect 26148 23112 26200 23118
rect 26148 23054 26200 23060
rect 25976 20182 26096 20210
rect 25780 19848 25832 19854
rect 25778 19816 25780 19825
rect 25832 19816 25834 19825
rect 25778 19751 25834 19760
rect 25778 19408 25834 19417
rect 25976 19378 26004 20182
rect 26056 20052 26108 20058
rect 26056 19994 26108 20000
rect 26068 19961 26096 19994
rect 26054 19952 26110 19961
rect 26054 19887 26110 19896
rect 26056 19848 26108 19854
rect 26056 19790 26108 19796
rect 26068 19718 26096 19790
rect 26056 19712 26108 19718
rect 26056 19654 26108 19660
rect 25778 19343 25780 19352
rect 25832 19343 25834 19352
rect 25964 19372 26016 19378
rect 25780 19314 25832 19320
rect 25964 19314 26016 19320
rect 26056 19372 26108 19378
rect 26056 19314 26108 19320
rect 25872 19168 25924 19174
rect 25872 19110 25924 19116
rect 25884 18970 25912 19110
rect 25872 18964 25924 18970
rect 25872 18906 25924 18912
rect 25964 17536 26016 17542
rect 25964 17478 26016 17484
rect 25780 17196 25832 17202
rect 25780 17138 25832 17144
rect 25792 16794 25820 17138
rect 25780 16788 25832 16794
rect 25780 16730 25832 16736
rect 25780 16108 25832 16114
rect 25780 16050 25832 16056
rect 25792 13462 25820 16050
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 25780 13456 25832 13462
rect 25780 13398 25832 13404
rect 25778 13016 25834 13025
rect 25778 12951 25834 12960
rect 25792 12646 25820 12951
rect 25780 12640 25832 12646
rect 25780 12582 25832 12588
rect 25778 12472 25834 12481
rect 25778 12407 25834 12416
rect 25792 12374 25820 12407
rect 25780 12368 25832 12374
rect 25780 12310 25832 12316
rect 25792 11762 25820 12310
rect 25780 11756 25832 11762
rect 25780 11698 25832 11704
rect 25688 11144 25740 11150
rect 25688 11086 25740 11092
rect 25686 10704 25742 10713
rect 25686 10639 25742 10648
rect 25700 10606 25728 10639
rect 25884 10606 25912 15302
rect 25976 14346 26004 17478
rect 26068 15162 26096 19314
rect 26160 18970 26188 23054
rect 26240 23044 26292 23050
rect 26240 22986 26292 22992
rect 26252 22681 26280 22986
rect 26238 22672 26294 22681
rect 26238 22607 26294 22616
rect 26344 22094 26372 26007
rect 26528 25362 26556 27474
rect 26792 27396 26844 27402
rect 26792 27338 26844 27344
rect 26804 25673 26832 27338
rect 26884 27328 26936 27334
rect 26884 27270 26936 27276
rect 26790 25664 26846 25673
rect 26790 25599 26846 25608
rect 26606 25392 26662 25401
rect 26516 25356 26568 25362
rect 26606 25327 26662 25336
rect 26516 25298 26568 25304
rect 26620 25294 26648 25327
rect 26608 25288 26660 25294
rect 26804 25265 26832 25599
rect 26608 25230 26660 25236
rect 26790 25256 26846 25265
rect 26516 25220 26568 25226
rect 26790 25191 26846 25200
rect 26516 25162 26568 25168
rect 26422 23352 26478 23361
rect 26422 23287 26424 23296
rect 26476 23287 26478 23296
rect 26424 23258 26476 23264
rect 26528 23186 26556 25162
rect 26792 25152 26844 25158
rect 26792 25094 26844 25100
rect 26804 24993 26832 25094
rect 26790 24984 26846 24993
rect 26790 24919 26846 24928
rect 26700 24880 26752 24886
rect 26700 24822 26752 24828
rect 26516 23180 26568 23186
rect 26516 23122 26568 23128
rect 26252 22066 26372 22094
rect 26252 19922 26280 22066
rect 26516 21480 26568 21486
rect 26516 21422 26568 21428
rect 26424 21072 26476 21078
rect 26424 21014 26476 21020
rect 26436 20942 26464 21014
rect 26424 20936 26476 20942
rect 26424 20878 26476 20884
rect 26436 20398 26464 20878
rect 26424 20392 26476 20398
rect 26424 20334 26476 20340
rect 26528 20233 26556 21422
rect 26608 21344 26660 21350
rect 26608 21286 26660 21292
rect 26620 20806 26648 21286
rect 26608 20800 26660 20806
rect 26608 20742 26660 20748
rect 26514 20224 26570 20233
rect 26514 20159 26570 20168
rect 26424 20052 26476 20058
rect 26424 19994 26476 20000
rect 26240 19916 26292 19922
rect 26240 19858 26292 19864
rect 26436 19854 26464 19994
rect 26424 19848 26476 19854
rect 26424 19790 26476 19796
rect 26422 19544 26478 19553
rect 26422 19479 26478 19488
rect 26436 19378 26464 19479
rect 26240 19372 26292 19378
rect 26240 19314 26292 19320
rect 26424 19372 26476 19378
rect 26424 19314 26476 19320
rect 26252 19174 26280 19314
rect 26240 19168 26292 19174
rect 26528 19145 26556 20159
rect 26240 19110 26292 19116
rect 26514 19136 26570 19145
rect 26514 19071 26570 19080
rect 26148 18964 26200 18970
rect 26148 18906 26200 18912
rect 26620 18465 26648 20742
rect 26712 20058 26740 24822
rect 26792 24812 26844 24818
rect 26792 24754 26844 24760
rect 26804 20505 26832 24754
rect 26790 20496 26846 20505
rect 26790 20431 26846 20440
rect 26896 20262 26924 27270
rect 26988 26994 27016 30738
rect 32312 30660 32364 30666
rect 32312 30602 32364 30608
rect 28264 30592 28316 30598
rect 28264 30534 28316 30540
rect 27250 29200 27306 29209
rect 27250 29135 27306 29144
rect 27066 27568 27122 27577
rect 27066 27503 27122 27512
rect 26976 26988 27028 26994
rect 26976 26930 27028 26936
rect 27080 26858 27108 27503
rect 27264 26994 27292 29135
rect 27344 27328 27396 27334
rect 27344 27270 27396 27276
rect 27252 26988 27304 26994
rect 27252 26930 27304 26936
rect 27068 26852 27120 26858
rect 27068 26794 27120 26800
rect 26976 26580 27028 26586
rect 26976 26522 27028 26528
rect 26988 26489 27016 26522
rect 26974 26480 27030 26489
rect 26974 26415 26976 26424
rect 27028 26415 27030 26424
rect 26976 26386 27028 26392
rect 27080 26314 27108 26794
rect 27160 26784 27212 26790
rect 27160 26726 27212 26732
rect 27172 26382 27200 26726
rect 27160 26376 27212 26382
rect 27160 26318 27212 26324
rect 27068 26308 27120 26314
rect 27068 26250 27120 26256
rect 27252 26240 27304 26246
rect 27252 26182 27304 26188
rect 27264 25945 27292 26182
rect 27250 25936 27306 25945
rect 27250 25871 27306 25880
rect 27160 23112 27212 23118
rect 27160 23054 27212 23060
rect 27068 22024 27120 22030
rect 27068 21966 27120 21972
rect 26976 21548 27028 21554
rect 26976 21490 27028 21496
rect 26988 21146 27016 21490
rect 27080 21146 27108 21966
rect 27172 21350 27200 23054
rect 27252 21548 27304 21554
rect 27252 21490 27304 21496
rect 27160 21344 27212 21350
rect 27160 21286 27212 21292
rect 26976 21140 27028 21146
rect 26976 21082 27028 21088
rect 27068 21140 27120 21146
rect 27068 21082 27120 21088
rect 26884 20256 26936 20262
rect 26884 20198 26936 20204
rect 26700 20052 26752 20058
rect 26700 19994 26752 20000
rect 26792 20052 26844 20058
rect 26792 19994 26844 20000
rect 26700 19916 26752 19922
rect 26700 19858 26752 19864
rect 26712 19689 26740 19858
rect 26698 19680 26754 19689
rect 26698 19615 26754 19624
rect 26804 19378 26832 19994
rect 26884 19984 26936 19990
rect 26884 19926 26936 19932
rect 26896 19446 26924 19926
rect 26884 19440 26936 19446
rect 26884 19382 26936 19388
rect 26792 19372 26844 19378
rect 27080 19334 27108 21082
rect 27172 20618 27200 21286
rect 27264 20777 27292 21490
rect 27250 20768 27306 20777
rect 27250 20703 27306 20712
rect 27172 20590 27292 20618
rect 26792 19314 26844 19320
rect 26606 18456 26662 18465
rect 26606 18391 26662 18400
rect 26148 18284 26200 18290
rect 26148 18226 26200 18232
rect 26160 17746 26188 18226
rect 26238 18184 26294 18193
rect 26238 18119 26294 18128
rect 26252 17746 26280 18119
rect 26700 18080 26752 18086
rect 26700 18022 26752 18028
rect 26712 17882 26740 18022
rect 26700 17876 26752 17882
rect 26700 17818 26752 17824
rect 26516 17808 26568 17814
rect 26514 17776 26516 17785
rect 26568 17776 26570 17785
rect 26148 17740 26200 17746
rect 26148 17682 26200 17688
rect 26240 17740 26292 17746
rect 26514 17711 26570 17720
rect 26240 17682 26292 17688
rect 26148 17604 26200 17610
rect 26148 17546 26200 17552
rect 26160 17202 26188 17546
rect 26700 17536 26752 17542
rect 26700 17478 26752 17484
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 26712 16590 26740 17478
rect 26700 16584 26752 16590
rect 26700 16526 26752 16532
rect 26424 16108 26476 16114
rect 26424 16050 26476 16056
rect 26332 16040 26384 16046
rect 26332 15982 26384 15988
rect 26056 15156 26108 15162
rect 26056 15098 26108 15104
rect 26056 14952 26108 14958
rect 26056 14894 26108 14900
rect 25964 14340 26016 14346
rect 25964 14282 26016 14288
rect 26068 13444 26096 14894
rect 26240 14340 26292 14346
rect 26240 14282 26292 14288
rect 26252 13938 26280 14282
rect 26240 13932 26292 13938
rect 26240 13874 26292 13880
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26252 13569 26280 13670
rect 26238 13560 26294 13569
rect 26238 13495 26294 13504
rect 26068 13416 26280 13444
rect 26056 13252 26108 13258
rect 26056 13194 26108 13200
rect 26068 12850 26096 13194
rect 26148 12912 26200 12918
rect 26148 12854 26200 12860
rect 26056 12844 26108 12850
rect 26056 12786 26108 12792
rect 25962 12336 26018 12345
rect 25962 12271 25964 12280
rect 26016 12271 26018 12280
rect 25964 12242 26016 12248
rect 25964 12164 26016 12170
rect 25964 12106 26016 12112
rect 25976 11626 26004 12106
rect 25964 11620 26016 11626
rect 25964 11562 26016 11568
rect 25964 11280 26016 11286
rect 25964 11222 26016 11228
rect 25688 10600 25740 10606
rect 25688 10542 25740 10548
rect 25872 10600 25924 10606
rect 25872 10542 25924 10548
rect 25976 10538 26004 11222
rect 26068 10826 26096 12786
rect 26160 12238 26188 12854
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 26252 11354 26280 13416
rect 26344 11393 26372 15982
rect 26436 14090 26464 16050
rect 26804 15978 26832 19314
rect 26988 19306 27108 19334
rect 26884 17196 26936 17202
rect 26884 17138 26936 17144
rect 26896 16658 26924 17138
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 26792 15972 26844 15978
rect 26792 15914 26844 15920
rect 26700 15904 26752 15910
rect 26700 15846 26752 15852
rect 26608 14272 26660 14278
rect 26608 14214 26660 14220
rect 26436 14062 26556 14090
rect 26424 14000 26476 14006
rect 26424 13942 26476 13948
rect 26330 11384 26386 11393
rect 26240 11348 26292 11354
rect 26330 11319 26386 11328
rect 26240 11290 26292 11296
rect 26332 11280 26384 11286
rect 26332 11222 26384 11228
rect 26068 10798 26280 10826
rect 26148 10736 26200 10742
rect 26148 10678 26200 10684
rect 25964 10532 26016 10538
rect 25964 10474 26016 10480
rect 26160 10470 26188 10678
rect 26252 10470 26280 10798
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 26148 10464 26200 10470
rect 26148 10406 26200 10412
rect 26240 10464 26292 10470
rect 26240 10406 26292 10412
rect 25964 9920 26016 9926
rect 25594 9888 25650 9897
rect 25964 9862 26016 9868
rect 25594 9823 25650 9832
rect 25502 9208 25558 9217
rect 25502 9143 25558 9152
rect 25608 8974 25636 9823
rect 25688 9444 25740 9450
rect 25688 9386 25740 9392
rect 25700 9178 25728 9386
rect 25688 9172 25740 9178
rect 25688 9114 25740 9120
rect 25700 8974 25728 9114
rect 25872 9104 25924 9110
rect 25778 9072 25834 9081
rect 25872 9046 25924 9052
rect 25778 9007 25834 9016
rect 25792 8974 25820 9007
rect 25596 8968 25648 8974
rect 25596 8910 25648 8916
rect 25688 8968 25740 8974
rect 25688 8910 25740 8916
rect 25780 8968 25832 8974
rect 25780 8910 25832 8916
rect 25608 8820 25636 8910
rect 25884 8820 25912 9046
rect 25608 8792 25912 8820
rect 25778 8528 25834 8537
rect 25778 8463 25834 8472
rect 25424 8214 25544 8242
rect 25516 7954 25544 8214
rect 25792 8090 25820 8463
rect 25780 8084 25832 8090
rect 25780 8026 25832 8032
rect 25504 7948 25556 7954
rect 25240 7908 25360 7936
rect 25332 6798 25360 7908
rect 25504 7890 25556 7896
rect 25320 6792 25372 6798
rect 25320 6734 25372 6740
rect 25044 6316 25096 6322
rect 25044 6258 25096 6264
rect 25228 6316 25280 6322
rect 25228 6258 25280 6264
rect 25056 5846 25084 6258
rect 25240 6118 25268 6258
rect 25332 6202 25360 6734
rect 25792 6322 25820 8026
rect 25976 7410 26004 9862
rect 26240 9580 26292 9586
rect 26240 9522 26292 9528
rect 26056 9172 26108 9178
rect 26056 9114 26108 9120
rect 26068 8922 26096 9114
rect 26146 9072 26202 9081
rect 26146 9007 26148 9016
rect 26200 9007 26202 9016
rect 26148 8978 26200 8984
rect 26068 8906 26188 8922
rect 26068 8900 26200 8906
rect 26068 8894 26148 8900
rect 26148 8842 26200 8848
rect 26056 7744 26108 7750
rect 26056 7686 26108 7692
rect 25964 7404 26016 7410
rect 25964 7346 26016 7352
rect 26068 7206 26096 7686
rect 26056 7200 26108 7206
rect 26056 7142 26108 7148
rect 26148 6860 26200 6866
rect 26148 6802 26200 6808
rect 25962 6352 26018 6361
rect 25780 6316 25832 6322
rect 25962 6287 25964 6296
rect 25780 6258 25832 6264
rect 26016 6287 26018 6296
rect 25964 6258 26016 6264
rect 25504 6248 25556 6254
rect 25332 6196 25504 6202
rect 25332 6190 25556 6196
rect 25686 6216 25742 6225
rect 25332 6174 25544 6190
rect 25332 6118 25360 6174
rect 25686 6151 25742 6160
rect 25700 6118 25728 6151
rect 25976 6118 26004 6258
rect 25228 6112 25280 6118
rect 25228 6054 25280 6060
rect 25320 6112 25372 6118
rect 25320 6054 25372 6060
rect 25688 6112 25740 6118
rect 25688 6054 25740 6060
rect 25964 6112 26016 6118
rect 25964 6054 26016 6060
rect 25044 5840 25096 5846
rect 25044 5782 25096 5788
rect 25240 5778 25268 6054
rect 25228 5772 25280 5778
rect 25228 5714 25280 5720
rect 24780 5086 24992 5114
rect 25688 5160 25740 5166
rect 25688 5102 25740 5108
rect 24780 5030 24808 5086
rect 24768 5024 24820 5030
rect 24768 4966 24820 4972
rect 24952 5024 25004 5030
rect 24952 4966 25004 4972
rect 24964 4622 24992 4966
rect 24216 4616 24268 4622
rect 24216 4558 24268 4564
rect 24584 4616 24636 4622
rect 24584 4558 24636 4564
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 24952 4616 25004 4622
rect 24952 4558 25004 4564
rect 24872 4146 24900 4558
rect 25700 4486 25728 5102
rect 26160 4554 26188 6802
rect 26252 4826 26280 9522
rect 26344 9382 26372 11222
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 26436 6458 26464 13942
rect 26528 13870 26556 14062
rect 26620 13938 26648 14214
rect 26608 13932 26660 13938
rect 26608 13874 26660 13880
rect 26516 13864 26568 13870
rect 26514 13832 26516 13841
rect 26568 13832 26570 13841
rect 26514 13767 26570 13776
rect 26620 13410 26648 13874
rect 26712 13734 26740 15846
rect 26988 15552 27016 19306
rect 27160 17672 27212 17678
rect 27160 17614 27212 17620
rect 27068 17536 27120 17542
rect 27068 17478 27120 17484
rect 27080 15570 27108 17478
rect 27172 16794 27200 17614
rect 27264 17338 27292 20590
rect 27252 17332 27304 17338
rect 27252 17274 27304 17280
rect 27160 16788 27212 16794
rect 27160 16730 27212 16736
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 26896 15524 27016 15552
rect 27068 15564 27120 15570
rect 26792 14000 26844 14006
rect 26792 13942 26844 13948
rect 26804 13841 26832 13942
rect 26896 13938 26924 15524
rect 27068 15506 27120 15512
rect 26974 15464 27030 15473
rect 26974 15399 26976 15408
rect 27028 15399 27030 15408
rect 26976 15370 27028 15376
rect 27080 14618 27108 15506
rect 27068 14612 27120 14618
rect 27068 14554 27120 14560
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 27068 14408 27120 14414
rect 27068 14350 27120 14356
rect 26988 14074 27016 14350
rect 26976 14068 27028 14074
rect 26976 14010 27028 14016
rect 26884 13932 26936 13938
rect 26884 13874 26936 13880
rect 26790 13832 26846 13841
rect 26790 13767 26846 13776
rect 26976 13796 27028 13802
rect 26976 13738 27028 13744
rect 26700 13728 26752 13734
rect 26884 13728 26936 13734
rect 26700 13670 26752 13676
rect 26804 13688 26884 13716
rect 26528 13382 26648 13410
rect 26528 10062 26556 13382
rect 26608 12640 26660 12646
rect 26608 12582 26660 12588
rect 26620 12442 26648 12582
rect 26608 12436 26660 12442
rect 26804 12434 26832 13688
rect 26884 13670 26936 13676
rect 26884 12776 26936 12782
rect 26884 12718 26936 12724
rect 26896 12442 26924 12718
rect 26608 12378 26660 12384
rect 26712 12406 26832 12434
rect 26884 12436 26936 12442
rect 26608 12164 26660 12170
rect 26608 12106 26660 12112
rect 26620 11150 26648 12106
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 26608 11008 26660 11014
rect 26608 10950 26660 10956
rect 26620 10470 26648 10950
rect 26608 10464 26660 10470
rect 26608 10406 26660 10412
rect 26516 10056 26568 10062
rect 26516 9998 26568 10004
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26528 9110 26556 9318
rect 26608 9172 26660 9178
rect 26712 9160 26740 12406
rect 26884 12378 26936 12384
rect 26988 12322 27016 13738
rect 26896 12294 27016 12322
rect 26792 11552 26844 11558
rect 26792 11494 26844 11500
rect 26804 11354 26832 11494
rect 26792 11348 26844 11354
rect 26792 11290 26844 11296
rect 26792 11144 26844 11150
rect 26792 11086 26844 11092
rect 26804 10810 26832 11086
rect 26792 10804 26844 10810
rect 26792 10746 26844 10752
rect 26790 10704 26846 10713
rect 26790 10639 26792 10648
rect 26844 10639 26846 10648
rect 26792 10610 26844 10616
rect 26790 9480 26846 9489
rect 26790 9415 26846 9424
rect 26660 9132 26740 9160
rect 26608 9114 26660 9120
rect 26516 9104 26568 9110
rect 26516 9046 26568 9052
rect 26606 9072 26662 9081
rect 26804 9042 26832 9415
rect 26606 9007 26662 9016
rect 26792 9036 26844 9042
rect 26620 8974 26648 9007
rect 26792 8978 26844 8984
rect 26608 8968 26660 8974
rect 26608 8910 26660 8916
rect 26896 7886 26924 12294
rect 26976 11076 27028 11082
rect 26976 11018 27028 11024
rect 26988 10606 27016 11018
rect 27080 10810 27108 14350
rect 27172 13734 27200 16594
rect 27264 13938 27292 17274
rect 27356 15502 27384 27270
rect 28276 27130 28304 30534
rect 29000 29572 29052 29578
rect 29000 29514 29052 29520
rect 28264 27124 28316 27130
rect 28264 27066 28316 27072
rect 27436 26784 27488 26790
rect 27436 26726 27488 26732
rect 28356 26784 28408 26790
rect 28356 26726 28408 26732
rect 27448 26586 27476 26726
rect 27710 26616 27766 26625
rect 27436 26580 27488 26586
rect 28368 26586 28396 26726
rect 27710 26551 27766 26560
rect 27896 26580 27948 26586
rect 27436 26522 27488 26528
rect 27724 26382 27752 26551
rect 27896 26522 27948 26528
rect 28356 26580 28408 26586
rect 28356 26522 28408 26528
rect 27908 26450 27936 26522
rect 27896 26444 27948 26450
rect 27896 26386 27948 26392
rect 27712 26376 27764 26382
rect 27712 26318 27764 26324
rect 27436 25356 27488 25362
rect 27436 25298 27488 25304
rect 27448 21078 27476 25298
rect 28262 24848 28318 24857
rect 28080 24812 28132 24818
rect 28080 24754 28132 24760
rect 28172 24812 28224 24818
rect 28262 24783 28264 24792
rect 28172 24754 28224 24760
rect 28316 24783 28318 24792
rect 28264 24754 28316 24760
rect 28092 24410 28120 24754
rect 27896 24404 27948 24410
rect 27896 24346 27948 24352
rect 28080 24404 28132 24410
rect 28080 24346 28132 24352
rect 27712 24064 27764 24070
rect 27712 24006 27764 24012
rect 27804 24064 27856 24070
rect 27804 24006 27856 24012
rect 27620 22636 27672 22642
rect 27620 22578 27672 22584
rect 27632 21690 27660 22578
rect 27620 21684 27672 21690
rect 27620 21626 27672 21632
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 27540 21146 27568 21490
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27528 21140 27580 21146
rect 27528 21082 27580 21088
rect 27436 21072 27488 21078
rect 27436 21014 27488 21020
rect 27436 20936 27488 20942
rect 27434 20904 27436 20913
rect 27488 20904 27490 20913
rect 27434 20839 27490 20848
rect 27436 20256 27488 20262
rect 27436 20198 27488 20204
rect 27344 15496 27396 15502
rect 27344 15438 27396 15444
rect 27252 13932 27304 13938
rect 27252 13874 27304 13880
rect 27160 13728 27212 13734
rect 27160 13670 27212 13676
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 27172 12442 27200 12786
rect 27252 12776 27304 12782
rect 27252 12718 27304 12724
rect 27160 12436 27212 12442
rect 27160 12378 27212 12384
rect 27160 12300 27212 12306
rect 27160 12242 27212 12248
rect 27172 11830 27200 12242
rect 27264 12209 27292 12718
rect 27250 12200 27306 12209
rect 27250 12135 27306 12144
rect 27160 11824 27212 11830
rect 27160 11766 27212 11772
rect 27158 11384 27214 11393
rect 27158 11319 27214 11328
rect 27068 10804 27120 10810
rect 27068 10746 27120 10752
rect 27172 10690 27200 11319
rect 27356 11218 27384 15438
rect 27448 15434 27476 20198
rect 27528 19304 27580 19310
rect 27528 19246 27580 19252
rect 27540 18834 27568 19246
rect 27528 18828 27580 18834
rect 27528 18770 27580 18776
rect 27528 18284 27580 18290
rect 27528 18226 27580 18232
rect 27540 17202 27568 18226
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 27632 16810 27660 21422
rect 27724 18290 27752 24006
rect 27816 23866 27844 24006
rect 27804 23860 27856 23866
rect 27804 23802 27856 23808
rect 27908 23526 27936 24346
rect 27986 24168 28042 24177
rect 27986 24103 28042 24112
rect 28000 23746 28028 24103
rect 28092 23866 28120 24346
rect 28080 23860 28132 23866
rect 28080 23802 28132 23808
rect 28000 23718 28120 23746
rect 27804 23520 27856 23526
rect 27804 23462 27856 23468
rect 27896 23520 27948 23526
rect 27896 23462 27948 23468
rect 27816 22438 27844 23462
rect 27896 22704 27948 22710
rect 27896 22646 27948 22652
rect 27804 22432 27856 22438
rect 27804 22374 27856 22380
rect 27804 21684 27856 21690
rect 27804 21626 27856 21632
rect 27712 18284 27764 18290
rect 27712 18226 27764 18232
rect 27816 17882 27844 21626
rect 27908 20058 27936 22646
rect 27988 22636 28040 22642
rect 27988 22578 28040 22584
rect 28000 21690 28028 22578
rect 27988 21684 28040 21690
rect 27988 21626 28040 21632
rect 27988 21480 28040 21486
rect 27988 21422 28040 21428
rect 28000 21049 28028 21422
rect 27986 21040 28042 21049
rect 27986 20975 28042 20984
rect 27986 20496 28042 20505
rect 27986 20431 28042 20440
rect 27896 20052 27948 20058
rect 27896 19994 27948 20000
rect 28000 19854 28028 20431
rect 27988 19848 28040 19854
rect 27988 19790 28040 19796
rect 28092 19786 28120 23718
rect 28184 23497 28212 24754
rect 28264 24676 28316 24682
rect 28264 24618 28316 24624
rect 28276 24274 28304 24618
rect 28264 24268 28316 24274
rect 28264 24210 28316 24216
rect 28368 24154 28396 26522
rect 28448 26512 28500 26518
rect 28448 26454 28500 26460
rect 28276 24126 28396 24154
rect 28170 23488 28226 23497
rect 28170 23423 28226 23432
rect 28276 21350 28304 24126
rect 28356 23860 28408 23866
rect 28356 23802 28408 23808
rect 28368 21554 28396 23802
rect 28356 21548 28408 21554
rect 28356 21490 28408 21496
rect 28172 21344 28224 21350
rect 28172 21286 28224 21292
rect 28264 21344 28316 21350
rect 28264 21286 28316 21292
rect 28184 21162 28212 21286
rect 28184 21134 28304 21162
rect 28172 19916 28224 19922
rect 28172 19858 28224 19864
rect 28080 19780 28132 19786
rect 28080 19722 28132 19728
rect 28092 19378 28120 19722
rect 28184 19514 28212 19858
rect 28276 19689 28304 21134
rect 28356 20936 28408 20942
rect 28356 20878 28408 20884
rect 28262 19680 28318 19689
rect 28262 19615 28318 19624
rect 28172 19508 28224 19514
rect 28172 19450 28224 19456
rect 28080 19372 28132 19378
rect 28080 19314 28132 19320
rect 27896 19168 27948 19174
rect 27896 19110 27948 19116
rect 27908 18290 27936 19110
rect 28172 18624 28224 18630
rect 28172 18566 28224 18572
rect 27896 18284 27948 18290
rect 27896 18226 27948 18232
rect 27908 18170 27936 18226
rect 27908 18142 28028 18170
rect 27896 18080 27948 18086
rect 27896 18022 27948 18028
rect 27804 17876 27856 17882
rect 27804 17818 27856 17824
rect 27710 17368 27766 17377
rect 27710 17303 27766 17312
rect 27724 17134 27752 17303
rect 27712 17128 27764 17134
rect 27712 17070 27764 17076
rect 27804 17128 27856 17134
rect 27804 17070 27856 17076
rect 27632 16782 27752 16810
rect 27620 16720 27672 16726
rect 27620 16662 27672 16668
rect 27528 16652 27580 16658
rect 27528 16594 27580 16600
rect 27540 16250 27568 16594
rect 27528 16244 27580 16250
rect 27528 16186 27580 16192
rect 27632 16153 27660 16662
rect 27618 16144 27674 16153
rect 27618 16079 27674 16088
rect 27528 15700 27580 15706
rect 27724 15688 27752 16782
rect 27816 16658 27844 17070
rect 27804 16652 27856 16658
rect 27804 16594 27856 16600
rect 27580 15660 27752 15688
rect 27528 15642 27580 15648
rect 27540 15502 27568 15642
rect 27528 15496 27580 15502
rect 27528 15438 27580 15444
rect 27436 15428 27488 15434
rect 27436 15370 27488 15376
rect 27540 15314 27568 15438
rect 27448 15286 27568 15314
rect 27448 14414 27476 15286
rect 27618 15056 27674 15065
rect 27618 14991 27674 15000
rect 27528 14612 27580 14618
rect 27528 14554 27580 14560
rect 27436 14408 27488 14414
rect 27436 14350 27488 14356
rect 27436 14272 27488 14278
rect 27436 14214 27488 14220
rect 27448 14006 27476 14214
rect 27436 14000 27488 14006
rect 27436 13942 27488 13948
rect 27436 13864 27488 13870
rect 27434 13832 27436 13841
rect 27488 13832 27490 13841
rect 27434 13767 27490 13776
rect 27436 13728 27488 13734
rect 27436 13670 27488 13676
rect 27448 12850 27476 13670
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 27344 11212 27396 11218
rect 27344 11154 27396 11160
rect 27540 11098 27568 14554
rect 27632 14482 27660 14991
rect 27804 14544 27856 14550
rect 27804 14486 27856 14492
rect 27620 14476 27672 14482
rect 27620 14418 27672 14424
rect 27710 14376 27766 14385
rect 27620 14340 27672 14346
rect 27710 14311 27712 14320
rect 27620 14282 27672 14288
rect 27764 14311 27766 14320
rect 27712 14282 27764 14288
rect 27632 12434 27660 14282
rect 27816 14006 27844 14486
rect 27804 14000 27856 14006
rect 27804 13942 27856 13948
rect 27712 13728 27764 13734
rect 27712 13670 27764 13676
rect 27724 13190 27752 13670
rect 27816 13326 27844 13942
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 27712 13184 27764 13190
rect 27712 13126 27764 13132
rect 27804 12436 27856 12442
rect 27632 12406 27752 12434
rect 27080 10662 27200 10690
rect 27264 11070 27568 11098
rect 26976 10600 27028 10606
rect 26976 10542 27028 10548
rect 26884 7880 26936 7886
rect 26884 7822 26936 7828
rect 26516 6792 26568 6798
rect 26516 6734 26568 6740
rect 26424 6452 26476 6458
rect 26424 6394 26476 6400
rect 26528 6322 26556 6734
rect 26988 6458 27016 10542
rect 27080 9382 27108 10662
rect 27158 10024 27214 10033
rect 27158 9959 27160 9968
rect 27212 9959 27214 9968
rect 27160 9930 27212 9936
rect 27264 9874 27292 11070
rect 27436 11008 27488 11014
rect 27436 10950 27488 10956
rect 27344 10668 27396 10674
rect 27448 10656 27476 10950
rect 27396 10628 27476 10656
rect 27344 10610 27396 10616
rect 27172 9846 27292 9874
rect 27344 9920 27396 9926
rect 27344 9862 27396 9868
rect 27068 9376 27120 9382
rect 27068 9318 27120 9324
rect 27172 8838 27200 9846
rect 27356 9654 27384 9862
rect 27344 9648 27396 9654
rect 27344 9590 27396 9596
rect 27448 9518 27476 10628
rect 27724 10266 27752 12406
rect 27804 12378 27856 12384
rect 27816 12170 27844 12378
rect 27804 12164 27856 12170
rect 27804 12106 27856 12112
rect 27802 11112 27858 11121
rect 27802 11047 27804 11056
rect 27856 11047 27858 11056
rect 27804 11018 27856 11024
rect 27712 10260 27764 10266
rect 27712 10202 27764 10208
rect 27528 10056 27580 10062
rect 27528 9998 27580 10004
rect 27436 9512 27488 9518
rect 27436 9454 27488 9460
rect 27252 9444 27304 9450
rect 27252 9386 27304 9392
rect 27344 9444 27396 9450
rect 27344 9386 27396 9392
rect 27264 9110 27292 9386
rect 27252 9104 27304 9110
rect 27252 9046 27304 9052
rect 27356 8906 27384 9386
rect 27540 9042 27568 9998
rect 27724 9450 27752 10202
rect 27712 9444 27764 9450
rect 27712 9386 27764 9392
rect 27620 9172 27672 9178
rect 27620 9114 27672 9120
rect 27528 9036 27580 9042
rect 27632 9024 27660 9114
rect 27804 9036 27856 9042
rect 27632 8996 27804 9024
rect 27528 8978 27580 8984
rect 27804 8978 27856 8984
rect 27344 8900 27396 8906
rect 27344 8842 27396 8848
rect 27160 8832 27212 8838
rect 27160 8774 27212 8780
rect 27172 7954 27200 8774
rect 27356 8294 27384 8842
rect 27540 8838 27568 8978
rect 27528 8832 27580 8838
rect 27528 8774 27580 8780
rect 27620 8560 27672 8566
rect 27620 8502 27672 8508
rect 27344 8288 27396 8294
rect 27344 8230 27396 8236
rect 27160 7948 27212 7954
rect 27160 7890 27212 7896
rect 27632 7546 27660 8502
rect 27620 7540 27672 7546
rect 27620 7482 27672 7488
rect 27908 7478 27936 18022
rect 28000 14414 28028 18142
rect 28080 16992 28132 16998
rect 28080 16934 28132 16940
rect 28092 16794 28120 16934
rect 28080 16788 28132 16794
rect 28080 16730 28132 16736
rect 28092 16658 28120 16730
rect 28184 16674 28212 18566
rect 28262 18320 28318 18329
rect 28262 18255 28264 18264
rect 28316 18255 28318 18264
rect 28264 18226 28316 18232
rect 28080 16652 28132 16658
rect 28080 16594 28132 16600
rect 28184 16646 28304 16674
rect 28184 15473 28212 16646
rect 28276 16590 28304 16646
rect 28264 16584 28316 16590
rect 28264 16526 28316 16532
rect 28264 16448 28316 16454
rect 28264 16390 28316 16396
rect 28170 15464 28226 15473
rect 28170 15399 28226 15408
rect 28172 15360 28224 15366
rect 28172 15302 28224 15308
rect 28080 15020 28132 15026
rect 28080 14962 28132 14968
rect 27988 14408 28040 14414
rect 27988 14350 28040 14356
rect 27986 13696 28042 13705
rect 27986 13631 28042 13640
rect 28000 10962 28028 13631
rect 28092 12918 28120 14962
rect 28184 12918 28212 15302
rect 28276 13802 28304 16390
rect 28264 13796 28316 13802
rect 28264 13738 28316 13744
rect 28368 13682 28396 20878
rect 28460 17678 28488 26454
rect 28540 24744 28592 24750
rect 28540 24686 28592 24692
rect 28552 24070 28580 24686
rect 28816 24200 28868 24206
rect 28816 24142 28868 24148
rect 28540 24064 28592 24070
rect 28538 24032 28540 24041
rect 28592 24032 28594 24041
rect 28538 23967 28594 23976
rect 28828 23798 28856 24142
rect 28816 23792 28868 23798
rect 28816 23734 28868 23740
rect 29012 23526 29040 29514
rect 29920 29232 29972 29238
rect 29920 29174 29972 29180
rect 29092 28484 29144 28490
rect 29092 28426 29144 28432
rect 28724 23520 28776 23526
rect 28724 23462 28776 23468
rect 29000 23520 29052 23526
rect 29000 23462 29052 23468
rect 28736 21706 28764 23462
rect 28908 23112 28960 23118
rect 28908 23054 28960 23060
rect 28552 21678 28764 21706
rect 28448 17672 28500 17678
rect 28448 17614 28500 17620
rect 28552 17626 28580 21678
rect 28632 21548 28684 21554
rect 28632 21490 28684 21496
rect 28644 19786 28672 21490
rect 28816 21480 28868 21486
rect 28816 21422 28868 21428
rect 28724 21344 28776 21350
rect 28724 21286 28776 21292
rect 28736 20874 28764 21286
rect 28828 20942 28856 21422
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 28724 20868 28776 20874
rect 28724 20810 28776 20816
rect 28724 20460 28776 20466
rect 28724 20402 28776 20408
rect 28632 19780 28684 19786
rect 28632 19722 28684 19728
rect 28644 19242 28672 19722
rect 28736 19446 28764 20402
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 28724 19440 28776 19446
rect 28724 19382 28776 19388
rect 28632 19236 28684 19242
rect 28632 19178 28684 19184
rect 28828 18601 28856 19790
rect 28814 18592 28870 18601
rect 28814 18527 28870 18536
rect 28920 18426 28948 23054
rect 28998 22808 29054 22817
rect 28998 22743 29054 22752
rect 29012 20058 29040 22743
rect 29000 20052 29052 20058
rect 29000 19994 29052 20000
rect 29000 19712 29052 19718
rect 29000 19654 29052 19660
rect 29012 19378 29040 19654
rect 29000 19372 29052 19378
rect 29000 19314 29052 19320
rect 29000 19236 29052 19242
rect 29000 19178 29052 19184
rect 29012 18766 29040 19178
rect 29000 18760 29052 18766
rect 29000 18702 29052 18708
rect 28908 18420 28960 18426
rect 28908 18362 28960 18368
rect 28998 18048 29054 18057
rect 28998 17983 29054 17992
rect 28908 17672 28960 17678
rect 28552 17598 28856 17626
rect 28908 17614 28960 17620
rect 28632 17536 28684 17542
rect 28684 17484 28764 17490
rect 28632 17478 28764 17484
rect 28644 17462 28764 17478
rect 28448 17196 28500 17202
rect 28448 17138 28500 17144
rect 28540 17196 28592 17202
rect 28540 17138 28592 17144
rect 28460 15366 28488 17138
rect 28552 16794 28580 17138
rect 28736 16794 28764 17462
rect 28540 16788 28592 16794
rect 28540 16730 28592 16736
rect 28724 16788 28776 16794
rect 28724 16730 28776 16736
rect 28632 16448 28684 16454
rect 28632 16390 28684 16396
rect 28540 15428 28592 15434
rect 28540 15370 28592 15376
rect 28448 15360 28500 15366
rect 28448 15302 28500 15308
rect 28448 13796 28500 13802
rect 28448 13738 28500 13744
rect 28276 13654 28396 13682
rect 28080 12912 28132 12918
rect 28080 12854 28132 12860
rect 28172 12912 28224 12918
rect 28172 12854 28224 12860
rect 28092 12442 28120 12854
rect 28276 12764 28304 13654
rect 28356 13524 28408 13530
rect 28356 13466 28408 13472
rect 28184 12736 28304 12764
rect 28080 12436 28132 12442
rect 28080 12378 28132 12384
rect 28080 11756 28132 11762
rect 28080 11698 28132 11704
rect 28092 11354 28120 11698
rect 28080 11348 28132 11354
rect 28080 11290 28132 11296
rect 28000 10934 28120 10962
rect 27986 10840 28042 10849
rect 27986 10775 27988 10784
rect 28040 10775 28042 10784
rect 27988 10746 28040 10752
rect 28000 10062 28028 10746
rect 27988 10056 28040 10062
rect 27988 9998 28040 10004
rect 27896 7472 27948 7478
rect 27896 7414 27948 7420
rect 27802 7304 27858 7313
rect 27802 7239 27858 7248
rect 27816 7206 27844 7239
rect 27804 7200 27856 7206
rect 27804 7142 27856 7148
rect 27908 6662 27936 7414
rect 27896 6656 27948 6662
rect 27896 6598 27948 6604
rect 26976 6452 27028 6458
rect 26976 6394 27028 6400
rect 26516 6316 26568 6322
rect 26516 6258 26568 6264
rect 26240 4820 26292 4826
rect 26240 4762 26292 4768
rect 26148 4548 26200 4554
rect 26148 4490 26200 4496
rect 25688 4480 25740 4486
rect 25688 4422 25740 4428
rect 24124 4140 24176 4146
rect 24124 4082 24176 4088
rect 24860 4140 24912 4146
rect 24860 4082 24912 4088
rect 25228 4072 25280 4078
rect 25228 4014 25280 4020
rect 25240 3942 25268 4014
rect 25228 3936 25280 3942
rect 25228 3878 25280 3884
rect 24030 3496 24086 3505
rect 24030 3431 24086 3440
rect 25700 2446 25728 4422
rect 25872 4072 25924 4078
rect 25872 4014 25924 4020
rect 25884 2446 25912 4014
rect 28092 3126 28120 10934
rect 28184 9178 28212 12736
rect 28264 12300 28316 12306
rect 28264 12242 28316 12248
rect 28276 11218 28304 12242
rect 28264 11212 28316 11218
rect 28264 11154 28316 11160
rect 28264 11008 28316 11014
rect 28264 10950 28316 10956
rect 28276 10674 28304 10950
rect 28368 10810 28396 13466
rect 28460 13326 28488 13738
rect 28552 13326 28580 15370
rect 28644 13530 28672 16390
rect 28632 13524 28684 13530
rect 28632 13466 28684 13472
rect 28448 13320 28500 13326
rect 28448 13262 28500 13268
rect 28540 13320 28592 13326
rect 28540 13262 28592 13268
rect 28448 13184 28500 13190
rect 28448 13126 28500 13132
rect 28460 12594 28488 13126
rect 28644 12782 28672 13466
rect 28632 12776 28684 12782
rect 28632 12718 28684 12724
rect 28460 12566 28580 12594
rect 28446 12472 28502 12481
rect 28446 12407 28502 12416
rect 28460 12186 28488 12407
rect 28552 12306 28580 12566
rect 28540 12300 28592 12306
rect 28540 12242 28592 12248
rect 28460 12158 28580 12186
rect 28448 12096 28500 12102
rect 28448 12038 28500 12044
rect 28460 11558 28488 12038
rect 28552 11830 28580 12158
rect 28630 12064 28686 12073
rect 28630 11999 28686 12008
rect 28540 11824 28592 11830
rect 28540 11766 28592 11772
rect 28448 11552 28500 11558
rect 28448 11494 28500 11500
rect 28448 11212 28500 11218
rect 28448 11154 28500 11160
rect 28356 10804 28408 10810
rect 28356 10746 28408 10752
rect 28264 10668 28316 10674
rect 28264 10610 28316 10616
rect 28368 10130 28396 10746
rect 28356 10124 28408 10130
rect 28356 10066 28408 10072
rect 28356 9376 28408 9382
rect 28356 9318 28408 9324
rect 28172 9172 28224 9178
rect 28172 9114 28224 9120
rect 28184 7478 28212 9114
rect 28368 8974 28396 9318
rect 28356 8968 28408 8974
rect 28356 8910 28408 8916
rect 28172 7472 28224 7478
rect 28172 7414 28224 7420
rect 28460 3194 28488 11154
rect 28552 11150 28580 11766
rect 28644 11762 28672 11999
rect 28736 11762 28764 16730
rect 28828 15502 28856 17598
rect 28920 16658 28948 17614
rect 28908 16652 28960 16658
rect 28908 16594 28960 16600
rect 28816 15496 28868 15502
rect 28868 15456 28948 15484
rect 28816 15438 28868 15444
rect 28816 14340 28868 14346
rect 28816 14282 28868 14288
rect 28828 14074 28856 14282
rect 28816 14068 28868 14074
rect 28816 14010 28868 14016
rect 28920 13410 28948 15456
rect 29012 15201 29040 17983
rect 28998 15192 29054 15201
rect 28998 15127 29054 15136
rect 29000 14816 29052 14822
rect 29000 14758 29052 14764
rect 29012 14482 29040 14758
rect 29000 14476 29052 14482
rect 29000 14418 29052 14424
rect 28828 13382 28948 13410
rect 28828 12866 28856 13382
rect 29104 13376 29132 28426
rect 29736 27668 29788 27674
rect 29736 27610 29788 27616
rect 29366 27160 29422 27169
rect 29366 27095 29422 27104
rect 29276 26376 29328 26382
rect 29276 26318 29328 26324
rect 29184 24608 29236 24614
rect 29184 24550 29236 24556
rect 29196 24206 29224 24550
rect 29184 24200 29236 24206
rect 29184 24142 29236 24148
rect 29184 24064 29236 24070
rect 29184 24006 29236 24012
rect 29196 20330 29224 24006
rect 29184 20324 29236 20330
rect 29184 20266 29236 20272
rect 29184 19780 29236 19786
rect 29184 19722 29236 19728
rect 29196 19378 29224 19722
rect 29184 19372 29236 19378
rect 29184 19314 29236 19320
rect 29196 18766 29224 19314
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 29184 18624 29236 18630
rect 29184 18566 29236 18572
rect 29196 14414 29224 18566
rect 29288 18222 29316 26318
rect 29380 25140 29408 27095
rect 29644 25900 29696 25906
rect 29644 25842 29696 25848
rect 29460 25764 29512 25770
rect 29460 25706 29512 25712
rect 29472 25294 29500 25706
rect 29656 25498 29684 25842
rect 29552 25492 29604 25498
rect 29552 25434 29604 25440
rect 29644 25492 29696 25498
rect 29644 25434 29696 25440
rect 29460 25288 29512 25294
rect 29460 25230 29512 25236
rect 29380 25112 29500 25140
rect 29368 24812 29420 24818
rect 29368 24754 29420 24760
rect 29380 24274 29408 24754
rect 29368 24268 29420 24274
rect 29368 24210 29420 24216
rect 29368 24064 29420 24070
rect 29368 24006 29420 24012
rect 29380 23798 29408 24006
rect 29368 23792 29420 23798
rect 29368 23734 29420 23740
rect 29472 23610 29500 25112
rect 29380 23582 29500 23610
rect 29380 19938 29408 23582
rect 29460 23520 29512 23526
rect 29460 23462 29512 23468
rect 29472 20262 29500 23462
rect 29564 21690 29592 25434
rect 29644 25288 29696 25294
rect 29644 25230 29696 25236
rect 29656 24682 29684 25230
rect 29644 24676 29696 24682
rect 29644 24618 29696 24624
rect 29644 24200 29696 24206
rect 29644 24142 29696 24148
rect 29552 21684 29604 21690
rect 29552 21626 29604 21632
rect 29460 20256 29512 20262
rect 29460 20198 29512 20204
rect 29380 19910 29592 19938
rect 29368 19848 29420 19854
rect 29368 19790 29420 19796
rect 29380 19514 29408 19790
rect 29368 19508 29420 19514
rect 29368 19450 29420 19456
rect 29460 19440 29512 19446
rect 29460 19382 29512 19388
rect 29368 19168 29420 19174
rect 29368 19110 29420 19116
rect 29276 18216 29328 18222
rect 29276 18158 29328 18164
rect 29380 16794 29408 19110
rect 29368 16788 29420 16794
rect 29368 16730 29420 16736
rect 29472 16522 29500 19382
rect 29460 16516 29512 16522
rect 29460 16458 29512 16464
rect 29368 16448 29420 16454
rect 29368 16390 29420 16396
rect 29276 16040 29328 16046
rect 29276 15982 29328 15988
rect 29288 15434 29316 15982
rect 29276 15428 29328 15434
rect 29276 15370 29328 15376
rect 29184 14408 29236 14414
rect 29184 14350 29236 14356
rect 29276 13864 29328 13870
rect 29276 13806 29328 13812
rect 29184 13796 29236 13802
rect 29184 13738 29236 13744
rect 29012 13348 29132 13376
rect 28908 13320 28960 13326
rect 28908 13262 28960 13268
rect 28920 12986 28948 13262
rect 28908 12980 28960 12986
rect 28908 12922 28960 12928
rect 28828 12838 28948 12866
rect 28814 12744 28870 12753
rect 28814 12679 28870 12688
rect 28632 11756 28684 11762
rect 28632 11698 28684 11704
rect 28724 11756 28776 11762
rect 28724 11698 28776 11704
rect 28632 11280 28684 11286
rect 28632 11222 28684 11228
rect 28540 11144 28592 11150
rect 28540 11086 28592 11092
rect 28644 10198 28672 11222
rect 28632 10192 28684 10198
rect 28632 10134 28684 10140
rect 28828 9042 28856 12679
rect 28920 12374 28948 12838
rect 28908 12368 28960 12374
rect 28908 12310 28960 12316
rect 29012 11642 29040 13348
rect 29196 11898 29224 13738
rect 29288 11937 29316 13806
rect 29274 11928 29330 11937
rect 29184 11892 29236 11898
rect 29274 11863 29330 11872
rect 29184 11834 29236 11840
rect 29380 11830 29408 16390
rect 29472 15910 29500 16458
rect 29460 15904 29512 15910
rect 29460 15846 29512 15852
rect 29472 15706 29500 15846
rect 29460 15700 29512 15706
rect 29460 15642 29512 15648
rect 29460 15428 29512 15434
rect 29460 15370 29512 15376
rect 29472 15042 29500 15370
rect 29564 15162 29592 19910
rect 29656 19378 29684 24142
rect 29748 20398 29776 27610
rect 29932 27062 29960 29174
rect 30380 29028 30432 29034
rect 30380 28970 30432 28976
rect 29920 27056 29972 27062
rect 29920 26998 29972 27004
rect 29828 26852 29880 26858
rect 29828 26794 29880 26800
rect 29840 23610 29868 26794
rect 29932 25974 29960 26998
rect 30392 26926 30420 28970
rect 32034 27976 32090 27985
rect 32034 27911 32090 27920
rect 30932 26988 30984 26994
rect 30932 26930 30984 26936
rect 31300 26988 31352 26994
rect 31300 26930 31352 26936
rect 30380 26920 30432 26926
rect 30380 26862 30432 26868
rect 30104 26036 30156 26042
rect 30392 26024 30420 26862
rect 30944 26353 30972 26930
rect 31312 26586 31340 26930
rect 31392 26784 31444 26790
rect 31392 26726 31444 26732
rect 31668 26784 31720 26790
rect 31668 26726 31720 26732
rect 31300 26580 31352 26586
rect 31300 26522 31352 26528
rect 30930 26344 30986 26353
rect 30930 26279 30986 26288
rect 30932 26240 30984 26246
rect 30932 26182 30984 26188
rect 30156 25996 30512 26024
rect 30104 25978 30156 25984
rect 29920 25968 29972 25974
rect 29920 25910 29972 25916
rect 29932 24342 29960 25910
rect 30484 24750 30512 25996
rect 30944 25906 30972 26182
rect 30932 25900 30984 25906
rect 30932 25842 30984 25848
rect 30932 25696 30984 25702
rect 30932 25638 30984 25644
rect 30944 25362 30972 25638
rect 30932 25356 30984 25362
rect 30932 25298 30984 25304
rect 30840 25152 30892 25158
rect 30840 25094 30892 25100
rect 30472 24744 30524 24750
rect 30472 24686 30524 24692
rect 29920 24336 29972 24342
rect 29920 24278 29972 24284
rect 29932 23712 29960 24278
rect 30484 24256 30512 24686
rect 30852 24585 30880 25094
rect 30838 24576 30894 24585
rect 30838 24511 30894 24520
rect 30392 24228 30512 24256
rect 30288 24064 30340 24070
rect 30288 24006 30340 24012
rect 30300 23730 30328 24006
rect 30196 23724 30248 23730
rect 29932 23684 30196 23712
rect 30196 23666 30248 23672
rect 30288 23724 30340 23730
rect 30288 23666 30340 23672
rect 29840 23582 29960 23610
rect 30392 23594 30420 24228
rect 30944 24206 30972 25298
rect 31404 25294 31432 26726
rect 31680 25945 31708 26726
rect 31760 26376 31812 26382
rect 31760 26318 31812 26324
rect 31666 25936 31722 25945
rect 31666 25871 31722 25880
rect 31772 25838 31800 26318
rect 31760 25832 31812 25838
rect 31760 25774 31812 25780
rect 31760 25696 31812 25702
rect 31680 25644 31760 25650
rect 31680 25638 31812 25644
rect 31680 25622 31800 25638
rect 31392 25288 31444 25294
rect 31392 25230 31444 25236
rect 31576 24812 31628 24818
rect 31576 24754 31628 24760
rect 30656 24200 30708 24206
rect 30656 24142 30708 24148
rect 30932 24200 30984 24206
rect 30932 24142 30984 24148
rect 30472 24132 30524 24138
rect 30472 24074 30524 24080
rect 30484 23866 30512 24074
rect 30472 23860 30524 23866
rect 30472 23802 30524 23808
rect 30668 23730 30696 24142
rect 30656 23724 30708 23730
rect 30656 23666 30708 23672
rect 29828 22976 29880 22982
rect 29828 22918 29880 22924
rect 29840 22642 29868 22918
rect 29828 22636 29880 22642
rect 29828 22578 29880 22584
rect 29828 22432 29880 22438
rect 29828 22374 29880 22380
rect 29840 22234 29868 22374
rect 29828 22228 29880 22234
rect 29828 22170 29880 22176
rect 29736 20392 29788 20398
rect 29736 20334 29788 20340
rect 29828 20324 29880 20330
rect 29828 20266 29880 20272
rect 29736 20256 29788 20262
rect 29736 20198 29788 20204
rect 29644 19372 29696 19378
rect 29644 19314 29696 19320
rect 29748 18873 29776 20198
rect 29840 19174 29868 20266
rect 29828 19168 29880 19174
rect 29828 19110 29880 19116
rect 29828 18964 29880 18970
rect 29828 18906 29880 18912
rect 29734 18864 29790 18873
rect 29734 18799 29790 18808
rect 29644 18080 29696 18086
rect 29644 18022 29696 18028
rect 29656 16114 29684 18022
rect 29840 16538 29868 18906
rect 29748 16510 29868 16538
rect 29644 16108 29696 16114
rect 29644 16050 29696 16056
rect 29552 15156 29604 15162
rect 29552 15098 29604 15104
rect 29472 15014 29592 15042
rect 29460 13456 29512 13462
rect 29460 13398 29512 13404
rect 29472 12442 29500 13398
rect 29564 12986 29592 15014
rect 29552 12980 29604 12986
rect 29552 12922 29604 12928
rect 29460 12436 29512 12442
rect 29460 12378 29512 12384
rect 29368 11824 29420 11830
rect 29368 11766 29420 11772
rect 29012 11614 29224 11642
rect 29092 11552 29144 11558
rect 29092 11494 29144 11500
rect 29000 9648 29052 9654
rect 29000 9590 29052 9596
rect 28816 9036 28868 9042
rect 28816 8978 28868 8984
rect 28814 7984 28870 7993
rect 28814 7919 28870 7928
rect 28828 7886 28856 7919
rect 28816 7880 28868 7886
rect 28816 7822 28868 7828
rect 29012 7818 29040 9590
rect 29104 8974 29132 11494
rect 29092 8968 29144 8974
rect 29092 8910 29144 8916
rect 29196 7970 29224 11614
rect 29552 10600 29604 10606
rect 29552 10542 29604 10548
rect 29276 9580 29328 9586
rect 29276 9522 29328 9528
rect 29288 9178 29316 9522
rect 29276 9172 29328 9178
rect 29276 9114 29328 9120
rect 29564 8634 29592 10542
rect 29656 10266 29684 16050
rect 29748 15434 29776 16510
rect 29828 16040 29880 16046
rect 29828 15982 29880 15988
rect 29840 15570 29868 15982
rect 29828 15564 29880 15570
rect 29828 15506 29880 15512
rect 29736 15428 29788 15434
rect 29736 15370 29788 15376
rect 29736 14816 29788 14822
rect 29736 14758 29788 14764
rect 29748 13818 29776 14758
rect 29840 14482 29868 15506
rect 29828 14476 29880 14482
rect 29828 14418 29880 14424
rect 29828 14272 29880 14278
rect 29828 14214 29880 14220
rect 29840 13938 29868 14214
rect 29828 13932 29880 13938
rect 29828 13874 29880 13880
rect 29748 13790 29868 13818
rect 29736 13252 29788 13258
rect 29736 13194 29788 13200
rect 29748 10606 29776 13194
rect 29736 10600 29788 10606
rect 29736 10542 29788 10548
rect 29736 10464 29788 10470
rect 29736 10406 29788 10412
rect 29644 10260 29696 10266
rect 29644 10202 29696 10208
rect 29748 9994 29776 10406
rect 29736 9988 29788 9994
rect 29736 9930 29788 9936
rect 29748 9654 29776 9930
rect 29736 9648 29788 9654
rect 29736 9590 29788 9596
rect 29552 8628 29604 8634
rect 29552 8570 29604 8576
rect 29104 7942 29224 7970
rect 29000 7812 29052 7818
rect 29000 7754 29052 7760
rect 29012 6730 29040 7754
rect 29104 6905 29132 7942
rect 29184 7880 29236 7886
rect 29184 7822 29236 7828
rect 29552 7880 29604 7886
rect 29552 7822 29604 7828
rect 29196 7546 29224 7822
rect 29184 7540 29236 7546
rect 29184 7482 29236 7488
rect 29090 6896 29146 6905
rect 29564 6866 29592 7822
rect 29090 6831 29146 6840
rect 29552 6860 29604 6866
rect 29552 6802 29604 6808
rect 29000 6724 29052 6730
rect 29000 6666 29052 6672
rect 29840 5234 29868 13790
rect 29932 13462 29960 23582
rect 30380 23588 30432 23594
rect 30380 23530 30432 23536
rect 30564 23520 30616 23526
rect 30564 23462 30616 23468
rect 30104 22976 30156 22982
rect 30104 22918 30156 22924
rect 30116 22642 30144 22918
rect 30104 22636 30156 22642
rect 30104 22578 30156 22584
rect 30380 22568 30432 22574
rect 30380 22510 30432 22516
rect 30392 22137 30420 22510
rect 30378 22128 30434 22137
rect 30378 22063 30434 22072
rect 30392 21622 30420 22063
rect 30380 21616 30432 21622
rect 30380 21558 30432 21564
rect 30288 21548 30340 21554
rect 30288 21490 30340 21496
rect 30012 20800 30064 20806
rect 30012 20742 30064 20748
rect 30024 20262 30052 20742
rect 30102 20632 30158 20641
rect 30102 20567 30158 20576
rect 30116 20398 30144 20567
rect 30196 20460 30248 20466
rect 30196 20402 30248 20408
rect 30104 20392 30156 20398
rect 30104 20334 30156 20340
rect 30012 20256 30064 20262
rect 30012 20198 30064 20204
rect 30104 20256 30156 20262
rect 30104 20198 30156 20204
rect 30116 19718 30144 20198
rect 30104 19712 30156 19718
rect 30104 19654 30156 19660
rect 30208 19530 30236 20402
rect 30116 19502 30236 19530
rect 30116 18816 30144 19502
rect 30300 19258 30328 21490
rect 30472 21004 30524 21010
rect 30472 20946 30524 20952
rect 30380 20460 30432 20466
rect 30380 20402 30432 20408
rect 30392 20369 30420 20402
rect 30378 20360 30434 20369
rect 30378 20295 30434 20304
rect 30380 19848 30432 19854
rect 30380 19790 30432 19796
rect 30392 19514 30420 19790
rect 30380 19508 30432 19514
rect 30380 19450 30432 19456
rect 30208 19230 30328 19258
rect 30208 18970 30236 19230
rect 30196 18964 30248 18970
rect 30196 18906 30248 18912
rect 30288 18964 30340 18970
rect 30288 18906 30340 18912
rect 30116 18788 30236 18816
rect 30104 18692 30156 18698
rect 30104 18634 30156 18640
rect 30012 16108 30064 16114
rect 30012 16050 30064 16056
rect 30024 15434 30052 16050
rect 30012 15428 30064 15434
rect 30012 15370 30064 15376
rect 30012 14544 30064 14550
rect 30012 14486 30064 14492
rect 30024 13870 30052 14486
rect 30012 13864 30064 13870
rect 30012 13806 30064 13812
rect 29920 13456 29972 13462
rect 29920 13398 29972 13404
rect 30116 13258 30144 18634
rect 30208 16250 30236 18788
rect 30300 18290 30328 18906
rect 30288 18284 30340 18290
rect 30288 18226 30340 18232
rect 30392 17678 30420 19450
rect 30484 19446 30512 20946
rect 30576 20058 30604 23462
rect 30668 23186 30696 23666
rect 30656 23180 30708 23186
rect 30656 23122 30708 23128
rect 30564 20052 30616 20058
rect 30564 19994 30616 20000
rect 30564 19712 30616 19718
rect 30564 19654 30616 19660
rect 30472 19440 30524 19446
rect 30472 19382 30524 19388
rect 30484 18426 30512 19382
rect 30576 19378 30604 19654
rect 30564 19372 30616 19378
rect 30564 19314 30616 19320
rect 30472 18420 30524 18426
rect 30472 18362 30524 18368
rect 30380 17672 30432 17678
rect 30380 17614 30432 17620
rect 30484 17610 30512 18362
rect 30472 17604 30524 17610
rect 30472 17546 30524 17552
rect 30288 16992 30340 16998
rect 30288 16934 30340 16940
rect 30300 16590 30328 16934
rect 30288 16584 30340 16590
rect 30288 16526 30340 16532
rect 30380 16448 30432 16454
rect 30380 16390 30432 16396
rect 30196 16244 30248 16250
rect 30196 16186 30248 16192
rect 30196 16108 30248 16114
rect 30196 16050 30248 16056
rect 30208 15706 30236 16050
rect 30196 15700 30248 15706
rect 30196 15642 30248 15648
rect 30196 15156 30248 15162
rect 30196 15098 30248 15104
rect 30104 13252 30156 13258
rect 30104 13194 30156 13200
rect 30104 12980 30156 12986
rect 30104 12922 30156 12928
rect 29918 12336 29974 12345
rect 29918 12271 29920 12280
rect 29972 12271 29974 12280
rect 29920 12242 29972 12248
rect 30012 11552 30064 11558
rect 30012 11494 30064 11500
rect 29920 9920 29972 9926
rect 29920 9862 29972 9868
rect 29932 8294 29960 9862
rect 30024 8498 30052 11494
rect 30116 10062 30144 12922
rect 30208 12434 30236 15098
rect 30392 15094 30420 16390
rect 30576 16250 30604 19314
rect 30668 18834 30696 23122
rect 31484 23044 31536 23050
rect 31484 22986 31536 22992
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 30748 22228 30800 22234
rect 30748 22170 30800 22176
rect 30760 22030 30788 22170
rect 30748 22024 30800 22030
rect 30748 21966 30800 21972
rect 30748 21888 30800 21894
rect 30748 21830 30800 21836
rect 30760 21078 30788 21830
rect 30748 21072 30800 21078
rect 30748 21014 30800 21020
rect 30840 21072 30892 21078
rect 30840 21014 30892 21020
rect 30748 20936 30800 20942
rect 30748 20878 30800 20884
rect 30760 20602 30788 20878
rect 30748 20596 30800 20602
rect 30748 20538 30800 20544
rect 30852 20534 30880 21014
rect 30944 20534 30972 22578
rect 31024 22432 31076 22438
rect 31024 22374 31076 22380
rect 31036 21078 31064 22374
rect 31496 22234 31524 22986
rect 31484 22228 31536 22234
rect 31484 22170 31536 22176
rect 31208 21956 31260 21962
rect 31208 21898 31260 21904
rect 31116 21616 31168 21622
rect 31116 21558 31168 21564
rect 31024 21072 31076 21078
rect 31024 21014 31076 21020
rect 31024 20868 31076 20874
rect 31024 20810 31076 20816
rect 30840 20528 30892 20534
rect 30840 20470 30892 20476
rect 30932 20528 30984 20534
rect 30932 20470 30984 20476
rect 30748 20460 30800 20466
rect 30748 20402 30800 20408
rect 30760 19378 30788 20402
rect 30944 20058 30972 20470
rect 30932 20052 30984 20058
rect 30932 19994 30984 20000
rect 31036 19514 31064 20810
rect 31128 19854 31156 21558
rect 31220 20874 31248 21898
rect 31300 21548 31352 21554
rect 31300 21490 31352 21496
rect 31312 21146 31340 21490
rect 31300 21140 31352 21146
rect 31300 21082 31352 21088
rect 31208 20868 31260 20874
rect 31208 20810 31260 20816
rect 31208 20256 31260 20262
rect 31208 20198 31260 20204
rect 31220 19854 31248 20198
rect 31298 20088 31354 20097
rect 31298 20023 31354 20032
rect 31116 19848 31168 19854
rect 31116 19790 31168 19796
rect 31208 19848 31260 19854
rect 31208 19790 31260 19796
rect 31024 19508 31076 19514
rect 31024 19450 31076 19456
rect 30748 19372 30800 19378
rect 30748 19314 30800 19320
rect 30930 18864 30986 18873
rect 30656 18828 30708 18834
rect 30930 18799 30986 18808
rect 30656 18770 30708 18776
rect 30668 18290 30696 18770
rect 30944 18766 30972 18799
rect 30932 18760 30984 18766
rect 30932 18702 30984 18708
rect 30656 18284 30708 18290
rect 30656 18226 30708 18232
rect 30668 17202 30696 18226
rect 31036 17882 31064 19450
rect 31024 17876 31076 17882
rect 31024 17818 31076 17824
rect 31036 17678 31064 17818
rect 30932 17672 30984 17678
rect 30932 17614 30984 17620
rect 31024 17672 31076 17678
rect 31024 17614 31076 17620
rect 30944 17338 30972 17614
rect 30932 17332 30984 17338
rect 30932 17274 30984 17280
rect 30656 17196 30708 17202
rect 30656 17138 30708 17144
rect 30564 16244 30616 16250
rect 30564 16186 30616 16192
rect 30576 16114 30604 16186
rect 30564 16108 30616 16114
rect 30564 16050 30616 16056
rect 30564 15972 30616 15978
rect 30564 15914 30616 15920
rect 30472 15904 30524 15910
rect 30472 15846 30524 15852
rect 30380 15088 30432 15094
rect 30300 15036 30380 15042
rect 30300 15030 30432 15036
rect 30300 15014 30420 15030
rect 30300 14618 30328 15014
rect 30380 14952 30432 14958
rect 30380 14894 30432 14900
rect 30288 14612 30340 14618
rect 30288 14554 30340 14560
rect 30288 14272 30340 14278
rect 30288 14214 30340 14220
rect 30300 13938 30328 14214
rect 30288 13932 30340 13938
rect 30288 13874 30340 13880
rect 30392 13530 30420 14894
rect 30484 14822 30512 15846
rect 30576 15706 30604 15914
rect 30564 15700 30616 15706
rect 30564 15642 30616 15648
rect 30668 15570 30696 17138
rect 30932 16516 30984 16522
rect 30932 16458 30984 16464
rect 30748 16176 30800 16182
rect 30748 16118 30800 16124
rect 30656 15564 30708 15570
rect 30656 15506 30708 15512
rect 30564 15360 30616 15366
rect 30564 15302 30616 15308
rect 30472 14816 30524 14822
rect 30472 14758 30524 14764
rect 30576 14618 30604 15302
rect 30656 14816 30708 14822
rect 30656 14758 30708 14764
rect 30564 14612 30616 14618
rect 30564 14554 30616 14560
rect 30576 13954 30604 14554
rect 30668 14464 30696 14758
rect 30760 14618 30788 16118
rect 30840 16108 30892 16114
rect 30840 16050 30892 16056
rect 30852 15178 30880 16050
rect 30944 15366 30972 16458
rect 30932 15360 30984 15366
rect 30932 15302 30984 15308
rect 30852 15150 30972 15178
rect 30840 15020 30892 15026
rect 30840 14962 30892 14968
rect 30852 14822 30880 14962
rect 30840 14816 30892 14822
rect 30838 14784 30840 14793
rect 30892 14784 30894 14793
rect 30838 14719 30894 14728
rect 30944 14618 30972 15150
rect 31022 15056 31078 15065
rect 31022 14991 31024 15000
rect 31076 14991 31078 15000
rect 31024 14962 31076 14968
rect 30748 14612 30800 14618
rect 30748 14554 30800 14560
rect 30932 14612 30984 14618
rect 30932 14554 30984 14560
rect 30668 14436 30880 14464
rect 30852 14396 30880 14436
rect 30932 14408 30984 14414
rect 30852 14368 30932 14396
rect 30932 14350 30984 14356
rect 31024 14272 31076 14278
rect 31024 14214 31076 14220
rect 30932 14068 30984 14074
rect 30932 14010 30984 14016
rect 30576 13926 30696 13954
rect 30564 13864 30616 13870
rect 30564 13806 30616 13812
rect 30380 13524 30432 13530
rect 30380 13466 30432 13472
rect 30576 13394 30604 13806
rect 30564 13388 30616 13394
rect 30564 13330 30616 13336
rect 30288 13320 30340 13326
rect 30288 13262 30340 13268
rect 30300 12850 30328 13262
rect 30576 12918 30604 13330
rect 30668 13258 30696 13926
rect 30944 13326 30972 14010
rect 30932 13320 30984 13326
rect 30932 13262 30984 13268
rect 30656 13252 30708 13258
rect 30656 13194 30708 13200
rect 30840 13252 30892 13258
rect 30840 13194 30892 13200
rect 30564 12912 30616 12918
rect 30564 12854 30616 12860
rect 30288 12844 30340 12850
rect 30288 12786 30340 12792
rect 30208 12406 30328 12434
rect 30196 11144 30248 11150
rect 30196 11086 30248 11092
rect 30208 10742 30236 11086
rect 30196 10736 30248 10742
rect 30196 10678 30248 10684
rect 30104 10056 30156 10062
rect 30104 9998 30156 10004
rect 30012 8492 30064 8498
rect 30012 8434 30064 8440
rect 30104 8356 30156 8362
rect 30104 8298 30156 8304
rect 29920 8288 29972 8294
rect 29920 8230 29972 8236
rect 30116 6798 30144 8298
rect 30300 7585 30328 12406
rect 30380 12164 30432 12170
rect 30380 12106 30432 12112
rect 30392 11150 30420 12106
rect 30472 12096 30524 12102
rect 30472 12038 30524 12044
rect 30484 11626 30512 12038
rect 30576 11694 30604 12854
rect 30656 12844 30708 12850
rect 30656 12786 30708 12792
rect 30668 12102 30696 12786
rect 30852 12170 30880 13194
rect 30932 12640 30984 12646
rect 30932 12582 30984 12588
rect 30944 12238 30972 12582
rect 30932 12232 30984 12238
rect 30932 12174 30984 12180
rect 30840 12164 30892 12170
rect 30840 12106 30892 12112
rect 30656 12096 30708 12102
rect 30656 12038 30708 12044
rect 30564 11688 30616 11694
rect 30564 11630 30616 11636
rect 30472 11620 30524 11626
rect 30472 11562 30524 11568
rect 30840 11552 30892 11558
rect 30840 11494 30892 11500
rect 30852 11150 30880 11494
rect 30380 11144 30432 11150
rect 30380 11086 30432 11092
rect 30564 11144 30616 11150
rect 30564 11086 30616 11092
rect 30840 11144 30892 11150
rect 30840 11086 30892 11092
rect 30576 10810 30604 11086
rect 30564 10804 30616 10810
rect 30564 10746 30616 10752
rect 30472 10668 30524 10674
rect 30392 10628 30472 10656
rect 30286 7576 30342 7585
rect 30286 7511 30342 7520
rect 30104 6792 30156 6798
rect 30104 6734 30156 6740
rect 30392 5302 30420 10628
rect 30472 10610 30524 10616
rect 30564 10464 30616 10470
rect 30564 10406 30616 10412
rect 30472 9988 30524 9994
rect 30472 9930 30524 9936
rect 30484 9722 30512 9930
rect 30472 9716 30524 9722
rect 30472 9658 30524 9664
rect 30484 7750 30512 9658
rect 30576 8566 30604 10406
rect 30656 9988 30708 9994
rect 30656 9930 30708 9936
rect 30668 9654 30696 9930
rect 30748 9920 30800 9926
rect 30748 9862 30800 9868
rect 30656 9648 30708 9654
rect 30656 9590 30708 9596
rect 30760 8906 30788 9862
rect 30852 9382 30880 11086
rect 31036 10674 31064 14214
rect 31024 10668 31076 10674
rect 31024 10610 31076 10616
rect 31128 9466 31156 19790
rect 31208 19168 31260 19174
rect 31208 19110 31260 19116
rect 31220 18766 31248 19110
rect 31208 18760 31260 18766
rect 31208 18702 31260 18708
rect 31208 15904 31260 15910
rect 31208 15846 31260 15852
rect 31220 15502 31248 15846
rect 31208 15496 31260 15502
rect 31208 15438 31260 15444
rect 31208 15088 31260 15094
rect 31208 15030 31260 15036
rect 31220 13326 31248 15030
rect 31208 13320 31260 13326
rect 31208 13262 31260 13268
rect 31220 12850 31248 13262
rect 31208 12844 31260 12850
rect 31208 12786 31260 12792
rect 31208 12164 31260 12170
rect 31208 12106 31260 12112
rect 31220 11082 31248 12106
rect 31208 11076 31260 11082
rect 31208 11018 31260 11024
rect 31036 9438 31156 9466
rect 30840 9376 30892 9382
rect 30840 9318 30892 9324
rect 30748 8900 30800 8906
rect 30748 8842 30800 8848
rect 30564 8560 30616 8566
rect 30564 8502 30616 8508
rect 30472 7744 30524 7750
rect 30472 7686 30524 7692
rect 30748 7744 30800 7750
rect 30748 7686 30800 7692
rect 30932 7744 30984 7750
rect 30932 7686 30984 7692
rect 30760 6798 30788 7686
rect 30944 7342 30972 7686
rect 30932 7336 30984 7342
rect 30932 7278 30984 7284
rect 30840 7200 30892 7206
rect 30840 7142 30892 7148
rect 30852 6798 30880 7142
rect 30748 6792 30800 6798
rect 30748 6734 30800 6740
rect 30840 6792 30892 6798
rect 30840 6734 30892 6740
rect 30380 5296 30432 5302
rect 30380 5238 30432 5244
rect 29828 5228 29880 5234
rect 29828 5170 29880 5176
rect 31036 4010 31064 9438
rect 31116 9376 31168 9382
rect 31116 9318 31168 9324
rect 31128 8974 31156 9318
rect 31116 8968 31168 8974
rect 31116 8910 31168 8916
rect 31128 7886 31156 8910
rect 31312 8378 31340 20023
rect 31588 19334 31616 24754
rect 31680 23905 31708 25622
rect 31852 25220 31904 25226
rect 31852 25162 31904 25168
rect 31864 24818 31892 25162
rect 31942 25120 31998 25129
rect 31942 25055 31998 25064
rect 31852 24812 31904 24818
rect 31852 24754 31904 24760
rect 31666 23896 31722 23905
rect 31864 23866 31892 24754
rect 31666 23831 31722 23840
rect 31852 23860 31904 23866
rect 31852 23802 31904 23808
rect 31760 23112 31812 23118
rect 31760 23054 31812 23060
rect 31772 22438 31800 23054
rect 31760 22432 31812 22438
rect 31760 22374 31812 22380
rect 31772 20466 31800 22374
rect 31852 20936 31904 20942
rect 31852 20878 31904 20884
rect 31760 20460 31812 20466
rect 31760 20402 31812 20408
rect 31404 19306 31616 19334
rect 31404 18630 31432 19306
rect 31864 18970 31892 20878
rect 31852 18964 31904 18970
rect 31852 18906 31904 18912
rect 31392 18624 31444 18630
rect 31392 18566 31444 18572
rect 31392 18284 31444 18290
rect 31392 18226 31444 18232
rect 31404 17882 31432 18226
rect 31392 17876 31444 17882
rect 31392 17818 31444 17824
rect 31576 17196 31628 17202
rect 31576 17138 31628 17144
rect 31588 16794 31616 17138
rect 31576 16788 31628 16794
rect 31576 16730 31628 16736
rect 31760 16244 31812 16250
rect 31760 16186 31812 16192
rect 31392 14816 31444 14822
rect 31392 14758 31444 14764
rect 31404 14414 31432 14758
rect 31772 14482 31800 16186
rect 31760 14476 31812 14482
rect 31760 14418 31812 14424
rect 31392 14408 31444 14414
rect 31392 14350 31444 14356
rect 31668 14408 31720 14414
rect 31668 14350 31720 14356
rect 31404 10742 31432 14350
rect 31680 12986 31708 14350
rect 31852 14272 31904 14278
rect 31852 14214 31904 14220
rect 31760 13932 31812 13938
rect 31760 13874 31812 13880
rect 31772 13530 31800 13874
rect 31760 13524 31812 13530
rect 31760 13466 31812 13472
rect 31668 12980 31720 12986
rect 31668 12922 31720 12928
rect 31484 12096 31536 12102
rect 31484 12038 31536 12044
rect 31496 11830 31524 12038
rect 31484 11824 31536 11830
rect 31484 11766 31536 11772
rect 31392 10736 31444 10742
rect 31392 10678 31444 10684
rect 31484 10668 31536 10674
rect 31484 10610 31536 10616
rect 31496 10062 31524 10610
rect 31576 10464 31628 10470
rect 31576 10406 31628 10412
rect 31588 10062 31616 10406
rect 31484 10056 31536 10062
rect 31484 9998 31536 10004
rect 31576 10056 31628 10062
rect 31864 10010 31892 14214
rect 31576 9998 31628 10004
rect 31496 9722 31524 9998
rect 31484 9716 31536 9722
rect 31484 9658 31536 9664
rect 31312 8350 31432 8378
rect 31208 8288 31260 8294
rect 31208 8230 31260 8236
rect 31300 8288 31352 8294
rect 31300 8230 31352 8236
rect 31220 7886 31248 8230
rect 31312 8090 31340 8230
rect 31300 8084 31352 8090
rect 31300 8026 31352 8032
rect 31116 7880 31168 7886
rect 31116 7822 31168 7828
rect 31208 7880 31260 7886
rect 31208 7822 31260 7828
rect 31024 4004 31076 4010
rect 31024 3946 31076 3952
rect 31404 3738 31432 8350
rect 31588 5370 31616 9998
rect 31772 9982 31892 10010
rect 31772 8294 31800 9982
rect 31852 9920 31904 9926
rect 31852 9862 31904 9868
rect 31864 9586 31892 9862
rect 31852 9580 31904 9586
rect 31852 9522 31904 9528
rect 31864 8566 31892 9522
rect 31852 8560 31904 8566
rect 31852 8502 31904 8508
rect 31760 8288 31812 8294
rect 31760 8230 31812 8236
rect 31666 7576 31722 7585
rect 31666 7511 31722 7520
rect 31680 6458 31708 7511
rect 31956 6914 31984 25055
rect 32048 11529 32076 27911
rect 32128 25900 32180 25906
rect 32128 25842 32180 25848
rect 32140 24274 32168 25842
rect 32220 25764 32272 25770
rect 32220 25706 32272 25712
rect 32232 24818 32260 25706
rect 32220 24812 32272 24818
rect 32220 24754 32272 24760
rect 32128 24268 32180 24274
rect 32128 24210 32180 24216
rect 32220 22636 32272 22642
rect 32220 22578 32272 22584
rect 32232 21690 32260 22578
rect 32220 21684 32272 21690
rect 32220 21626 32272 21632
rect 32128 21548 32180 21554
rect 32128 21490 32180 21496
rect 32140 20398 32168 21490
rect 32232 21010 32260 21626
rect 32220 21004 32272 21010
rect 32220 20946 32272 20952
rect 32128 20392 32180 20398
rect 32128 20334 32180 20340
rect 32126 19408 32182 19417
rect 32126 19343 32182 19352
rect 32220 19372 32272 19378
rect 32140 14278 32168 19343
rect 32220 19314 32272 19320
rect 32232 18426 32260 19314
rect 32220 18420 32272 18426
rect 32220 18362 32272 18368
rect 32232 17746 32260 18362
rect 32220 17740 32272 17746
rect 32220 17682 32272 17688
rect 32324 17626 32352 30602
rect 32496 26988 32548 26994
rect 32496 26930 32548 26936
rect 32508 26382 32536 26930
rect 32496 26376 32548 26382
rect 32496 26318 32548 26324
rect 32508 25498 32536 26318
rect 32496 25492 32548 25498
rect 32496 25434 32548 25440
rect 32496 24608 32548 24614
rect 32496 24550 32548 24556
rect 32404 23520 32456 23526
rect 32404 23462 32456 23468
rect 32416 22545 32444 23462
rect 32508 23225 32536 24550
rect 32588 23724 32640 23730
rect 32588 23666 32640 23672
rect 32494 23216 32550 23225
rect 32494 23151 32550 23160
rect 32600 22982 32628 23666
rect 32680 23316 32732 23322
rect 32680 23258 32732 23264
rect 32588 22976 32640 22982
rect 32588 22918 32640 22924
rect 32402 22536 32458 22545
rect 32402 22471 32458 22480
rect 32496 22432 32548 22438
rect 32496 22374 32548 22380
rect 32404 21344 32456 21350
rect 32404 21286 32456 21292
rect 32416 20505 32444 21286
rect 32508 21185 32536 22374
rect 32600 22098 32628 22918
rect 32588 22092 32640 22098
rect 32588 22034 32640 22040
rect 32692 21978 32720 23258
rect 32600 21950 32720 21978
rect 32494 21176 32550 21185
rect 32494 21111 32550 21120
rect 32402 20496 32458 20505
rect 32402 20431 32458 20440
rect 32496 20392 32548 20398
rect 32496 20334 32548 20340
rect 32404 20256 32456 20262
rect 32404 20198 32456 20204
rect 32416 19825 32444 20198
rect 32508 20058 32536 20334
rect 32496 20052 32548 20058
rect 32496 19994 32548 20000
rect 32402 19816 32458 19825
rect 32402 19751 32458 19760
rect 32404 19508 32456 19514
rect 32404 19450 32456 19456
rect 32416 19145 32444 19450
rect 32402 19136 32458 19145
rect 32402 19071 32458 19080
rect 32404 18080 32456 18086
rect 32404 18022 32456 18028
rect 32416 17785 32444 18022
rect 32402 17776 32458 17785
rect 32402 17711 32458 17720
rect 32232 17598 32352 17626
rect 32232 16266 32260 17598
rect 32312 17196 32364 17202
rect 32312 17138 32364 17144
rect 32324 16658 32352 17138
rect 32402 17096 32458 17105
rect 32402 17031 32404 17040
rect 32456 17031 32458 17040
rect 32404 17002 32456 17008
rect 32312 16652 32364 16658
rect 32312 16594 32364 16600
rect 32232 16238 32352 16266
rect 32220 16108 32272 16114
rect 32220 16050 32272 16056
rect 32232 15706 32260 16050
rect 32220 15700 32272 15706
rect 32220 15642 32272 15648
rect 32220 15020 32272 15026
rect 32220 14962 32272 14968
rect 32128 14272 32180 14278
rect 32128 14214 32180 14220
rect 32232 14074 32260 14962
rect 32220 14068 32272 14074
rect 32220 14010 32272 14016
rect 32128 13932 32180 13938
rect 32128 13874 32180 13880
rect 32034 11520 32090 11529
rect 32034 11455 32090 11464
rect 32140 11354 32168 13874
rect 32232 13394 32260 14010
rect 32220 13388 32272 13394
rect 32220 13330 32272 13336
rect 32220 12232 32272 12238
rect 32220 12174 32272 12180
rect 32232 11898 32260 12174
rect 32220 11892 32272 11898
rect 32220 11834 32272 11840
rect 32232 11762 32260 11834
rect 32220 11756 32272 11762
rect 32220 11698 32272 11704
rect 32128 11348 32180 11354
rect 32128 11290 32180 11296
rect 32140 10606 32168 11290
rect 32128 10600 32180 10606
rect 32128 10542 32180 10548
rect 32324 9738 32352 16238
rect 32404 15904 32456 15910
rect 32404 15846 32456 15852
rect 32416 15745 32444 15846
rect 32402 15736 32458 15745
rect 32402 15671 32458 15680
rect 32404 15156 32456 15162
rect 32404 15098 32456 15104
rect 32416 15065 32444 15098
rect 32402 15056 32458 15065
rect 32402 14991 32458 15000
rect 32404 14068 32456 14074
rect 32404 14010 32456 14016
rect 32416 13705 32444 14010
rect 32402 13696 32458 13705
rect 32402 13631 32458 13640
rect 32494 13016 32550 13025
rect 32494 12951 32550 12960
rect 32508 12850 32536 12951
rect 32496 12844 32548 12850
rect 32496 12786 32548 12792
rect 32402 11656 32458 11665
rect 32402 11591 32404 11600
rect 32456 11591 32458 11600
rect 32404 11562 32456 11568
rect 32404 10464 32456 10470
rect 32600 10441 32628 21950
rect 32678 17232 32734 17241
rect 32678 17167 32734 17176
rect 32404 10406 32456 10412
rect 32586 10432 32642 10441
rect 32416 10305 32444 10406
rect 32586 10367 32642 10376
rect 32402 10296 32458 10305
rect 32402 10231 32458 10240
rect 32496 10056 32548 10062
rect 32496 9998 32548 10004
rect 32140 9710 32352 9738
rect 32140 9625 32168 9710
rect 32126 9616 32182 9625
rect 32126 9551 32182 9560
rect 32310 9616 32366 9625
rect 32508 9586 32536 9998
rect 32310 9551 32366 9560
rect 32496 9580 32548 9586
rect 32324 9450 32352 9551
rect 32496 9522 32548 9528
rect 32312 9444 32364 9450
rect 32312 9386 32364 9392
rect 32508 9178 32536 9522
rect 32496 9172 32548 9178
rect 32496 9114 32548 9120
rect 32220 8492 32272 8498
rect 32220 8434 32272 8440
rect 32232 8090 32260 8434
rect 32404 8356 32456 8362
rect 32404 8298 32456 8304
rect 32416 8265 32444 8298
rect 32402 8256 32458 8265
rect 32402 8191 32458 8200
rect 32220 8084 32272 8090
rect 32220 8026 32272 8032
rect 32496 7404 32548 7410
rect 32496 7346 32548 7352
rect 32220 7336 32272 7342
rect 32220 7278 32272 7284
rect 31772 6886 31984 6914
rect 31668 6452 31720 6458
rect 31668 6394 31720 6400
rect 31772 5710 31800 6886
rect 32232 6322 32260 7278
rect 32312 7200 32364 7206
rect 32312 7142 32364 7148
rect 32324 6905 32352 7142
rect 32508 7002 32536 7346
rect 32496 6996 32548 7002
rect 32496 6938 32548 6944
rect 32310 6896 32366 6905
rect 32310 6831 32366 6840
rect 32220 6316 32272 6322
rect 32220 6258 32272 6264
rect 31760 5704 31812 5710
rect 31760 5646 31812 5652
rect 32692 5545 32720 17167
rect 32678 5536 32734 5545
rect 32678 5471 32734 5480
rect 31576 5364 31628 5370
rect 31576 5306 31628 5312
rect 31392 3732 31444 3738
rect 31392 3674 31444 3680
rect 28448 3188 28500 3194
rect 28448 3130 28500 3136
rect 28080 3120 28132 3126
rect 28080 3062 28132 3068
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 19708 2440 19760 2446
rect 19708 2382 19760 2388
rect 21364 2440 21416 2446
rect 21364 2382 21416 2388
rect 23572 2440 23624 2446
rect 23572 2382 23624 2388
rect 25688 2440 25740 2446
rect 25688 2382 25740 2388
rect 25872 2440 25924 2446
rect 25872 2382 25924 2388
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 17420 800 17448 2246
rect 19352 800 19380 2246
rect 21284 800 21312 2246
rect 22572 800 22600 2246
rect 24504 800 24532 2246
rect 25792 800 25820 2246
rect 29656 800 29684 2382
rect 17406 0 17462 800
rect 19338 0 19394 800
rect 21270 0 21326 800
rect 22558 0 22614 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 29642 0 29698 800
<< via2 >>
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 13726 30776 13782 30832
rect 1122 30232 1178 30288
rect 846 25744 902 25800
rect 386 24656 442 24712
rect 754 24112 810 24168
rect 478 23160 534 23216
rect 570 20848 626 20904
rect 662 14048 718 14104
rect 846 23976 902 24032
rect 846 18808 902 18864
rect 1030 20712 1086 20768
rect 938 17584 994 17640
rect 846 16532 848 16552
rect 848 16532 900 16552
rect 900 16532 902 16552
rect 846 16496 902 16532
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 6826 30368 6882 30424
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 1398 28600 1454 28656
rect 1490 27920 1546 27976
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 3330 28364 3332 28384
rect 3332 28364 3384 28384
rect 3384 28364 3386 28384
rect 3330 28328 3386 28364
rect 2594 26868 2596 26888
rect 2596 26868 2648 26888
rect 2648 26868 2650 26888
rect 2594 26832 2650 26868
rect 2134 25744 2190 25800
rect 3698 28872 3754 28928
rect 4250 28960 4306 29008
rect 4250 28952 4252 28960
rect 4252 28952 4304 28960
rect 4304 28952 4306 28960
rect 1766 25064 1822 25120
rect 1398 21548 1454 21584
rect 1398 21528 1400 21548
rect 1400 21528 1452 21548
rect 1452 21528 1454 21548
rect 1306 19080 1362 19136
rect 1122 15408 1178 15464
rect 846 14456 902 14512
rect 938 10784 994 10840
rect 386 7928 442 7984
rect 1858 19624 1914 19680
rect 2226 20576 2282 20632
rect 3698 27548 3700 27568
rect 3700 27548 3752 27568
rect 3752 27548 3754 27568
rect 3698 27512 3754 27548
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4618 28056 4674 28112
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4710 26988 4766 27024
rect 4710 26968 4712 26988
rect 4712 26968 4764 26988
rect 4764 26968 4766 26988
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 5354 27104 5410 27160
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4986 25900 5042 25936
rect 4986 25880 4988 25900
rect 4988 25880 5040 25900
rect 5040 25880 5042 25900
rect 5354 26152 5410 26208
rect 3146 23568 3202 23624
rect 3146 22480 3202 22536
rect 3514 23568 3570 23624
rect 5078 25608 5134 25664
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4342 24792 4398 24848
rect 3882 23704 3938 23760
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 5262 24248 5318 24304
rect 5538 27240 5594 27296
rect 5630 27104 5686 27160
rect 5538 26424 5594 26480
rect 5722 26188 5724 26208
rect 5724 26188 5776 26208
rect 5776 26188 5778 26208
rect 5722 26152 5778 26188
rect 6734 28328 6790 28384
rect 5906 26016 5962 26072
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 3514 21664 3570 21720
rect 3422 20984 3478 21040
rect 3330 20440 3386 20496
rect 2502 19760 2558 19816
rect 2042 16224 2098 16280
rect 2870 19488 2926 19544
rect 2686 17196 2742 17232
rect 2686 17176 2688 17196
rect 2688 17176 2740 17196
rect 2740 17176 2742 17196
rect 3790 21392 3846 21448
rect 3514 18672 3570 18728
rect 3146 17176 3202 17232
rect 3054 16360 3110 16416
rect 2778 15952 2834 16008
rect 2502 15272 2558 15328
rect 1398 10920 1454 10976
rect 2318 13368 2374 13424
rect 2226 11092 2228 11112
rect 2228 11092 2280 11112
rect 2280 11092 2282 11112
rect 2226 11056 2282 11092
rect 2318 5616 2374 5672
rect 2042 5072 2098 5128
rect 3054 15408 3110 15464
rect 3054 15156 3110 15192
rect 3054 15136 3056 15156
rect 3056 15136 3108 15156
rect 3108 15136 3110 15156
rect 3238 15952 3294 16008
rect 3054 13776 3110 13832
rect 3146 13232 3202 13288
rect 3146 13096 3202 13152
rect 2962 12144 3018 12200
rect 2502 9016 2558 9072
rect 2870 11228 2872 11248
rect 2872 11228 2924 11248
rect 2924 11228 2926 11248
rect 2870 11192 2926 11228
rect 2870 11092 2872 11112
rect 2872 11092 2924 11112
rect 2924 11092 2926 11112
rect 2870 11056 2926 11092
rect 3790 20748 3792 20768
rect 3792 20748 3844 20768
rect 3844 20748 3846 20768
rect 3790 20712 3846 20748
rect 4342 21936 4398 21992
rect 4066 21800 4122 21856
rect 4526 22072 4582 22128
rect 4526 21836 4528 21856
rect 4528 21836 4580 21856
rect 4580 21836 4582 21856
rect 4526 21800 4582 21836
rect 3790 20440 3846 20496
rect 4250 21392 4306 21448
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4250 20984 4306 21040
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 3422 17856 3478 17912
rect 4066 19624 4122 19680
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 5906 25608 5962 25664
rect 6182 26560 6238 26616
rect 6090 26152 6146 26208
rect 5722 23976 5778 24032
rect 4986 23160 5042 23216
rect 4894 23024 4950 23080
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 5354 22888 5410 22944
rect 5354 22752 5410 22808
rect 4710 22208 4766 22264
rect 4710 20576 4766 20632
rect 5078 22480 5134 22536
rect 4986 22344 5042 22400
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 5538 23432 5594 23488
rect 5722 22480 5778 22536
rect 5538 21936 5594 21992
rect 5354 21392 5410 21448
rect 4894 21140 4950 21176
rect 4894 21120 4896 21140
rect 4896 21120 4948 21140
rect 4948 21120 4950 21140
rect 5446 20884 5448 20904
rect 5448 20884 5500 20904
rect 5500 20884 5502 20904
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4802 20304 4858 20360
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4710 19488 4766 19544
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 3882 17060 3938 17096
rect 3882 17040 3884 17060
rect 3884 17040 3936 17060
rect 3936 17040 3938 17060
rect 3882 16496 3938 16552
rect 3882 15544 3938 15600
rect 4802 17720 4858 17776
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4342 16496 4398 16552
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 5170 17040 5226 17096
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4434 15544 4490 15600
rect 3882 14456 3938 14512
rect 3790 14320 3846 14376
rect 4434 15272 4490 15328
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 5170 15816 5226 15872
rect 5446 20848 5502 20884
rect 5722 20440 5778 20496
rect 5538 19080 5594 19136
rect 5354 18672 5410 18728
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 3606 12844 3662 12880
rect 3606 12824 3608 12844
rect 3608 12824 3660 12844
rect 3660 12824 3662 12844
rect 3790 12960 3846 13016
rect 4710 14612 4766 14648
rect 4710 14592 4712 14612
rect 4712 14592 4764 14612
rect 4764 14592 4766 14612
rect 4894 14764 4896 14784
rect 4896 14764 4948 14784
rect 4948 14764 4950 14784
rect 4894 14728 4950 14764
rect 4250 14320 4306 14376
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4434 13388 4490 13424
rect 4434 13368 4436 13388
rect 4436 13368 4488 13388
rect 4488 13368 4490 13388
rect 4342 13268 4344 13288
rect 4344 13268 4396 13288
rect 4396 13268 4398 13288
rect 4342 13232 4398 13268
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4894 13812 4896 13832
rect 4896 13812 4948 13832
rect 4948 13812 4950 13832
rect 4894 13776 4950 13812
rect 4802 13504 4858 13560
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4342 11892 4398 11928
rect 4342 11872 4344 11892
rect 4344 11872 4396 11892
rect 4396 11872 4398 11892
rect 4710 12960 4766 13016
rect 4894 13252 4950 13288
rect 4894 13232 4896 13252
rect 4896 13232 4948 13252
rect 4948 13232 4950 13252
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 5630 18400 5686 18456
rect 5538 16360 5594 16416
rect 5906 24112 5962 24168
rect 5998 23976 6054 24032
rect 5906 23432 5962 23488
rect 5906 23024 5962 23080
rect 5906 22208 5962 22264
rect 5906 22108 5908 22128
rect 5908 22108 5960 22128
rect 5960 22108 5962 22128
rect 5906 22072 5962 22108
rect 6090 23296 6146 23352
rect 6090 22752 6146 22808
rect 6734 27648 6790 27704
rect 6918 28736 6974 28792
rect 7470 29552 7526 29608
rect 7194 28500 7196 28520
rect 7196 28500 7248 28520
rect 7248 28500 7250 28520
rect 7194 28464 7250 28500
rect 7194 28364 7196 28384
rect 7196 28364 7248 28384
rect 7248 28364 7250 28384
rect 7194 28328 7250 28364
rect 7010 27512 7066 27568
rect 6826 27376 6882 27432
rect 7470 27784 7526 27840
rect 6826 27104 6882 27160
rect 6366 26832 6422 26888
rect 7194 27376 7250 27432
rect 7010 27240 7066 27296
rect 6642 26188 6644 26208
rect 6644 26188 6696 26208
rect 6696 26188 6698 26208
rect 6642 26152 6698 26188
rect 6366 23724 6422 23760
rect 6366 23704 6368 23724
rect 6368 23704 6420 23724
rect 6420 23704 6422 23724
rect 6366 23588 6422 23624
rect 6366 23568 6368 23588
rect 6368 23568 6420 23588
rect 6420 23568 6422 23588
rect 6182 21664 6238 21720
rect 6090 21256 6146 21312
rect 5906 21120 5962 21176
rect 5998 20304 6054 20360
rect 6826 25064 6882 25120
rect 6550 23976 6606 24032
rect 6550 22752 6606 22808
rect 7102 25780 7104 25800
rect 7104 25780 7156 25800
rect 7156 25780 7158 25800
rect 7102 25744 7158 25780
rect 7746 27920 7802 27976
rect 8022 27648 8078 27704
rect 7930 27276 7932 27296
rect 7932 27276 7984 27296
rect 7984 27276 7986 27296
rect 7930 27240 7986 27276
rect 7746 26016 7802 26072
rect 7378 23296 7434 23352
rect 6918 23060 6920 23080
rect 6920 23060 6972 23080
rect 6972 23060 6974 23080
rect 6918 23024 6974 23060
rect 6918 22752 6974 22808
rect 6550 22208 6606 22264
rect 6274 20848 6330 20904
rect 7286 23180 7342 23216
rect 7286 23160 7288 23180
rect 7288 23160 7340 23180
rect 7340 23160 7342 23180
rect 7194 22888 7250 22944
rect 6642 20304 6698 20360
rect 6550 18808 6606 18864
rect 5630 15680 5686 15736
rect 5446 14864 5502 14920
rect 5354 13776 5410 13832
rect 5078 12708 5134 12744
rect 5722 14900 5724 14920
rect 5724 14900 5776 14920
rect 5776 14900 5778 14920
rect 5722 14864 5778 14900
rect 5630 14456 5686 14512
rect 5906 15136 5962 15192
rect 5722 14320 5778 14376
rect 6458 17856 6514 17912
rect 6826 20440 6882 20496
rect 6642 17312 6698 17368
rect 6642 17196 6698 17232
rect 6642 17176 6644 17196
rect 6644 17176 6696 17196
rect 6696 17176 6698 17196
rect 5722 14068 5778 14104
rect 5722 14048 5724 14068
rect 5724 14048 5776 14068
rect 5776 14048 5778 14068
rect 5538 13096 5594 13152
rect 5078 12688 5080 12708
rect 5080 12688 5132 12708
rect 5132 12688 5134 12708
rect 5262 12588 5264 12608
rect 5264 12588 5316 12608
rect 5316 12588 5318 12608
rect 5262 12552 5318 12588
rect 5262 12416 5318 12472
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4158 11600 4214 11656
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 5170 11464 5226 11520
rect 4434 10648 4490 10704
rect 5354 11328 5410 11384
rect 4710 10784 4766 10840
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4802 10376 4858 10432
rect 4710 10240 4766 10296
rect 4158 10004 4160 10024
rect 4160 10004 4212 10024
rect 4212 10004 4214 10024
rect 4158 9968 4214 10004
rect 4434 9560 4490 9616
rect 3882 9424 3938 9480
rect 4986 10104 5042 10160
rect 5354 10920 5410 10976
rect 5354 10140 5356 10160
rect 5356 10140 5408 10160
rect 5408 10140 5410 10160
rect 5354 10104 5410 10140
rect 5538 12688 5594 12744
rect 5722 12280 5778 12336
rect 7010 18944 7066 19000
rect 7010 18808 7066 18864
rect 6826 16904 6882 16960
rect 6734 16108 6790 16144
rect 6734 16088 6736 16108
rect 6736 16088 6788 16108
rect 6788 16088 6790 16108
rect 6734 15700 6790 15736
rect 6734 15680 6736 15700
rect 6736 15680 6788 15700
rect 6788 15680 6790 15700
rect 6642 15544 6698 15600
rect 6550 15272 6606 15328
rect 6182 12824 6238 12880
rect 6090 12416 6146 12472
rect 5722 12008 5778 12064
rect 5630 11892 5686 11928
rect 5630 11872 5632 11892
rect 5632 11872 5684 11892
rect 5684 11872 5686 11892
rect 5630 11756 5686 11792
rect 5630 11736 5632 11756
rect 5632 11736 5684 11756
rect 5684 11736 5686 11756
rect 5630 11092 5632 11112
rect 5632 11092 5684 11112
rect 5684 11092 5686 11112
rect 5630 11056 5686 11092
rect 5998 11328 6054 11384
rect 5906 10920 5962 10976
rect 5538 10784 5594 10840
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3790 7384 3846 7440
rect 4894 9288 4950 9344
rect 5078 8880 5134 8936
rect 5814 9696 5870 9752
rect 6458 12824 6514 12880
rect 6826 14492 6828 14512
rect 6828 14492 6880 14512
rect 6880 14492 6882 14512
rect 6826 14456 6882 14492
rect 6734 13132 6736 13152
rect 6736 13132 6788 13152
rect 6788 13132 6790 13152
rect 6734 13096 6790 13132
rect 6642 12552 6698 12608
rect 6826 12824 6882 12880
rect 6826 12708 6882 12744
rect 6826 12688 6828 12708
rect 6828 12688 6880 12708
rect 6880 12688 6882 12708
rect 7010 15952 7066 16008
rect 7010 15000 7066 15056
rect 7654 23296 7710 23352
rect 7562 23060 7564 23080
rect 7564 23060 7616 23080
rect 7616 23060 7618 23080
rect 7562 23024 7618 23060
rect 7654 22344 7710 22400
rect 7562 19932 7564 19952
rect 7564 19932 7616 19952
rect 7616 19932 7618 19952
rect 7562 19896 7618 19932
rect 7562 19352 7618 19408
rect 7470 18572 7472 18592
rect 7472 18572 7524 18592
rect 7524 18572 7526 18592
rect 7470 18536 7526 18572
rect 7470 17992 7526 18048
rect 7838 23160 7894 23216
rect 9126 29144 9182 29200
rect 9678 29688 9734 29744
rect 8482 26732 8484 26752
rect 8484 26732 8536 26752
rect 8536 26732 8538 26752
rect 8482 26696 8538 26732
rect 8574 26152 8630 26208
rect 8206 25064 8262 25120
rect 8114 24792 8170 24848
rect 8666 25200 8722 25256
rect 9862 29008 9918 29064
rect 9402 28872 9458 28928
rect 9126 27940 9182 27976
rect 9126 27920 9128 27940
rect 9128 27920 9180 27940
rect 9180 27920 9182 27940
rect 9126 27276 9128 27296
rect 9128 27276 9180 27296
rect 9180 27276 9182 27296
rect 9126 27240 9182 27276
rect 9586 28328 9642 28384
rect 10138 28328 10194 28384
rect 9586 26560 9642 26616
rect 9770 26560 9826 26616
rect 8114 22888 8170 22944
rect 7930 20984 7986 21040
rect 7838 20712 7894 20768
rect 7654 18572 7656 18592
rect 7656 18572 7708 18592
rect 7708 18572 7710 18592
rect 7654 18536 7710 18572
rect 7746 18284 7802 18320
rect 7930 20032 7986 20088
rect 7746 18264 7748 18284
rect 7748 18264 7800 18284
rect 7800 18264 7802 18284
rect 7746 17992 7802 18048
rect 7194 16088 7250 16144
rect 7378 16496 7434 16552
rect 7286 15000 7342 15056
rect 7194 14592 7250 14648
rect 7470 14728 7526 14784
rect 7378 14048 7434 14104
rect 7286 13404 7288 13424
rect 7288 13404 7340 13424
rect 7340 13404 7342 13424
rect 7286 13368 7342 13404
rect 7194 13096 7250 13152
rect 6550 11872 6606 11928
rect 6734 11872 6790 11928
rect 6458 11620 6514 11656
rect 6458 11600 6460 11620
rect 6460 11600 6512 11620
rect 6512 11600 6514 11620
rect 6366 11092 6368 11112
rect 6368 11092 6420 11112
rect 6420 11092 6422 11112
rect 6366 11056 6422 11092
rect 6366 10920 6422 10976
rect 5262 8744 5318 8800
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4802 8472 4858 8528
rect 4986 8472 5042 8528
rect 4618 8200 4674 8256
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4250 7404 4306 7440
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4250 7384 4252 7404
rect 4252 7384 4304 7404
rect 4304 7384 4306 7404
rect 4986 7404 5042 7440
rect 4986 7384 4988 7404
rect 4988 7384 5040 7404
rect 5040 7384 5042 7404
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 5446 8336 5502 8392
rect 6090 9152 6146 9208
rect 5814 8336 5870 8392
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 6090 8200 6146 8256
rect 6274 9696 6330 9752
rect 6642 11192 6698 11248
rect 6642 10920 6698 10976
rect 6918 12280 6974 12336
rect 7010 11892 7066 11928
rect 7010 11872 7012 11892
rect 7012 11872 7064 11892
rect 7064 11872 7066 11892
rect 7010 11600 7066 11656
rect 7010 11464 7066 11520
rect 8298 22480 8354 22536
rect 8206 19760 8262 19816
rect 8666 24520 8722 24576
rect 9034 24384 9090 24440
rect 8850 24248 8906 24304
rect 9218 24792 9274 24848
rect 9586 25372 9588 25392
rect 9588 25372 9640 25392
rect 9640 25372 9642 25392
rect 9586 25336 9642 25372
rect 10138 27784 10194 27840
rect 10230 27648 10286 27704
rect 10230 27240 10286 27296
rect 9402 25064 9458 25120
rect 9494 24556 9496 24576
rect 9496 24556 9548 24576
rect 9548 24556 9550 24576
rect 9494 24520 9550 24556
rect 9034 23024 9090 23080
rect 8666 21972 8668 21992
rect 8668 21972 8720 21992
rect 8720 21972 8722 21992
rect 8666 21936 8722 21972
rect 8574 21120 8630 21176
rect 8942 21800 8998 21856
rect 8942 20712 8998 20768
rect 8942 20576 8998 20632
rect 8298 17040 8354 17096
rect 7746 16496 7802 16552
rect 8022 15952 8078 16008
rect 7654 14048 7710 14104
rect 7746 13948 7748 13968
rect 7748 13948 7800 13968
rect 7800 13948 7802 13968
rect 7746 13912 7802 13948
rect 7654 13812 7656 13832
rect 7656 13812 7708 13832
rect 7708 13812 7710 13832
rect 7654 13776 7710 13812
rect 7930 14592 7986 14648
rect 7838 12688 7894 12744
rect 7654 12416 7710 12472
rect 7654 12144 7710 12200
rect 7562 12008 7618 12064
rect 7470 11212 7526 11248
rect 7470 11192 7472 11212
rect 7472 11192 7524 11212
rect 7524 11192 7526 11212
rect 6734 10376 6790 10432
rect 7102 10376 7158 10432
rect 6734 10260 6790 10296
rect 6734 10240 6736 10260
rect 6736 10240 6788 10260
rect 6788 10240 6790 10260
rect 6918 10140 6920 10160
rect 6920 10140 6972 10160
rect 6972 10140 6974 10160
rect 6550 9832 6606 9888
rect 6458 9696 6514 9752
rect 6918 10104 6974 10140
rect 6918 10004 6920 10024
rect 6920 10004 6972 10024
rect 6972 10004 6974 10024
rect 6918 9968 6974 10004
rect 6642 9152 6698 9208
rect 6642 8780 6644 8800
rect 6644 8780 6696 8800
rect 6696 8780 6698 8800
rect 6642 8744 6698 8780
rect 6366 8608 6422 8664
rect 6734 8336 6790 8392
rect 7654 11600 7710 11656
rect 7930 12588 7932 12608
rect 7932 12588 7984 12608
rect 7984 12588 7986 12608
rect 7930 12552 7986 12588
rect 7654 10920 7710 10976
rect 7378 10648 7434 10704
rect 7470 9560 7526 9616
rect 7470 9152 7526 9208
rect 8482 15408 8538 15464
rect 8666 17076 8668 17096
rect 8668 17076 8720 17096
rect 8720 17076 8722 17096
rect 8666 17040 8722 17076
rect 8666 15408 8722 15464
rect 8666 15272 8722 15328
rect 9770 25200 9826 25256
rect 9862 24928 9918 24984
rect 9770 24520 9826 24576
rect 9678 24384 9734 24440
rect 9678 24112 9734 24168
rect 9126 22500 9182 22536
rect 9126 22480 9128 22500
rect 9128 22480 9180 22500
rect 9180 22480 9182 22500
rect 9034 18264 9090 18320
rect 9310 21392 9366 21448
rect 9218 21140 9274 21176
rect 9218 21120 9220 21140
rect 9220 21120 9272 21140
rect 9272 21120 9274 21140
rect 9310 20984 9366 21040
rect 9218 20576 9274 20632
rect 8942 16768 8998 16824
rect 8114 12008 8170 12064
rect 8666 14728 8722 14784
rect 8574 14456 8630 14512
rect 8666 11600 8722 11656
rect 8574 11464 8630 11520
rect 8666 11328 8722 11384
rect 8574 11192 8630 11248
rect 8666 10784 8722 10840
rect 8574 10240 8630 10296
rect 8574 9560 8630 9616
rect 8482 9288 8538 9344
rect 8390 8880 8446 8936
rect 8114 8336 8170 8392
rect 6918 6296 6974 6352
rect 7378 6296 7434 6352
rect 7102 6024 7158 6080
rect 8206 8200 8262 8256
rect 8390 8200 8446 8256
rect 8206 7520 8262 7576
rect 8206 6704 8262 6760
rect 8942 13096 8998 13152
rect 9126 11736 9182 11792
rect 8758 9424 8814 9480
rect 8942 9596 8944 9616
rect 8944 9596 8996 9616
rect 8996 9596 8998 9616
rect 8942 9560 8998 9596
rect 8850 9288 8906 9344
rect 8758 9016 8814 9072
rect 8758 8472 8814 8528
rect 9494 21800 9550 21856
rect 9954 22344 10010 22400
rect 9862 20712 9918 20768
rect 9586 20168 9642 20224
rect 9310 13776 9366 13832
rect 9310 13640 9366 13696
rect 9678 19488 9734 19544
rect 9678 19216 9734 19272
rect 9678 17176 9734 17232
rect 10138 24792 10194 24848
rect 10598 27784 10654 27840
rect 10506 26152 10562 26208
rect 10506 24928 10562 24984
rect 10782 28076 10838 28112
rect 10782 28056 10784 28076
rect 10784 28056 10836 28076
rect 10836 28056 10838 28076
rect 10782 27784 10838 27840
rect 11058 28464 11114 28520
rect 11334 28328 11390 28384
rect 11150 27784 11206 27840
rect 10782 26560 10838 26616
rect 10690 25064 10746 25120
rect 10414 23840 10470 23896
rect 11058 27512 11114 27568
rect 11058 26832 11114 26888
rect 10966 25744 11022 25800
rect 9862 18536 9918 18592
rect 10230 19916 10286 19952
rect 10230 19896 10232 19916
rect 10232 19896 10284 19916
rect 10284 19896 10286 19916
rect 10414 23160 10470 23216
rect 10506 22752 10562 22808
rect 10414 21664 10470 21720
rect 10414 21528 10470 21584
rect 10506 20324 10562 20360
rect 10506 20304 10508 20324
rect 10508 20304 10560 20324
rect 10560 20304 10562 20324
rect 10506 18964 10562 19000
rect 10506 18944 10508 18964
rect 10508 18944 10560 18964
rect 10560 18944 10562 18964
rect 10966 23432 11022 23488
rect 11426 27648 11482 27704
rect 11334 27104 11390 27160
rect 11242 26832 11298 26888
rect 11150 23840 11206 23896
rect 10690 19896 10746 19952
rect 10506 17992 10562 18048
rect 10506 17620 10508 17640
rect 10508 17620 10560 17640
rect 10560 17620 10562 17640
rect 10506 17584 10562 17620
rect 9954 16904 10010 16960
rect 9494 15272 9550 15328
rect 9494 14728 9550 14784
rect 9494 14592 9550 14648
rect 9770 15680 9826 15736
rect 10230 16904 10286 16960
rect 10506 16768 10562 16824
rect 9954 15272 10010 15328
rect 9862 15136 9918 15192
rect 10138 15272 10194 15328
rect 9862 14592 9918 14648
rect 9494 13812 9496 13832
rect 9496 13812 9548 13832
rect 9548 13812 9550 13832
rect 9494 13776 9550 13812
rect 9586 13640 9642 13696
rect 10138 14320 10194 14376
rect 9862 14184 9918 14240
rect 9862 13776 9918 13832
rect 9310 13096 9366 13152
rect 9494 13096 9550 13152
rect 9310 12724 9312 12744
rect 9312 12724 9364 12744
rect 9364 12724 9366 12744
rect 9310 12688 9366 12724
rect 9678 12688 9734 12744
rect 9862 12688 9918 12744
rect 9770 12552 9826 12608
rect 9586 12008 9642 12064
rect 9494 11600 9550 11656
rect 9402 10648 9458 10704
rect 9126 9560 9182 9616
rect 9494 9968 9550 10024
rect 9402 9288 9458 9344
rect 9402 8900 9458 8936
rect 9402 8880 9404 8900
rect 9404 8880 9456 8900
rect 9456 8880 9458 8900
rect 9034 8336 9090 8392
rect 9218 8200 9274 8256
rect 10046 12844 10102 12880
rect 10046 12824 10048 12844
rect 10048 12824 10100 12844
rect 10100 12824 10102 12844
rect 10138 12552 10194 12608
rect 10046 11600 10102 11656
rect 10230 11092 10232 11112
rect 10232 11092 10284 11112
rect 10284 11092 10286 11112
rect 10230 11056 10286 11092
rect 10230 9968 10286 10024
rect 10414 14320 10470 14376
rect 10966 21548 11022 21584
rect 10966 21528 10968 21548
rect 10968 21528 11020 21548
rect 11020 21528 11022 21548
rect 10874 21256 10930 21312
rect 10874 19216 10930 19272
rect 11058 20712 11114 20768
rect 12530 28872 12586 28928
rect 12346 28600 12402 28656
rect 11886 27784 11942 27840
rect 11794 27648 11850 27704
rect 12070 23704 12126 23760
rect 11794 23568 11850 23624
rect 11518 23044 11574 23080
rect 11518 23024 11520 23044
rect 11520 23024 11572 23044
rect 11572 23024 11574 23044
rect 11886 23160 11942 23216
rect 11978 22888 12034 22944
rect 11702 22208 11758 22264
rect 11610 21972 11612 21992
rect 11612 21972 11664 21992
rect 11664 21972 11666 21992
rect 11610 21936 11666 21972
rect 12254 27648 12310 27704
rect 12530 28600 12586 28656
rect 12346 27412 12348 27432
rect 12348 27412 12400 27432
rect 12400 27412 12402 27432
rect 12346 27376 12402 27412
rect 12254 27240 12310 27296
rect 12806 27412 12808 27432
rect 12808 27412 12860 27432
rect 12860 27412 12862 27432
rect 12806 27376 12862 27412
rect 12254 25880 12310 25936
rect 12714 27104 12770 27160
rect 12438 25336 12494 25392
rect 12346 24656 12402 24712
rect 12346 23160 12402 23216
rect 11150 19252 11152 19272
rect 11152 19252 11204 19272
rect 11204 19252 11206 19272
rect 11150 19216 11206 19252
rect 11886 21800 11942 21856
rect 11794 21548 11850 21584
rect 11794 21528 11796 21548
rect 11796 21528 11848 21548
rect 11848 21528 11850 21548
rect 11794 21120 11850 21176
rect 11886 20848 11942 20904
rect 11794 20168 11850 20224
rect 11610 19896 11666 19952
rect 11058 18128 11114 18184
rect 11058 17448 11114 17504
rect 11058 17196 11114 17232
rect 11058 17176 11060 17196
rect 11060 17176 11112 17196
rect 11112 17176 11114 17196
rect 10598 15272 10654 15328
rect 11058 16496 11114 16552
rect 11242 17312 11298 17368
rect 12346 21528 12402 21584
rect 11886 19896 11942 19952
rect 12990 26560 13046 26616
rect 13174 28636 13176 28656
rect 13176 28636 13228 28656
rect 13228 28636 13230 28656
rect 13174 28600 13230 28636
rect 13174 26988 13230 27024
rect 13174 26968 13176 26988
rect 13176 26968 13228 26988
rect 13228 26968 13230 26988
rect 12898 24384 12954 24440
rect 12530 23568 12586 23624
rect 12806 23432 12862 23488
rect 12530 22344 12586 22400
rect 13358 28212 13414 28248
rect 13358 28192 13360 28212
rect 13360 28192 13412 28212
rect 13412 28192 13414 28212
rect 14002 29144 14058 29200
rect 13726 27376 13782 27432
rect 13450 26288 13506 26344
rect 13358 26016 13414 26072
rect 13266 24928 13322 24984
rect 13266 24656 13322 24712
rect 13082 23432 13138 23488
rect 13082 22752 13138 22808
rect 13450 24520 13506 24576
rect 13450 23296 13506 23352
rect 12806 22344 12862 22400
rect 12622 22072 12678 22128
rect 12438 21392 12494 21448
rect 12622 21428 12624 21448
rect 12624 21428 12676 21448
rect 12676 21428 12678 21448
rect 12622 21392 12678 21428
rect 12806 21664 12862 21720
rect 13174 22072 13230 22128
rect 13082 21936 13138 21992
rect 12898 21392 12954 21448
rect 12806 20712 12862 20768
rect 12898 20576 12954 20632
rect 12530 19624 12586 19680
rect 12438 19488 12494 19544
rect 11426 17312 11482 17368
rect 11150 15852 11152 15872
rect 11152 15852 11204 15872
rect 11204 15852 11206 15872
rect 11150 15816 11206 15852
rect 11242 15136 11298 15192
rect 10598 14048 10654 14104
rect 10506 12688 10562 12744
rect 10414 11600 10470 11656
rect 11058 14728 11114 14784
rect 10874 14048 10930 14104
rect 10874 13776 10930 13832
rect 11242 13776 11298 13832
rect 11886 18964 11942 19000
rect 11886 18944 11888 18964
rect 11888 18944 11940 18964
rect 11940 18944 11942 18964
rect 12162 18944 12218 19000
rect 12530 19216 12586 19272
rect 12806 19216 12862 19272
rect 12530 19080 12586 19136
rect 11794 18536 11850 18592
rect 11702 17196 11758 17232
rect 11702 17176 11704 17196
rect 11704 17176 11756 17196
rect 11756 17176 11758 17196
rect 11610 17040 11666 17096
rect 11794 16496 11850 16552
rect 11610 16224 11666 16280
rect 11518 15952 11574 16008
rect 12162 18420 12218 18456
rect 12162 18400 12164 18420
rect 12164 18400 12216 18420
rect 12216 18400 12218 18420
rect 12346 18400 12402 18456
rect 12162 18128 12218 18184
rect 11886 16224 11942 16280
rect 11978 15952 12034 16008
rect 11518 15272 11574 15328
rect 12162 17076 12164 17096
rect 12164 17076 12216 17096
rect 12216 17076 12218 17096
rect 12162 17040 12218 17076
rect 12714 18264 12770 18320
rect 12530 16496 12586 16552
rect 12438 16396 12440 16416
rect 12440 16396 12492 16416
rect 12492 16396 12494 16416
rect 12438 16360 12494 16396
rect 12254 15272 12310 15328
rect 11518 14068 11574 14104
rect 11518 14048 11520 14068
rect 11520 14048 11572 14068
rect 11572 14048 11574 14068
rect 10506 10376 10562 10432
rect 9586 8472 9642 8528
rect 10046 8744 10102 8800
rect 9954 8472 10010 8528
rect 9494 7520 9550 7576
rect 9310 6840 9366 6896
rect 9494 6840 9550 6896
rect 9310 6024 9366 6080
rect 9954 4564 9956 4584
rect 9956 4564 10008 4584
rect 10008 4564 10010 4584
rect 9954 4528 10010 4564
rect 10874 12008 10930 12064
rect 11150 12824 11206 12880
rect 11426 12844 11482 12880
rect 11426 12824 11428 12844
rect 11428 12824 11480 12844
rect 11480 12824 11482 12844
rect 11334 12552 11390 12608
rect 11426 12180 11428 12200
rect 11428 12180 11480 12200
rect 11480 12180 11482 12200
rect 11426 12144 11482 12180
rect 11058 12008 11114 12064
rect 11242 12008 11298 12064
rect 10874 11600 10930 11656
rect 10874 11092 10876 11112
rect 10876 11092 10928 11112
rect 10928 11092 10930 11112
rect 10874 11056 10930 11092
rect 11242 9968 11298 10024
rect 11242 9696 11298 9752
rect 11150 9152 11206 9208
rect 11058 8744 11114 8800
rect 11058 8508 11060 8528
rect 11060 8508 11112 8528
rect 11112 8508 11114 8528
rect 11058 8472 11114 8508
rect 11426 8356 11482 8392
rect 11426 8336 11428 8356
rect 11428 8336 11480 8356
rect 11480 8336 11482 8356
rect 11702 14048 11758 14104
rect 11702 12960 11758 13016
rect 11978 13948 11980 13968
rect 11980 13948 12032 13968
rect 12032 13948 12034 13968
rect 12254 14900 12256 14920
rect 12256 14900 12308 14920
rect 12308 14900 12310 14920
rect 12254 14864 12310 14900
rect 12254 14592 12310 14648
rect 11978 13912 12034 13948
rect 11978 13776 12034 13832
rect 12162 13812 12164 13832
rect 12164 13812 12216 13832
rect 12216 13812 12218 13832
rect 12162 13776 12218 13812
rect 13174 20712 13230 20768
rect 13082 18400 13138 18456
rect 12990 17856 13046 17912
rect 12990 17312 13046 17368
rect 12898 17040 12954 17096
rect 13358 21120 13414 21176
rect 13358 20884 13360 20904
rect 13360 20884 13412 20904
rect 13412 20884 13414 20904
rect 13358 20848 13414 20884
rect 13358 19624 13414 19680
rect 13266 17856 13322 17912
rect 13266 16768 13322 16824
rect 12806 15272 12862 15328
rect 12714 14728 12770 14784
rect 13266 15544 13322 15600
rect 12622 14184 12678 14240
rect 12438 13932 12494 13968
rect 12438 13912 12440 13932
rect 12440 13912 12492 13932
rect 12492 13912 12494 13932
rect 11794 12688 11850 12744
rect 11702 12144 11758 12200
rect 12070 12688 12126 12744
rect 12346 12280 12402 12336
rect 11794 12008 11850 12064
rect 11702 10668 11758 10704
rect 11702 10648 11704 10668
rect 11704 10648 11756 10668
rect 11756 10648 11758 10668
rect 11702 9152 11758 9208
rect 12070 11464 12126 11520
rect 12070 10240 12126 10296
rect 11978 9424 12034 9480
rect 11702 8628 11758 8664
rect 11702 8608 11704 8628
rect 11704 8608 11756 8628
rect 11756 8608 11758 8628
rect 11978 8608 12034 8664
rect 11518 7112 11574 7168
rect 10782 6568 10838 6624
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 11150 6568 11206 6624
rect 11058 6160 11114 6216
rect 11978 8064 12034 8120
rect 12254 9424 12310 9480
rect 12530 10376 12586 10432
rect 12806 13932 12862 13968
rect 12806 13912 12808 13932
rect 12808 13912 12860 13932
rect 12860 13912 12862 13932
rect 13266 13912 13322 13968
rect 12990 13232 13046 13288
rect 13082 12960 13138 13016
rect 13082 12688 13138 12744
rect 12714 10240 12770 10296
rect 12622 9696 12678 9752
rect 12254 8492 12310 8528
rect 12254 8472 12256 8492
rect 12256 8472 12308 8492
rect 12308 8472 12310 8492
rect 12438 8472 12494 8528
rect 11242 5888 11298 5944
rect 11334 5752 11390 5808
rect 11150 5616 11206 5672
rect 11794 6568 11850 6624
rect 11978 6060 11980 6080
rect 11980 6060 12032 6080
rect 12032 6060 12034 6080
rect 11978 6024 12034 6060
rect 12622 7384 12678 7440
rect 12622 7148 12624 7168
rect 12624 7148 12676 7168
rect 12676 7148 12678 7168
rect 12622 7112 12678 7148
rect 13910 27648 13966 27704
rect 13818 26968 13874 27024
rect 14554 28328 14610 28384
rect 13726 25356 13782 25392
rect 13726 25336 13728 25356
rect 13728 25336 13780 25356
rect 13780 25336 13782 25356
rect 15014 30504 15070 30560
rect 15934 30096 15990 30152
rect 14646 27820 14648 27840
rect 14648 27820 14700 27840
rect 14700 27820 14702 27840
rect 14646 27784 14702 27820
rect 15014 27920 15070 27976
rect 14370 26968 14426 27024
rect 14278 26696 14334 26752
rect 14186 25100 14188 25120
rect 14188 25100 14240 25120
rect 14240 25100 14242 25120
rect 14186 25064 14242 25100
rect 13818 21936 13874 21992
rect 13634 21664 13690 21720
rect 13818 21684 13874 21720
rect 13818 21664 13820 21684
rect 13820 21664 13872 21684
rect 13872 21664 13874 21684
rect 13542 21392 13598 21448
rect 13542 20848 13598 20904
rect 13634 20712 13690 20768
rect 14462 26696 14518 26752
rect 15198 27668 15254 27704
rect 15198 27648 15200 27668
rect 15200 27648 15252 27668
rect 15252 27648 15254 27668
rect 15106 27104 15162 27160
rect 14646 26016 14702 26072
rect 14462 25472 14518 25528
rect 14278 24384 14334 24440
rect 14554 24792 14610 24848
rect 14002 23976 14058 24032
rect 14002 20848 14058 20904
rect 14278 21664 14334 21720
rect 14094 20304 14150 20360
rect 14278 20168 14334 20224
rect 13910 19352 13966 19408
rect 13726 18572 13728 18592
rect 13728 18572 13780 18592
rect 13780 18572 13782 18592
rect 13726 18536 13782 18572
rect 13634 15000 13690 15056
rect 14554 23432 14610 23488
rect 15014 26580 15070 26616
rect 15290 27376 15346 27432
rect 15014 26560 15016 26580
rect 15016 26560 15068 26580
rect 15068 26560 15070 26580
rect 14830 26152 14886 26208
rect 14922 25336 14978 25392
rect 14830 25200 14886 25256
rect 14738 21528 14794 21584
rect 14646 21120 14702 21176
rect 14462 20340 14464 20360
rect 14464 20340 14516 20360
rect 14516 20340 14518 20360
rect 14462 20304 14518 20340
rect 15198 25236 15200 25256
rect 15200 25236 15252 25256
rect 15252 25236 15254 25256
rect 15198 25200 15254 25236
rect 15106 23976 15162 24032
rect 15382 24928 15438 24984
rect 15474 24792 15530 24848
rect 15290 23568 15346 23624
rect 15014 20984 15070 21040
rect 15198 20984 15254 21040
rect 15014 20576 15070 20632
rect 14646 19896 14702 19952
rect 14554 19760 14610 19816
rect 14370 18536 14426 18592
rect 14094 17856 14150 17912
rect 14002 15680 14058 15736
rect 13910 15408 13966 15464
rect 13818 14592 13874 14648
rect 13726 14184 13782 14240
rect 12898 8608 12954 8664
rect 12806 8200 12862 8256
rect 12714 6840 12770 6896
rect 12162 5480 12218 5536
rect 12622 4700 12624 4720
rect 12624 4700 12676 4720
rect 12676 4700 12678 4720
rect 12622 4664 12678 4700
rect 13174 8880 13230 8936
rect 13818 13096 13874 13152
rect 13818 11872 13874 11928
rect 13818 11464 13874 11520
rect 13358 7520 13414 7576
rect 13634 7520 13690 7576
rect 12898 3712 12954 3768
rect 13634 6704 13690 6760
rect 14278 17040 14334 17096
rect 14278 16632 14334 16688
rect 14186 15000 14242 15056
rect 14094 8608 14150 8664
rect 14094 7112 14150 7168
rect 14278 14728 14334 14784
rect 14278 14592 14334 14648
rect 14278 13096 14334 13152
rect 14370 12960 14426 13016
rect 14370 12416 14426 12472
rect 14646 18536 14702 18592
rect 14922 19352 14978 19408
rect 14738 17992 14794 18048
rect 14830 17584 14886 17640
rect 14646 13912 14702 13968
rect 15658 23724 15714 23760
rect 15658 23704 15660 23724
rect 15660 23704 15712 23724
rect 15712 23704 15714 23724
rect 16026 27668 16082 27704
rect 16026 27648 16028 27668
rect 16028 27648 16080 27668
rect 16080 27648 16082 27668
rect 16118 27104 16174 27160
rect 16026 26424 16082 26480
rect 15934 25880 15990 25936
rect 15842 24792 15898 24848
rect 15106 19116 15108 19136
rect 15108 19116 15160 19136
rect 15160 19116 15162 19136
rect 15106 19080 15162 19116
rect 15290 18944 15346 19000
rect 15106 17720 15162 17776
rect 15474 17312 15530 17368
rect 15658 18400 15714 18456
rect 15566 16768 15622 16824
rect 15198 16532 15200 16552
rect 15200 16532 15252 16552
rect 15252 16532 15254 16552
rect 15014 16360 15070 16416
rect 15198 16496 15254 16532
rect 15014 15444 15016 15464
rect 15016 15444 15068 15464
rect 15068 15444 15070 15464
rect 15014 15408 15070 15444
rect 15198 15000 15254 15056
rect 15106 14456 15162 14512
rect 14830 13912 14886 13968
rect 14554 12416 14610 12472
rect 14830 12960 14886 13016
rect 15290 14764 15292 14784
rect 15292 14764 15344 14784
rect 15344 14764 15346 14784
rect 15290 14728 15346 14764
rect 15382 13096 15438 13152
rect 15290 12960 15346 13016
rect 14554 12280 14610 12336
rect 14462 11872 14518 11928
rect 14462 11736 14518 11792
rect 14462 10240 14518 10296
rect 14278 9424 14334 9480
rect 14278 9152 14334 9208
rect 14554 9172 14610 9208
rect 14554 9152 14556 9172
rect 14556 9152 14608 9172
rect 14608 9152 14610 9172
rect 14278 8880 14334 8936
rect 14554 8336 14610 8392
rect 14554 7948 14610 7984
rect 14554 7928 14556 7948
rect 14556 7928 14608 7948
rect 14608 7928 14610 7948
rect 13726 5344 13782 5400
rect 14370 5244 14372 5264
rect 14372 5244 14424 5264
rect 14424 5244 14426 5264
rect 14370 5208 14426 5244
rect 14738 11736 14794 11792
rect 15014 11600 15070 11656
rect 15106 10920 15162 10976
rect 15106 9560 15162 9616
rect 15014 8608 15070 8664
rect 15014 8472 15070 8528
rect 15198 8492 15254 8528
rect 15198 8472 15200 8492
rect 15200 8472 15252 8492
rect 15252 8472 15254 8492
rect 15014 8336 15070 8392
rect 15474 11872 15530 11928
rect 16302 26424 16358 26480
rect 15934 19488 15990 19544
rect 16210 20576 16266 20632
rect 16946 27396 17002 27432
rect 16946 27376 16948 27396
rect 16948 27376 17000 27396
rect 17000 27376 17002 27396
rect 16762 26016 16818 26072
rect 16946 25900 17002 25936
rect 16946 25880 16948 25900
rect 16948 25880 17000 25900
rect 17000 25880 17002 25900
rect 16854 25608 16910 25664
rect 16762 25064 16818 25120
rect 17038 25608 17094 25664
rect 16578 23316 16634 23352
rect 16578 23296 16580 23316
rect 16580 23296 16632 23316
rect 16632 23296 16634 23316
rect 16026 18944 16082 19000
rect 16026 18672 16082 18728
rect 16026 18400 16082 18456
rect 15934 16496 15990 16552
rect 15934 15680 15990 15736
rect 15934 15544 15990 15600
rect 16118 15952 16174 16008
rect 16578 20032 16634 20088
rect 16946 24656 17002 24712
rect 17038 23704 17094 23760
rect 16762 22888 16818 22944
rect 16946 22752 17002 22808
rect 16854 22072 16910 22128
rect 16762 21120 16818 21176
rect 16394 19080 16450 19136
rect 16302 17740 16358 17776
rect 16302 17720 16304 17740
rect 16304 17720 16356 17740
rect 16356 17720 16358 17740
rect 16946 21256 17002 21312
rect 17222 23296 17278 23352
rect 15842 12280 15898 12336
rect 15842 12008 15898 12064
rect 15566 9580 15622 9616
rect 15566 9560 15568 9580
rect 15568 9560 15620 9580
rect 15620 9560 15622 9580
rect 15474 9424 15530 9480
rect 15382 8356 15438 8392
rect 15382 8336 15384 8356
rect 15384 8336 15436 8356
rect 15436 8336 15438 8356
rect 15382 8200 15438 8256
rect 15198 6840 15254 6896
rect 16762 15700 16818 15736
rect 16762 15680 16764 15700
rect 16764 15680 16816 15700
rect 16816 15680 16818 15700
rect 16762 14864 16818 14920
rect 16762 14728 16818 14784
rect 17130 20324 17186 20360
rect 17130 20304 17132 20324
rect 17132 20304 17184 20324
rect 17184 20304 17186 20324
rect 18142 29028 18198 29064
rect 18142 29008 18144 29028
rect 18144 29008 18196 29028
rect 18196 29008 18198 29028
rect 17498 25608 17554 25664
rect 17498 24792 17554 24848
rect 17406 24556 17408 24576
rect 17408 24556 17460 24576
rect 17460 24556 17462 24576
rect 17406 24520 17462 24556
rect 17498 23976 17554 24032
rect 18142 28056 18198 28112
rect 17958 27376 18014 27432
rect 17774 26288 17830 26344
rect 17590 23044 17646 23080
rect 18418 28192 18474 28248
rect 23110 31184 23166 31240
rect 23018 30232 23074 30288
rect 20166 29280 20222 29336
rect 19522 28736 19578 28792
rect 18602 27648 18658 27704
rect 19338 28328 19394 28384
rect 19154 27512 19210 27568
rect 20166 28872 20222 28928
rect 19614 28600 19670 28656
rect 18510 27376 18566 27432
rect 18602 27240 18658 27296
rect 18510 26696 18566 26752
rect 17958 24656 18014 24712
rect 17590 23024 17592 23044
rect 17592 23024 17644 23044
rect 17644 23024 17646 23044
rect 17498 22636 17554 22672
rect 17498 22616 17500 22636
rect 17500 22616 17552 22636
rect 17552 22616 17554 22636
rect 17406 21664 17462 21720
rect 17314 18264 17370 18320
rect 17130 16768 17186 16824
rect 17038 16360 17094 16416
rect 16946 15408 17002 15464
rect 17222 14048 17278 14104
rect 17038 12960 17094 13016
rect 16302 11328 16358 11384
rect 16578 11464 16634 11520
rect 16486 11328 16542 11384
rect 15842 10512 15898 10568
rect 16026 10512 16082 10568
rect 16026 9016 16082 9072
rect 15658 7928 15714 7984
rect 15934 8236 15936 8256
rect 15936 8236 15988 8256
rect 15988 8236 15990 8256
rect 15934 8200 15990 8236
rect 16302 10412 16304 10432
rect 16304 10412 16356 10432
rect 16356 10412 16358 10432
rect 16302 10376 16358 10412
rect 16486 11192 16542 11248
rect 16762 10784 16818 10840
rect 16762 10104 16818 10160
rect 16394 9832 16450 9888
rect 16302 9424 16358 9480
rect 16302 9016 16358 9072
rect 15842 3984 15898 4040
rect 15106 3576 15162 3632
rect 16670 9560 16726 9616
rect 16670 7520 16726 7576
rect 17314 12688 17370 12744
rect 17222 12008 17278 12064
rect 17130 11600 17186 11656
rect 16946 11092 16948 11112
rect 16948 11092 17000 11112
rect 17000 11092 17002 11112
rect 16946 11056 17002 11092
rect 17130 8880 17186 8936
rect 17958 23432 18014 23488
rect 17866 22752 17922 22808
rect 17682 21392 17738 21448
rect 17682 21292 17684 21312
rect 17684 21292 17736 21312
rect 17736 21292 17738 21312
rect 17682 21256 17738 21292
rect 17682 20984 17738 21040
rect 17866 20712 17922 20768
rect 17774 19080 17830 19136
rect 18234 22616 18290 22672
rect 18234 20848 18290 20904
rect 18786 26696 18842 26752
rect 18418 23160 18474 23216
rect 18326 20032 18382 20088
rect 18142 19896 18198 19952
rect 18142 18264 18198 18320
rect 18142 17992 18198 18048
rect 18234 17312 18290 17368
rect 17590 15000 17646 15056
rect 17866 15000 17922 15056
rect 17682 14592 17738 14648
rect 17590 13368 17646 13424
rect 17590 11056 17646 11112
rect 16854 7248 16910 7304
rect 17222 7248 17278 7304
rect 17222 6568 17278 6624
rect 17498 10784 17554 10840
rect 17406 10104 17462 10160
rect 17590 8880 17646 8936
rect 17038 5636 17094 5672
rect 17038 5616 17040 5636
rect 17040 5616 17092 5636
rect 17092 5616 17094 5636
rect 13542 3304 13598 3360
rect 17774 12416 17830 12472
rect 17958 13912 18014 13968
rect 17958 13640 18014 13696
rect 17866 11872 17922 11928
rect 19614 27376 19670 27432
rect 19154 26968 19210 27024
rect 19154 26288 19210 26344
rect 19154 25472 19210 25528
rect 19338 25472 19394 25528
rect 19706 27276 19708 27296
rect 19708 27276 19760 27296
rect 19760 27276 19762 27296
rect 19706 27240 19762 27276
rect 19982 27512 20038 27568
rect 19890 27240 19946 27296
rect 19522 26016 19578 26072
rect 19614 25900 19670 25936
rect 19614 25880 19616 25900
rect 19616 25880 19668 25900
rect 19668 25880 19670 25900
rect 19706 24928 19762 24984
rect 19246 24656 19302 24712
rect 18694 23432 18750 23488
rect 18970 23160 19026 23216
rect 18878 22616 18934 22672
rect 18878 22344 18934 22400
rect 18418 16360 18474 16416
rect 18142 12416 18198 12472
rect 18694 16632 18750 16688
rect 18970 16496 19026 16552
rect 18602 14592 18658 14648
rect 18878 15136 18934 15192
rect 18786 14884 18842 14920
rect 18786 14864 18788 14884
rect 18788 14864 18840 14884
rect 18840 14864 18842 14884
rect 18786 14592 18842 14648
rect 18878 14456 18934 14512
rect 18786 13932 18842 13968
rect 18786 13912 18788 13932
rect 18788 13912 18840 13932
rect 18840 13912 18842 13932
rect 18786 12724 18788 12744
rect 18788 12724 18840 12744
rect 18840 12724 18842 12744
rect 18786 12688 18842 12724
rect 18970 12960 19026 13016
rect 18970 12688 19026 12744
rect 19154 22072 19210 22128
rect 19430 24656 19486 24712
rect 19890 25900 19946 25936
rect 19890 25880 19892 25900
rect 19892 25880 19944 25900
rect 19944 25880 19946 25900
rect 19798 24656 19854 24712
rect 19430 23024 19486 23080
rect 19338 22888 19394 22944
rect 19338 22344 19394 22400
rect 19430 22208 19486 22264
rect 19338 22072 19394 22128
rect 19246 21800 19302 21856
rect 19338 21684 19394 21720
rect 19338 21664 19340 21684
rect 19340 21664 19392 21684
rect 19392 21664 19394 21684
rect 19246 20984 19302 21040
rect 19614 22092 19670 22128
rect 19614 22072 19616 22092
rect 19616 22072 19668 22092
rect 19668 22072 19670 22092
rect 19522 20984 19578 21040
rect 19338 20848 19394 20904
rect 19522 20848 19578 20904
rect 19430 19624 19486 19680
rect 19246 17992 19302 18048
rect 19890 21548 19946 21584
rect 19890 21528 19892 21548
rect 19892 21528 19944 21548
rect 19944 21528 19946 21548
rect 19706 21392 19762 21448
rect 19982 21392 20038 21448
rect 19706 20984 19762 21040
rect 19706 20712 19762 20768
rect 19706 20032 19762 20088
rect 19430 17992 19486 18048
rect 19154 14592 19210 14648
rect 19338 16768 19394 16824
rect 19706 16124 19708 16144
rect 19708 16124 19760 16144
rect 19760 16124 19762 16144
rect 19706 16088 19762 16124
rect 19706 15680 19762 15736
rect 19522 15136 19578 15192
rect 19614 15020 19670 15056
rect 19614 15000 19616 15020
rect 19616 15000 19668 15020
rect 19668 15000 19670 15020
rect 19522 14456 19578 14512
rect 19890 20032 19946 20088
rect 20350 28328 20406 28384
rect 20534 28328 20590 28384
rect 20442 28056 20498 28112
rect 20166 27376 20222 27432
rect 20166 26832 20222 26888
rect 20258 26152 20314 26208
rect 20258 25336 20314 25392
rect 20258 24928 20314 24984
rect 20442 26016 20498 26072
rect 20626 26832 20682 26888
rect 21178 26308 21234 26344
rect 21178 26288 21180 26308
rect 21180 26288 21232 26308
rect 21232 26288 21234 26308
rect 20994 25744 21050 25800
rect 20534 25336 20590 25392
rect 20534 24112 20590 24168
rect 20166 22888 20222 22944
rect 20166 22092 20222 22128
rect 20166 22072 20168 22092
rect 20168 22072 20220 22092
rect 20220 22072 20222 22092
rect 21914 29008 21970 29064
rect 22190 29008 22246 29064
rect 21822 27940 21878 27976
rect 21822 27920 21824 27940
rect 21824 27920 21876 27940
rect 21876 27920 21878 27940
rect 22098 27784 22154 27840
rect 22098 27648 22154 27704
rect 22006 27376 22062 27432
rect 22558 28464 22614 28520
rect 22190 27512 22246 27568
rect 22098 27104 22154 27160
rect 21822 26968 21878 27024
rect 21362 25744 21418 25800
rect 21454 24928 21510 24984
rect 20810 23704 20866 23760
rect 20902 23432 20958 23488
rect 20258 21664 20314 21720
rect 20258 21392 20314 21448
rect 20718 22888 20774 22944
rect 20718 22344 20774 22400
rect 20350 20712 20406 20768
rect 20166 19252 20168 19272
rect 20168 19252 20220 19272
rect 20220 19252 20222 19272
rect 20166 19216 20222 19252
rect 19982 16632 20038 16688
rect 20074 15000 20130 15056
rect 18510 11056 18566 11112
rect 17774 8900 17830 8936
rect 17774 8880 17776 8900
rect 17776 8880 17828 8900
rect 17828 8880 17830 8900
rect 18050 8472 18106 8528
rect 17774 6840 17830 6896
rect 17590 6432 17646 6488
rect 17774 6060 17776 6080
rect 17776 6060 17828 6080
rect 17828 6060 17830 6080
rect 17774 6024 17830 6060
rect 17958 5752 18014 5808
rect 17406 3168 17462 3224
rect 10874 2624 10930 2680
rect 18786 10920 18842 10976
rect 18786 10512 18842 10568
rect 18602 9424 18658 9480
rect 18418 6296 18474 6352
rect 18418 5888 18474 5944
rect 18694 8880 18750 8936
rect 18786 7792 18842 7848
rect 19338 13640 19394 13696
rect 19614 12280 19670 12336
rect 19430 12164 19486 12200
rect 19430 12144 19432 12164
rect 19432 12144 19484 12164
rect 19484 12144 19486 12164
rect 19430 11872 19486 11928
rect 19338 11328 19394 11384
rect 19246 10920 19302 10976
rect 19614 11192 19670 11248
rect 19246 9832 19302 9888
rect 19430 9696 19486 9752
rect 19614 9696 19670 9752
rect 19338 9560 19394 9616
rect 19522 9424 19578 9480
rect 19430 8508 19432 8528
rect 19432 8508 19484 8528
rect 19484 8508 19486 8528
rect 19430 8472 19486 8508
rect 19338 7420 19340 7440
rect 19340 7420 19392 7440
rect 19392 7420 19394 7440
rect 19338 7384 19394 7420
rect 19890 13948 19892 13968
rect 19892 13948 19944 13968
rect 19944 13948 19946 13968
rect 19890 13912 19946 13948
rect 19798 13368 19854 13424
rect 19890 11076 19946 11112
rect 19890 11056 19892 11076
rect 19892 11056 19944 11076
rect 19944 11056 19946 11076
rect 19798 10512 19854 10568
rect 19890 8628 19946 8664
rect 19890 8608 19892 8628
rect 19892 8608 19944 8628
rect 19944 8608 19946 8628
rect 20442 19372 20498 19408
rect 20442 19352 20444 19372
rect 20444 19352 20496 19372
rect 20496 19352 20498 19372
rect 20258 16668 20260 16688
rect 20260 16668 20312 16688
rect 20312 16668 20314 16688
rect 20258 16632 20314 16668
rect 21362 24520 21418 24576
rect 21270 24112 21326 24168
rect 20810 21564 20812 21584
rect 20812 21564 20864 21584
rect 20864 21564 20866 21584
rect 20810 21528 20866 21564
rect 20810 19624 20866 19680
rect 20626 19488 20682 19544
rect 20718 19352 20774 19408
rect 20258 15680 20314 15736
rect 20810 16360 20866 16416
rect 20718 16108 20774 16144
rect 20718 16088 20720 16108
rect 20720 16088 20772 16108
rect 20772 16088 20774 16108
rect 20718 15952 20774 16008
rect 21086 20032 21142 20088
rect 20718 15272 20774 15328
rect 20350 14456 20406 14512
rect 20626 15000 20682 15056
rect 20442 14184 20498 14240
rect 20350 13912 20406 13968
rect 20350 11600 20406 11656
rect 20810 13640 20866 13696
rect 20350 11056 20406 11112
rect 20350 10804 20406 10840
rect 20350 10784 20352 10804
rect 20352 10784 20404 10804
rect 20404 10784 20406 10804
rect 20534 10804 20590 10840
rect 20534 10784 20536 10804
rect 20536 10784 20588 10804
rect 20588 10784 20590 10804
rect 20626 10240 20682 10296
rect 20350 9560 20406 9616
rect 20350 9152 20406 9208
rect 20350 8608 20406 8664
rect 20258 6860 20314 6896
rect 20258 6840 20260 6860
rect 20260 6840 20312 6860
rect 20312 6840 20314 6860
rect 19522 5616 19578 5672
rect 20534 6704 20590 6760
rect 20534 6432 20590 6488
rect 20718 5616 20774 5672
rect 21270 18808 21326 18864
rect 21638 24112 21694 24168
rect 21914 26152 21970 26208
rect 21914 25236 21916 25256
rect 21916 25236 21968 25256
rect 21968 25236 21970 25256
rect 21914 25200 21970 25236
rect 21914 24248 21970 24304
rect 21914 24112 21970 24168
rect 21822 23432 21878 23488
rect 21638 20984 21694 21040
rect 21454 19080 21510 19136
rect 20902 11056 20958 11112
rect 20902 10920 20958 10976
rect 22098 24520 22154 24576
rect 22282 24656 22338 24712
rect 22282 23160 22338 23216
rect 22742 26696 22798 26752
rect 22742 26288 22798 26344
rect 22650 25236 22652 25256
rect 22652 25236 22704 25256
rect 22704 25236 22706 25256
rect 22650 25200 22706 25236
rect 22006 20984 22062 21040
rect 21730 19216 21786 19272
rect 22006 18672 22062 18728
rect 22006 17992 22062 18048
rect 21546 15952 21602 16008
rect 21454 14184 21510 14240
rect 21454 13776 21510 13832
rect 22742 23160 22798 23216
rect 22742 22924 22744 22944
rect 22744 22924 22796 22944
rect 22796 22924 22798 22944
rect 22742 22888 22798 22924
rect 22650 22480 22706 22536
rect 22742 22208 22798 22264
rect 22558 20460 22614 20496
rect 22558 20440 22560 20460
rect 22560 20440 22612 20460
rect 22612 20440 22614 20460
rect 22558 19896 22614 19952
rect 22742 21664 22798 21720
rect 22742 20848 22798 20904
rect 22466 18964 22522 19000
rect 22466 18944 22468 18964
rect 22468 18944 22520 18964
rect 22520 18944 22522 18964
rect 22466 18708 22468 18728
rect 22468 18708 22520 18728
rect 22520 18708 22522 18728
rect 22466 18672 22522 18708
rect 22558 18128 22614 18184
rect 21546 13640 21602 13696
rect 21454 12280 21510 12336
rect 21086 10920 21142 10976
rect 21178 10512 21234 10568
rect 20994 7656 21050 7712
rect 21730 13232 21786 13288
rect 21822 12960 21878 13016
rect 22006 15680 22062 15736
rect 22742 17584 22798 17640
rect 22098 13232 22154 13288
rect 22650 15272 22706 15328
rect 23570 30912 23626 30968
rect 23202 29416 23258 29472
rect 23294 28600 23350 28656
rect 23478 27784 23534 27840
rect 23570 27648 23626 27704
rect 23478 25744 23534 25800
rect 23846 27396 23902 27432
rect 23846 27376 23848 27396
rect 23848 27376 23900 27396
rect 23900 27376 23902 27396
rect 23018 24656 23074 24712
rect 23386 24656 23442 24712
rect 23386 23840 23442 23896
rect 22926 15680 22982 15736
rect 23294 19352 23350 19408
rect 23754 25336 23810 25392
rect 23662 23976 23718 24032
rect 23754 23568 23810 23624
rect 24214 27512 24270 27568
rect 24306 24928 24362 24984
rect 23570 23432 23626 23488
rect 23846 23468 23848 23488
rect 23848 23468 23900 23488
rect 23900 23468 23902 23488
rect 23846 23432 23902 23468
rect 24030 23568 24086 23624
rect 23202 17196 23258 17232
rect 23202 17176 23204 17196
rect 23204 17176 23256 17196
rect 23256 17176 23258 17196
rect 22374 14592 22430 14648
rect 22282 14184 22338 14240
rect 21362 10512 21418 10568
rect 21546 9460 21548 9480
rect 21548 9460 21600 9480
rect 21600 9460 21602 9480
rect 21546 9424 21602 9460
rect 21454 8744 21510 8800
rect 22098 12552 22154 12608
rect 21822 11464 21878 11520
rect 22190 12044 22192 12064
rect 22192 12044 22244 12064
rect 22244 12044 22246 12064
rect 22190 12008 22246 12044
rect 22374 13640 22430 13696
rect 22006 10668 22062 10704
rect 22006 10648 22008 10668
rect 22008 10648 22060 10668
rect 22060 10648 22062 10668
rect 22282 9424 22338 9480
rect 22006 8916 22008 8936
rect 22008 8916 22060 8936
rect 22060 8916 22062 8936
rect 22006 8880 22062 8916
rect 21362 5616 21418 5672
rect 22282 9152 22338 9208
rect 22650 13232 22706 13288
rect 22926 13912 22982 13968
rect 22650 12552 22706 12608
rect 22650 11092 22652 11112
rect 22652 11092 22704 11112
rect 22704 11092 22706 11112
rect 22650 11056 22706 11092
rect 22742 10784 22798 10840
rect 22650 10240 22706 10296
rect 23662 17448 23718 17504
rect 23478 16244 23534 16280
rect 23478 16224 23480 16244
rect 23480 16224 23532 16244
rect 23532 16224 23534 16244
rect 23662 15544 23718 15600
rect 23386 13776 23442 13832
rect 23294 13232 23350 13288
rect 23018 11192 23074 11248
rect 23202 12416 23258 12472
rect 23018 10240 23074 10296
rect 22558 9324 22560 9344
rect 22560 9324 22612 9344
rect 22612 9324 22614 9344
rect 22558 9288 22614 9324
rect 22834 8084 22890 8120
rect 22834 8064 22836 8084
rect 22836 8064 22888 8084
rect 22888 8064 22890 8084
rect 22742 5344 22798 5400
rect 20718 4528 20774 4584
rect 22926 6704 22982 6760
rect 23110 8064 23166 8120
rect 23202 6160 23258 6216
rect 23846 21292 23848 21312
rect 23848 21292 23900 21312
rect 23900 21292 23902 21312
rect 23846 21256 23902 21292
rect 25594 28192 25650 28248
rect 24490 24384 24546 24440
rect 25502 27820 25504 27840
rect 25504 27820 25556 27840
rect 25556 27820 25558 27840
rect 25502 27784 25558 27820
rect 25134 25744 25190 25800
rect 24674 23704 24730 23760
rect 24582 22208 24638 22264
rect 23846 20440 23902 20496
rect 23846 19760 23902 19816
rect 23938 16904 23994 16960
rect 23662 14320 23718 14376
rect 23938 15816 23994 15872
rect 23570 10240 23626 10296
rect 23478 8608 23534 8664
rect 23386 7384 23442 7440
rect 23754 8236 23756 8256
rect 23756 8236 23808 8256
rect 23808 8236 23810 8256
rect 23754 8200 23810 8236
rect 23938 13812 23940 13832
rect 23940 13812 23992 13832
rect 23992 13812 23994 13832
rect 23938 13776 23994 13812
rect 23938 13640 23994 13696
rect 23938 12316 23940 12336
rect 23940 12316 23992 12336
rect 23992 12316 23994 12336
rect 23938 12280 23994 12316
rect 23938 11736 23994 11792
rect 24490 20712 24546 20768
rect 24214 17196 24270 17232
rect 24214 17176 24216 17196
rect 24216 17176 24268 17196
rect 24268 17176 24270 17196
rect 24306 16360 24362 16416
rect 24306 14456 24362 14512
rect 24122 13676 24124 13696
rect 24124 13676 24176 13696
rect 24176 13676 24178 13696
rect 24122 13640 24178 13676
rect 24122 13268 24124 13288
rect 24124 13268 24176 13288
rect 24176 13268 24178 13288
rect 24122 13232 24178 13268
rect 24582 17992 24638 18048
rect 25134 25064 25190 25120
rect 24950 23024 25006 23080
rect 24766 20052 24822 20088
rect 24766 20032 24768 20052
rect 24768 20032 24820 20052
rect 24820 20032 24822 20052
rect 24950 19624 25006 19680
rect 25226 22344 25282 22400
rect 25134 21392 25190 21448
rect 24950 19080 25006 19136
rect 25594 26424 25650 26480
rect 25962 28056 26018 28112
rect 26330 26016 26386 26072
rect 26238 25220 26294 25256
rect 26238 25200 26240 25220
rect 26240 25200 26292 25220
rect 26292 25200 26294 25220
rect 25134 16768 25190 16824
rect 24950 14900 24952 14920
rect 24952 14900 25004 14920
rect 25004 14900 25006 14920
rect 24950 14864 25006 14900
rect 24490 14320 24546 14376
rect 24490 13368 24546 13424
rect 24214 11092 24216 11112
rect 24216 11092 24268 11112
rect 24268 11092 24270 11112
rect 24214 11056 24270 11092
rect 23938 10784 23994 10840
rect 24306 10920 24362 10976
rect 24122 10668 24178 10704
rect 24122 10648 24124 10668
rect 24124 10648 24176 10668
rect 24176 10648 24178 10668
rect 24122 10240 24178 10296
rect 24122 9832 24178 9888
rect 23478 5636 23534 5672
rect 23478 5616 23480 5636
rect 23480 5616 23532 5636
rect 23532 5616 23534 5636
rect 23202 5208 23258 5264
rect 22834 3848 22890 3904
rect 24122 7384 24178 7440
rect 24306 9696 24362 9752
rect 24766 12844 24822 12880
rect 24766 12824 24768 12844
rect 24768 12824 24820 12844
rect 24820 12824 24822 12844
rect 24950 12436 25006 12472
rect 24950 12416 24952 12436
rect 24952 12416 25004 12436
rect 25004 12416 25006 12436
rect 24950 12280 25006 12336
rect 24766 8628 24822 8664
rect 25226 15816 25282 15872
rect 25502 21936 25558 21992
rect 25686 21956 25742 21992
rect 25686 21936 25688 21956
rect 25688 21936 25740 21956
rect 25740 21936 25742 21956
rect 25594 17992 25650 18048
rect 25502 15952 25558 16008
rect 25410 12416 25466 12472
rect 24766 8608 24768 8628
rect 24768 8608 24820 8628
rect 24820 8608 24822 8628
rect 24582 8336 24638 8392
rect 24582 5344 24638 5400
rect 25594 14764 25596 14784
rect 25596 14764 25648 14784
rect 25648 14764 25650 14784
rect 25594 14728 25650 14764
rect 25594 12008 25650 12064
rect 25410 10376 25466 10432
rect 25870 20712 25926 20768
rect 25778 19796 25780 19816
rect 25780 19796 25832 19816
rect 25832 19796 25834 19816
rect 25778 19760 25834 19796
rect 25778 19372 25834 19408
rect 26054 19896 26110 19952
rect 25778 19352 25780 19372
rect 25780 19352 25832 19372
rect 25832 19352 25834 19372
rect 25778 12960 25834 13016
rect 25778 12416 25834 12472
rect 25686 10648 25742 10704
rect 26238 22616 26294 22672
rect 26790 25608 26846 25664
rect 26606 25336 26662 25392
rect 26790 25200 26846 25256
rect 26422 23316 26478 23352
rect 26422 23296 26424 23316
rect 26424 23296 26476 23316
rect 26476 23296 26478 23316
rect 26790 24928 26846 24984
rect 26514 20168 26570 20224
rect 26422 19488 26478 19544
rect 26514 19080 26570 19136
rect 26790 20440 26846 20496
rect 27250 29144 27306 29200
rect 27066 27512 27122 27568
rect 26974 26444 27030 26480
rect 26974 26424 26976 26444
rect 26976 26424 27028 26444
rect 27028 26424 27030 26444
rect 27250 25880 27306 25936
rect 26698 19624 26754 19680
rect 27250 20712 27306 20768
rect 26606 18400 26662 18456
rect 26238 18128 26294 18184
rect 26514 17756 26516 17776
rect 26516 17756 26568 17776
rect 26568 17756 26570 17776
rect 26514 17720 26570 17756
rect 26238 13504 26294 13560
rect 25962 12300 26018 12336
rect 25962 12280 25964 12300
rect 25964 12280 26016 12300
rect 26016 12280 26018 12300
rect 26330 11328 26386 11384
rect 25594 9832 25650 9888
rect 25502 9152 25558 9208
rect 25778 9016 25834 9072
rect 25778 8472 25834 8528
rect 26146 9036 26202 9072
rect 26146 9016 26148 9036
rect 26148 9016 26200 9036
rect 26200 9016 26202 9036
rect 25962 6316 26018 6352
rect 25962 6296 25964 6316
rect 25964 6296 26016 6316
rect 26016 6296 26018 6316
rect 25686 6160 25742 6216
rect 26514 13812 26516 13832
rect 26516 13812 26568 13832
rect 26568 13812 26570 13832
rect 26514 13776 26570 13812
rect 26974 15428 27030 15464
rect 26974 15408 26976 15428
rect 26976 15408 27028 15428
rect 27028 15408 27030 15428
rect 26790 13776 26846 13832
rect 26790 10668 26846 10704
rect 26790 10648 26792 10668
rect 26792 10648 26844 10668
rect 26844 10648 26846 10668
rect 26790 9424 26846 9480
rect 26606 9016 26662 9072
rect 27710 26560 27766 26616
rect 28262 24812 28318 24848
rect 28262 24792 28264 24812
rect 28264 24792 28316 24812
rect 28316 24792 28318 24812
rect 27434 20884 27436 20904
rect 27436 20884 27488 20904
rect 27488 20884 27490 20904
rect 27434 20848 27490 20884
rect 27250 12144 27306 12200
rect 27158 11328 27214 11384
rect 27986 24112 28042 24168
rect 27986 20984 28042 21040
rect 27986 20440 28042 20496
rect 28170 23432 28226 23488
rect 28262 19624 28318 19680
rect 27710 17312 27766 17368
rect 27618 16088 27674 16144
rect 27618 15000 27674 15056
rect 27434 13812 27436 13832
rect 27436 13812 27488 13832
rect 27488 13812 27490 13832
rect 27434 13776 27490 13812
rect 27710 14340 27766 14376
rect 27710 14320 27712 14340
rect 27712 14320 27764 14340
rect 27764 14320 27766 14340
rect 27158 9988 27214 10024
rect 27158 9968 27160 9988
rect 27160 9968 27212 9988
rect 27212 9968 27214 9988
rect 27802 11076 27858 11112
rect 27802 11056 27804 11076
rect 27804 11056 27856 11076
rect 27856 11056 27858 11076
rect 28262 18284 28318 18320
rect 28262 18264 28264 18284
rect 28264 18264 28316 18284
rect 28316 18264 28318 18284
rect 28170 15408 28226 15464
rect 27986 13640 28042 13696
rect 28538 24012 28540 24032
rect 28540 24012 28592 24032
rect 28592 24012 28594 24032
rect 28538 23976 28594 24012
rect 28814 18536 28870 18592
rect 28998 22752 29054 22808
rect 28998 17992 29054 18048
rect 27986 10804 28042 10840
rect 27986 10784 27988 10804
rect 27988 10784 28040 10804
rect 28040 10784 28042 10804
rect 27802 7248 27858 7304
rect 24030 3440 24086 3496
rect 28446 12416 28502 12472
rect 28630 12008 28686 12064
rect 28998 15136 29054 15192
rect 29366 27104 29422 27160
rect 28814 12688 28870 12744
rect 29274 11872 29330 11928
rect 32034 27920 32090 27976
rect 30930 26288 30986 26344
rect 30838 24520 30894 24576
rect 31666 25880 31722 25936
rect 29734 18808 29790 18864
rect 28814 7928 28870 7984
rect 29090 6840 29146 6896
rect 30378 22072 30434 22128
rect 30102 20576 30158 20632
rect 30378 20304 30434 20360
rect 29918 12300 29974 12336
rect 29918 12280 29920 12300
rect 29920 12280 29972 12300
rect 29972 12280 29974 12300
rect 31298 20032 31354 20088
rect 30930 18808 30986 18864
rect 30838 14764 30840 14784
rect 30840 14764 30892 14784
rect 30892 14764 30894 14784
rect 30838 14728 30894 14764
rect 31022 15020 31078 15056
rect 31022 15000 31024 15020
rect 31024 15000 31076 15020
rect 31076 15000 31078 15020
rect 30286 7520 30342 7576
rect 31942 25064 31998 25120
rect 31666 23840 31722 23896
rect 31666 7520 31722 7576
rect 32126 19352 32182 19408
rect 32494 23160 32550 23216
rect 32402 22480 32458 22536
rect 32494 21120 32550 21176
rect 32402 20440 32458 20496
rect 32402 19760 32458 19816
rect 32402 19080 32458 19136
rect 32402 17720 32458 17776
rect 32402 17060 32458 17096
rect 32402 17040 32404 17060
rect 32404 17040 32456 17060
rect 32456 17040 32458 17060
rect 32034 11464 32090 11520
rect 32402 15680 32458 15736
rect 32402 15000 32458 15056
rect 32402 13640 32458 13696
rect 32494 12960 32550 13016
rect 32402 11620 32458 11656
rect 32402 11600 32404 11620
rect 32404 11600 32456 11620
rect 32456 11600 32458 11620
rect 32678 17176 32734 17232
rect 32586 10376 32642 10432
rect 32402 10240 32458 10296
rect 32126 9560 32182 9616
rect 32310 9560 32366 9616
rect 32402 8200 32458 8256
rect 32310 6840 32366 6896
rect 32678 5480 32734 5536
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 974 31316 980 31380
rect 1044 31378 1050 31380
rect 20662 31378 20668 31380
rect 1044 31318 20668 31378
rect 1044 31316 1050 31318
rect 20662 31316 20668 31318
rect 20732 31316 20738 31380
rect 2078 31180 2084 31244
rect 2148 31242 2154 31244
rect 23105 31242 23171 31245
rect 2148 31240 23171 31242
rect 2148 31184 23110 31240
rect 23166 31184 23171 31240
rect 2148 31182 23171 31184
rect 2148 31180 2154 31182
rect 23105 31179 23171 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 14406 30908 14412 30972
rect 14476 30970 14482 30972
rect 23565 30970 23631 30973
rect 14476 30968 23631 30970
rect 14476 30912 23570 30968
rect 23626 30912 23631 30968
rect 14476 30910 23631 30912
rect 14476 30908 14482 30910
rect 23565 30907 23631 30910
rect 13721 30834 13787 30837
rect 30414 30834 30420 30836
rect 13721 30832 30420 30834
rect 13721 30776 13726 30832
rect 13782 30776 30420 30832
rect 13721 30774 30420 30776
rect 13721 30771 13787 30774
rect 30414 30772 30420 30774
rect 30484 30772 30490 30836
rect 15009 30562 15075 30565
rect 30598 30562 30604 30564
rect 15009 30560 30604 30562
rect 15009 30504 15014 30560
rect 15070 30504 30604 30560
rect 15009 30502 30604 30504
rect 15009 30499 15075 30502
rect 30598 30500 30604 30502
rect 30668 30500 30674 30564
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 6821 30426 6887 30429
rect 17902 30426 17908 30428
rect 6821 30424 17908 30426
rect 6821 30368 6826 30424
rect 6882 30368 17908 30424
rect 6821 30366 17908 30368
rect 6821 30363 6887 30366
rect 17902 30364 17908 30366
rect 17972 30364 17978 30428
rect 1117 30290 1183 30293
rect 23013 30290 23079 30293
rect 1117 30288 23079 30290
rect 1117 30232 1122 30288
rect 1178 30232 23018 30288
rect 23074 30232 23079 30288
rect 1117 30230 23079 30232
rect 1117 30227 1183 30230
rect 23013 30227 23079 30230
rect 606 30092 612 30156
rect 676 30154 682 30156
rect 15929 30154 15995 30157
rect 676 30152 15995 30154
rect 676 30096 15934 30152
rect 15990 30096 15995 30152
rect 676 30094 15995 30096
rect 676 30092 682 30094
rect 15929 30091 15995 30094
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 2630 29684 2636 29748
rect 2700 29746 2706 29748
rect 9673 29746 9739 29749
rect 2700 29744 9739 29746
rect 2700 29688 9678 29744
rect 9734 29688 9739 29744
rect 2700 29686 9739 29688
rect 2700 29684 2706 29686
rect 9673 29683 9739 29686
rect 1158 29548 1164 29612
rect 1228 29610 1234 29612
rect 7465 29610 7531 29613
rect 1228 29608 7531 29610
rect 1228 29552 7470 29608
rect 7526 29552 7531 29608
rect 1228 29550 7531 29552
rect 1228 29548 1234 29550
rect 7465 29547 7531 29550
rect 5390 29412 5396 29476
rect 5460 29474 5466 29476
rect 23197 29474 23263 29477
rect 5460 29472 23263 29474
rect 5460 29416 23202 29472
rect 23258 29416 23263 29472
rect 5460 29414 23263 29416
rect 5460 29412 5466 29414
rect 23197 29411 23263 29414
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 20161 29338 20227 29341
rect 29310 29338 29316 29340
rect 20161 29336 29316 29338
rect 20161 29280 20166 29336
rect 20222 29280 29316 29336
rect 20161 29278 29316 29280
rect 20161 29275 20227 29278
rect 29310 29276 29316 29278
rect 29380 29276 29386 29340
rect 2446 29140 2452 29204
rect 2516 29202 2522 29204
rect 9121 29202 9187 29205
rect 2516 29200 9187 29202
rect 2516 29144 9126 29200
rect 9182 29144 9187 29200
rect 2516 29142 9187 29144
rect 2516 29140 2522 29142
rect 9121 29139 9187 29142
rect 13997 29202 14063 29205
rect 27245 29202 27311 29205
rect 13997 29200 27311 29202
rect 13997 29144 14002 29200
rect 14058 29144 27250 29200
rect 27306 29144 27311 29200
rect 13997 29142 27311 29144
rect 13997 29139 14063 29142
rect 27245 29139 27311 29142
rect 4245 29010 4311 29013
rect 4064 29008 4311 29010
rect 4064 28952 4250 29008
rect 4306 28952 4311 29008
rect 8150 29004 8156 29068
rect 8220 29066 8226 29068
rect 9857 29066 9923 29069
rect 8220 29064 9923 29066
rect 8220 29008 9862 29064
rect 9918 29008 9923 29064
rect 8220 29006 9923 29008
rect 8220 29004 8226 29006
rect 9857 29003 9923 29006
rect 18137 29066 18203 29069
rect 18270 29066 18276 29068
rect 18137 29064 18276 29066
rect 18137 29008 18142 29064
rect 18198 29008 18276 29064
rect 18137 29006 18276 29008
rect 18137 29003 18203 29006
rect 18270 29004 18276 29006
rect 18340 29004 18346 29068
rect 21909 29066 21975 29069
rect 22185 29066 22251 29069
rect 21909 29064 22251 29066
rect 21909 29008 21914 29064
rect 21970 29008 22190 29064
rect 22246 29008 22251 29064
rect 21909 29006 22251 29008
rect 21909 29003 21975 29006
rect 22185 29003 22251 29006
rect 4064 28950 4311 28952
rect 3693 28930 3759 28933
rect 4064 28930 4124 28950
rect 4245 28947 4311 28950
rect 3693 28928 4124 28930
rect 3693 28872 3698 28928
rect 3754 28872 4124 28928
rect 3693 28870 4124 28872
rect 3693 28867 3759 28870
rect 6310 28868 6316 28932
rect 6380 28930 6386 28932
rect 9397 28930 9463 28933
rect 6380 28928 9463 28930
rect 6380 28872 9402 28928
rect 9458 28872 9463 28928
rect 6380 28870 9463 28872
rect 6380 28868 6386 28870
rect 9397 28867 9463 28870
rect 12525 28930 12591 28933
rect 20161 28930 20227 28933
rect 12525 28928 20227 28930
rect 12525 28872 12530 28928
rect 12586 28872 20166 28928
rect 20222 28872 20227 28928
rect 12525 28870 20227 28872
rect 12525 28867 12591 28870
rect 20161 28867 20227 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 6913 28794 6979 28797
rect 12934 28794 12940 28796
rect 6913 28792 12940 28794
rect 6913 28736 6918 28792
rect 6974 28736 12940 28792
rect 6913 28734 12940 28736
rect 6913 28731 6979 28734
rect 12934 28732 12940 28734
rect 13004 28794 13010 28796
rect 19517 28794 19583 28797
rect 13004 28792 19583 28794
rect 13004 28736 19522 28792
rect 19578 28736 19583 28792
rect 13004 28734 19583 28736
rect 13004 28732 13010 28734
rect 19517 28731 19583 28734
rect 0 28658 800 28688
rect 1393 28658 1459 28661
rect 0 28656 1459 28658
rect 0 28600 1398 28656
rect 1454 28600 1459 28656
rect 0 28598 1459 28600
rect 0 28568 800 28598
rect 1393 28595 1459 28598
rect 7414 28596 7420 28660
rect 7484 28658 7490 28660
rect 12341 28658 12407 28661
rect 7484 28656 12407 28658
rect 7484 28600 12346 28656
rect 12402 28600 12407 28656
rect 7484 28598 12407 28600
rect 7484 28596 7490 28598
rect 12341 28595 12407 28598
rect 12525 28658 12591 28661
rect 13169 28658 13235 28661
rect 12525 28656 13235 28658
rect 12525 28600 12530 28656
rect 12586 28600 13174 28656
rect 13230 28600 13235 28656
rect 12525 28598 13235 28600
rect 12525 28595 12591 28598
rect 13169 28595 13235 28598
rect 19609 28658 19675 28661
rect 23289 28658 23355 28661
rect 19609 28656 23355 28658
rect 19609 28600 19614 28656
rect 19670 28600 23294 28656
rect 23350 28600 23355 28656
rect 19609 28598 23355 28600
rect 19609 28595 19675 28598
rect 23289 28595 23355 28598
rect 7189 28522 7255 28525
rect 3374 28520 7255 28522
rect 3374 28464 7194 28520
rect 7250 28464 7255 28520
rect 3374 28462 7255 28464
rect 3374 28389 3434 28462
rect 7189 28459 7255 28462
rect 11053 28522 11119 28525
rect 22553 28522 22619 28525
rect 11053 28520 22619 28522
rect 11053 28464 11058 28520
rect 11114 28464 22558 28520
rect 22614 28464 22619 28520
rect 11053 28462 22619 28464
rect 11053 28459 11119 28462
rect 22553 28459 22619 28462
rect 3325 28388 3434 28389
rect 3325 28386 3372 28388
rect 3280 28384 3372 28386
rect 3280 28328 3330 28384
rect 3280 28326 3372 28328
rect 3325 28324 3372 28326
rect 3436 28324 3442 28388
rect 6494 28324 6500 28388
rect 6564 28386 6570 28388
rect 6729 28386 6795 28389
rect 6564 28384 6795 28386
rect 6564 28328 6734 28384
rect 6790 28328 6795 28384
rect 6564 28326 6795 28328
rect 6564 28324 6570 28326
rect 3325 28323 3391 28324
rect 6729 28323 6795 28326
rect 7189 28386 7255 28389
rect 9581 28386 9647 28389
rect 10133 28388 10199 28389
rect 10133 28386 10180 28388
rect 7189 28384 9647 28386
rect 7189 28328 7194 28384
rect 7250 28328 9586 28384
rect 9642 28328 9647 28384
rect 7189 28326 9647 28328
rect 10088 28384 10180 28386
rect 10088 28328 10138 28384
rect 10088 28326 10180 28328
rect 7189 28323 7255 28326
rect 9581 28323 9647 28326
rect 10133 28324 10180 28326
rect 10244 28324 10250 28388
rect 11329 28386 11395 28389
rect 14549 28386 14615 28389
rect 11329 28384 14615 28386
rect 11329 28328 11334 28384
rect 11390 28328 14554 28384
rect 14610 28328 14615 28384
rect 11329 28326 14615 28328
rect 10133 28323 10199 28324
rect 11329 28323 11395 28326
rect 14549 28323 14615 28326
rect 19333 28386 19399 28389
rect 20345 28386 20411 28389
rect 19333 28384 20411 28386
rect 19333 28328 19338 28384
rect 19394 28328 20350 28384
rect 20406 28328 20411 28384
rect 19333 28326 20411 28328
rect 19333 28323 19399 28326
rect 20345 28323 20411 28326
rect 20529 28386 20595 28389
rect 21030 28386 21036 28388
rect 20529 28384 21036 28386
rect 20529 28328 20534 28384
rect 20590 28328 21036 28384
rect 20529 28326 21036 28328
rect 20529 28323 20595 28326
rect 21030 28324 21036 28326
rect 21100 28324 21106 28388
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 11094 28188 11100 28252
rect 11164 28250 11170 28252
rect 13353 28250 13419 28253
rect 11164 28248 13419 28250
rect 11164 28192 13358 28248
rect 13414 28192 13419 28248
rect 11164 28190 13419 28192
rect 11164 28188 11170 28190
rect 13353 28187 13419 28190
rect 13486 28188 13492 28252
rect 13556 28250 13562 28252
rect 18413 28250 18479 28253
rect 25589 28250 25655 28253
rect 13556 28248 18479 28250
rect 13556 28192 18418 28248
rect 18474 28192 18479 28248
rect 13556 28190 18479 28192
rect 13556 28188 13562 28190
rect 18413 28187 18479 28190
rect 19290 28248 25655 28250
rect 19290 28192 25594 28248
rect 25650 28192 25655 28248
rect 19290 28190 25655 28192
rect 4613 28116 4679 28117
rect 4613 28112 4660 28116
rect 4724 28114 4730 28116
rect 10777 28114 10843 28117
rect 18137 28114 18203 28117
rect 4613 28056 4618 28112
rect 4613 28052 4660 28056
rect 4724 28054 4770 28114
rect 10777 28112 18203 28114
rect 10777 28056 10782 28112
rect 10838 28056 18142 28112
rect 18198 28056 18203 28112
rect 10777 28054 18203 28056
rect 4724 28052 4730 28054
rect 4613 28051 4679 28052
rect 10777 28051 10843 28054
rect 18137 28051 18203 28054
rect 0 27978 800 28008
rect 1485 27978 1551 27981
rect 0 27976 1551 27978
rect 0 27920 1490 27976
rect 1546 27920 1551 27976
rect 0 27918 1551 27920
rect 0 27888 800 27918
rect 1485 27915 1551 27918
rect 6862 27916 6868 27980
rect 6932 27978 6938 27980
rect 7741 27978 7807 27981
rect 6932 27976 7807 27978
rect 6932 27920 7746 27976
rect 7802 27920 7807 27976
rect 6932 27918 7807 27920
rect 6932 27916 6938 27918
rect 7741 27915 7807 27918
rect 9121 27978 9187 27981
rect 15009 27978 15075 27981
rect 19290 27978 19350 28190
rect 25589 28187 25655 28190
rect 20437 28114 20503 28117
rect 25957 28114 26023 28117
rect 20437 28112 26023 28114
rect 20437 28056 20442 28112
rect 20498 28056 25962 28112
rect 26018 28056 26023 28112
rect 20437 28054 26023 28056
rect 20437 28051 20503 28054
rect 25957 28051 26023 28054
rect 9121 27976 19350 27978
rect 9121 27920 9126 27976
rect 9182 27920 15014 27976
rect 15070 27920 19350 27976
rect 9121 27918 19350 27920
rect 21817 27978 21883 27981
rect 32029 27978 32095 27981
rect 21817 27976 32095 27978
rect 21817 27920 21822 27976
rect 21878 27920 32034 27976
rect 32090 27920 32095 27976
rect 21817 27918 32095 27920
rect 9121 27915 9187 27918
rect 15009 27915 15075 27918
rect 21817 27915 21883 27918
rect 32029 27915 32095 27918
rect 7465 27842 7531 27845
rect 9438 27842 9444 27844
rect 7465 27840 9444 27842
rect 7465 27784 7470 27840
rect 7526 27784 9444 27840
rect 7465 27782 9444 27784
rect 7465 27779 7531 27782
rect 9438 27780 9444 27782
rect 9508 27842 9514 27844
rect 10133 27842 10199 27845
rect 9508 27840 10199 27842
rect 9508 27784 10138 27840
rect 10194 27784 10199 27840
rect 9508 27782 10199 27784
rect 9508 27780 9514 27782
rect 10133 27779 10199 27782
rect 10593 27842 10659 27845
rect 10777 27842 10843 27845
rect 10593 27840 10843 27842
rect 10593 27784 10598 27840
rect 10654 27784 10782 27840
rect 10838 27784 10843 27840
rect 10593 27782 10843 27784
rect 10593 27779 10659 27782
rect 10777 27779 10843 27782
rect 11145 27842 11211 27845
rect 11278 27842 11284 27844
rect 11145 27840 11284 27842
rect 11145 27784 11150 27840
rect 11206 27784 11284 27840
rect 11145 27782 11284 27784
rect 11145 27779 11211 27782
rect 11278 27780 11284 27782
rect 11348 27780 11354 27844
rect 11881 27842 11947 27845
rect 12750 27842 12756 27844
rect 11881 27840 12756 27842
rect 11881 27784 11886 27840
rect 11942 27784 12756 27840
rect 11881 27782 12756 27784
rect 11881 27779 11947 27782
rect 12750 27780 12756 27782
rect 12820 27780 12826 27844
rect 14641 27842 14707 27845
rect 22093 27842 22159 27845
rect 23473 27842 23539 27845
rect 14641 27840 23539 27842
rect 14641 27784 14646 27840
rect 14702 27784 22098 27840
rect 22154 27784 23478 27840
rect 23534 27784 23539 27840
rect 14641 27782 23539 27784
rect 14641 27779 14707 27782
rect 22093 27779 22159 27782
rect 23473 27779 23539 27782
rect 25497 27842 25563 27845
rect 27838 27842 27844 27844
rect 25497 27840 27844 27842
rect 25497 27784 25502 27840
rect 25558 27784 27844 27840
rect 25497 27782 27844 27784
rect 25497 27779 25563 27782
rect 27838 27780 27844 27782
rect 27908 27780 27914 27844
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 6729 27706 6795 27709
rect 8017 27706 8083 27709
rect 6729 27704 8083 27706
rect 6729 27648 6734 27704
rect 6790 27648 8022 27704
rect 8078 27648 8083 27704
rect 6729 27646 8083 27648
rect 6729 27643 6795 27646
rect 8017 27643 8083 27646
rect 10225 27706 10291 27709
rect 11421 27706 11487 27709
rect 10225 27704 11487 27706
rect 10225 27648 10230 27704
rect 10286 27648 11426 27704
rect 11482 27648 11487 27704
rect 10225 27646 11487 27648
rect 10225 27643 10291 27646
rect 11421 27643 11487 27646
rect 11789 27706 11855 27709
rect 12249 27706 12315 27709
rect 11789 27704 12315 27706
rect 11789 27648 11794 27704
rect 11850 27648 12254 27704
rect 12310 27648 12315 27704
rect 11789 27646 12315 27648
rect 11789 27643 11855 27646
rect 12249 27643 12315 27646
rect 12566 27644 12572 27708
rect 12636 27706 12642 27708
rect 13905 27706 13971 27709
rect 15193 27708 15259 27709
rect 15142 27706 15148 27708
rect 12636 27704 13971 27706
rect 12636 27648 13910 27704
rect 13966 27648 13971 27704
rect 12636 27646 13971 27648
rect 15102 27646 15148 27706
rect 15212 27704 15259 27708
rect 15254 27648 15259 27704
rect 12636 27644 12642 27646
rect 13905 27643 13971 27646
rect 15142 27644 15148 27646
rect 15212 27644 15259 27648
rect 15193 27643 15259 27644
rect 16021 27708 16087 27709
rect 16021 27704 16068 27708
rect 16132 27706 16138 27708
rect 18597 27706 18663 27709
rect 20478 27706 20484 27708
rect 16021 27648 16026 27704
rect 16021 27644 16068 27648
rect 16132 27646 16178 27706
rect 18597 27704 20484 27706
rect 18597 27648 18602 27704
rect 18658 27648 20484 27704
rect 18597 27646 20484 27648
rect 16132 27644 16138 27646
rect 16021 27643 16087 27644
rect 18597 27643 18663 27646
rect 20478 27644 20484 27646
rect 20548 27644 20554 27708
rect 22093 27706 22159 27709
rect 22093 27704 22754 27706
rect 22093 27648 22098 27704
rect 22154 27648 22754 27704
rect 22093 27646 22754 27648
rect 22093 27643 22159 27646
rect 3693 27570 3759 27573
rect 7005 27570 7071 27573
rect 3693 27568 7071 27570
rect 3693 27512 3698 27568
rect 3754 27512 7010 27568
rect 7066 27512 7071 27568
rect 3693 27510 7071 27512
rect 3693 27507 3759 27510
rect 7005 27507 7071 27510
rect 11053 27570 11119 27573
rect 19149 27570 19215 27573
rect 11053 27568 19215 27570
rect 11053 27512 11058 27568
rect 11114 27512 19154 27568
rect 19210 27512 19215 27568
rect 11053 27510 19215 27512
rect 11053 27507 11119 27510
rect 19149 27507 19215 27510
rect 19374 27508 19380 27572
rect 19444 27570 19450 27572
rect 19977 27570 20043 27573
rect 19444 27568 20043 27570
rect 19444 27512 19982 27568
rect 20038 27512 20043 27568
rect 19444 27510 20043 27512
rect 19444 27508 19450 27510
rect 19977 27507 20043 27510
rect 22185 27570 22251 27573
rect 22502 27570 22508 27572
rect 22185 27568 22508 27570
rect 22185 27512 22190 27568
rect 22246 27512 22508 27568
rect 22185 27510 22508 27512
rect 22185 27507 22251 27510
rect 22502 27508 22508 27510
rect 22572 27508 22578 27572
rect 22694 27570 22754 27646
rect 23422 27644 23428 27708
rect 23492 27706 23498 27708
rect 23565 27706 23631 27709
rect 23492 27704 23631 27706
rect 23492 27648 23570 27704
rect 23626 27648 23631 27704
rect 23492 27646 23631 27648
rect 23492 27644 23498 27646
rect 23565 27643 23631 27646
rect 23982 27646 24778 27706
rect 23982 27570 24042 27646
rect 22694 27510 24042 27570
rect 24209 27570 24275 27573
rect 24526 27570 24532 27572
rect 24209 27568 24532 27570
rect 24209 27512 24214 27568
rect 24270 27512 24532 27568
rect 24209 27510 24532 27512
rect 24209 27507 24275 27510
rect 24526 27508 24532 27510
rect 24596 27508 24602 27572
rect 24718 27570 24778 27646
rect 27061 27570 27127 27573
rect 24718 27568 27127 27570
rect 24718 27512 27066 27568
rect 27122 27512 27127 27568
rect 24718 27510 27127 27512
rect 27061 27507 27127 27510
rect 6821 27434 6887 27437
rect 2730 27432 6887 27434
rect 2730 27376 6826 27432
rect 6882 27376 6887 27432
rect 2730 27374 6887 27376
rect 0 27298 800 27328
rect 2730 27298 2790 27374
rect 6821 27371 6887 27374
rect 7189 27436 7255 27437
rect 7189 27432 7236 27436
rect 7300 27434 7306 27436
rect 12341 27434 12407 27437
rect 12801 27434 12867 27437
rect 7189 27376 7194 27432
rect 7189 27372 7236 27376
rect 7300 27374 7346 27434
rect 12341 27432 12867 27434
rect 12341 27376 12346 27432
rect 12402 27376 12806 27432
rect 12862 27376 12867 27432
rect 12341 27374 12867 27376
rect 7300 27372 7306 27374
rect 7189 27371 7255 27372
rect 12341 27371 12407 27374
rect 12801 27371 12867 27374
rect 13721 27434 13787 27437
rect 15285 27434 15351 27437
rect 13721 27432 15351 27434
rect 13721 27376 13726 27432
rect 13782 27376 15290 27432
rect 15346 27376 15351 27432
rect 13721 27374 15351 27376
rect 13721 27371 13787 27374
rect 15285 27371 15351 27374
rect 16941 27434 17007 27437
rect 17953 27434 18019 27437
rect 16941 27432 18019 27434
rect 16941 27376 16946 27432
rect 17002 27376 17958 27432
rect 18014 27376 18019 27432
rect 16941 27374 18019 27376
rect 16941 27371 17007 27374
rect 17953 27371 18019 27374
rect 18505 27434 18571 27437
rect 19609 27434 19675 27437
rect 18505 27432 19675 27434
rect 18505 27376 18510 27432
rect 18566 27376 19614 27432
rect 19670 27376 19675 27432
rect 18505 27374 19675 27376
rect 18505 27371 18571 27374
rect 19609 27371 19675 27374
rect 19926 27372 19932 27436
rect 19996 27434 20002 27436
rect 20161 27434 20227 27437
rect 19996 27432 20227 27434
rect 19996 27376 20166 27432
rect 20222 27376 20227 27432
rect 19996 27374 20227 27376
rect 19996 27372 20002 27374
rect 20161 27371 20227 27374
rect 22001 27434 22067 27437
rect 23841 27434 23907 27437
rect 22001 27432 23907 27434
rect 22001 27376 22006 27432
rect 22062 27376 23846 27432
rect 23902 27376 23907 27432
rect 22001 27374 23907 27376
rect 22001 27371 22067 27374
rect 23841 27371 23907 27374
rect 0 27238 2790 27298
rect 5533 27298 5599 27301
rect 7005 27300 7071 27301
rect 7925 27300 7991 27301
rect 5533 27296 5826 27298
rect 5533 27240 5538 27296
rect 5594 27240 5826 27296
rect 5533 27238 5826 27240
rect 0 27208 800 27238
rect 5533 27235 5599 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 5349 27162 5415 27165
rect 5625 27162 5691 27165
rect 5349 27160 5691 27162
rect 5349 27104 5354 27160
rect 5410 27104 5630 27160
rect 5686 27104 5691 27160
rect 5349 27102 5691 27104
rect 5349 27099 5415 27102
rect 5625 27099 5691 27102
rect 4705 27026 4771 27029
rect 5766 27026 5826 27238
rect 7005 27296 7052 27300
rect 7116 27298 7122 27300
rect 7925 27298 7972 27300
rect 7005 27240 7010 27296
rect 7005 27236 7052 27240
rect 7116 27238 7162 27298
rect 7880 27296 7972 27298
rect 7880 27240 7930 27296
rect 7880 27238 7972 27240
rect 7116 27236 7122 27238
rect 7925 27236 7972 27238
rect 8036 27236 8042 27300
rect 9121 27298 9187 27301
rect 10225 27298 10291 27301
rect 9121 27296 10291 27298
rect 9121 27240 9126 27296
rect 9182 27240 10230 27296
rect 10286 27240 10291 27296
rect 9121 27238 10291 27240
rect 7005 27235 7071 27236
rect 7925 27235 7991 27236
rect 9121 27235 9187 27238
rect 10225 27235 10291 27238
rect 12249 27298 12315 27301
rect 18597 27298 18663 27301
rect 12249 27296 18663 27298
rect 12249 27240 12254 27296
rect 12310 27240 18602 27296
rect 18658 27240 18663 27296
rect 12249 27238 18663 27240
rect 12249 27235 12315 27238
rect 18597 27235 18663 27238
rect 18822 27236 18828 27300
rect 18892 27298 18898 27300
rect 19701 27298 19767 27301
rect 18892 27296 19767 27298
rect 18892 27240 19706 27296
rect 19762 27240 19767 27296
rect 18892 27238 19767 27240
rect 18892 27236 18898 27238
rect 19701 27235 19767 27238
rect 19885 27298 19951 27301
rect 19885 27296 27630 27298
rect 19885 27240 19890 27296
rect 19946 27240 27630 27296
rect 19885 27238 27630 27240
rect 19885 27235 19951 27238
rect 6821 27162 6887 27165
rect 11329 27162 11395 27165
rect 12709 27162 12775 27165
rect 15101 27162 15167 27165
rect 6821 27160 11395 27162
rect 6821 27104 6826 27160
rect 6882 27104 11334 27160
rect 11390 27104 11395 27160
rect 6821 27102 11395 27104
rect 6821 27099 6887 27102
rect 11329 27099 11395 27102
rect 11470 27160 12775 27162
rect 11470 27104 12714 27160
rect 12770 27104 12775 27160
rect 11470 27102 12775 27104
rect 4705 27024 5826 27026
rect 4705 26968 4710 27024
rect 4766 26968 5826 27024
rect 4705 26966 5826 26968
rect 4705 26963 4771 26966
rect 6126 26964 6132 27028
rect 6196 27026 6202 27028
rect 11470 27026 11530 27102
rect 12709 27099 12775 27102
rect 12988 27160 15167 27162
rect 12988 27104 15106 27160
rect 15162 27104 15167 27160
rect 12988 27102 15167 27104
rect 12988 27026 13048 27102
rect 15101 27099 15167 27102
rect 16113 27162 16179 27165
rect 22093 27162 22159 27165
rect 16113 27160 22159 27162
rect 16113 27104 16118 27160
rect 16174 27104 22098 27160
rect 22154 27104 22159 27160
rect 16113 27102 22159 27104
rect 27570 27162 27630 27238
rect 29361 27162 29427 27165
rect 27570 27160 29427 27162
rect 27570 27104 29366 27160
rect 29422 27104 29427 27160
rect 27570 27102 29427 27104
rect 16113 27099 16179 27102
rect 22093 27099 22159 27102
rect 29361 27099 29427 27102
rect 6196 26966 11530 27026
rect 12620 26966 13048 27026
rect 13169 27026 13235 27029
rect 13813 27026 13879 27029
rect 13169 27024 13879 27026
rect 13169 26968 13174 27024
rect 13230 26968 13818 27024
rect 13874 26968 13879 27024
rect 13169 26966 13879 26968
rect 6196 26964 6202 26966
rect 2589 26890 2655 26893
rect 6361 26890 6427 26893
rect 2589 26888 6427 26890
rect 2589 26832 2594 26888
rect 2650 26832 6366 26888
rect 6422 26832 6427 26888
rect 2589 26830 6427 26832
rect 2589 26827 2655 26830
rect 6361 26827 6427 26830
rect 9254 26828 9260 26892
rect 9324 26890 9330 26892
rect 11053 26890 11119 26893
rect 9324 26888 11119 26890
rect 9324 26832 11058 26888
rect 11114 26832 11119 26888
rect 9324 26830 11119 26832
rect 9324 26828 9330 26830
rect 11053 26827 11119 26830
rect 11237 26890 11303 26893
rect 12620 26890 12680 26966
rect 13169 26963 13235 26966
rect 13813 26963 13879 26966
rect 14365 27026 14431 27029
rect 19006 27026 19012 27028
rect 14365 27024 19012 27026
rect 14365 26968 14370 27024
rect 14426 26968 19012 27024
rect 14365 26966 19012 26968
rect 14365 26963 14431 26966
rect 19006 26964 19012 26966
rect 19076 26964 19082 27028
rect 19149 27026 19215 27029
rect 21817 27026 21883 27029
rect 29862 27026 29868 27028
rect 19149 27024 21883 27026
rect 19149 26968 19154 27024
rect 19210 26968 21822 27024
rect 21878 26968 21883 27024
rect 19149 26966 21883 26968
rect 19149 26963 19215 26966
rect 21817 26963 21883 26966
rect 22510 26966 29868 27026
rect 11237 26888 12680 26890
rect 11237 26832 11242 26888
rect 11298 26832 12680 26888
rect 11237 26830 12680 26832
rect 11237 26827 11303 26830
rect 12750 26828 12756 26892
rect 12820 26890 12826 26892
rect 18822 26890 18828 26892
rect 12820 26830 18828 26890
rect 12820 26828 12826 26830
rect 18822 26828 18828 26830
rect 18892 26828 18898 26892
rect 20161 26890 20227 26893
rect 19428 26888 20227 26890
rect 19428 26832 20166 26888
rect 20222 26832 20227 26888
rect 19428 26830 20227 26832
rect 8477 26754 8543 26757
rect 14273 26754 14339 26757
rect 8477 26752 14339 26754
rect 8477 26696 8482 26752
rect 8538 26696 14278 26752
rect 14334 26696 14339 26752
rect 8477 26694 14339 26696
rect 8477 26691 8543 26694
rect 14273 26691 14339 26694
rect 14457 26754 14523 26757
rect 18505 26754 18571 26757
rect 14457 26752 18571 26754
rect 14457 26696 14462 26752
rect 14518 26696 18510 26752
rect 18566 26696 18571 26752
rect 14457 26694 18571 26696
rect 14457 26691 14523 26694
rect 18505 26691 18571 26694
rect 18781 26754 18847 26757
rect 19428 26754 19488 26830
rect 20161 26827 20227 26830
rect 20621 26890 20687 26893
rect 21398 26890 21404 26892
rect 20621 26888 21404 26890
rect 20621 26832 20626 26888
rect 20682 26832 21404 26888
rect 20621 26830 21404 26832
rect 20621 26827 20687 26830
rect 21398 26828 21404 26830
rect 21468 26828 21474 26892
rect 18781 26752 19488 26754
rect 18781 26696 18786 26752
rect 18842 26696 19488 26752
rect 18781 26694 19488 26696
rect 18781 26691 18847 26694
rect 19558 26692 19564 26756
rect 19628 26754 19634 26756
rect 22510 26754 22570 26966
rect 29862 26964 29868 26966
rect 29932 26964 29938 27028
rect 19628 26694 22570 26754
rect 22737 26754 22803 26757
rect 30782 26754 30788 26756
rect 22737 26752 30788 26754
rect 22737 26696 22742 26752
rect 22798 26696 30788 26752
rect 22737 26694 30788 26696
rect 19628 26692 19634 26694
rect 22737 26691 22803 26694
rect 30782 26692 30788 26694
rect 30852 26692 30858 26756
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 6177 26618 6243 26621
rect 9581 26618 9647 26621
rect 6177 26616 9647 26618
rect 6177 26560 6182 26616
rect 6238 26560 9586 26616
rect 9642 26560 9647 26616
rect 6177 26558 9647 26560
rect 6177 26555 6243 26558
rect 9581 26555 9647 26558
rect 9765 26618 9831 26621
rect 10777 26618 10843 26621
rect 9765 26616 10843 26618
rect 9765 26560 9770 26616
rect 9826 26560 10782 26616
rect 10838 26560 10843 26616
rect 9765 26558 10843 26560
rect 9765 26555 9831 26558
rect 10777 26555 10843 26558
rect 12985 26618 13051 26621
rect 13302 26618 13308 26620
rect 12985 26616 13308 26618
rect 12985 26560 12990 26616
rect 13046 26560 13308 26616
rect 12985 26558 13308 26560
rect 12985 26555 13051 26558
rect 13302 26556 13308 26558
rect 13372 26618 13378 26620
rect 15009 26618 15075 26621
rect 27705 26618 27771 26621
rect 13372 26616 27771 26618
rect 13372 26560 15014 26616
rect 15070 26560 27710 26616
rect 27766 26560 27771 26616
rect 13372 26558 27771 26560
rect 13372 26556 13378 26558
rect 15009 26555 15075 26558
rect 27705 26555 27771 26558
rect 5533 26484 5599 26485
rect 5533 26482 5580 26484
rect 5488 26480 5580 26482
rect 5488 26424 5538 26480
rect 5488 26422 5580 26424
rect 5533 26420 5580 26422
rect 5644 26420 5650 26484
rect 5942 26420 5948 26484
rect 6012 26482 6018 26484
rect 16021 26482 16087 26485
rect 6012 26480 16087 26482
rect 6012 26424 16026 26480
rect 16082 26424 16087 26480
rect 6012 26422 16087 26424
rect 6012 26420 6018 26422
rect 5533 26419 5599 26420
rect 16021 26419 16087 26422
rect 16297 26482 16363 26485
rect 25589 26482 25655 26485
rect 26969 26484 27035 26485
rect 16297 26480 25655 26482
rect 16297 26424 16302 26480
rect 16358 26424 25594 26480
rect 25650 26424 25655 26480
rect 16297 26422 25655 26424
rect 16297 26419 16363 26422
rect 25589 26419 25655 26422
rect 26918 26420 26924 26484
rect 26988 26482 27035 26484
rect 26988 26480 27080 26482
rect 27030 26424 27080 26480
rect 26988 26422 27080 26424
rect 26988 26420 27035 26422
rect 26969 26419 27035 26420
rect 13445 26346 13511 26349
rect 17769 26348 17835 26349
rect 17718 26346 17724 26348
rect 8710 26344 13511 26346
rect 8710 26288 13450 26344
rect 13506 26288 13511 26344
rect 8710 26286 13511 26288
rect 17678 26286 17724 26346
rect 17788 26344 17835 26348
rect 17830 26288 17835 26344
rect 5349 26210 5415 26213
rect 5717 26210 5783 26213
rect 5349 26208 5783 26210
rect 5349 26152 5354 26208
rect 5410 26152 5722 26208
rect 5778 26152 5783 26208
rect 5349 26150 5783 26152
rect 5349 26147 5415 26150
rect 5717 26147 5783 26150
rect 6085 26210 6151 26213
rect 6637 26210 6703 26213
rect 6085 26208 6703 26210
rect 6085 26152 6090 26208
rect 6146 26152 6642 26208
rect 6698 26152 6703 26208
rect 6085 26150 6703 26152
rect 6085 26147 6151 26150
rect 6637 26147 6703 26150
rect 8569 26210 8635 26213
rect 8710 26212 8770 26286
rect 13445 26283 13511 26286
rect 17718 26284 17724 26286
rect 17788 26284 17835 26288
rect 17769 26283 17835 26284
rect 19149 26346 19215 26349
rect 21173 26348 21239 26349
rect 19149 26344 21098 26346
rect 19149 26288 19154 26344
rect 19210 26288 21098 26344
rect 19149 26286 21098 26288
rect 19149 26283 19215 26286
rect 8702 26210 8708 26212
rect 8569 26208 8708 26210
rect 8569 26152 8574 26208
rect 8630 26152 8708 26208
rect 8569 26150 8708 26152
rect 8569 26147 8635 26150
rect 8702 26148 8708 26150
rect 8772 26148 8778 26212
rect 10174 26148 10180 26212
rect 10244 26210 10250 26212
rect 10501 26210 10567 26213
rect 10244 26208 10567 26210
rect 10244 26152 10506 26208
rect 10562 26152 10567 26208
rect 10244 26150 10567 26152
rect 10244 26148 10250 26150
rect 10501 26147 10567 26150
rect 14825 26210 14891 26213
rect 20253 26210 20319 26213
rect 14825 26208 20319 26210
rect 14825 26152 14830 26208
rect 14886 26152 20258 26208
rect 20314 26152 20319 26208
rect 14825 26150 20319 26152
rect 21038 26210 21098 26286
rect 21173 26344 21220 26348
rect 21284 26346 21290 26348
rect 22737 26346 22803 26349
rect 21173 26288 21178 26344
rect 21173 26284 21220 26288
rect 21284 26286 21330 26346
rect 21406 26344 22803 26346
rect 21406 26288 22742 26344
rect 22798 26288 22803 26344
rect 21406 26286 22803 26288
rect 21284 26284 21290 26286
rect 21173 26283 21239 26284
rect 21406 26210 21466 26286
rect 22737 26283 22803 26286
rect 24894 26284 24900 26348
rect 24964 26346 24970 26348
rect 30925 26346 30991 26349
rect 24964 26344 30991 26346
rect 24964 26288 30930 26344
rect 30986 26288 30991 26344
rect 24964 26286 30991 26288
rect 24964 26284 24970 26286
rect 30925 26283 30991 26286
rect 21038 26150 21466 26210
rect 21909 26210 21975 26213
rect 26182 26210 26188 26212
rect 21909 26208 26188 26210
rect 21909 26152 21914 26208
rect 21970 26152 26188 26208
rect 21909 26150 26188 26152
rect 14825 26147 14891 26150
rect 20253 26147 20319 26150
rect 21909 26147 21975 26150
rect 26182 26148 26188 26150
rect 26252 26148 26258 26212
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 5901 26074 5967 26077
rect 5398 26072 5967 26074
rect 5398 26016 5906 26072
rect 5962 26016 5967 26072
rect 5398 26014 5967 26016
rect 0 25938 800 25968
rect 4981 25938 5047 25941
rect 5398 25938 5458 26014
rect 5901 26011 5967 26014
rect 7741 26074 7807 26077
rect 13353 26074 13419 26077
rect 7741 26072 13419 26074
rect 7741 26016 7746 26072
rect 7802 26016 13358 26072
rect 13414 26016 13419 26072
rect 7741 26014 13419 26016
rect 7741 26011 7807 26014
rect 13353 26011 13419 26014
rect 14641 26074 14707 26077
rect 16757 26074 16823 26077
rect 14641 26072 16823 26074
rect 14641 26016 14646 26072
rect 14702 26016 16762 26072
rect 16818 26016 16823 26072
rect 14641 26014 16823 26016
rect 14641 26011 14707 26014
rect 16757 26011 16823 26014
rect 19517 26074 19583 26077
rect 20437 26074 20503 26077
rect 26325 26074 26391 26077
rect 19517 26072 26391 26074
rect 19517 26016 19522 26072
rect 19578 26016 20442 26072
rect 20498 26016 26330 26072
rect 26386 26016 26391 26072
rect 19517 26014 26391 26016
rect 19517 26011 19583 26014
rect 20437 26011 20503 26014
rect 26325 26011 26391 26014
rect 0 25848 858 25938
rect 4981 25936 5458 25938
rect 4981 25880 4986 25936
rect 5042 25880 5458 25936
rect 4981 25878 5458 25880
rect 12249 25938 12315 25941
rect 15929 25938 15995 25941
rect 12249 25936 15995 25938
rect 12249 25880 12254 25936
rect 12310 25880 15934 25936
rect 15990 25880 15995 25936
rect 12249 25878 15995 25880
rect 4981 25875 5047 25878
rect 12249 25875 12315 25878
rect 15929 25875 15995 25878
rect 16941 25938 17007 25941
rect 19374 25938 19380 25940
rect 16941 25936 19380 25938
rect 16941 25880 16946 25936
rect 17002 25880 19380 25936
rect 16941 25878 19380 25880
rect 16941 25875 17007 25878
rect 19374 25876 19380 25878
rect 19444 25876 19450 25940
rect 19609 25938 19675 25941
rect 19742 25938 19748 25940
rect 19609 25936 19748 25938
rect 19609 25880 19614 25936
rect 19670 25880 19748 25936
rect 19609 25878 19748 25880
rect 19609 25875 19675 25878
rect 19742 25876 19748 25878
rect 19812 25876 19818 25940
rect 19885 25938 19951 25941
rect 25814 25938 25820 25940
rect 19885 25936 25820 25938
rect 19885 25880 19890 25936
rect 19946 25880 25820 25936
rect 19885 25878 25820 25880
rect 19885 25875 19951 25878
rect 25814 25876 25820 25878
rect 25884 25938 25890 25940
rect 27245 25938 27311 25941
rect 25884 25936 27311 25938
rect 25884 25880 27250 25936
rect 27306 25880 27311 25936
rect 25884 25878 27311 25880
rect 25884 25876 25890 25878
rect 27245 25875 27311 25878
rect 31661 25938 31727 25941
rect 33200 25938 34000 25968
rect 31661 25936 34000 25938
rect 31661 25880 31666 25936
rect 31722 25880 34000 25936
rect 31661 25878 34000 25880
rect 31661 25875 31727 25878
rect 33200 25848 34000 25878
rect 798 25805 858 25848
rect 798 25800 907 25805
rect 798 25744 846 25800
rect 902 25744 907 25800
rect 798 25742 907 25744
rect 841 25739 907 25742
rect 2129 25802 2195 25805
rect 7097 25802 7163 25805
rect 2129 25800 7163 25802
rect 2129 25744 2134 25800
rect 2190 25744 7102 25800
rect 7158 25744 7163 25800
rect 2129 25742 7163 25744
rect 2129 25739 2195 25742
rect 7097 25739 7163 25742
rect 10961 25802 11027 25805
rect 20989 25802 21055 25805
rect 10961 25800 21055 25802
rect 10961 25744 10966 25800
rect 11022 25744 20994 25800
rect 21050 25744 21055 25800
rect 10961 25742 21055 25744
rect 10961 25739 11027 25742
rect 20989 25739 21055 25742
rect 21357 25802 21423 25805
rect 21766 25802 21772 25804
rect 21357 25800 21772 25802
rect 21357 25744 21362 25800
rect 21418 25744 21772 25800
rect 21357 25742 21772 25744
rect 21357 25739 21423 25742
rect 21766 25740 21772 25742
rect 21836 25740 21842 25804
rect 23473 25802 23539 25805
rect 25129 25802 25195 25805
rect 23473 25800 25195 25802
rect 23473 25744 23478 25800
rect 23534 25744 25134 25800
rect 25190 25744 25195 25800
rect 23473 25742 25195 25744
rect 23473 25739 23539 25742
rect 25129 25739 25195 25742
rect 5073 25666 5139 25669
rect 5758 25666 5764 25668
rect 5073 25664 5764 25666
rect 5073 25608 5078 25664
rect 5134 25608 5764 25664
rect 5073 25606 5764 25608
rect 5073 25603 5139 25606
rect 5758 25604 5764 25606
rect 5828 25666 5834 25668
rect 5901 25666 5967 25669
rect 7230 25666 7236 25668
rect 5828 25664 7236 25666
rect 5828 25608 5906 25664
rect 5962 25608 7236 25664
rect 5828 25606 7236 25608
rect 5828 25604 5834 25606
rect 5901 25603 5967 25606
rect 7230 25604 7236 25606
rect 7300 25604 7306 25668
rect 16849 25666 16915 25669
rect 12390 25664 16915 25666
rect 12390 25608 16854 25664
rect 16910 25608 16915 25664
rect 12390 25606 16915 25608
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 12390 25532 12450 25606
rect 16849 25603 16915 25606
rect 17033 25666 17099 25669
rect 17493 25666 17559 25669
rect 17033 25664 17559 25666
rect 17033 25608 17038 25664
rect 17094 25608 17498 25664
rect 17554 25608 17559 25664
rect 17033 25606 17559 25608
rect 17033 25603 17099 25606
rect 17493 25603 17559 25606
rect 19374 25604 19380 25668
rect 19444 25666 19450 25668
rect 26785 25666 26851 25669
rect 19444 25664 26851 25666
rect 19444 25608 26790 25664
rect 26846 25608 26851 25664
rect 19444 25606 26851 25608
rect 19444 25604 19450 25606
rect 26785 25603 26851 25606
rect 12382 25530 12388 25532
rect 4662 25470 12388 25530
rect 1761 25122 1827 25125
rect 4662 25122 4722 25470
rect 12382 25468 12388 25470
rect 12452 25468 12458 25532
rect 14457 25530 14523 25533
rect 19149 25530 19215 25533
rect 14457 25528 19215 25530
rect 14457 25472 14462 25528
rect 14518 25472 19154 25528
rect 19210 25472 19215 25528
rect 14457 25470 19215 25472
rect 14457 25467 14523 25470
rect 19149 25467 19215 25470
rect 19333 25530 19399 25533
rect 28942 25530 28948 25532
rect 19333 25528 28948 25530
rect 19333 25472 19338 25528
rect 19394 25472 28948 25528
rect 19333 25470 28948 25472
rect 19333 25467 19399 25470
rect 28942 25468 28948 25470
rect 29012 25468 29018 25532
rect 9581 25394 9647 25397
rect 12433 25394 12499 25397
rect 13721 25396 13787 25397
rect 9581 25392 12499 25394
rect 9581 25336 9586 25392
rect 9642 25336 12438 25392
rect 12494 25336 12499 25392
rect 9581 25334 12499 25336
rect 9581 25331 9647 25334
rect 12433 25331 12499 25334
rect 13670 25332 13676 25396
rect 13740 25394 13787 25396
rect 14917 25394 14983 25397
rect 16982 25394 16988 25396
rect 13740 25392 13832 25394
rect 13782 25336 13832 25392
rect 13740 25334 13832 25336
rect 14917 25392 16988 25394
rect 14917 25336 14922 25392
rect 14978 25336 16988 25392
rect 14917 25334 16988 25336
rect 13740 25332 13787 25334
rect 13721 25331 13787 25332
rect 14917 25331 14983 25334
rect 16982 25332 16988 25334
rect 17052 25394 17058 25396
rect 20253 25394 20319 25397
rect 17052 25392 20319 25394
rect 17052 25336 20258 25392
rect 20314 25336 20319 25392
rect 17052 25334 20319 25336
rect 17052 25332 17058 25334
rect 20253 25331 20319 25334
rect 20529 25394 20595 25397
rect 23749 25394 23815 25397
rect 26601 25394 26667 25397
rect 20529 25392 26667 25394
rect 20529 25336 20534 25392
rect 20590 25336 23754 25392
rect 23810 25336 26606 25392
rect 26662 25336 26667 25392
rect 20529 25334 26667 25336
rect 20529 25331 20595 25334
rect 23749 25331 23815 25334
rect 26601 25331 26667 25334
rect 8661 25258 8727 25261
rect 9765 25258 9831 25261
rect 8661 25256 9831 25258
rect 8661 25200 8666 25256
rect 8722 25200 9770 25256
rect 9826 25200 9831 25256
rect 8661 25198 9831 25200
rect 8661 25195 8727 25198
rect 9765 25195 9831 25198
rect 10542 25196 10548 25260
rect 10612 25258 10618 25260
rect 14825 25258 14891 25261
rect 10612 25256 14891 25258
rect 10612 25200 14830 25256
rect 14886 25200 14891 25256
rect 10612 25198 14891 25200
rect 10612 25196 10618 25198
rect 14825 25195 14891 25198
rect 15193 25258 15259 25261
rect 21909 25258 21975 25261
rect 15193 25256 21975 25258
rect 15193 25200 15198 25256
rect 15254 25200 21914 25256
rect 21970 25200 21975 25256
rect 15193 25198 21975 25200
rect 15193 25195 15259 25198
rect 21909 25195 21975 25198
rect 22645 25258 22711 25261
rect 26233 25258 26299 25261
rect 22645 25256 26299 25258
rect 22645 25200 22650 25256
rect 22706 25200 26238 25256
rect 26294 25200 26299 25256
rect 22645 25198 26299 25200
rect 22645 25195 22711 25198
rect 26233 25195 26299 25198
rect 26366 25196 26372 25260
rect 26436 25258 26442 25260
rect 26785 25258 26851 25261
rect 26436 25256 26851 25258
rect 26436 25200 26790 25256
rect 26846 25200 26851 25256
rect 26436 25198 26851 25200
rect 26436 25196 26442 25198
rect 26785 25195 26851 25198
rect 1761 25120 4722 25122
rect 1761 25064 1766 25120
rect 1822 25064 4722 25120
rect 1761 25062 4722 25064
rect 6821 25122 6887 25125
rect 8201 25122 8267 25125
rect 6821 25120 8267 25122
rect 6821 25064 6826 25120
rect 6882 25064 8206 25120
rect 8262 25064 8267 25120
rect 6821 25062 8267 25064
rect 1761 25059 1827 25062
rect 6821 25059 6887 25062
rect 8201 25059 8267 25062
rect 9397 25122 9463 25125
rect 10685 25122 10751 25125
rect 9397 25120 10751 25122
rect 9397 25064 9402 25120
rect 9458 25064 10690 25120
rect 10746 25064 10751 25120
rect 9397 25062 10751 25064
rect 9397 25059 9463 25062
rect 10685 25059 10751 25062
rect 14181 25122 14247 25125
rect 16614 25122 16620 25124
rect 14181 25120 16620 25122
rect 14181 25064 14186 25120
rect 14242 25064 16620 25120
rect 14181 25062 16620 25064
rect 14181 25059 14247 25062
rect 16614 25060 16620 25062
rect 16684 25060 16690 25124
rect 16757 25122 16823 25125
rect 25129 25122 25195 25125
rect 31937 25122 32003 25125
rect 16757 25120 25195 25122
rect 16757 25064 16762 25120
rect 16818 25064 25134 25120
rect 25190 25064 25195 25120
rect 16757 25062 25195 25064
rect 16757 25059 16823 25062
rect 25129 25059 25195 25062
rect 25270 25120 32003 25122
rect 25270 25064 31942 25120
rect 31998 25064 32003 25120
rect 25270 25062 32003 25064
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 9438 24924 9444 24988
rect 9508 24986 9514 24988
rect 9857 24986 9923 24989
rect 10501 24986 10567 24989
rect 9508 24984 10567 24986
rect 9508 24928 9862 24984
rect 9918 24928 10506 24984
rect 10562 24928 10567 24984
rect 9508 24926 10567 24928
rect 9508 24924 9514 24926
rect 9857 24923 9923 24926
rect 10501 24923 10567 24926
rect 11094 24924 11100 24988
rect 11164 24986 11170 24988
rect 13261 24986 13327 24989
rect 11164 24984 13327 24986
rect 11164 24928 13266 24984
rect 13322 24928 13327 24984
rect 11164 24926 13327 24928
rect 11164 24924 11170 24926
rect 13261 24923 13327 24926
rect 15377 24986 15443 24989
rect 15878 24986 15884 24988
rect 15377 24984 15884 24986
rect 15377 24928 15382 24984
rect 15438 24928 15884 24984
rect 15377 24926 15884 24928
rect 15377 24923 15443 24926
rect 15878 24924 15884 24926
rect 15948 24924 15954 24988
rect 19701 24986 19767 24989
rect 16024 24984 19767 24986
rect 16024 24928 19706 24984
rect 19762 24928 19767 24984
rect 16024 24926 19767 24928
rect 3734 24788 3740 24852
rect 3804 24850 3810 24852
rect 4337 24850 4403 24853
rect 8109 24850 8175 24853
rect 3804 24848 8175 24850
rect 3804 24792 4342 24848
rect 4398 24792 8114 24848
rect 8170 24792 8175 24848
rect 3804 24790 8175 24792
rect 3804 24788 3810 24790
rect 4337 24787 4403 24790
rect 8109 24787 8175 24790
rect 9213 24850 9279 24853
rect 9806 24850 9812 24852
rect 9213 24848 9812 24850
rect 9213 24792 9218 24848
rect 9274 24792 9812 24848
rect 9213 24790 9812 24792
rect 9213 24787 9279 24790
rect 9806 24788 9812 24790
rect 9876 24788 9882 24852
rect 10133 24850 10199 24853
rect 14549 24850 14615 24853
rect 10133 24848 14615 24850
rect 10133 24792 10138 24848
rect 10194 24792 14554 24848
rect 14610 24792 14615 24848
rect 10133 24790 14615 24792
rect 10133 24787 10199 24790
rect 14549 24787 14615 24790
rect 15469 24850 15535 24853
rect 15837 24850 15903 24853
rect 16024 24850 16084 24926
rect 19701 24923 19767 24926
rect 20253 24986 20319 24989
rect 20662 24986 20668 24988
rect 20253 24984 20668 24986
rect 20253 24928 20258 24984
rect 20314 24928 20668 24984
rect 20253 24926 20668 24928
rect 20253 24923 20319 24926
rect 20662 24924 20668 24926
rect 20732 24924 20738 24988
rect 20846 24924 20852 24988
rect 20916 24986 20922 24988
rect 21449 24986 21515 24989
rect 20916 24984 21515 24986
rect 20916 24928 21454 24984
rect 21510 24928 21515 24984
rect 20916 24926 21515 24928
rect 20916 24924 20922 24926
rect 21449 24923 21515 24926
rect 24301 24986 24367 24989
rect 25270 24986 25330 25062
rect 31937 25059 32003 25062
rect 24301 24984 25330 24986
rect 24301 24928 24306 24984
rect 24362 24928 25330 24984
rect 24301 24926 25330 24928
rect 26785 24986 26851 24989
rect 28574 24986 28580 24988
rect 26785 24984 28580 24986
rect 26785 24928 26790 24984
rect 26846 24928 28580 24984
rect 26785 24926 28580 24928
rect 24301 24923 24367 24926
rect 26785 24923 26851 24926
rect 28574 24924 28580 24926
rect 28644 24924 28650 24988
rect 15469 24848 16084 24850
rect 15469 24792 15474 24848
rect 15530 24792 15842 24848
rect 15898 24792 16084 24848
rect 15469 24790 16084 24792
rect 17493 24850 17559 24853
rect 28257 24850 28323 24853
rect 17493 24848 28323 24850
rect 17493 24792 17498 24848
rect 17554 24792 28262 24848
rect 28318 24792 28323 24848
rect 17493 24790 28323 24792
rect 15469 24787 15535 24790
rect 15837 24787 15903 24790
rect 17493 24787 17559 24790
rect 28257 24787 28323 24790
rect 381 24714 447 24717
rect 12341 24714 12407 24717
rect 381 24712 12407 24714
rect 381 24656 386 24712
rect 442 24656 12346 24712
rect 12402 24656 12407 24712
rect 381 24654 12407 24656
rect 381 24651 447 24654
rect 12341 24651 12407 24654
rect 13261 24714 13327 24717
rect 16941 24714 17007 24717
rect 17953 24714 18019 24717
rect 13261 24712 17007 24714
rect 13261 24656 13266 24712
rect 13322 24656 16946 24712
rect 17002 24656 17007 24712
rect 13261 24654 17007 24656
rect 13261 24651 13327 24654
rect 16941 24651 17007 24654
rect 17128 24712 18019 24714
rect 17128 24656 17958 24712
rect 18014 24656 18019 24712
rect 17128 24654 18019 24656
rect 8661 24578 8727 24581
rect 9489 24578 9555 24581
rect 8661 24576 9555 24578
rect 8661 24520 8666 24576
rect 8722 24520 9494 24576
rect 9550 24520 9555 24576
rect 8661 24518 9555 24520
rect 8661 24515 8727 24518
rect 9489 24515 9555 24518
rect 9765 24578 9831 24581
rect 13445 24578 13511 24581
rect 17128 24578 17188 24654
rect 17953 24651 18019 24654
rect 19241 24712 19307 24717
rect 19241 24656 19246 24712
rect 19302 24656 19307 24712
rect 19241 24651 19307 24656
rect 19425 24714 19491 24717
rect 19558 24714 19564 24716
rect 19425 24712 19564 24714
rect 19425 24656 19430 24712
rect 19486 24656 19564 24712
rect 19425 24654 19564 24656
rect 19425 24651 19491 24654
rect 19558 24652 19564 24654
rect 19628 24652 19634 24716
rect 19793 24714 19859 24717
rect 22277 24714 22343 24717
rect 19793 24712 22343 24714
rect 19793 24656 19798 24712
rect 19854 24656 22282 24712
rect 22338 24656 22343 24712
rect 19793 24654 22343 24656
rect 19793 24651 19859 24654
rect 22277 24651 22343 24654
rect 23013 24714 23079 24717
rect 23381 24714 23447 24717
rect 23013 24712 23447 24714
rect 23013 24656 23018 24712
rect 23074 24656 23386 24712
rect 23442 24656 23447 24712
rect 23013 24654 23447 24656
rect 23013 24651 23079 24654
rect 23381 24651 23447 24654
rect 9765 24576 13511 24578
rect 9765 24520 9770 24576
rect 9826 24520 13450 24576
rect 13506 24520 13511 24576
rect 9765 24518 13511 24520
rect 9765 24515 9831 24518
rect 13445 24515 13511 24518
rect 13678 24518 17188 24578
rect 17401 24578 17467 24581
rect 19244 24578 19304 24651
rect 20662 24578 20668 24580
rect 17401 24576 20668 24578
rect 17401 24520 17406 24576
rect 17462 24520 20668 24576
rect 17401 24518 20668 24520
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 9029 24442 9095 24445
rect 9673 24442 9739 24445
rect 9029 24440 9739 24442
rect 9029 24384 9034 24440
rect 9090 24384 9678 24440
rect 9734 24384 9739 24440
rect 9029 24382 9739 24384
rect 9029 24379 9095 24382
rect 9673 24379 9739 24382
rect 12893 24442 12959 24445
rect 13678 24442 13738 24518
rect 17401 24515 17467 24518
rect 20662 24516 20668 24518
rect 20732 24516 20738 24580
rect 21357 24578 21423 24581
rect 22093 24578 22159 24581
rect 21357 24576 22159 24578
rect 21357 24520 21362 24576
rect 21418 24520 22098 24576
rect 22154 24520 22159 24576
rect 21357 24518 22159 24520
rect 21357 24515 21423 24518
rect 22093 24515 22159 24518
rect 30833 24578 30899 24581
rect 33200 24578 34000 24608
rect 30833 24576 34000 24578
rect 30833 24520 30838 24576
rect 30894 24520 34000 24576
rect 30833 24518 34000 24520
rect 30833 24515 30899 24518
rect 33200 24488 34000 24518
rect 12893 24440 13738 24442
rect 12893 24384 12898 24440
rect 12954 24384 13738 24440
rect 12893 24382 13738 24384
rect 14273 24442 14339 24445
rect 24485 24442 24551 24445
rect 14273 24440 24551 24442
rect 14273 24384 14278 24440
rect 14334 24384 24490 24440
rect 24546 24384 24551 24440
rect 14273 24382 24551 24384
rect 12893 24379 12959 24382
rect 14273 24379 14339 24382
rect 24485 24379 24551 24382
rect 5257 24306 5323 24309
rect 7414 24306 7420 24308
rect 5257 24304 7420 24306
rect 5257 24248 5262 24304
rect 5318 24248 7420 24304
rect 5257 24246 7420 24248
rect 5257 24243 5323 24246
rect 7414 24244 7420 24246
rect 7484 24244 7490 24308
rect 8845 24306 8911 24309
rect 13118 24306 13124 24308
rect 8845 24304 13124 24306
rect 8845 24248 8850 24304
rect 8906 24248 13124 24304
rect 8845 24246 13124 24248
rect 8845 24243 8911 24246
rect 13118 24244 13124 24246
rect 13188 24306 13194 24308
rect 20846 24306 20852 24308
rect 13188 24246 20852 24306
rect 13188 24244 13194 24246
rect 20846 24244 20852 24246
rect 20916 24244 20922 24308
rect 21909 24306 21975 24309
rect 21636 24304 21975 24306
rect 21636 24248 21914 24304
rect 21970 24248 21975 24304
rect 21636 24246 21975 24248
rect 21636 24173 21696 24246
rect 21909 24243 21975 24246
rect 749 24170 815 24173
rect 5901 24170 5967 24173
rect 749 24168 5967 24170
rect 749 24112 754 24168
rect 810 24112 5906 24168
rect 5962 24112 5967 24168
rect 749 24110 5967 24112
rect 749 24107 815 24110
rect 5901 24107 5967 24110
rect 9673 24170 9739 24173
rect 20529 24170 20595 24173
rect 20846 24170 20852 24172
rect 9673 24168 18522 24170
rect 9673 24112 9678 24168
rect 9734 24112 18522 24168
rect 9673 24110 18522 24112
rect 9673 24107 9739 24110
rect 841 24034 907 24037
rect 798 24032 907 24034
rect 798 23976 846 24032
rect 902 23976 907 24032
rect 798 23971 907 23976
rect 5717 24034 5783 24037
rect 5993 24034 6059 24037
rect 5717 24032 6059 24034
rect 5717 23976 5722 24032
rect 5778 23976 5998 24032
rect 6054 23976 6059 24032
rect 5717 23974 6059 23976
rect 5717 23971 5783 23974
rect 5993 23971 6059 23974
rect 6310 23972 6316 24036
rect 6380 24034 6386 24036
rect 6545 24034 6611 24037
rect 6380 24032 6611 24034
rect 6380 23976 6550 24032
rect 6606 23976 6611 24032
rect 6380 23974 6611 23976
rect 6380 23972 6386 23974
rect 6545 23971 6611 23974
rect 10910 23972 10916 24036
rect 10980 24034 10986 24036
rect 13302 24034 13308 24036
rect 10980 23974 13308 24034
rect 10980 23972 10986 23974
rect 13302 23972 13308 23974
rect 13372 23972 13378 24036
rect 13997 24034 14063 24037
rect 15101 24034 15167 24037
rect 13997 24032 15167 24034
rect 13997 23976 14002 24032
rect 14058 23976 15106 24032
rect 15162 23976 15167 24032
rect 13997 23974 15167 23976
rect 13997 23971 14063 23974
rect 15101 23971 15167 23974
rect 16798 23972 16804 24036
rect 16868 24034 16874 24036
rect 17493 24034 17559 24037
rect 16868 24032 17559 24034
rect 16868 23976 17498 24032
rect 17554 23976 17559 24032
rect 16868 23974 17559 23976
rect 18462 24034 18522 24110
rect 20529 24168 20852 24170
rect 20529 24112 20534 24168
rect 20590 24112 20852 24168
rect 20529 24110 20852 24112
rect 20529 24107 20595 24110
rect 20846 24108 20852 24110
rect 20916 24108 20922 24172
rect 21265 24170 21331 24173
rect 21222 24168 21331 24170
rect 21222 24112 21270 24168
rect 21326 24112 21331 24168
rect 21222 24107 21331 24112
rect 21633 24168 21699 24173
rect 21633 24112 21638 24168
rect 21694 24112 21699 24168
rect 21633 24107 21699 24112
rect 21909 24170 21975 24173
rect 27981 24170 28047 24173
rect 21909 24168 28047 24170
rect 21909 24112 21914 24168
rect 21970 24112 27986 24168
rect 28042 24112 28047 24168
rect 21909 24110 28047 24112
rect 21909 24107 21975 24110
rect 27981 24107 28047 24110
rect 21222 24034 21282 24107
rect 23657 24034 23723 24037
rect 18462 24032 23723 24034
rect 18462 23976 23662 24032
rect 23718 23976 23723 24032
rect 18462 23974 23723 23976
rect 16868 23972 16874 23974
rect 17493 23971 17559 23974
rect 23657 23971 23723 23974
rect 28390 23972 28396 24036
rect 28460 24034 28466 24036
rect 28533 24034 28599 24037
rect 28460 24032 28599 24034
rect 28460 23976 28538 24032
rect 28594 23976 28599 24032
rect 28460 23974 28599 23976
rect 28460 23972 28466 23974
rect 28533 23971 28599 23974
rect 798 23928 858 23971
rect 0 23838 858 23928
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 10409 23898 10475 23901
rect 11145 23898 11211 23901
rect 23381 23898 23447 23901
rect 10409 23896 23447 23898
rect 10409 23840 10414 23896
rect 10470 23840 11150 23896
rect 11206 23840 23386 23896
rect 23442 23840 23447 23896
rect 10409 23838 23447 23840
rect 0 23808 800 23838
rect 10409 23835 10475 23838
rect 11145 23835 11211 23838
rect 23381 23835 23447 23838
rect 31661 23898 31727 23901
rect 33200 23898 34000 23928
rect 31661 23896 34000 23898
rect 31661 23840 31666 23896
rect 31722 23840 34000 23896
rect 31661 23838 34000 23840
rect 31661 23835 31727 23838
rect 33200 23808 34000 23838
rect 3877 23762 3943 23765
rect 6361 23762 6427 23765
rect 3877 23760 6427 23762
rect 3877 23704 3882 23760
rect 3938 23704 6366 23760
rect 6422 23704 6427 23760
rect 3877 23702 6427 23704
rect 3877 23699 3943 23702
rect 6361 23699 6427 23702
rect 12065 23762 12131 23765
rect 15653 23762 15719 23765
rect 17033 23762 17099 23765
rect 12065 23760 17099 23762
rect 12065 23704 12070 23760
rect 12126 23704 15658 23760
rect 15714 23704 17038 23760
rect 17094 23704 17099 23760
rect 12065 23702 17099 23704
rect 12065 23699 12131 23702
rect 15653 23699 15719 23702
rect 17033 23699 17099 23702
rect 20805 23762 20871 23765
rect 24669 23762 24735 23765
rect 20805 23760 24735 23762
rect 20805 23704 20810 23760
rect 20866 23704 24674 23760
rect 24730 23704 24735 23760
rect 20805 23702 24735 23704
rect 20805 23699 20871 23702
rect 24669 23699 24735 23702
rect 3141 23626 3207 23629
rect 3509 23626 3575 23629
rect 6361 23626 6427 23629
rect 3141 23624 6427 23626
rect 3141 23568 3146 23624
rect 3202 23568 3514 23624
rect 3570 23568 6366 23624
rect 6422 23568 6427 23624
rect 3141 23566 6427 23568
rect 3141 23563 3207 23566
rect 3509 23563 3575 23566
rect 6361 23563 6427 23566
rect 11462 23564 11468 23628
rect 11532 23626 11538 23628
rect 11789 23626 11855 23629
rect 11532 23624 11855 23626
rect 11532 23568 11794 23624
rect 11850 23568 11855 23624
rect 11532 23566 11855 23568
rect 11532 23564 11538 23566
rect 11789 23563 11855 23566
rect 12525 23626 12591 23629
rect 15285 23626 15351 23629
rect 23749 23626 23815 23629
rect 24025 23626 24091 23629
rect 12525 23624 15351 23626
rect 12525 23568 12530 23624
rect 12586 23568 15290 23624
rect 15346 23568 15351 23624
rect 12525 23566 15351 23568
rect 12525 23563 12591 23566
rect 15285 23563 15351 23566
rect 16990 23624 24091 23626
rect 16990 23568 23754 23624
rect 23810 23568 24030 23624
rect 24086 23568 24091 23624
rect 16990 23566 24091 23568
rect 4654 23428 4660 23492
rect 4724 23490 4730 23492
rect 5533 23490 5599 23493
rect 4724 23488 5599 23490
rect 4724 23432 5538 23488
rect 5594 23432 5599 23488
rect 4724 23430 5599 23432
rect 4724 23428 4730 23430
rect 5533 23427 5599 23430
rect 5901 23490 5967 23493
rect 6494 23490 6500 23492
rect 5901 23488 6500 23490
rect 5901 23432 5906 23488
rect 5962 23432 6500 23488
rect 5901 23430 6500 23432
rect 5901 23427 5967 23430
rect 6494 23428 6500 23430
rect 6564 23428 6570 23492
rect 10961 23490 11027 23493
rect 12801 23490 12867 23493
rect 10961 23488 12867 23490
rect 10961 23432 10966 23488
rect 11022 23432 12806 23488
rect 12862 23432 12867 23488
rect 10961 23430 12867 23432
rect 10961 23427 11027 23430
rect 12801 23427 12867 23430
rect 13077 23490 13143 23493
rect 14549 23492 14615 23493
rect 13077 23488 14474 23490
rect 13077 23432 13082 23488
rect 13138 23432 14474 23488
rect 13077 23430 14474 23432
rect 13077 23427 13143 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 6085 23354 6151 23357
rect 7373 23354 7439 23357
rect 6085 23352 7439 23354
rect 6085 23296 6090 23352
rect 6146 23296 7378 23352
rect 7434 23296 7439 23352
rect 6085 23294 7439 23296
rect 6085 23291 6151 23294
rect 7373 23291 7439 23294
rect 7649 23354 7715 23357
rect 11094 23354 11100 23356
rect 7649 23352 11100 23354
rect 7649 23296 7654 23352
rect 7710 23296 11100 23352
rect 7649 23294 11100 23296
rect 7649 23291 7715 23294
rect 11094 23292 11100 23294
rect 11164 23292 11170 23356
rect 12382 23292 12388 23356
rect 12452 23354 12458 23356
rect 13445 23354 13511 23357
rect 12452 23352 13511 23354
rect 12452 23296 13450 23352
rect 13506 23296 13511 23352
rect 12452 23294 13511 23296
rect 14414 23354 14474 23430
rect 14549 23488 14596 23492
rect 14660 23490 14666 23492
rect 16990 23490 17050 23566
rect 23749 23563 23815 23566
rect 24025 23563 24091 23566
rect 17953 23492 18019 23493
rect 17902 23490 17908 23492
rect 14549 23432 14554 23488
rect 14549 23428 14596 23432
rect 14660 23430 14706 23490
rect 14782 23430 17050 23490
rect 17862 23430 17908 23490
rect 17972 23488 18019 23492
rect 18014 23432 18019 23488
rect 14660 23428 14666 23430
rect 14549 23427 14615 23428
rect 14782 23354 14842 23430
rect 17902 23428 17908 23430
rect 17972 23428 18019 23432
rect 17953 23427 18019 23428
rect 18689 23490 18755 23493
rect 20897 23490 20963 23493
rect 18689 23488 20963 23490
rect 18689 23432 18694 23488
rect 18750 23432 20902 23488
rect 20958 23432 20963 23488
rect 18689 23430 20963 23432
rect 18689 23427 18755 23430
rect 20897 23427 20963 23430
rect 21817 23490 21883 23493
rect 21950 23490 21956 23492
rect 21817 23488 21956 23490
rect 21817 23432 21822 23488
rect 21878 23432 21956 23488
rect 21817 23430 21956 23432
rect 21817 23427 21883 23430
rect 21950 23428 21956 23430
rect 22020 23428 22026 23492
rect 22134 23428 22140 23492
rect 22204 23490 22210 23492
rect 23565 23490 23631 23493
rect 22204 23488 23631 23490
rect 22204 23432 23570 23488
rect 23626 23432 23631 23488
rect 22204 23430 23631 23432
rect 22204 23428 22210 23430
rect 23565 23427 23631 23430
rect 23841 23490 23907 23493
rect 28165 23492 28231 23493
rect 23974 23490 23980 23492
rect 23841 23488 23980 23490
rect 23841 23432 23846 23488
rect 23902 23432 23980 23488
rect 23841 23430 23980 23432
rect 23841 23427 23907 23430
rect 23974 23428 23980 23430
rect 24044 23428 24050 23492
rect 28165 23488 28212 23492
rect 28276 23490 28282 23492
rect 28165 23432 28170 23488
rect 28165 23428 28212 23432
rect 28276 23430 28322 23490
rect 28276 23428 28282 23430
rect 28165 23427 28231 23428
rect 14414 23294 14842 23354
rect 16573 23354 16639 23357
rect 17217 23354 17283 23357
rect 26417 23354 26483 23357
rect 16573 23352 26483 23354
rect 16573 23296 16578 23352
rect 16634 23296 17222 23352
rect 17278 23296 26422 23352
rect 26478 23296 26483 23352
rect 16573 23294 26483 23296
rect 12452 23292 12458 23294
rect 13445 23291 13511 23294
rect 16573 23291 16639 23294
rect 17217 23291 17283 23294
rect 26417 23291 26483 23294
rect 473 23218 539 23221
rect 4981 23218 5047 23221
rect 7281 23218 7347 23221
rect 7414 23218 7420 23220
rect 473 23216 2790 23218
rect 473 23160 478 23216
rect 534 23160 2790 23216
rect 473 23158 2790 23160
rect 473 23155 539 23158
rect 2730 22674 2790 23158
rect 4981 23216 5826 23218
rect 4981 23160 4986 23216
rect 5042 23160 5826 23216
rect 4981 23158 5826 23160
rect 4981 23155 5047 23158
rect 4654 23020 4660 23084
rect 4724 23082 4730 23084
rect 4889 23082 4955 23085
rect 5766 23084 5826 23158
rect 7281 23216 7420 23218
rect 7281 23160 7286 23216
rect 7342 23160 7420 23216
rect 7281 23158 7420 23160
rect 7281 23155 7347 23158
rect 7414 23156 7420 23158
rect 7484 23156 7490 23220
rect 7833 23218 7899 23221
rect 10409 23218 10475 23221
rect 11278 23218 11284 23220
rect 7833 23216 8034 23218
rect 7833 23160 7838 23216
rect 7894 23160 8034 23216
rect 7833 23158 8034 23160
rect 7833 23155 7899 23158
rect 5390 23082 5396 23084
rect 4724 23080 5396 23082
rect 4724 23024 4894 23080
rect 4950 23024 5396 23080
rect 4724 23022 5396 23024
rect 4724 23020 4730 23022
rect 4889 23019 4955 23022
rect 5390 23020 5396 23022
rect 5460 23020 5466 23084
rect 5758 23020 5764 23084
rect 5828 23082 5834 23084
rect 5901 23082 5967 23085
rect 5828 23080 5967 23082
rect 5828 23024 5906 23080
rect 5962 23024 5967 23080
rect 5828 23022 5967 23024
rect 5828 23020 5834 23022
rect 5901 23019 5967 23022
rect 6913 23082 6979 23085
rect 7557 23082 7623 23085
rect 6913 23080 7623 23082
rect 6913 23024 6918 23080
rect 6974 23024 7562 23080
rect 7618 23024 7623 23080
rect 6913 23022 7623 23024
rect 6913 23019 6979 23022
rect 7557 23019 7623 23022
rect 5349 22946 5415 22949
rect 7189 22946 7255 22949
rect 5349 22944 7255 22946
rect 5349 22888 5354 22944
rect 5410 22888 7194 22944
rect 7250 22888 7255 22944
rect 5349 22886 7255 22888
rect 7974 22946 8034 23158
rect 10409 23216 11284 23218
rect 10409 23160 10414 23216
rect 10470 23160 11284 23216
rect 10409 23158 11284 23160
rect 10409 23155 10475 23158
rect 11278 23156 11284 23158
rect 11348 23218 11354 23220
rect 11881 23218 11947 23221
rect 11348 23216 11947 23218
rect 11348 23160 11886 23216
rect 11942 23160 11947 23216
rect 11348 23158 11947 23160
rect 11348 23156 11354 23158
rect 11881 23155 11947 23158
rect 12341 23218 12407 23221
rect 18413 23218 18479 23221
rect 12341 23216 18479 23218
rect 12341 23160 12346 23216
rect 12402 23160 18418 23216
rect 18474 23160 18479 23216
rect 12341 23158 18479 23160
rect 12341 23155 12407 23158
rect 18413 23155 18479 23158
rect 18965 23218 19031 23221
rect 22277 23218 22343 23221
rect 18965 23216 22343 23218
rect 18965 23160 18970 23216
rect 19026 23160 22282 23216
rect 22338 23160 22343 23216
rect 18965 23158 22343 23160
rect 18965 23155 19031 23158
rect 22277 23155 22343 23158
rect 22737 23218 22803 23221
rect 22870 23218 22876 23220
rect 22737 23216 22876 23218
rect 22737 23160 22742 23216
rect 22798 23160 22876 23216
rect 22737 23158 22876 23160
rect 22737 23155 22803 23158
rect 22870 23156 22876 23158
rect 22940 23156 22946 23220
rect 32489 23218 32555 23221
rect 33200 23218 34000 23248
rect 32489 23216 34000 23218
rect 32489 23160 32494 23216
rect 32550 23160 34000 23216
rect 32489 23158 34000 23160
rect 32489 23155 32555 23158
rect 33200 23128 34000 23158
rect 9029 23082 9095 23085
rect 11513 23082 11579 23085
rect 17585 23082 17651 23085
rect 9029 23080 11579 23082
rect 9029 23024 9034 23080
rect 9090 23024 11518 23080
rect 11574 23024 11579 23080
rect 9029 23022 11579 23024
rect 9029 23019 9095 23022
rect 11513 23019 11579 23022
rect 11654 23080 17651 23082
rect 11654 23024 17590 23080
rect 17646 23024 17651 23080
rect 11654 23022 17651 23024
rect 8109 22946 8175 22949
rect 7974 22944 8175 22946
rect 7974 22888 8114 22944
rect 8170 22888 8175 22944
rect 7974 22886 8175 22888
rect 5349 22883 5415 22886
rect 7189 22883 7255 22886
rect 8109 22883 8175 22886
rect 8518 22884 8524 22948
rect 8588 22946 8594 22948
rect 11654 22946 11714 23022
rect 17585 23019 17651 23022
rect 19425 23082 19491 23085
rect 19558 23082 19564 23084
rect 19425 23080 19564 23082
rect 19425 23024 19430 23080
rect 19486 23024 19564 23080
rect 19425 23022 19564 23024
rect 19425 23019 19491 23022
rect 19558 23020 19564 23022
rect 19628 23082 19634 23084
rect 24945 23082 25011 23085
rect 19628 23080 25011 23082
rect 19628 23024 24950 23080
rect 25006 23024 25011 23080
rect 19628 23022 25011 23024
rect 19628 23020 19634 23022
rect 24945 23019 25011 23022
rect 8588 22886 11714 22946
rect 11973 22946 12039 22949
rect 16757 22946 16823 22949
rect 11973 22944 16823 22946
rect 11973 22888 11978 22944
rect 12034 22888 16762 22944
rect 16818 22888 16823 22944
rect 11973 22886 16823 22888
rect 8588 22884 8594 22886
rect 11973 22883 12039 22886
rect 16757 22883 16823 22886
rect 19333 22948 19399 22949
rect 20161 22948 20227 22949
rect 19333 22944 19380 22948
rect 19444 22946 19450 22948
rect 20110 22946 20116 22948
rect 19333 22888 19338 22944
rect 19333 22884 19380 22888
rect 19444 22886 19490 22946
rect 20070 22886 20116 22946
rect 20180 22946 20227 22948
rect 20713 22946 20779 22949
rect 20180 22944 20779 22946
rect 20222 22888 20718 22944
rect 20774 22888 20779 22944
rect 19444 22884 19450 22886
rect 20110 22884 20116 22886
rect 20180 22886 20779 22888
rect 20180 22884 20227 22886
rect 19333 22883 19399 22884
rect 20161 22883 20227 22884
rect 20713 22883 20779 22886
rect 22737 22946 22803 22949
rect 25262 22946 25268 22948
rect 22737 22944 25268 22946
rect 22737 22888 22742 22944
rect 22798 22888 25268 22944
rect 22737 22886 25268 22888
rect 22737 22883 22803 22886
rect 25262 22884 25268 22886
rect 25332 22884 25338 22948
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 5349 22810 5415 22813
rect 6085 22810 6151 22813
rect 5349 22808 6151 22810
rect 5349 22752 5354 22808
rect 5410 22752 6090 22808
rect 6146 22752 6151 22808
rect 5349 22750 6151 22752
rect 5349 22747 5415 22750
rect 6085 22747 6151 22750
rect 6545 22810 6611 22813
rect 6913 22810 6979 22813
rect 6545 22808 6979 22810
rect 6545 22752 6550 22808
rect 6606 22752 6918 22808
rect 6974 22752 6979 22808
rect 6545 22750 6979 22752
rect 6545 22747 6611 22750
rect 6913 22747 6979 22750
rect 10501 22810 10567 22813
rect 13077 22810 13143 22813
rect 10501 22808 13143 22810
rect 10501 22752 10506 22808
rect 10562 22752 13082 22808
rect 13138 22752 13143 22808
rect 10501 22750 13143 22752
rect 10501 22747 10567 22750
rect 13077 22747 13143 22750
rect 16941 22810 17007 22813
rect 17861 22810 17927 22813
rect 20294 22810 20300 22812
rect 16941 22808 20300 22810
rect 16941 22752 16946 22808
rect 17002 22752 17866 22808
rect 17922 22752 20300 22808
rect 16941 22750 20300 22752
rect 16941 22747 17007 22750
rect 17861 22747 17927 22750
rect 20294 22748 20300 22750
rect 20364 22748 20370 22812
rect 20662 22748 20668 22812
rect 20732 22810 20738 22812
rect 28993 22810 29059 22813
rect 20732 22808 29059 22810
rect 20732 22752 28998 22808
rect 29054 22752 29059 22808
rect 20732 22750 29059 22752
rect 20732 22748 20738 22750
rect 28993 22747 29059 22750
rect 17493 22674 17559 22677
rect 2730 22672 17559 22674
rect 2730 22616 17498 22672
rect 17554 22616 17559 22672
rect 2730 22614 17559 22616
rect 17493 22611 17559 22614
rect 18229 22674 18295 22677
rect 18454 22674 18460 22676
rect 18229 22672 18460 22674
rect 18229 22616 18234 22672
rect 18290 22616 18460 22672
rect 18229 22614 18460 22616
rect 18229 22611 18295 22614
rect 18454 22612 18460 22614
rect 18524 22612 18530 22676
rect 18873 22674 18939 22677
rect 26233 22674 26299 22677
rect 18873 22672 26299 22674
rect 18873 22616 18878 22672
rect 18934 22616 26238 22672
rect 26294 22616 26299 22672
rect 18873 22614 26299 22616
rect 18873 22611 18939 22614
rect 26233 22611 26299 22614
rect 3141 22538 3207 22541
rect 5073 22538 5139 22541
rect 5717 22538 5783 22541
rect 8293 22538 8359 22541
rect 3141 22536 4722 22538
rect 3141 22480 3146 22536
rect 3202 22480 4722 22536
rect 3141 22478 4722 22480
rect 3141 22475 3207 22478
rect 4662 22402 4722 22478
rect 5073 22536 8359 22538
rect 5073 22480 5078 22536
rect 5134 22480 5722 22536
rect 5778 22480 8298 22536
rect 8354 22480 8359 22536
rect 5073 22478 8359 22480
rect 5073 22475 5139 22478
rect 5717 22475 5783 22478
rect 8293 22475 8359 22478
rect 9121 22538 9187 22541
rect 22645 22538 22711 22541
rect 9121 22536 22711 22538
rect 9121 22480 9126 22536
rect 9182 22480 22650 22536
rect 22706 22480 22711 22536
rect 9121 22478 22711 22480
rect 9121 22475 9187 22478
rect 22645 22475 22711 22478
rect 32397 22538 32463 22541
rect 33200 22538 34000 22568
rect 32397 22536 34000 22538
rect 32397 22480 32402 22536
rect 32458 22480 34000 22536
rect 32397 22478 34000 22480
rect 32397 22475 32463 22478
rect 33200 22448 34000 22478
rect 4981 22402 5047 22405
rect 7649 22402 7715 22405
rect 4662 22400 7715 22402
rect 4662 22344 4986 22400
rect 5042 22344 7654 22400
rect 7710 22344 7715 22400
rect 4662 22342 7715 22344
rect 4981 22339 5047 22342
rect 7649 22339 7715 22342
rect 9949 22402 10015 22405
rect 12525 22402 12591 22405
rect 9949 22400 12591 22402
rect 9949 22344 9954 22400
rect 10010 22344 12530 22400
rect 12586 22344 12591 22400
rect 9949 22342 12591 22344
rect 9949 22339 10015 22342
rect 12525 22339 12591 22342
rect 12801 22402 12867 22405
rect 18873 22402 18939 22405
rect 12801 22400 18939 22402
rect 12801 22344 12806 22400
rect 12862 22344 18878 22400
rect 18934 22344 18939 22400
rect 12801 22342 18939 22344
rect 12801 22339 12867 22342
rect 18873 22339 18939 22342
rect 19333 22402 19399 22405
rect 20713 22402 20779 22405
rect 19333 22400 20779 22402
rect 19333 22344 19338 22400
rect 19394 22344 20718 22400
rect 20774 22344 20779 22400
rect 19333 22342 20779 22344
rect 19333 22339 19399 22342
rect 20713 22339 20779 22342
rect 25078 22340 25084 22404
rect 25148 22402 25154 22404
rect 25221 22402 25287 22405
rect 25148 22400 25287 22402
rect 25148 22344 25226 22400
rect 25282 22344 25287 22400
rect 25148 22342 25287 22344
rect 25148 22340 25154 22342
rect 25221 22339 25287 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 4705 22266 4771 22269
rect 5901 22266 5967 22269
rect 6545 22268 6611 22269
rect 4705 22264 5967 22266
rect 4705 22208 4710 22264
rect 4766 22208 5906 22264
rect 5962 22208 5967 22264
rect 4705 22206 5967 22208
rect 4705 22203 4771 22206
rect 5901 22203 5967 22206
rect 6494 22204 6500 22268
rect 6564 22266 6611 22268
rect 11697 22266 11763 22269
rect 12014 22266 12020 22268
rect 6564 22264 6656 22266
rect 6606 22208 6656 22264
rect 6564 22206 6656 22208
rect 11697 22264 12020 22266
rect 11697 22208 11702 22264
rect 11758 22208 12020 22264
rect 11697 22206 12020 22208
rect 6564 22204 6611 22206
rect 6545 22203 6611 22204
rect 11697 22203 11763 22206
rect 12014 22204 12020 22206
rect 12084 22204 12090 22268
rect 12198 22204 12204 22268
rect 12268 22266 12274 22268
rect 19425 22266 19491 22269
rect 12268 22264 19491 22266
rect 12268 22208 19430 22264
rect 19486 22208 19491 22264
rect 12268 22206 19491 22208
rect 12268 22204 12274 22206
rect 19425 22203 19491 22206
rect 20294 22204 20300 22268
rect 20364 22266 20370 22268
rect 22737 22266 22803 22269
rect 20364 22264 22803 22266
rect 20364 22208 22742 22264
rect 22798 22208 22803 22264
rect 20364 22206 22803 22208
rect 20364 22204 20370 22206
rect 22737 22203 22803 22206
rect 24577 22266 24643 22269
rect 24710 22266 24716 22268
rect 24577 22264 24716 22266
rect 24577 22208 24582 22264
rect 24638 22208 24716 22264
rect 24577 22206 24716 22208
rect 24577 22203 24643 22206
rect 24710 22204 24716 22206
rect 24780 22204 24786 22268
rect 4521 22130 4587 22133
rect 5574 22130 5580 22132
rect 4521 22128 5580 22130
rect 4521 22072 4526 22128
rect 4582 22072 5580 22128
rect 4521 22070 5580 22072
rect 4521 22067 4587 22070
rect 5574 22068 5580 22070
rect 5644 22068 5650 22132
rect 5901 22130 5967 22133
rect 6126 22130 6132 22132
rect 5901 22128 6132 22130
rect 5901 22072 5906 22128
rect 5962 22072 6132 22128
rect 5901 22070 6132 22072
rect 5901 22067 5967 22070
rect 6126 22068 6132 22070
rect 6196 22068 6202 22132
rect 6862 22068 6868 22132
rect 6932 22130 6938 22132
rect 12617 22130 12683 22133
rect 6932 22128 12683 22130
rect 6932 22072 12622 22128
rect 12678 22072 12683 22128
rect 6932 22070 12683 22072
rect 6932 22068 6938 22070
rect 12617 22067 12683 22070
rect 13169 22130 13235 22133
rect 16849 22130 16915 22133
rect 13169 22128 16915 22130
rect 13169 22072 13174 22128
rect 13230 22072 16854 22128
rect 16910 22072 16915 22128
rect 13169 22070 16915 22072
rect 13169 22067 13235 22070
rect 16849 22067 16915 22070
rect 19149 22130 19215 22133
rect 19333 22130 19399 22133
rect 19149 22128 19399 22130
rect 19149 22072 19154 22128
rect 19210 22072 19338 22128
rect 19394 22072 19399 22128
rect 19149 22070 19399 22072
rect 19149 22067 19215 22070
rect 19333 22067 19399 22070
rect 19609 22130 19675 22133
rect 19742 22130 19748 22132
rect 19609 22128 19748 22130
rect 19609 22072 19614 22128
rect 19670 22072 19748 22128
rect 19609 22070 19748 22072
rect 19609 22067 19675 22070
rect 19742 22068 19748 22070
rect 19812 22068 19818 22132
rect 20161 22130 20227 22133
rect 21398 22130 21404 22132
rect 20161 22128 21404 22130
rect 20161 22072 20166 22128
rect 20222 22072 21404 22128
rect 20161 22070 21404 22072
rect 20161 22067 20227 22070
rect 21398 22068 21404 22070
rect 21468 22130 21474 22132
rect 30373 22130 30439 22133
rect 21468 22128 30439 22130
rect 21468 22072 30378 22128
rect 30434 22072 30439 22128
rect 21468 22070 30439 22072
rect 21468 22068 21474 22070
rect 30373 22067 30439 22070
rect 4337 21994 4403 21997
rect 5533 21996 5599 21997
rect 4337 21992 5458 21994
rect 4337 21936 4342 21992
rect 4398 21936 5458 21992
rect 4337 21934 5458 21936
rect 4337 21931 4403 21934
rect 3550 21796 3556 21860
rect 3620 21858 3626 21860
rect 4061 21858 4127 21861
rect 4521 21858 4587 21861
rect 3620 21856 4587 21858
rect 3620 21800 4066 21856
rect 4122 21800 4526 21856
rect 4582 21800 4587 21856
rect 3620 21798 4587 21800
rect 3620 21796 3626 21798
rect 4061 21795 4127 21798
rect 4521 21795 4587 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 2262 21660 2268 21724
rect 2332 21722 2338 21724
rect 3509 21722 3575 21725
rect 2332 21720 3575 21722
rect 2332 21664 3514 21720
rect 3570 21664 3575 21720
rect 2332 21662 3575 21664
rect 5398 21722 5458 21934
rect 5533 21992 5580 21996
rect 5644 21994 5650 21996
rect 8661 21994 8727 21997
rect 11605 21994 11671 21997
rect 12382 21994 12388 21996
rect 5533 21936 5538 21992
rect 5533 21932 5580 21936
rect 5644 21934 5690 21994
rect 8661 21992 8770 21994
rect 8661 21936 8666 21992
rect 8722 21936 8770 21992
rect 5644 21932 5650 21934
rect 5533 21931 5599 21932
rect 8661 21931 8770 21936
rect 11605 21992 12388 21994
rect 11605 21936 11610 21992
rect 11666 21936 12388 21992
rect 11605 21934 12388 21936
rect 11605 21931 11671 21934
rect 12382 21932 12388 21934
rect 12452 21932 12458 21996
rect 13077 21994 13143 21997
rect 13486 21994 13492 21996
rect 13077 21992 13492 21994
rect 13077 21936 13082 21992
rect 13138 21936 13492 21992
rect 13077 21934 13492 21936
rect 13077 21931 13143 21934
rect 13486 21932 13492 21934
rect 13556 21932 13562 21996
rect 13813 21994 13879 21997
rect 25497 21994 25563 21997
rect 13813 21992 25563 21994
rect 13813 21936 13818 21992
rect 13874 21936 25502 21992
rect 25558 21936 25563 21992
rect 13813 21934 25563 21936
rect 13813 21931 13879 21934
rect 25497 21931 25563 21934
rect 25681 21994 25747 21997
rect 25814 21994 25820 21996
rect 25681 21992 25820 21994
rect 25681 21936 25686 21992
rect 25742 21936 25820 21992
rect 25681 21934 25820 21936
rect 25681 21931 25747 21934
rect 25814 21932 25820 21934
rect 25884 21932 25890 21996
rect 8710 21858 8770 21931
rect 8937 21858 9003 21861
rect 8710 21856 9003 21858
rect 8710 21800 8942 21856
rect 8998 21800 9003 21856
rect 8710 21798 9003 21800
rect 8937 21795 9003 21798
rect 9489 21858 9555 21861
rect 11881 21858 11947 21861
rect 14222 21858 14228 21860
rect 9489 21856 14228 21858
rect 9489 21800 9494 21856
rect 9550 21800 11886 21856
rect 11942 21800 14228 21856
rect 9489 21798 14228 21800
rect 9489 21795 9555 21798
rect 11881 21795 11947 21798
rect 14222 21796 14228 21798
rect 14292 21796 14298 21860
rect 19241 21858 19307 21861
rect 22686 21858 22692 21860
rect 19241 21856 22692 21858
rect 19241 21800 19246 21856
rect 19302 21800 22692 21856
rect 19241 21798 22692 21800
rect 19241 21795 19307 21798
rect 22686 21796 22692 21798
rect 22756 21796 22762 21860
rect 6177 21722 6243 21725
rect 10409 21722 10475 21725
rect 12801 21722 12867 21725
rect 13302 21722 13308 21724
rect 5398 21720 10475 21722
rect 5398 21664 6182 21720
rect 6238 21664 10414 21720
rect 10470 21664 10475 21720
rect 5398 21662 10475 21664
rect 2332 21660 2338 21662
rect 3509 21659 3575 21662
rect 6177 21659 6243 21662
rect 10409 21659 10475 21662
rect 12022 21720 13308 21722
rect 12022 21664 12806 21720
rect 12862 21664 13308 21720
rect 12022 21662 13308 21664
rect 1393 21586 1459 21589
rect 10409 21586 10475 21589
rect 1393 21584 10475 21586
rect 1393 21528 1398 21584
rect 1454 21528 10414 21584
rect 10470 21528 10475 21584
rect 1393 21526 10475 21528
rect 1393 21523 1459 21526
rect 10409 21523 10475 21526
rect 10726 21524 10732 21588
rect 10796 21586 10802 21588
rect 10961 21586 11027 21589
rect 10796 21584 11027 21586
rect 10796 21528 10966 21584
rect 11022 21528 11027 21584
rect 10796 21526 11027 21528
rect 10796 21524 10802 21526
rect 10961 21523 11027 21526
rect 11789 21586 11855 21589
rect 12022 21586 12082 21662
rect 12801 21659 12867 21662
rect 13302 21660 13308 21662
rect 13372 21660 13378 21724
rect 13486 21660 13492 21724
rect 13556 21722 13562 21724
rect 13629 21722 13695 21725
rect 13556 21720 13695 21722
rect 13556 21664 13634 21720
rect 13690 21664 13695 21720
rect 13556 21662 13695 21664
rect 13556 21660 13562 21662
rect 13629 21659 13695 21662
rect 13813 21722 13879 21725
rect 14038 21722 14044 21724
rect 13813 21720 14044 21722
rect 13813 21664 13818 21720
rect 13874 21664 14044 21720
rect 13813 21662 14044 21664
rect 13813 21659 13879 21662
rect 14038 21660 14044 21662
rect 14108 21660 14114 21724
rect 14273 21722 14339 21725
rect 17401 21722 17467 21725
rect 14273 21720 17467 21722
rect 14273 21664 14278 21720
rect 14334 21664 17406 21720
rect 17462 21664 17467 21720
rect 14273 21662 17467 21664
rect 14273 21659 14339 21662
rect 17401 21659 17467 21662
rect 19333 21722 19399 21725
rect 20253 21722 20319 21725
rect 19333 21720 20319 21722
rect 19333 21664 19338 21720
rect 19394 21664 20258 21720
rect 20314 21664 20319 21720
rect 19333 21662 20319 21664
rect 19333 21659 19399 21662
rect 20253 21659 20319 21662
rect 22737 21722 22803 21725
rect 22870 21722 22876 21724
rect 22737 21720 22876 21722
rect 22737 21664 22742 21720
rect 22798 21664 22876 21720
rect 22737 21662 22876 21664
rect 22737 21659 22803 21662
rect 22870 21660 22876 21662
rect 22940 21660 22946 21724
rect 23422 21660 23428 21724
rect 23492 21722 23498 21724
rect 24342 21722 24348 21724
rect 23492 21662 24348 21722
rect 23492 21660 23498 21662
rect 24342 21660 24348 21662
rect 24412 21660 24418 21724
rect 11789 21584 12082 21586
rect 11789 21528 11794 21584
rect 11850 21528 12082 21584
rect 11789 21526 12082 21528
rect 12341 21586 12407 21589
rect 14733 21586 14799 21589
rect 18086 21586 18092 21588
rect 12341 21584 18092 21586
rect 12341 21528 12346 21584
rect 12402 21528 14738 21584
rect 14794 21528 18092 21584
rect 12341 21526 18092 21528
rect 11789 21523 11855 21526
rect 12341 21523 12407 21526
rect 14733 21523 14799 21526
rect 18086 21524 18092 21526
rect 18156 21524 18162 21588
rect 19885 21586 19951 21589
rect 20294 21586 20300 21588
rect 19885 21584 20300 21586
rect 19885 21528 19890 21584
rect 19946 21528 20300 21584
rect 19885 21526 20300 21528
rect 19885 21523 19951 21526
rect 20294 21524 20300 21526
rect 20364 21524 20370 21588
rect 20478 21524 20484 21588
rect 20548 21586 20554 21588
rect 20805 21586 20871 21589
rect 23422 21586 23428 21588
rect 20548 21584 23428 21586
rect 20548 21528 20810 21584
rect 20866 21528 23428 21584
rect 20548 21526 23428 21528
rect 20548 21524 20554 21526
rect 20805 21523 20871 21526
rect 23422 21524 23428 21526
rect 23492 21524 23498 21588
rect 3785 21450 3851 21453
rect 4245 21450 4311 21453
rect 5349 21452 5415 21453
rect 5349 21450 5396 21452
rect 3785 21448 4768 21450
rect 3785 21392 3790 21448
rect 3846 21392 4250 21448
rect 4306 21392 4768 21448
rect 3785 21390 4768 21392
rect 5304 21448 5396 21450
rect 5304 21392 5354 21448
rect 5304 21390 5396 21392
rect 3785 21387 3851 21390
rect 4245 21387 4311 21390
rect 4708 21314 4768 21390
rect 5349 21388 5396 21390
rect 5460 21388 5466 21452
rect 9305 21450 9371 21453
rect 9990 21450 9996 21452
rect 9305 21448 9996 21450
rect 9305 21392 9310 21448
rect 9366 21392 9996 21448
rect 9305 21390 9996 21392
rect 5349 21387 5415 21388
rect 9305 21387 9371 21390
rect 9990 21388 9996 21390
rect 10060 21388 10066 21452
rect 11792 21450 11852 21523
rect 12433 21452 12499 21453
rect 12382 21450 12388 21452
rect 10136 21390 11852 21450
rect 12342 21390 12388 21450
rect 12452 21448 12499 21452
rect 12494 21392 12499 21448
rect 5758 21314 5764 21316
rect 4708 21254 5764 21314
rect 5758 21252 5764 21254
rect 5828 21314 5834 21316
rect 6085 21314 6151 21317
rect 5828 21312 6151 21314
rect 5828 21256 6090 21312
rect 6146 21256 6151 21312
rect 5828 21254 6151 21256
rect 5828 21252 5834 21254
rect 6085 21251 6151 21254
rect 7414 21252 7420 21316
rect 7484 21314 7490 21316
rect 10136 21314 10196 21390
rect 12382 21388 12388 21390
rect 12452 21388 12499 21392
rect 12433 21387 12499 21388
rect 12617 21450 12683 21453
rect 12893 21452 12959 21453
rect 12750 21450 12756 21452
rect 12617 21448 12756 21450
rect 12617 21392 12622 21448
rect 12678 21392 12756 21448
rect 12617 21390 12756 21392
rect 12617 21387 12683 21390
rect 12750 21388 12756 21390
rect 12820 21388 12826 21452
rect 12893 21448 12940 21452
rect 13004 21450 13010 21452
rect 13537 21450 13603 21453
rect 17677 21450 17743 21453
rect 19701 21450 19767 21453
rect 19977 21452 20043 21453
rect 19926 21450 19932 21452
rect 12893 21392 12898 21448
rect 12893 21388 12940 21392
rect 13004 21390 13050 21450
rect 13310 21448 17234 21450
rect 13310 21392 13542 21448
rect 13598 21392 17234 21448
rect 13310 21390 17234 21392
rect 13004 21388 13010 21390
rect 12893 21387 12959 21388
rect 7484 21254 10196 21314
rect 10869 21314 10935 21317
rect 13310 21314 13370 21390
rect 13537 21387 13603 21390
rect 10869 21312 13370 21314
rect 10869 21256 10874 21312
rect 10930 21256 13370 21312
rect 10869 21254 13370 21256
rect 7484 21252 7490 21254
rect 10869 21251 10935 21254
rect 13486 21252 13492 21316
rect 13556 21314 13562 21316
rect 16941 21314 17007 21317
rect 13556 21312 17007 21314
rect 13556 21256 16946 21312
rect 17002 21256 17007 21312
rect 13556 21254 17007 21256
rect 17174 21314 17234 21390
rect 17677 21448 19767 21450
rect 17677 21392 17682 21448
rect 17738 21392 19706 21448
rect 19762 21392 19767 21448
rect 17677 21390 19767 21392
rect 19886 21390 19932 21450
rect 19996 21450 20043 21452
rect 20253 21450 20319 21453
rect 19996 21448 20319 21450
rect 20038 21392 20258 21448
rect 20314 21392 20319 21448
rect 17677 21387 17743 21390
rect 19701 21387 19767 21390
rect 19926 21388 19932 21390
rect 19996 21390 20319 21392
rect 19996 21388 20043 21390
rect 19977 21387 20043 21388
rect 20253 21387 20319 21390
rect 20846 21388 20852 21452
rect 20916 21450 20922 21452
rect 25129 21450 25195 21453
rect 20916 21448 25195 21450
rect 20916 21392 25134 21448
rect 25190 21392 25195 21448
rect 20916 21390 25195 21392
rect 20916 21388 20922 21390
rect 25129 21387 25195 21390
rect 17677 21314 17743 21317
rect 22134 21314 22140 21316
rect 17174 21312 22140 21314
rect 17174 21256 17682 21312
rect 17738 21256 22140 21312
rect 17174 21254 22140 21256
rect 13556 21252 13562 21254
rect 16941 21251 17007 21254
rect 17677 21251 17743 21254
rect 22134 21252 22140 21254
rect 22204 21252 22210 21316
rect 23841 21314 23907 21317
rect 31150 21314 31156 21316
rect 23841 21312 31156 21314
rect 23841 21256 23846 21312
rect 23902 21256 31156 21312
rect 23841 21254 31156 21256
rect 23841 21251 23907 21254
rect 31150 21252 31156 21254
rect 31220 21252 31226 21316
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 4889 21178 4955 21181
rect 5901 21178 5967 21181
rect 4889 21176 5967 21178
rect 4889 21120 4894 21176
rect 4950 21120 5906 21176
rect 5962 21120 5967 21176
rect 4889 21118 5967 21120
rect 4889 21115 4955 21118
rect 5901 21115 5967 21118
rect 8569 21178 8635 21181
rect 9213 21178 9279 21181
rect 8569 21176 9279 21178
rect 8569 21120 8574 21176
rect 8630 21120 9218 21176
rect 9274 21120 9279 21176
rect 8569 21118 9279 21120
rect 8569 21115 8635 21118
rect 9213 21115 9279 21118
rect 11789 21178 11855 21181
rect 13353 21178 13419 21181
rect 11789 21176 13419 21178
rect 11789 21120 11794 21176
rect 11850 21120 13358 21176
rect 13414 21120 13419 21176
rect 11789 21118 13419 21120
rect 11789 21115 11855 21118
rect 13353 21115 13419 21118
rect 14641 21178 14707 21181
rect 14774 21178 14780 21180
rect 14641 21176 14780 21178
rect 14641 21120 14646 21176
rect 14702 21120 14780 21176
rect 14641 21118 14780 21120
rect 14641 21115 14707 21118
rect 14774 21116 14780 21118
rect 14844 21116 14850 21180
rect 16757 21178 16823 21181
rect 23054 21178 23060 21180
rect 16757 21176 23060 21178
rect 16757 21120 16762 21176
rect 16818 21120 23060 21176
rect 16757 21118 23060 21120
rect 16757 21115 16823 21118
rect 23054 21116 23060 21118
rect 23124 21116 23130 21180
rect 32489 21178 32555 21181
rect 33200 21178 34000 21208
rect 32489 21176 34000 21178
rect 32489 21120 32494 21176
rect 32550 21120 34000 21176
rect 32489 21118 34000 21120
rect 32489 21115 32555 21118
rect 33200 21088 34000 21118
rect 3417 21042 3483 21045
rect 4245 21042 4311 21045
rect 7925 21042 7991 21045
rect 3417 21040 7991 21042
rect 3417 20984 3422 21040
rect 3478 20984 4250 21040
rect 4306 20984 7930 21040
rect 7986 20984 7991 21040
rect 3417 20982 7991 20984
rect 3417 20979 3483 20982
rect 4245 20979 4311 20982
rect 7925 20979 7991 20982
rect 9305 21042 9371 21045
rect 15009 21042 15075 21045
rect 9305 21040 15075 21042
rect 9305 20984 9310 21040
rect 9366 20984 15014 21040
rect 15070 20984 15075 21040
rect 9305 20982 15075 20984
rect 9305 20979 9371 20982
rect 15009 20979 15075 20982
rect 15193 21042 15259 21045
rect 17677 21042 17743 21045
rect 15193 21040 17743 21042
rect 15193 20984 15198 21040
rect 15254 20984 17682 21040
rect 17738 20984 17743 21040
rect 15193 20982 17743 20984
rect 15193 20979 15259 20982
rect 17677 20979 17743 20982
rect 17902 20980 17908 21044
rect 17972 21042 17978 21044
rect 19241 21042 19307 21045
rect 19517 21044 19583 21045
rect 19517 21042 19564 21044
rect 17972 21040 19307 21042
rect 17972 20984 19246 21040
rect 19302 20984 19307 21040
rect 17972 20982 19307 20984
rect 19472 21040 19564 21042
rect 19472 20984 19522 21040
rect 19472 20982 19564 20984
rect 17972 20980 17978 20982
rect 19241 20979 19307 20982
rect 19517 20980 19564 20982
rect 19628 20980 19634 21044
rect 19701 21042 19767 21045
rect 21633 21044 21699 21045
rect 21582 21042 21588 21044
rect 19701 21040 21588 21042
rect 21652 21042 21699 21044
rect 22001 21042 22067 21045
rect 27981 21042 28047 21045
rect 21652 21040 21744 21042
rect 19701 20984 19706 21040
rect 19762 20984 21588 21040
rect 21694 20984 21744 21040
rect 19701 20982 21588 20984
rect 19517 20979 19583 20980
rect 19701 20979 19767 20982
rect 21582 20980 21588 20982
rect 21652 20982 21744 20984
rect 22001 21040 28047 21042
rect 22001 20984 22006 21040
rect 22062 20984 27986 21040
rect 28042 20984 28047 21040
rect 22001 20982 28047 20984
rect 21652 20980 21699 20982
rect 21633 20979 21699 20980
rect 22001 20979 22067 20982
rect 27981 20979 28047 20982
rect 565 20906 631 20909
rect 5441 20906 5507 20909
rect 565 20904 5507 20906
rect 565 20848 570 20904
rect 626 20848 5446 20904
rect 5502 20848 5507 20904
rect 565 20846 5507 20848
rect 565 20843 631 20846
rect 5441 20843 5507 20846
rect 6269 20906 6335 20909
rect 11881 20906 11947 20909
rect 13353 20906 13419 20909
rect 6269 20904 11947 20906
rect 6269 20848 6274 20904
rect 6330 20848 11886 20904
rect 11942 20848 11947 20904
rect 6269 20846 11947 20848
rect 6269 20843 6335 20846
rect 11881 20843 11947 20846
rect 12022 20904 13419 20906
rect 12022 20848 13358 20904
rect 13414 20848 13419 20904
rect 12022 20846 13419 20848
rect 790 20708 796 20772
rect 860 20770 866 20772
rect 1025 20770 1091 20773
rect 860 20768 1091 20770
rect 860 20712 1030 20768
rect 1086 20712 1091 20768
rect 860 20710 1091 20712
rect 860 20708 866 20710
rect 1025 20707 1091 20710
rect 3785 20770 3851 20773
rect 3918 20770 3924 20772
rect 3785 20768 3924 20770
rect 3785 20712 3790 20768
rect 3846 20712 3924 20768
rect 3785 20710 3924 20712
rect 3785 20707 3851 20710
rect 3918 20708 3924 20710
rect 3988 20708 3994 20772
rect 7046 20708 7052 20772
rect 7116 20770 7122 20772
rect 7833 20770 7899 20773
rect 8937 20770 9003 20773
rect 7116 20768 7899 20770
rect 7116 20712 7838 20768
rect 7894 20712 7899 20768
rect 7116 20710 7899 20712
rect 7116 20708 7122 20710
rect 7833 20707 7899 20710
rect 8526 20768 9003 20770
rect 8526 20712 8942 20768
rect 8998 20712 9003 20768
rect 8526 20710 9003 20712
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 2221 20634 2287 20637
rect 4705 20634 4771 20637
rect 8526 20634 8586 20710
rect 8937 20707 9003 20710
rect 9857 20770 9923 20773
rect 11053 20770 11119 20773
rect 12022 20770 12082 20846
rect 13353 20843 13419 20846
rect 13537 20906 13603 20909
rect 13997 20908 14063 20909
rect 13670 20906 13676 20908
rect 13537 20904 13676 20906
rect 13537 20848 13542 20904
rect 13598 20848 13676 20904
rect 13537 20846 13676 20848
rect 13537 20843 13603 20846
rect 13670 20844 13676 20846
rect 13740 20844 13746 20908
rect 13997 20906 14044 20908
rect 13952 20904 14044 20906
rect 13952 20848 14002 20904
rect 13952 20846 14044 20848
rect 13997 20844 14044 20846
rect 14108 20844 14114 20908
rect 15510 20844 15516 20908
rect 15580 20906 15586 20908
rect 18229 20906 18295 20909
rect 15580 20904 18295 20906
rect 15580 20848 18234 20904
rect 18290 20848 18295 20904
rect 15580 20846 18295 20848
rect 15580 20844 15586 20846
rect 13997 20843 14063 20844
rect 18229 20843 18295 20846
rect 19333 20906 19399 20909
rect 19517 20906 19583 20909
rect 22737 20906 22803 20909
rect 27429 20906 27495 20909
rect 19333 20904 20868 20906
rect 19333 20848 19338 20904
rect 19394 20848 19522 20904
rect 19578 20848 20868 20904
rect 19333 20846 20868 20848
rect 19333 20843 19399 20846
rect 19517 20843 19583 20846
rect 12801 20770 12867 20773
rect 9857 20768 12082 20770
rect 9857 20712 9862 20768
rect 9918 20712 11058 20768
rect 11114 20712 12082 20768
rect 9857 20710 12082 20712
rect 12160 20768 12867 20770
rect 12160 20712 12806 20768
rect 12862 20712 12867 20768
rect 12160 20710 12867 20712
rect 9857 20707 9923 20710
rect 11053 20707 11119 20710
rect 2221 20632 4771 20634
rect 2221 20576 2226 20632
rect 2282 20576 4710 20632
rect 4766 20576 4771 20632
rect 2221 20574 4771 20576
rect 2221 20571 2287 20574
rect 4705 20571 4771 20574
rect 6686 20574 8586 20634
rect 3325 20498 3391 20501
rect 3785 20498 3851 20501
rect 5717 20498 5783 20501
rect 3325 20496 5783 20498
rect 3325 20440 3330 20496
rect 3386 20440 3790 20496
rect 3846 20440 5722 20496
rect 5778 20440 5783 20496
rect 3325 20438 5783 20440
rect 3325 20435 3391 20438
rect 3785 20435 3851 20438
rect 5717 20435 5783 20438
rect 6686 20365 6746 20574
rect 8702 20572 8708 20636
rect 8772 20634 8778 20636
rect 8937 20634 9003 20637
rect 8772 20632 9003 20634
rect 8772 20576 8942 20632
rect 8998 20576 9003 20632
rect 8772 20574 9003 20576
rect 8772 20572 8778 20574
rect 8937 20571 9003 20574
rect 9213 20634 9279 20637
rect 12160 20634 12220 20710
rect 12801 20707 12867 20710
rect 12934 20708 12940 20772
rect 13004 20770 13010 20772
rect 13169 20770 13235 20773
rect 13004 20768 13235 20770
rect 13004 20712 13174 20768
rect 13230 20712 13235 20768
rect 13004 20710 13235 20712
rect 13004 20708 13010 20710
rect 13169 20707 13235 20710
rect 13629 20770 13695 20773
rect 17861 20770 17927 20773
rect 13629 20768 17927 20770
rect 13629 20712 13634 20768
rect 13690 20712 17866 20768
rect 17922 20712 17927 20768
rect 13629 20710 17927 20712
rect 13629 20707 13695 20710
rect 17861 20707 17927 20710
rect 18086 20708 18092 20772
rect 18156 20770 18162 20772
rect 19701 20770 19767 20773
rect 18156 20768 19767 20770
rect 18156 20712 19706 20768
rect 19762 20712 19767 20768
rect 18156 20710 19767 20712
rect 18156 20708 18162 20710
rect 19701 20707 19767 20710
rect 20345 20770 20411 20773
rect 20662 20770 20668 20772
rect 20345 20768 20668 20770
rect 20345 20712 20350 20768
rect 20406 20712 20668 20768
rect 20345 20710 20668 20712
rect 20345 20707 20411 20710
rect 20662 20708 20668 20710
rect 20732 20708 20738 20772
rect 20808 20770 20868 20846
rect 22737 20904 27495 20906
rect 22737 20848 22742 20904
rect 22798 20848 27434 20904
rect 27490 20848 27495 20904
rect 22737 20846 27495 20848
rect 22737 20843 22803 20846
rect 27429 20843 27495 20846
rect 24485 20770 24551 20773
rect 20808 20768 24551 20770
rect 20808 20712 24490 20768
rect 24546 20712 24551 20768
rect 20808 20710 24551 20712
rect 24485 20707 24551 20710
rect 25446 20708 25452 20772
rect 25516 20770 25522 20772
rect 25865 20770 25931 20773
rect 25516 20768 25931 20770
rect 25516 20712 25870 20768
rect 25926 20712 25931 20768
rect 25516 20710 25931 20712
rect 25516 20708 25522 20710
rect 25865 20707 25931 20710
rect 26550 20708 26556 20772
rect 26620 20770 26626 20772
rect 27245 20770 27311 20773
rect 26620 20768 27311 20770
rect 26620 20712 27250 20768
rect 27306 20712 27311 20768
rect 26620 20710 27311 20712
rect 26620 20708 26626 20710
rect 27245 20707 27311 20710
rect 9213 20632 12220 20634
rect 9213 20576 9218 20632
rect 9274 20576 12220 20632
rect 9213 20574 12220 20576
rect 12893 20634 12959 20637
rect 15009 20634 15075 20637
rect 12893 20632 15075 20634
rect 12893 20576 12898 20632
rect 12954 20576 15014 20632
rect 15070 20576 15075 20632
rect 12893 20574 15075 20576
rect 9213 20571 9279 20574
rect 12893 20571 12959 20574
rect 15009 20571 15075 20574
rect 16205 20634 16271 20637
rect 30097 20634 30163 20637
rect 16205 20632 30163 20634
rect 16205 20576 16210 20632
rect 16266 20576 30102 20632
rect 30158 20576 30163 20632
rect 16205 20574 30163 20576
rect 16205 20571 16271 20574
rect 30097 20571 30163 20574
rect 6821 20498 6887 20501
rect 22553 20498 22619 20501
rect 6821 20496 22619 20498
rect 6821 20440 6826 20496
rect 6882 20440 22558 20496
rect 22614 20440 22619 20496
rect 6821 20438 22619 20440
rect 6821 20435 6887 20438
rect 22553 20435 22619 20438
rect 23841 20498 23907 20501
rect 26785 20498 26851 20501
rect 23841 20496 26851 20498
rect 23841 20440 23846 20496
rect 23902 20440 26790 20496
rect 26846 20440 26851 20496
rect 23841 20438 26851 20440
rect 23841 20435 23907 20438
rect 26785 20435 26851 20438
rect 27981 20498 28047 20501
rect 30414 20498 30420 20500
rect 27981 20496 30420 20498
rect 27981 20440 27986 20496
rect 28042 20440 30420 20496
rect 27981 20438 30420 20440
rect 27981 20435 28047 20438
rect 30414 20436 30420 20438
rect 30484 20436 30490 20500
rect 32397 20498 32463 20501
rect 33200 20498 34000 20528
rect 32397 20496 34000 20498
rect 32397 20440 32402 20496
rect 32458 20440 34000 20496
rect 32397 20438 34000 20440
rect 32397 20435 32463 20438
rect 33200 20408 34000 20438
rect 3182 20300 3188 20364
rect 3252 20362 3258 20364
rect 4797 20362 4863 20365
rect 5993 20362 6059 20365
rect 3252 20302 4722 20362
rect 3252 20300 3258 20302
rect 4662 20226 4722 20302
rect 4797 20360 6059 20362
rect 4797 20304 4802 20360
rect 4858 20304 5998 20360
rect 6054 20304 6059 20360
rect 4797 20302 6059 20304
rect 4797 20299 4863 20302
rect 5993 20299 6059 20302
rect 6637 20360 6746 20365
rect 6637 20304 6642 20360
rect 6698 20304 6746 20360
rect 6637 20302 6746 20304
rect 10501 20362 10567 20365
rect 12198 20362 12204 20364
rect 10501 20360 12204 20362
rect 10501 20304 10506 20360
rect 10562 20304 12204 20360
rect 10501 20302 12204 20304
rect 6637 20299 6703 20302
rect 10501 20299 10567 20302
rect 12198 20300 12204 20302
rect 12268 20300 12274 20364
rect 14089 20362 14155 20365
rect 14457 20362 14523 20365
rect 14089 20360 14523 20362
rect 14089 20304 14094 20360
rect 14150 20304 14462 20360
rect 14518 20304 14523 20360
rect 14089 20302 14523 20304
rect 14089 20299 14155 20302
rect 14457 20299 14523 20302
rect 17125 20362 17191 20365
rect 30373 20362 30439 20365
rect 17125 20360 30439 20362
rect 17125 20304 17130 20360
rect 17186 20304 30378 20360
rect 30434 20304 30439 20360
rect 17125 20302 30439 20304
rect 17125 20299 17191 20302
rect 30373 20299 30439 20302
rect 9581 20226 9647 20229
rect 11789 20228 11855 20229
rect 11789 20226 11836 20228
rect 4662 20166 7850 20226
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 1894 19892 1900 19956
rect 1964 19954 1970 19956
rect 7557 19954 7623 19957
rect 1964 19952 7623 19954
rect 1964 19896 7562 19952
rect 7618 19896 7623 19952
rect 1964 19894 7623 19896
rect 1964 19892 1970 19894
rect 7557 19891 7623 19894
rect 2497 19818 2563 19821
rect 5942 19818 5948 19820
rect 2497 19816 5948 19818
rect 2497 19760 2502 19816
rect 2558 19760 5948 19816
rect 2497 19758 5948 19760
rect 2497 19755 2563 19758
rect 5942 19756 5948 19758
rect 6012 19756 6018 19820
rect 1853 19682 1919 19685
rect 2262 19682 2268 19684
rect 1853 19680 2268 19682
rect 1853 19624 1858 19680
rect 1914 19624 2268 19680
rect 1853 19622 2268 19624
rect 1853 19619 1919 19622
rect 2262 19620 2268 19622
rect 2332 19620 2338 19684
rect 3366 19620 3372 19684
rect 3436 19682 3442 19684
rect 4061 19682 4127 19685
rect 3436 19680 4127 19682
rect 3436 19624 4066 19680
rect 4122 19624 4127 19680
rect 3436 19622 4127 19624
rect 7790 19682 7850 20166
rect 9581 20224 11836 20226
rect 11900 20226 11906 20228
rect 9581 20168 9586 20224
rect 9642 20168 11794 20224
rect 9581 20166 11836 20168
rect 9581 20163 9647 20166
rect 11789 20164 11836 20166
rect 11900 20166 11982 20226
rect 11900 20164 11906 20166
rect 12198 20164 12204 20228
rect 12268 20226 12274 20228
rect 14273 20226 14339 20229
rect 12268 20224 14339 20226
rect 12268 20168 14278 20224
rect 14334 20168 14339 20224
rect 12268 20166 14339 20168
rect 14460 20226 14520 20299
rect 26509 20226 26575 20229
rect 14460 20224 26575 20226
rect 14460 20168 26514 20224
rect 26570 20168 26575 20224
rect 14460 20166 26575 20168
rect 12268 20164 12274 20166
rect 11789 20163 11855 20164
rect 14273 20163 14339 20166
rect 26509 20163 26575 20166
rect 7925 20090 7991 20093
rect 16573 20090 16639 20093
rect 7925 20088 16639 20090
rect 7925 20032 7930 20088
rect 7986 20032 16578 20088
rect 16634 20032 16639 20088
rect 7925 20030 16639 20032
rect 7925 20027 7991 20030
rect 16573 20027 16639 20030
rect 18086 20028 18092 20092
rect 18156 20090 18162 20092
rect 18321 20090 18387 20093
rect 18156 20088 18387 20090
rect 18156 20032 18326 20088
rect 18382 20032 18387 20088
rect 18156 20030 18387 20032
rect 18156 20028 18162 20030
rect 18321 20027 18387 20030
rect 19374 20028 19380 20092
rect 19444 20090 19450 20092
rect 19701 20090 19767 20093
rect 19444 20088 19767 20090
rect 19444 20032 19706 20088
rect 19762 20032 19767 20088
rect 19444 20030 19767 20032
rect 19444 20028 19450 20030
rect 19701 20027 19767 20030
rect 19885 20090 19951 20093
rect 21081 20090 21147 20093
rect 19885 20088 21147 20090
rect 19885 20032 19890 20088
rect 19946 20032 21086 20088
rect 21142 20032 21147 20088
rect 19885 20030 21147 20032
rect 19885 20027 19951 20030
rect 21081 20027 21147 20030
rect 24761 20090 24827 20093
rect 24894 20090 24900 20092
rect 24761 20088 24900 20090
rect 24761 20032 24766 20088
rect 24822 20032 24900 20088
rect 24761 20030 24900 20032
rect 24761 20027 24827 20030
rect 24894 20028 24900 20030
rect 24964 20028 24970 20092
rect 31293 20090 31359 20093
rect 25086 20088 31359 20090
rect 25086 20032 31298 20088
rect 31354 20032 31359 20088
rect 25086 20030 31359 20032
rect 10225 19954 10291 19957
rect 10685 19954 10751 19957
rect 10225 19952 10751 19954
rect 10225 19896 10230 19952
rect 10286 19896 10690 19952
rect 10746 19896 10751 19952
rect 10225 19894 10751 19896
rect 10225 19891 10291 19894
rect 10685 19891 10751 19894
rect 11605 19956 11671 19957
rect 11605 19952 11652 19956
rect 11716 19954 11722 19956
rect 11881 19954 11947 19957
rect 13670 19954 13676 19956
rect 11605 19896 11610 19952
rect 11605 19892 11652 19896
rect 11716 19894 11762 19954
rect 11881 19952 13676 19954
rect 11881 19896 11886 19952
rect 11942 19896 13676 19952
rect 11881 19894 13676 19896
rect 11716 19892 11722 19894
rect 11605 19891 11671 19892
rect 11881 19891 11947 19894
rect 13670 19892 13676 19894
rect 13740 19892 13746 19956
rect 14641 19954 14707 19957
rect 18137 19954 18203 19957
rect 14276 19952 18203 19954
rect 14276 19896 14646 19952
rect 14702 19896 18142 19952
rect 18198 19896 18203 19952
rect 14276 19894 18203 19896
rect 8201 19818 8267 19821
rect 14276 19818 14336 19894
rect 14641 19891 14707 19894
rect 18137 19891 18203 19894
rect 21766 19892 21772 19956
rect 21836 19954 21842 19956
rect 22553 19954 22619 19957
rect 25086 19954 25146 20030
rect 31293 20027 31359 20030
rect 26049 19956 26115 19957
rect 21836 19952 25146 19954
rect 21836 19896 22558 19952
rect 22614 19896 25146 19952
rect 21836 19894 25146 19896
rect 21836 19892 21842 19894
rect 22553 19891 22619 19894
rect 25998 19892 26004 19956
rect 26068 19954 26115 19956
rect 26068 19952 26160 19954
rect 26110 19896 26160 19952
rect 26068 19894 26160 19896
rect 26068 19892 26115 19894
rect 26049 19891 26115 19892
rect 8201 19816 14336 19818
rect 8201 19760 8206 19816
rect 8262 19760 14336 19816
rect 8201 19758 14336 19760
rect 14549 19818 14615 19821
rect 23841 19818 23907 19821
rect 25773 19820 25839 19821
rect 14549 19816 23907 19818
rect 14549 19760 14554 19816
rect 14610 19760 23846 19816
rect 23902 19760 23907 19816
rect 14549 19758 23907 19760
rect 8201 19755 8267 19758
rect 14549 19755 14615 19758
rect 23841 19755 23907 19758
rect 25262 19756 25268 19820
rect 25332 19818 25338 19820
rect 25773 19818 25820 19820
rect 25332 19816 25820 19818
rect 25332 19760 25778 19816
rect 25332 19758 25820 19760
rect 25332 19756 25338 19758
rect 25773 19756 25820 19758
rect 25884 19756 25890 19820
rect 32397 19818 32463 19821
rect 33200 19818 34000 19848
rect 32397 19816 34000 19818
rect 32397 19760 32402 19816
rect 32458 19760 34000 19816
rect 32397 19758 34000 19760
rect 25773 19755 25839 19756
rect 32397 19755 32463 19758
rect 33200 19728 34000 19758
rect 12525 19682 12591 19685
rect 13353 19682 13419 19685
rect 7790 19622 12082 19682
rect 3436 19620 3442 19622
rect 4061 19619 4127 19622
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 2262 19484 2268 19548
rect 2332 19546 2338 19548
rect 2865 19546 2931 19549
rect 4705 19546 4771 19549
rect 2332 19486 2790 19546
rect 2332 19484 2338 19486
rect 2078 19348 2084 19412
rect 2148 19348 2154 19412
rect 2730 19410 2790 19486
rect 2865 19544 4771 19546
rect 2865 19488 2870 19544
rect 2926 19488 4710 19544
rect 4766 19488 4771 19544
rect 2865 19486 4771 19488
rect 2865 19483 2931 19486
rect 4705 19483 4771 19486
rect 9673 19546 9739 19549
rect 9806 19546 9812 19548
rect 9673 19544 9812 19546
rect 9673 19488 9678 19544
rect 9734 19488 9812 19544
rect 9673 19486 9812 19488
rect 9673 19483 9739 19486
rect 9806 19484 9812 19486
rect 9876 19484 9882 19548
rect 7557 19410 7623 19413
rect 2730 19408 7623 19410
rect 2730 19352 7562 19408
rect 7618 19352 7623 19408
rect 2730 19350 7623 19352
rect 2086 19274 2146 19348
rect 7557 19347 7623 19350
rect 9438 19348 9444 19412
rect 9508 19410 9514 19412
rect 10542 19410 10548 19412
rect 9508 19350 10548 19410
rect 9508 19348 9514 19350
rect 10542 19348 10548 19350
rect 10612 19348 10618 19412
rect 12022 19410 12082 19622
rect 12525 19680 13419 19682
rect 12525 19624 12530 19680
rect 12586 19624 13358 19680
rect 13414 19624 13419 19680
rect 12525 19622 13419 19624
rect 12525 19619 12591 19622
rect 13353 19619 13419 19622
rect 13670 19620 13676 19684
rect 13740 19682 13746 19684
rect 19425 19682 19491 19685
rect 13740 19680 19491 19682
rect 13740 19624 19430 19680
rect 19486 19624 19491 19680
rect 13740 19622 19491 19624
rect 13740 19620 13746 19622
rect 19425 19619 19491 19622
rect 20805 19682 20871 19685
rect 21030 19682 21036 19684
rect 20805 19680 21036 19682
rect 20805 19624 20810 19680
rect 20866 19624 21036 19680
rect 20805 19622 21036 19624
rect 20805 19619 20871 19622
rect 21030 19620 21036 19622
rect 21100 19620 21106 19684
rect 24945 19682 25011 19685
rect 26693 19682 26759 19685
rect 28257 19682 28323 19685
rect 24945 19680 28323 19682
rect 24945 19624 24950 19680
rect 25006 19624 26698 19680
rect 26754 19624 28262 19680
rect 28318 19624 28323 19680
rect 24945 19622 28323 19624
rect 24945 19619 25011 19622
rect 26693 19619 26759 19622
rect 28257 19619 28323 19622
rect 12433 19546 12499 19549
rect 15929 19546 15995 19549
rect 20621 19546 20687 19549
rect 26417 19546 26483 19549
rect 12433 19544 15995 19546
rect 12433 19488 12438 19544
rect 12494 19488 15934 19544
rect 15990 19488 15995 19544
rect 12433 19486 15995 19488
rect 12433 19483 12499 19486
rect 15929 19483 15995 19486
rect 19290 19544 26483 19546
rect 19290 19488 20626 19544
rect 20682 19488 26422 19544
rect 26478 19488 26483 19544
rect 19290 19486 26483 19488
rect 13905 19410 13971 19413
rect 12022 19408 13971 19410
rect 12022 19352 13910 19408
rect 13966 19352 13971 19408
rect 12022 19350 13971 19352
rect 13905 19347 13971 19350
rect 14774 19348 14780 19412
rect 14844 19410 14850 19412
rect 14917 19410 14983 19413
rect 14844 19408 14983 19410
rect 14844 19352 14922 19408
rect 14978 19352 14983 19408
rect 14844 19350 14983 19352
rect 14844 19348 14850 19350
rect 14917 19347 14983 19350
rect 9673 19274 9739 19277
rect 2086 19272 9739 19274
rect 2086 19216 9678 19272
rect 9734 19216 9739 19272
rect 2086 19214 9739 19216
rect 9673 19211 9739 19214
rect 10869 19276 10935 19277
rect 10869 19272 10916 19276
rect 10980 19274 10986 19276
rect 11145 19274 11211 19277
rect 12525 19274 12591 19277
rect 10869 19216 10874 19272
rect 10869 19212 10916 19216
rect 10980 19214 11026 19274
rect 11145 19272 12591 19274
rect 11145 19216 11150 19272
rect 11206 19216 12530 19272
rect 12586 19216 12591 19272
rect 11145 19214 12591 19216
rect 10980 19212 10986 19214
rect 10869 19211 10935 19212
rect 11145 19211 11211 19214
rect 12525 19211 12591 19214
rect 12801 19274 12867 19277
rect 13118 19274 13124 19276
rect 12801 19272 13124 19274
rect 12801 19216 12806 19272
rect 12862 19216 13124 19272
rect 12801 19214 13124 19216
rect 12801 19211 12867 19214
rect 13118 19212 13124 19214
rect 13188 19212 13194 19276
rect 13670 19212 13676 19276
rect 13740 19274 13746 19276
rect 13740 19214 18154 19274
rect 13740 19212 13746 19214
rect 0 19138 800 19168
rect 1301 19138 1367 19141
rect 0 19136 1367 19138
rect 0 19080 1306 19136
rect 1362 19080 1367 19136
rect 0 19078 1367 19080
rect 0 19048 800 19078
rect 1301 19075 1367 19078
rect 5533 19138 5599 19141
rect 7966 19138 7972 19140
rect 5533 19136 7972 19138
rect 5533 19080 5538 19136
rect 5594 19080 7972 19136
rect 5533 19078 7972 19080
rect 5533 19075 5599 19078
rect 7966 19076 7972 19078
rect 8036 19076 8042 19140
rect 12525 19138 12591 19141
rect 13486 19138 13492 19140
rect 12525 19136 13492 19138
rect 12525 19080 12530 19136
rect 12586 19080 13492 19136
rect 12525 19078 13492 19080
rect 12525 19075 12591 19078
rect 13486 19076 13492 19078
rect 13556 19076 13562 19140
rect 15101 19138 15167 19141
rect 16246 19138 16252 19140
rect 15101 19136 16252 19138
rect 15101 19080 15106 19136
rect 15162 19080 16252 19136
rect 15101 19078 16252 19080
rect 15101 19075 15167 19078
rect 16246 19076 16252 19078
rect 16316 19076 16322 19140
rect 16389 19138 16455 19141
rect 17769 19138 17835 19141
rect 16389 19136 17835 19138
rect 16389 19080 16394 19136
rect 16450 19080 17774 19136
rect 17830 19080 17835 19136
rect 16389 19078 17835 19080
rect 18094 19138 18154 19214
rect 19290 19138 19350 19486
rect 20621 19483 20687 19486
rect 26417 19483 26483 19486
rect 20110 19348 20116 19412
rect 20180 19410 20186 19412
rect 20437 19410 20503 19413
rect 20180 19408 20503 19410
rect 20180 19352 20442 19408
rect 20498 19352 20503 19408
rect 20180 19350 20503 19352
rect 20180 19348 20186 19350
rect 20437 19347 20503 19350
rect 20713 19410 20779 19413
rect 21214 19410 21220 19412
rect 20713 19408 21220 19410
rect 20713 19352 20718 19408
rect 20774 19352 21220 19408
rect 20713 19350 21220 19352
rect 20713 19347 20779 19350
rect 21214 19348 21220 19350
rect 21284 19348 21290 19412
rect 22318 19348 22324 19412
rect 22388 19410 22394 19412
rect 23289 19410 23355 19413
rect 22388 19408 23355 19410
rect 22388 19352 23294 19408
rect 23350 19352 23355 19408
rect 22388 19350 23355 19352
rect 22388 19348 22394 19350
rect 23289 19347 23355 19350
rect 25773 19410 25839 19413
rect 32121 19410 32187 19413
rect 25773 19408 32187 19410
rect 25773 19352 25778 19408
rect 25834 19352 32126 19408
rect 32182 19352 32187 19408
rect 25773 19350 32187 19352
rect 25773 19347 25839 19350
rect 32121 19347 32187 19350
rect 20161 19274 20227 19277
rect 21725 19274 21791 19277
rect 28390 19274 28396 19276
rect 20161 19272 21650 19274
rect 20161 19216 20166 19272
rect 20222 19216 21650 19272
rect 20161 19214 21650 19216
rect 20161 19211 20227 19214
rect 18094 19078 19350 19138
rect 16389 19075 16455 19078
rect 17769 19075 17835 19078
rect 20846 19076 20852 19140
rect 20916 19138 20922 19140
rect 21449 19138 21515 19141
rect 20916 19136 21515 19138
rect 20916 19080 21454 19136
rect 21510 19080 21515 19136
rect 20916 19078 21515 19080
rect 21590 19138 21650 19214
rect 21725 19272 28396 19274
rect 21725 19216 21730 19272
rect 21786 19216 28396 19272
rect 21725 19214 28396 19216
rect 21725 19211 21791 19214
rect 28390 19212 28396 19214
rect 28460 19212 28466 19276
rect 24710 19138 24716 19140
rect 21590 19078 24716 19138
rect 20916 19076 20922 19078
rect 21449 19075 21515 19078
rect 24710 19076 24716 19078
rect 24780 19138 24786 19140
rect 24945 19138 25011 19141
rect 24780 19136 25011 19138
rect 24780 19080 24950 19136
rect 25006 19080 25011 19136
rect 24780 19078 25011 19080
rect 24780 19076 24786 19078
rect 24945 19075 25011 19078
rect 26509 19138 26575 19141
rect 29678 19138 29684 19140
rect 26509 19136 29684 19138
rect 26509 19080 26514 19136
rect 26570 19080 29684 19136
rect 26509 19078 29684 19080
rect 26509 19075 26575 19078
rect 29678 19076 29684 19078
rect 29748 19076 29754 19140
rect 32397 19138 32463 19141
rect 33200 19138 34000 19168
rect 32397 19136 34000 19138
rect 32397 19080 32402 19136
rect 32458 19080 34000 19136
rect 32397 19078 34000 19080
rect 32397 19075 32463 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 33200 19048 34000 19078
rect 4210 19007 4526 19008
rect 6310 18940 6316 19004
rect 6380 19002 6386 19004
rect 7005 19002 7071 19005
rect 6380 19000 7071 19002
rect 6380 18944 7010 19000
rect 7066 18944 7071 19000
rect 6380 18942 7071 18944
rect 6380 18940 6386 18942
rect 7005 18939 7071 18942
rect 10501 19002 10567 19005
rect 11881 19002 11947 19005
rect 10501 19000 11947 19002
rect 10501 18944 10506 19000
rect 10562 18944 11886 19000
rect 11942 18944 11947 19000
rect 10501 18942 11947 18944
rect 10501 18939 10567 18942
rect 11881 18939 11947 18942
rect 12157 19002 12223 19005
rect 15285 19002 15351 19005
rect 12157 19000 15351 19002
rect 12157 18944 12162 19000
rect 12218 18944 15290 19000
rect 15346 18944 15351 19000
rect 12157 18942 15351 18944
rect 12157 18939 12223 18942
rect 15285 18939 15351 18942
rect 16021 19002 16087 19005
rect 22461 19004 22527 19005
rect 22134 19002 22140 19004
rect 16021 19000 22140 19002
rect 16021 18944 16026 19000
rect 16082 18944 22140 19000
rect 16021 18942 22140 18944
rect 16021 18939 16087 18942
rect 22134 18940 22140 18942
rect 22204 18940 22210 19004
rect 22461 19002 22508 19004
rect 22416 19000 22508 19002
rect 22416 18944 22466 19000
rect 22416 18942 22508 18944
rect 22461 18940 22508 18942
rect 22572 18940 22578 19004
rect 30414 19002 30420 19004
rect 26190 18942 30420 19002
rect 22461 18939 22527 18940
rect 841 18866 907 18869
rect 6545 18866 6611 18869
rect 841 18864 6611 18866
rect 841 18808 846 18864
rect 902 18808 6550 18864
rect 6606 18808 6611 18864
rect 841 18806 6611 18808
rect 841 18803 907 18806
rect 6545 18803 6611 18806
rect 7005 18866 7071 18869
rect 21265 18866 21331 18869
rect 26190 18866 26250 18942
rect 30414 18940 30420 18942
rect 30484 18940 30490 19004
rect 7005 18864 17418 18866
rect 7005 18808 7010 18864
rect 7066 18808 17418 18864
rect 7005 18806 17418 18808
rect 7005 18803 7071 18806
rect 3509 18730 3575 18733
rect 5349 18730 5415 18733
rect 16021 18730 16087 18733
rect 3509 18728 5415 18730
rect 3509 18672 3514 18728
rect 3570 18672 5354 18728
rect 5410 18672 5415 18728
rect 3509 18670 5415 18672
rect 3509 18667 3575 18670
rect 5349 18667 5415 18670
rect 7468 18728 16087 18730
rect 7468 18672 16026 18728
rect 16082 18672 16087 18728
rect 7468 18670 16087 18672
rect 17358 18730 17418 18806
rect 21265 18864 26250 18866
rect 21265 18808 21270 18864
rect 21326 18808 26250 18864
rect 21265 18806 26250 18808
rect 29729 18866 29795 18869
rect 30925 18868 30991 18869
rect 30925 18866 30972 18868
rect 29729 18864 30972 18866
rect 31036 18866 31042 18868
rect 29729 18808 29734 18864
rect 29790 18808 30930 18864
rect 29729 18806 30972 18808
rect 21265 18803 21331 18806
rect 29729 18803 29795 18806
rect 30925 18804 30972 18806
rect 31036 18806 31118 18866
rect 31036 18804 31042 18806
rect 30925 18803 30991 18804
rect 22001 18730 22067 18733
rect 17358 18728 22067 18730
rect 17358 18672 22006 18728
rect 22062 18672 22067 18728
rect 17358 18670 22067 18672
rect 7468 18597 7528 18670
rect 16021 18667 16087 18670
rect 22001 18667 22067 18670
rect 22134 18668 22140 18732
rect 22204 18730 22210 18732
rect 22461 18730 22527 18733
rect 30598 18730 30604 18732
rect 22204 18670 22386 18730
rect 22204 18668 22210 18670
rect 6678 18532 6684 18596
rect 6748 18594 6754 18596
rect 7465 18594 7531 18597
rect 7649 18596 7715 18597
rect 6748 18592 7531 18594
rect 6748 18536 7470 18592
rect 7526 18536 7531 18592
rect 6748 18534 7531 18536
rect 6748 18532 6754 18534
rect 7465 18531 7531 18534
rect 7598 18532 7604 18596
rect 7668 18594 7715 18596
rect 9857 18594 9923 18597
rect 10358 18594 10364 18596
rect 7668 18592 7760 18594
rect 7710 18536 7760 18592
rect 7668 18534 7760 18536
rect 9857 18592 10364 18594
rect 9857 18536 9862 18592
rect 9918 18536 10364 18592
rect 9857 18534 10364 18536
rect 7668 18532 7715 18534
rect 7649 18531 7715 18532
rect 9857 18531 9923 18534
rect 10358 18532 10364 18534
rect 10428 18532 10434 18596
rect 11094 18532 11100 18596
rect 11164 18594 11170 18596
rect 11789 18594 11855 18597
rect 13721 18594 13787 18597
rect 11164 18592 13787 18594
rect 11164 18536 11794 18592
rect 11850 18536 13726 18592
rect 13782 18536 13787 18592
rect 11164 18534 13787 18536
rect 11164 18532 11170 18534
rect 11789 18531 11855 18534
rect 13721 18531 13787 18534
rect 14222 18532 14228 18596
rect 14292 18594 14298 18596
rect 14365 18594 14431 18597
rect 14292 18592 14431 18594
rect 14292 18536 14370 18592
rect 14426 18536 14431 18592
rect 14292 18534 14431 18536
rect 14292 18532 14298 18534
rect 14365 18531 14431 18534
rect 14641 18594 14707 18597
rect 18270 18594 18276 18596
rect 14641 18592 18276 18594
rect 14641 18536 14646 18592
rect 14702 18536 18276 18592
rect 14641 18534 18276 18536
rect 14641 18531 14707 18534
rect 18270 18532 18276 18534
rect 18340 18594 18346 18596
rect 21030 18594 21036 18596
rect 18340 18534 21036 18594
rect 18340 18532 18346 18534
rect 21030 18532 21036 18534
rect 21100 18532 21106 18596
rect 22326 18594 22386 18670
rect 22461 18728 30604 18730
rect 22461 18672 22466 18728
rect 22522 18672 30604 18728
rect 22461 18670 30604 18672
rect 22461 18667 22527 18670
rect 30598 18668 30604 18670
rect 30668 18668 30674 18732
rect 25630 18594 25636 18596
rect 22326 18534 25636 18594
rect 25630 18532 25636 18534
rect 25700 18594 25706 18596
rect 28809 18594 28875 18597
rect 25700 18592 28875 18594
rect 25700 18536 28814 18592
rect 28870 18536 28875 18592
rect 25700 18534 28875 18536
rect 25700 18532 25706 18534
rect 28809 18531 28875 18534
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 5625 18458 5691 18461
rect 5758 18458 5764 18460
rect 5625 18456 5764 18458
rect 5625 18400 5630 18456
rect 5686 18400 5764 18456
rect 5625 18398 5764 18400
rect 5625 18395 5691 18398
rect 5758 18396 5764 18398
rect 5828 18396 5834 18460
rect 12014 18396 12020 18460
rect 12084 18458 12090 18460
rect 12157 18458 12223 18461
rect 12084 18456 12223 18458
rect 12084 18400 12162 18456
rect 12218 18400 12223 18456
rect 12084 18398 12223 18400
rect 12084 18396 12090 18398
rect 12157 18395 12223 18398
rect 12341 18458 12407 18461
rect 12934 18458 12940 18460
rect 12341 18456 12940 18458
rect 12341 18400 12346 18456
rect 12402 18400 12940 18456
rect 12341 18398 12940 18400
rect 12341 18395 12407 18398
rect 12934 18396 12940 18398
rect 13004 18396 13010 18460
rect 13077 18458 13143 18461
rect 15653 18458 15719 18461
rect 13077 18456 15719 18458
rect 13077 18400 13082 18456
rect 13138 18400 15658 18456
rect 15714 18400 15719 18456
rect 13077 18398 15719 18400
rect 13077 18395 13143 18398
rect 15653 18395 15719 18398
rect 16021 18458 16087 18461
rect 26601 18458 26667 18461
rect 16021 18456 26667 18458
rect 16021 18400 16026 18456
rect 16082 18400 26606 18456
rect 26662 18400 26667 18456
rect 16021 18398 26667 18400
rect 16021 18395 16087 18398
rect 26601 18395 26667 18398
rect 606 18260 612 18324
rect 676 18322 682 18324
rect 7741 18322 7807 18325
rect 9029 18324 9095 18325
rect 9029 18322 9076 18324
rect 676 18320 7807 18322
rect 676 18264 7746 18320
rect 7802 18264 7807 18320
rect 676 18262 7807 18264
rect 8948 18320 9076 18322
rect 9140 18322 9146 18324
rect 12709 18322 12775 18325
rect 17309 18322 17375 18325
rect 8948 18264 9034 18320
rect 8948 18262 9076 18264
rect 676 18260 682 18262
rect 7741 18259 7807 18262
rect 9029 18260 9076 18262
rect 9140 18262 12450 18322
rect 9140 18260 9146 18262
rect 9029 18259 9095 18260
rect 11053 18186 11119 18189
rect 2730 18184 11119 18186
rect 2730 18128 11058 18184
rect 11114 18128 11119 18184
rect 2730 18126 11119 18128
rect 2730 18050 2790 18126
rect 11053 18123 11119 18126
rect 11646 18124 11652 18188
rect 11716 18186 11722 18188
rect 12157 18186 12223 18189
rect 11716 18184 12223 18186
rect 11716 18128 12162 18184
rect 12218 18128 12223 18184
rect 11716 18126 12223 18128
rect 12390 18186 12450 18262
rect 12709 18320 17375 18322
rect 12709 18264 12714 18320
rect 12770 18264 17314 18320
rect 17370 18264 17375 18320
rect 12709 18262 17375 18264
rect 12709 18259 12775 18262
rect 17309 18259 17375 18262
rect 18137 18322 18203 18325
rect 28257 18322 28323 18325
rect 18137 18320 28323 18322
rect 18137 18264 18142 18320
rect 18198 18264 28262 18320
rect 28318 18264 28323 18320
rect 18137 18262 28323 18264
rect 18137 18259 18203 18262
rect 28257 18259 28323 18262
rect 22553 18186 22619 18189
rect 12390 18184 22619 18186
rect 12390 18128 22558 18184
rect 22614 18128 22619 18184
rect 12390 18126 22619 18128
rect 11716 18124 11722 18126
rect 12157 18123 12223 18126
rect 22553 18123 22619 18126
rect 23422 18124 23428 18188
rect 23492 18186 23498 18188
rect 26233 18186 26299 18189
rect 23492 18184 26299 18186
rect 23492 18128 26238 18184
rect 26294 18128 26299 18184
rect 23492 18126 26299 18128
rect 23492 18124 23498 18126
rect 26233 18123 26299 18126
rect 2086 17990 2790 18050
rect 7465 18050 7531 18053
rect 7741 18050 7807 18053
rect 10501 18052 10567 18053
rect 10501 18050 10548 18052
rect 7465 18048 7807 18050
rect 7465 17992 7470 18048
rect 7526 17992 7746 18048
rect 7802 17992 7807 18048
rect 7465 17990 7807 17992
rect 10456 18048 10548 18050
rect 10456 17992 10506 18048
rect 10456 17990 10548 17992
rect 2086 17916 2146 17990
rect 7465 17987 7531 17990
rect 7741 17987 7807 17990
rect 10501 17988 10548 17990
rect 10612 17988 10618 18052
rect 11462 17988 11468 18052
rect 11532 18050 11538 18052
rect 14733 18050 14799 18053
rect 14958 18050 14964 18052
rect 11532 17990 14658 18050
rect 11532 17988 11538 17990
rect 10501 17987 10567 17988
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 2078 17852 2084 17916
rect 2148 17852 2154 17916
rect 2446 17852 2452 17916
rect 2516 17914 2522 17916
rect 3417 17914 3483 17917
rect 2516 17912 3483 17914
rect 2516 17856 3422 17912
rect 3478 17856 3483 17912
rect 2516 17854 3483 17856
rect 2516 17852 2522 17854
rect 3417 17851 3483 17854
rect 6453 17916 6519 17917
rect 6453 17912 6500 17916
rect 6564 17914 6570 17916
rect 6453 17856 6458 17912
rect 6453 17852 6500 17856
rect 6564 17854 6610 17914
rect 6564 17852 6570 17854
rect 8150 17852 8156 17916
rect 8220 17914 8226 17916
rect 8886 17914 8892 17916
rect 8220 17854 8892 17914
rect 8220 17852 8226 17854
rect 8886 17852 8892 17854
rect 8956 17852 8962 17916
rect 12198 17852 12204 17916
rect 12268 17914 12274 17916
rect 12985 17914 13051 17917
rect 12268 17912 13051 17914
rect 12268 17856 12990 17912
rect 13046 17856 13051 17912
rect 12268 17854 13051 17856
rect 12268 17852 12274 17854
rect 6453 17851 6519 17852
rect 12985 17851 13051 17854
rect 13261 17914 13327 17917
rect 14089 17914 14155 17917
rect 13261 17912 14155 17914
rect 13261 17856 13266 17912
rect 13322 17856 14094 17912
rect 14150 17856 14155 17912
rect 13261 17854 14155 17856
rect 14598 17914 14658 17990
rect 14733 18048 14964 18050
rect 14733 17992 14738 18048
rect 14794 17992 14964 18048
rect 14733 17990 14964 17992
rect 14733 17987 14799 17990
rect 14958 17988 14964 17990
rect 15028 17988 15034 18052
rect 18137 18050 18203 18053
rect 15150 18048 18203 18050
rect 15150 17992 18142 18048
rect 18198 17992 18203 18048
rect 15150 17990 18203 17992
rect 15150 17914 15210 17990
rect 18137 17987 18203 17990
rect 18822 17988 18828 18052
rect 18892 18050 18898 18052
rect 19241 18050 19307 18053
rect 18892 18048 19307 18050
rect 18892 17992 19246 18048
rect 19302 17992 19307 18048
rect 18892 17990 19307 17992
rect 18892 17988 18898 17990
rect 19241 17987 19307 17990
rect 19425 18048 19491 18053
rect 19425 17992 19430 18048
rect 19486 17992 19491 18048
rect 19425 17987 19491 17992
rect 22001 18050 22067 18053
rect 24577 18050 24643 18053
rect 22001 18048 24643 18050
rect 22001 17992 22006 18048
rect 22062 17992 24582 18048
rect 24638 17992 24643 18048
rect 22001 17990 24643 17992
rect 22001 17987 22067 17990
rect 24577 17987 24643 17990
rect 25589 18050 25655 18053
rect 28993 18052 29059 18053
rect 27654 18050 27660 18052
rect 25589 18048 27660 18050
rect 25589 17992 25594 18048
rect 25650 17992 27660 18048
rect 25589 17990 27660 17992
rect 25589 17987 25655 17990
rect 27654 17988 27660 17990
rect 27724 17988 27730 18052
rect 28942 18050 28948 18052
rect 28902 17990 28948 18050
rect 29012 18048 29059 18052
rect 29054 17992 29059 18048
rect 28942 17988 28948 17990
rect 29012 17988 29059 17992
rect 28993 17987 29059 17988
rect 14598 17854 15210 17914
rect 19428 17914 19488 17987
rect 23238 17914 23244 17916
rect 19428 17854 23244 17914
rect 13261 17851 13327 17854
rect 14089 17851 14155 17854
rect 23238 17852 23244 17854
rect 23308 17852 23314 17916
rect 2630 17716 2636 17780
rect 2700 17778 2706 17780
rect 4797 17778 4863 17781
rect 2700 17776 4863 17778
rect 2700 17720 4802 17776
rect 4858 17720 4863 17776
rect 2700 17718 4863 17720
rect 2700 17716 2706 17718
rect 4797 17715 4863 17718
rect 9990 17716 9996 17780
rect 10060 17778 10066 17780
rect 15101 17778 15167 17781
rect 10060 17776 15167 17778
rect 10060 17720 15106 17776
rect 15162 17720 15167 17776
rect 10060 17718 15167 17720
rect 10060 17716 10066 17718
rect 15101 17715 15167 17718
rect 16297 17778 16363 17781
rect 26509 17778 26575 17781
rect 16297 17776 26575 17778
rect 16297 17720 16302 17776
rect 16358 17720 26514 17776
rect 26570 17720 26575 17776
rect 16297 17718 26575 17720
rect 16297 17715 16363 17718
rect 26509 17715 26575 17718
rect 32397 17778 32463 17781
rect 33200 17778 34000 17808
rect 32397 17776 34000 17778
rect 32397 17720 32402 17776
rect 32458 17720 34000 17776
rect 32397 17718 34000 17720
rect 32397 17715 32463 17718
rect 33200 17688 34000 17718
rect 933 17642 999 17645
rect 7782 17642 7788 17644
rect 933 17640 7788 17642
rect 933 17584 938 17640
rect 994 17584 7788 17640
rect 933 17582 7788 17584
rect 933 17579 999 17582
rect 7782 17580 7788 17582
rect 7852 17580 7858 17644
rect 10501 17642 10567 17645
rect 14406 17642 14412 17644
rect 10501 17640 14412 17642
rect 10501 17584 10506 17640
rect 10562 17584 14412 17640
rect 10501 17582 14412 17584
rect 10501 17579 10567 17582
rect 14406 17580 14412 17582
rect 14476 17580 14482 17644
rect 14825 17642 14891 17645
rect 22737 17642 22803 17645
rect 14825 17640 22803 17642
rect 14825 17584 14830 17640
rect 14886 17584 22742 17640
rect 22798 17584 22803 17640
rect 14825 17582 22803 17584
rect 14825 17579 14891 17582
rect 22737 17579 22803 17582
rect 11053 17506 11119 17509
rect 23657 17506 23723 17509
rect 11053 17504 23723 17506
rect 11053 17448 11058 17504
rect 11114 17448 23662 17504
rect 23718 17448 23723 17504
rect 11053 17446 23723 17448
rect 11053 17443 11119 17446
rect 23657 17443 23723 17446
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 6637 17370 6703 17373
rect 11237 17370 11303 17373
rect 6502 17368 6703 17370
rect 6502 17312 6642 17368
rect 6698 17312 6703 17368
rect 6502 17310 6703 17312
rect 2681 17234 2747 17237
rect 3141 17234 3207 17237
rect 6502 17234 6562 17310
rect 6637 17307 6703 17310
rect 6870 17368 11303 17370
rect 6870 17312 11242 17368
rect 11298 17312 11303 17368
rect 6870 17310 11303 17312
rect 2681 17232 3207 17234
rect 2681 17176 2686 17232
rect 2742 17176 3146 17232
rect 3202 17176 3207 17232
rect 2681 17174 3207 17176
rect 2681 17171 2747 17174
rect 3141 17171 3207 17174
rect 3742 17174 6562 17234
rect 6637 17234 6703 17237
rect 6870 17234 6930 17310
rect 11237 17307 11303 17310
rect 11421 17368 11487 17373
rect 11421 17312 11426 17368
rect 11482 17312 11487 17368
rect 11421 17307 11487 17312
rect 12985 17370 13051 17373
rect 15142 17370 15148 17372
rect 12985 17368 15148 17370
rect 12985 17312 12990 17368
rect 13046 17312 15148 17368
rect 12985 17310 15148 17312
rect 12985 17307 13051 17310
rect 15142 17308 15148 17310
rect 15212 17308 15218 17372
rect 15469 17370 15535 17373
rect 15878 17370 15884 17372
rect 15469 17368 15884 17370
rect 15469 17312 15474 17368
rect 15530 17312 15884 17368
rect 15469 17310 15884 17312
rect 15469 17307 15535 17310
rect 15878 17308 15884 17310
rect 15948 17370 15954 17372
rect 18229 17370 18295 17373
rect 15948 17368 18295 17370
rect 15948 17312 18234 17368
rect 18290 17312 18295 17368
rect 15948 17310 18295 17312
rect 15948 17308 15954 17310
rect 18229 17307 18295 17310
rect 23974 17308 23980 17372
rect 24044 17370 24050 17372
rect 24710 17370 24716 17372
rect 24044 17310 24716 17370
rect 24044 17308 24050 17310
rect 24710 17308 24716 17310
rect 24780 17370 24786 17372
rect 27705 17370 27771 17373
rect 24780 17368 27771 17370
rect 24780 17312 27710 17368
rect 27766 17312 27771 17368
rect 24780 17310 27771 17312
rect 24780 17308 24786 17310
rect 27705 17307 27771 17310
rect 6637 17232 6930 17234
rect 6637 17176 6642 17232
rect 6698 17176 6930 17232
rect 6637 17174 6930 17176
rect 9673 17234 9739 17237
rect 11053 17234 11119 17237
rect 11424 17234 11484 17307
rect 9673 17232 11484 17234
rect 9673 17176 9678 17232
rect 9734 17176 11058 17232
rect 11114 17176 11484 17232
rect 9673 17174 11484 17176
rect 11697 17234 11763 17237
rect 21766 17234 21772 17236
rect 11697 17232 21772 17234
rect 11697 17176 11702 17232
rect 11758 17176 21772 17232
rect 11697 17174 21772 17176
rect 841 16554 907 16557
rect 798 16552 907 16554
rect 798 16496 846 16552
rect 902 16496 907 16552
rect 798 16491 907 16496
rect 798 16448 858 16491
rect 0 16358 858 16448
rect 3049 16418 3115 16421
rect 3742 16418 3802 17174
rect 6637 17171 6703 17174
rect 9673 17171 9739 17174
rect 11053 17171 11119 17174
rect 11697 17171 11763 17174
rect 21766 17172 21772 17174
rect 21836 17172 21842 17236
rect 23054 17172 23060 17236
rect 23124 17234 23130 17236
rect 23197 17234 23263 17237
rect 23124 17232 23263 17234
rect 23124 17176 23202 17232
rect 23258 17176 23263 17232
rect 23124 17174 23263 17176
rect 23124 17172 23130 17174
rect 23197 17171 23263 17174
rect 24209 17234 24275 17237
rect 25078 17234 25084 17236
rect 24209 17232 25084 17234
rect 24209 17176 24214 17232
rect 24270 17176 25084 17232
rect 24209 17174 25084 17176
rect 24209 17171 24275 17174
rect 25078 17172 25084 17174
rect 25148 17172 25154 17236
rect 25998 17172 26004 17236
rect 26068 17234 26074 17236
rect 32673 17234 32739 17237
rect 26068 17232 32739 17234
rect 26068 17176 32678 17232
rect 32734 17176 32739 17232
rect 26068 17174 32739 17176
rect 26068 17172 26074 17174
rect 32673 17171 32739 17174
rect 3877 17098 3943 17101
rect 5165 17098 5231 17101
rect 8293 17098 8359 17101
rect 3877 17096 5090 17098
rect 3877 17040 3882 17096
rect 3938 17040 5090 17096
rect 3877 17038 5090 17040
rect 3877 17035 3943 17038
rect 5030 16962 5090 17038
rect 5165 17096 8359 17098
rect 5165 17040 5170 17096
rect 5226 17040 8298 17096
rect 8354 17040 8359 17096
rect 5165 17038 8359 17040
rect 5165 17035 5231 17038
rect 8293 17035 8359 17038
rect 8661 17098 8727 17101
rect 11605 17098 11671 17101
rect 8661 17096 11671 17098
rect 8661 17040 8666 17096
rect 8722 17040 11610 17096
rect 11666 17040 11671 17096
rect 8661 17038 11671 17040
rect 8661 17035 8727 17038
rect 11605 17035 11671 17038
rect 12157 17098 12223 17101
rect 12893 17098 12959 17101
rect 12157 17096 12959 17098
rect 12157 17040 12162 17096
rect 12218 17040 12898 17096
rect 12954 17040 12959 17096
rect 12157 17038 12959 17040
rect 12157 17035 12223 17038
rect 12893 17035 12959 17038
rect 14273 17098 14339 17101
rect 32397 17098 32463 17101
rect 33200 17098 34000 17128
rect 14273 17096 22110 17098
rect 14273 17040 14278 17096
rect 14334 17040 22110 17096
rect 14273 17038 22110 17040
rect 14273 17035 14339 17038
rect 6821 16962 6887 16965
rect 5030 16960 6887 16962
rect 5030 16904 6826 16960
rect 6882 16904 6887 16960
rect 5030 16902 6887 16904
rect 6821 16899 6887 16902
rect 9806 16900 9812 16964
rect 9876 16962 9882 16964
rect 9949 16962 10015 16965
rect 9876 16960 10015 16962
rect 9876 16904 9954 16960
rect 10010 16904 10015 16960
rect 9876 16902 10015 16904
rect 9876 16900 9882 16902
rect 9949 16899 10015 16902
rect 10225 16962 10291 16965
rect 14276 16962 14336 17035
rect 10225 16960 14336 16962
rect 10225 16904 10230 16960
rect 10286 16904 14336 16960
rect 10225 16902 14336 16904
rect 10225 16899 10291 16902
rect 14406 16900 14412 16964
rect 14476 16962 14482 16964
rect 17902 16962 17908 16964
rect 14476 16902 17908 16962
rect 14476 16900 14482 16902
rect 17902 16900 17908 16902
rect 17972 16900 17978 16964
rect 22050 16962 22110 17038
rect 32397 17096 34000 17098
rect 32397 17040 32402 17096
rect 32458 17040 34000 17096
rect 32397 17038 34000 17040
rect 32397 17035 32463 17038
rect 33200 17008 34000 17038
rect 23933 16962 23999 16965
rect 24158 16962 24164 16964
rect 22050 16960 24164 16962
rect 22050 16904 23938 16960
rect 23994 16904 24164 16960
rect 22050 16902 24164 16904
rect 23933 16899 23999 16902
rect 24158 16900 24164 16902
rect 24228 16900 24234 16964
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 8937 16826 9003 16829
rect 10501 16826 10567 16829
rect 13261 16826 13327 16829
rect 6456 16766 8770 16826
rect 4110 16630 4906 16690
rect 3877 16554 3943 16557
rect 4110 16554 4170 16630
rect 3877 16552 4170 16554
rect 3877 16496 3882 16552
rect 3938 16496 4170 16552
rect 3877 16494 4170 16496
rect 4337 16554 4403 16557
rect 4654 16554 4660 16556
rect 4337 16552 4660 16554
rect 4337 16496 4342 16552
rect 4398 16496 4660 16552
rect 4337 16494 4660 16496
rect 3877 16491 3943 16494
rect 4337 16491 4403 16494
rect 4654 16492 4660 16494
rect 4724 16492 4730 16556
rect 4846 16554 4906 16630
rect 5758 16628 5764 16692
rect 5828 16690 5834 16692
rect 6456 16690 6516 16766
rect 5828 16630 6516 16690
rect 8710 16690 8770 16766
rect 8937 16824 10567 16826
rect 8937 16768 8942 16824
rect 8998 16768 10506 16824
rect 10562 16768 10567 16824
rect 8937 16766 10567 16768
rect 8937 16763 9003 16766
rect 10501 16763 10567 16766
rect 12390 16824 13327 16826
rect 12390 16768 13266 16824
rect 13322 16768 13327 16824
rect 12390 16766 13327 16768
rect 12390 16690 12450 16766
rect 13261 16763 13327 16766
rect 15326 16764 15332 16828
rect 15396 16826 15402 16828
rect 15561 16826 15627 16829
rect 15396 16824 15627 16826
rect 15396 16768 15566 16824
rect 15622 16768 15627 16824
rect 15396 16766 15627 16768
rect 15396 16764 15402 16766
rect 15561 16763 15627 16766
rect 15694 16764 15700 16828
rect 15764 16826 15770 16828
rect 17125 16826 17191 16829
rect 15764 16824 17191 16826
rect 15764 16768 17130 16824
rect 17186 16768 17191 16824
rect 15764 16766 17191 16768
rect 15764 16764 15770 16766
rect 17125 16763 17191 16766
rect 19333 16826 19399 16829
rect 25129 16826 25195 16829
rect 19333 16824 25195 16826
rect 19333 16768 19338 16824
rect 19394 16768 25134 16824
rect 25190 16768 25195 16824
rect 19333 16766 25195 16768
rect 19333 16763 19399 16766
rect 25129 16763 25195 16766
rect 8710 16630 12450 16690
rect 5828 16628 5834 16630
rect 12566 16628 12572 16692
rect 12636 16690 12642 16692
rect 12934 16690 12940 16692
rect 12636 16630 12940 16690
rect 12636 16628 12642 16630
rect 12934 16628 12940 16630
rect 13004 16628 13010 16692
rect 14273 16690 14339 16693
rect 18689 16690 18755 16693
rect 14273 16688 18755 16690
rect 14273 16632 14278 16688
rect 14334 16632 18694 16688
rect 18750 16632 18755 16688
rect 14273 16630 18755 16632
rect 14273 16627 14339 16630
rect 18689 16627 18755 16630
rect 19742 16628 19748 16692
rect 19812 16690 19818 16692
rect 19977 16690 20043 16693
rect 19812 16688 20043 16690
rect 19812 16632 19982 16688
rect 20038 16632 20043 16688
rect 19812 16630 20043 16632
rect 19812 16628 19818 16630
rect 19977 16627 20043 16630
rect 20253 16690 20319 16693
rect 20253 16688 20362 16690
rect 20253 16632 20258 16688
rect 20314 16632 20362 16688
rect 20253 16627 20362 16632
rect 7373 16554 7439 16557
rect 4846 16552 7439 16554
rect 4846 16496 7378 16552
rect 7434 16496 7439 16552
rect 4846 16494 7439 16496
rect 7373 16491 7439 16494
rect 7741 16554 7807 16557
rect 9622 16554 9628 16556
rect 7741 16552 9628 16554
rect 7741 16496 7746 16552
rect 7802 16496 9628 16552
rect 7741 16494 9628 16496
rect 7741 16491 7807 16494
rect 9622 16492 9628 16494
rect 9692 16492 9698 16556
rect 10358 16492 10364 16556
rect 10428 16554 10434 16556
rect 11053 16554 11119 16557
rect 10428 16552 11119 16554
rect 10428 16496 11058 16552
rect 11114 16496 11119 16552
rect 10428 16494 11119 16496
rect 10428 16492 10434 16494
rect 11053 16491 11119 16494
rect 11278 16492 11284 16556
rect 11348 16554 11354 16556
rect 11789 16554 11855 16557
rect 12525 16556 12591 16557
rect 12525 16554 12572 16556
rect 11348 16552 11855 16554
rect 11348 16496 11794 16552
rect 11850 16496 11855 16552
rect 11348 16494 11855 16496
rect 12480 16552 12572 16554
rect 12480 16496 12530 16552
rect 12480 16494 12572 16496
rect 11348 16492 11354 16494
rect 11789 16491 11855 16494
rect 12525 16492 12572 16494
rect 12636 16492 12642 16556
rect 15193 16554 15259 16557
rect 12712 16552 15259 16554
rect 12712 16496 15198 16552
rect 15254 16496 15259 16552
rect 12712 16494 15259 16496
rect 12525 16491 12591 16492
rect 3049 16416 3802 16418
rect 3049 16360 3054 16416
rect 3110 16360 3802 16416
rect 3049 16358 3802 16360
rect 5533 16418 5599 16421
rect 12014 16418 12020 16420
rect 5533 16416 12020 16418
rect 5533 16360 5538 16416
rect 5594 16360 12020 16416
rect 5533 16358 12020 16360
rect 0 16328 800 16358
rect 3049 16355 3115 16358
rect 5533 16355 5599 16358
rect 12014 16356 12020 16358
rect 12084 16356 12090 16420
rect 12433 16418 12499 16421
rect 12712 16418 12772 16494
rect 15193 16491 15259 16494
rect 15929 16554 15995 16557
rect 16062 16554 16068 16556
rect 15929 16552 16068 16554
rect 15929 16496 15934 16552
rect 15990 16496 16068 16552
rect 15929 16494 16068 16496
rect 15929 16491 15995 16494
rect 16062 16492 16068 16494
rect 16132 16492 16138 16556
rect 18965 16554 19031 16557
rect 20302 16554 20362 16627
rect 25262 16554 25268 16556
rect 18965 16552 25268 16554
rect 18965 16496 18970 16552
rect 19026 16496 25268 16552
rect 18965 16494 25268 16496
rect 18965 16491 19031 16494
rect 25262 16492 25268 16494
rect 25332 16554 25338 16556
rect 26550 16554 26556 16556
rect 25332 16494 26556 16554
rect 25332 16492 25338 16494
rect 26550 16492 26556 16494
rect 26620 16492 26626 16556
rect 12433 16416 12772 16418
rect 12433 16360 12438 16416
rect 12494 16360 12772 16416
rect 12433 16358 12772 16360
rect 15009 16418 15075 16421
rect 17033 16418 17099 16421
rect 18413 16418 18479 16421
rect 15009 16416 18479 16418
rect 15009 16360 15014 16416
rect 15070 16360 17038 16416
rect 17094 16360 18418 16416
rect 18474 16360 18479 16416
rect 15009 16358 18479 16360
rect 12433 16355 12499 16358
rect 15009 16355 15075 16358
rect 17033 16355 17099 16358
rect 18413 16355 18479 16358
rect 19558 16356 19564 16420
rect 19628 16418 19634 16420
rect 20805 16418 20871 16421
rect 19628 16416 20871 16418
rect 19628 16360 20810 16416
rect 20866 16360 20871 16416
rect 19628 16358 20871 16360
rect 19628 16356 19634 16358
rect 20805 16355 20871 16358
rect 24301 16420 24367 16421
rect 24301 16416 24348 16420
rect 24412 16418 24418 16420
rect 24301 16360 24306 16416
rect 24301 16356 24348 16360
rect 24412 16358 24458 16418
rect 24412 16356 24418 16358
rect 24301 16355 24367 16356
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 2037 16282 2103 16285
rect 2037 16280 2790 16282
rect 2037 16224 2042 16280
rect 2098 16224 2790 16280
rect 2037 16222 2790 16224
rect 2037 16219 2103 16222
rect 2730 16146 2790 16222
rect 7230 16220 7236 16284
rect 7300 16282 7306 16284
rect 11605 16282 11671 16285
rect 7300 16280 11671 16282
rect 7300 16224 11610 16280
rect 11666 16224 11671 16280
rect 7300 16222 11671 16224
rect 7300 16220 7306 16222
rect 11605 16219 11671 16222
rect 11881 16282 11947 16285
rect 23473 16282 23539 16285
rect 11881 16280 23539 16282
rect 11881 16224 11886 16280
rect 11942 16224 23478 16280
rect 23534 16224 23539 16280
rect 11881 16222 23539 16224
rect 11881 16219 11947 16222
rect 23473 16219 23539 16222
rect 6729 16146 6795 16149
rect 2730 16144 6795 16146
rect 2730 16088 6734 16144
rect 6790 16088 6795 16144
rect 2730 16086 6795 16088
rect 6729 16083 6795 16086
rect 7189 16146 7255 16149
rect 19701 16146 19767 16149
rect 7189 16144 19767 16146
rect 7189 16088 7194 16144
rect 7250 16088 19706 16144
rect 19762 16088 19767 16144
rect 7189 16086 19767 16088
rect 7189 16083 7255 16086
rect 19701 16083 19767 16086
rect 20713 16146 20779 16149
rect 27613 16146 27679 16149
rect 20713 16144 27679 16146
rect 20713 16088 20718 16144
rect 20774 16088 27618 16144
rect 27674 16088 27679 16144
rect 20713 16086 27679 16088
rect 20713 16083 20779 16086
rect 27613 16083 27679 16086
rect 2773 16010 2839 16013
rect 3233 16010 3299 16013
rect 7005 16010 7071 16013
rect 2773 16008 7071 16010
rect 2773 15952 2778 16008
rect 2834 15952 3238 16008
rect 3294 15952 7010 16008
rect 7066 15952 7071 16008
rect 2773 15950 7071 15952
rect 2773 15947 2839 15950
rect 3233 15947 3299 15950
rect 7005 15947 7071 15950
rect 8017 16010 8083 16013
rect 11513 16010 11579 16013
rect 11973 16010 12039 16013
rect 8017 16008 12039 16010
rect 8017 15952 8022 16008
rect 8078 15952 11518 16008
rect 11574 15952 11978 16008
rect 12034 15952 12039 16008
rect 8017 15950 12039 15952
rect 8017 15947 8083 15950
rect 11513 15947 11579 15950
rect 11973 15947 12039 15950
rect 13118 15948 13124 16012
rect 13188 16010 13194 16012
rect 16113 16010 16179 16013
rect 13188 16008 16179 16010
rect 13188 15952 16118 16008
rect 16174 15952 16179 16008
rect 13188 15950 16179 15952
rect 13188 15948 13194 15950
rect 16113 15947 16179 15950
rect 20713 16010 20779 16013
rect 21541 16010 21607 16013
rect 25497 16010 25563 16013
rect 20713 16008 25563 16010
rect 20713 15952 20718 16008
rect 20774 15952 21546 16008
rect 21602 15952 25502 16008
rect 25558 15952 25563 16008
rect 20713 15950 25563 15952
rect 20713 15947 20779 15950
rect 21541 15947 21607 15950
rect 25497 15947 25563 15950
rect 5165 15874 5231 15877
rect 5390 15874 5396 15876
rect 5165 15872 5396 15874
rect 5165 15816 5170 15872
rect 5226 15816 5396 15872
rect 5165 15814 5396 15816
rect 5165 15811 5231 15814
rect 5390 15812 5396 15814
rect 5460 15812 5466 15876
rect 10910 15874 10916 15876
rect 6502 15814 10916 15874
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 4654 15676 4660 15740
rect 4724 15738 4730 15740
rect 5625 15738 5691 15741
rect 4724 15736 5691 15738
rect 4724 15680 5630 15736
rect 5686 15680 5691 15736
rect 4724 15678 5691 15680
rect 4724 15676 4730 15678
rect 5625 15675 5691 15678
rect 3877 15604 3943 15605
rect 3877 15602 3924 15604
rect 3832 15600 3924 15602
rect 3832 15544 3882 15600
rect 3832 15542 3924 15544
rect 3877 15540 3924 15542
rect 3988 15540 3994 15604
rect 4429 15602 4495 15605
rect 6502 15602 6562 15814
rect 10910 15812 10916 15814
rect 10980 15812 10986 15876
rect 11145 15874 11211 15877
rect 23933 15874 23999 15877
rect 25221 15874 25287 15877
rect 11145 15872 25287 15874
rect 11145 15816 11150 15872
rect 11206 15816 23938 15872
rect 23994 15816 25226 15872
rect 25282 15816 25287 15872
rect 11145 15814 25287 15816
rect 11145 15811 11211 15814
rect 23933 15811 23999 15814
rect 25221 15811 25287 15814
rect 6729 15738 6795 15741
rect 6862 15738 6868 15740
rect 6729 15736 6868 15738
rect 6729 15680 6734 15736
rect 6790 15680 6868 15736
rect 6729 15678 6868 15680
rect 6729 15675 6795 15678
rect 6862 15676 6868 15678
rect 6932 15676 6938 15740
rect 9765 15738 9831 15741
rect 13486 15738 13492 15740
rect 9765 15736 13492 15738
rect 9765 15680 9770 15736
rect 9826 15680 13492 15736
rect 9765 15678 13492 15680
rect 9765 15675 9831 15678
rect 13486 15676 13492 15678
rect 13556 15676 13562 15740
rect 13997 15738 14063 15741
rect 15929 15738 15995 15741
rect 16757 15740 16823 15741
rect 16757 15738 16804 15740
rect 13997 15736 15995 15738
rect 13997 15680 14002 15736
rect 14058 15680 15934 15736
rect 15990 15680 15995 15736
rect 13997 15678 15995 15680
rect 16712 15736 16804 15738
rect 16712 15680 16762 15736
rect 16712 15678 16804 15680
rect 13997 15675 14063 15678
rect 15929 15675 15995 15678
rect 16757 15676 16804 15678
rect 16868 15676 16874 15740
rect 19701 15738 19767 15741
rect 20253 15738 20319 15741
rect 22001 15740 22067 15741
rect 21950 15738 21956 15740
rect 19701 15736 20319 15738
rect 19701 15680 19706 15736
rect 19762 15680 20258 15736
rect 20314 15680 20319 15736
rect 19701 15678 20319 15680
rect 21910 15678 21956 15738
rect 22020 15736 22067 15740
rect 22062 15680 22067 15736
rect 16757 15675 16823 15676
rect 19701 15675 19767 15678
rect 20253 15675 20319 15678
rect 21950 15676 21956 15678
rect 22020 15676 22067 15680
rect 22001 15675 22067 15676
rect 22921 15738 22987 15741
rect 27838 15738 27844 15740
rect 22921 15736 27844 15738
rect 22921 15680 22926 15736
rect 22982 15680 27844 15736
rect 22921 15678 27844 15680
rect 22921 15675 22987 15678
rect 27838 15676 27844 15678
rect 27908 15676 27914 15740
rect 32397 15738 32463 15741
rect 33200 15738 34000 15768
rect 32397 15736 34000 15738
rect 32397 15680 32402 15736
rect 32458 15680 34000 15736
rect 32397 15678 34000 15680
rect 32397 15675 32463 15678
rect 33200 15648 34000 15678
rect 4429 15600 6562 15602
rect 4429 15544 4434 15600
rect 4490 15544 6562 15600
rect 4429 15542 6562 15544
rect 6637 15602 6703 15605
rect 13118 15602 13124 15604
rect 6637 15600 13124 15602
rect 6637 15544 6642 15600
rect 6698 15544 13124 15600
rect 6637 15542 13124 15544
rect 3877 15539 3943 15540
rect 4429 15539 4495 15542
rect 6637 15539 6703 15542
rect 13118 15540 13124 15542
rect 13188 15540 13194 15604
rect 13261 15602 13327 15605
rect 15929 15602 15995 15605
rect 23657 15602 23723 15605
rect 13261 15600 15210 15602
rect 13261 15544 13266 15600
rect 13322 15544 15210 15600
rect 13261 15542 15210 15544
rect 13261 15539 13327 15542
rect 1117 15466 1183 15469
rect 3049 15466 3115 15469
rect 1117 15464 3115 15466
rect 1117 15408 1122 15464
rect 1178 15408 3054 15464
rect 3110 15408 3115 15464
rect 1117 15406 3115 15408
rect 1117 15403 1183 15406
rect 3049 15403 3115 15406
rect 3550 15404 3556 15468
rect 3620 15466 3626 15468
rect 8477 15466 8543 15469
rect 3620 15464 8543 15466
rect 3620 15408 8482 15464
rect 8538 15408 8543 15464
rect 3620 15406 8543 15408
rect 3620 15404 3626 15406
rect 8477 15403 8543 15406
rect 8661 15466 8727 15469
rect 13905 15466 13971 15469
rect 15009 15466 15075 15469
rect 8661 15464 15075 15466
rect 8661 15408 8666 15464
rect 8722 15408 13910 15464
rect 13966 15408 15014 15464
rect 15070 15408 15075 15464
rect 8661 15406 15075 15408
rect 15150 15466 15210 15542
rect 15929 15600 23723 15602
rect 15929 15544 15934 15600
rect 15990 15544 23662 15600
rect 23718 15544 23723 15600
rect 15929 15542 23723 15544
rect 15929 15539 15995 15542
rect 23657 15539 23723 15542
rect 16941 15466 17007 15469
rect 15150 15464 17007 15466
rect 15150 15408 16946 15464
rect 17002 15408 17007 15464
rect 15150 15406 17007 15408
rect 8661 15403 8727 15406
rect 13905 15403 13971 15406
rect 15009 15403 15075 15406
rect 16941 15403 17007 15406
rect 18086 15404 18092 15468
rect 18156 15466 18162 15468
rect 26969 15466 27035 15469
rect 18156 15464 27035 15466
rect 18156 15408 26974 15464
rect 27030 15408 27035 15464
rect 18156 15406 27035 15408
rect 18156 15404 18162 15406
rect 26969 15403 27035 15406
rect 28165 15466 28231 15469
rect 28390 15466 28396 15468
rect 28165 15464 28396 15466
rect 28165 15408 28170 15464
rect 28226 15408 28396 15464
rect 28165 15406 28396 15408
rect 28165 15403 28231 15406
rect 28390 15404 28396 15406
rect 28460 15404 28466 15468
rect 2497 15330 2563 15333
rect 4429 15330 4495 15333
rect 2497 15328 4495 15330
rect 2497 15272 2502 15328
rect 2558 15272 4434 15328
rect 4490 15272 4495 15328
rect 2497 15270 4495 15272
rect 2497 15267 2563 15270
rect 4429 15267 4495 15270
rect 5942 15268 5948 15332
rect 6012 15330 6018 15332
rect 6545 15330 6611 15333
rect 6012 15328 6611 15330
rect 6012 15272 6550 15328
rect 6606 15272 6611 15328
rect 6012 15270 6611 15272
rect 6012 15268 6018 15270
rect 6545 15267 6611 15270
rect 8661 15330 8727 15333
rect 9489 15330 9555 15333
rect 9949 15330 10015 15333
rect 8661 15328 9555 15330
rect 8661 15272 8666 15328
rect 8722 15272 9494 15328
rect 9550 15272 9555 15328
rect 8661 15270 9555 15272
rect 8661 15267 8727 15270
rect 9489 15267 9555 15270
rect 9630 15328 10015 15330
rect 9630 15272 9954 15328
rect 10010 15272 10015 15328
rect 9630 15270 10015 15272
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 3049 15194 3115 15197
rect 3182 15194 3188 15196
rect 3049 15192 3188 15194
rect 3049 15136 3054 15192
rect 3110 15136 3188 15192
rect 3049 15134 3188 15136
rect 3049 15131 3115 15134
rect 3182 15132 3188 15134
rect 3252 15132 3258 15196
rect 5901 15194 5967 15197
rect 9630 15194 9690 15270
rect 9949 15267 10015 15270
rect 10133 15330 10199 15333
rect 10593 15330 10659 15333
rect 11513 15330 11579 15333
rect 12249 15330 12315 15333
rect 10133 15328 10426 15330
rect 10133 15272 10138 15328
rect 10194 15272 10426 15328
rect 10133 15270 10426 15272
rect 10133 15267 10199 15270
rect 5901 15192 9690 15194
rect 5901 15136 5906 15192
rect 5962 15136 9690 15192
rect 5901 15134 9690 15136
rect 9857 15194 9923 15197
rect 9990 15194 9996 15196
rect 9857 15192 9996 15194
rect 9857 15136 9862 15192
rect 9918 15136 9996 15192
rect 9857 15134 9996 15136
rect 5901 15131 5967 15134
rect 9857 15131 9923 15134
rect 9990 15132 9996 15134
rect 10060 15132 10066 15196
rect 10366 15194 10426 15270
rect 10593 15328 12315 15330
rect 10593 15272 10598 15328
rect 10654 15272 11518 15328
rect 11574 15272 12254 15328
rect 12310 15272 12315 15328
rect 10593 15270 12315 15272
rect 10593 15267 10659 15270
rect 11513 15267 11579 15270
rect 12249 15267 12315 15270
rect 12801 15330 12867 15333
rect 20713 15330 20779 15333
rect 12801 15328 20779 15330
rect 12801 15272 12806 15328
rect 12862 15272 20718 15328
rect 20774 15272 20779 15328
rect 12801 15270 20779 15272
rect 12801 15267 12867 15270
rect 20713 15267 20779 15270
rect 22645 15330 22711 15333
rect 23422 15330 23428 15332
rect 22645 15328 23428 15330
rect 22645 15272 22650 15328
rect 22706 15272 23428 15328
rect 22645 15270 23428 15272
rect 22645 15267 22711 15270
rect 23422 15268 23428 15270
rect 23492 15268 23498 15332
rect 11237 15194 11303 15197
rect 10366 15192 11303 15194
rect 10366 15136 11242 15192
rect 11298 15136 11303 15192
rect 10366 15134 11303 15136
rect 11237 15131 11303 15134
rect 11830 15132 11836 15196
rect 11900 15194 11906 15196
rect 18873 15194 18939 15197
rect 11900 15192 18939 15194
rect 11900 15136 18878 15192
rect 18934 15136 18939 15192
rect 11900 15134 18939 15136
rect 11900 15132 11906 15134
rect 18873 15131 18939 15134
rect 19517 15196 19583 15197
rect 19517 15192 19564 15196
rect 19628 15194 19634 15196
rect 28993 15194 29059 15197
rect 29126 15194 29132 15196
rect 19517 15136 19522 15192
rect 19517 15132 19564 15136
rect 19628 15134 19674 15194
rect 28993 15192 29132 15194
rect 28993 15136 28998 15192
rect 29054 15136 29132 15192
rect 28993 15134 29132 15136
rect 19628 15132 19634 15134
rect 19517 15131 19583 15132
rect 28993 15131 29059 15134
rect 29126 15132 29132 15134
rect 29196 15132 29202 15196
rect 974 14996 980 15060
rect 1044 15058 1050 15060
rect 7005 15058 7071 15061
rect 1044 15056 7071 15058
rect 1044 15000 7010 15056
rect 7066 15000 7071 15056
rect 1044 14998 7071 15000
rect 1044 14996 1050 14998
rect 7005 14995 7071 14998
rect 7281 15058 7347 15061
rect 12198 15058 12204 15060
rect 7281 15056 12204 15058
rect 7281 15000 7286 15056
rect 7342 15000 12204 15056
rect 7281 14998 12204 15000
rect 7281 14995 7347 14998
rect 12198 14996 12204 14998
rect 12268 14996 12274 15060
rect 13629 15058 13695 15061
rect 14181 15058 14247 15061
rect 13629 15056 14247 15058
rect 13629 15000 13634 15056
rect 13690 15000 14186 15056
rect 14242 15000 14247 15056
rect 13629 14998 14247 15000
rect 13629 14995 13695 14998
rect 14181 14995 14247 14998
rect 15193 15058 15259 15061
rect 17585 15058 17651 15061
rect 15193 15056 17651 15058
rect 15193 15000 15198 15056
rect 15254 15000 17590 15056
rect 17646 15000 17651 15056
rect 15193 14998 17651 15000
rect 15193 14995 15259 14998
rect 17585 14995 17651 14998
rect 17718 14996 17724 15060
rect 17788 15058 17794 15060
rect 17861 15058 17927 15061
rect 17788 15056 17927 15058
rect 17788 15000 17866 15056
rect 17922 15000 17927 15056
rect 17788 14998 17927 15000
rect 17788 14996 17794 14998
rect 17861 14995 17927 14998
rect 19609 15058 19675 15061
rect 20069 15058 20135 15061
rect 20621 15058 20687 15061
rect 19609 15056 20687 15058
rect 19609 15000 19614 15056
rect 19670 15000 20074 15056
rect 20130 15000 20626 15056
rect 20682 15000 20687 15056
rect 19609 14998 20687 15000
rect 19609 14995 19675 14998
rect 20069 14995 20135 14998
rect 20621 14995 20687 14998
rect 21214 14996 21220 15060
rect 21284 15058 21290 15060
rect 27613 15058 27679 15061
rect 31017 15060 31083 15061
rect 21284 15056 27679 15058
rect 21284 15000 27618 15056
rect 27674 15000 27679 15056
rect 21284 14998 27679 15000
rect 21284 14996 21290 14998
rect 27613 14995 27679 14998
rect 30966 14996 30972 15060
rect 31036 15058 31083 15060
rect 32397 15058 32463 15061
rect 33200 15058 34000 15088
rect 31036 15056 31128 15058
rect 31078 15000 31128 15056
rect 31036 14998 31128 15000
rect 32397 15056 34000 15058
rect 32397 15000 32402 15056
rect 32458 15000 34000 15056
rect 32397 14998 34000 15000
rect 31036 14996 31083 14998
rect 31017 14995 31083 14996
rect 32397 14995 32463 14998
rect 33200 14968 34000 14998
rect 5441 14922 5507 14925
rect 5574 14922 5580 14924
rect 5441 14920 5580 14922
rect 5441 14864 5446 14920
rect 5502 14864 5580 14920
rect 5441 14862 5580 14864
rect 5441 14859 5507 14862
rect 5574 14860 5580 14862
rect 5644 14860 5650 14924
rect 5717 14922 5783 14925
rect 8702 14922 8708 14924
rect 5717 14920 8708 14922
rect 5717 14864 5722 14920
rect 5778 14864 8708 14920
rect 5717 14862 8708 14864
rect 5717 14859 5783 14862
rect 8702 14860 8708 14862
rect 8772 14922 8778 14924
rect 12249 14922 12315 14925
rect 12382 14922 12388 14924
rect 8772 14862 11898 14922
rect 8772 14860 8778 14862
rect 4889 14786 4955 14789
rect 7465 14786 7531 14789
rect 4889 14784 7531 14786
rect 4889 14728 4894 14784
rect 4950 14728 7470 14784
rect 7526 14728 7531 14784
rect 4889 14726 7531 14728
rect 4889 14723 4955 14726
rect 7465 14723 7531 14726
rect 8661 14786 8727 14789
rect 9254 14786 9260 14788
rect 8661 14784 9260 14786
rect 8661 14728 8666 14784
rect 8722 14728 9260 14784
rect 8661 14726 9260 14728
rect 8661 14723 8727 14726
rect 9254 14724 9260 14726
rect 9324 14724 9330 14788
rect 9489 14786 9555 14789
rect 11053 14786 11119 14789
rect 9489 14784 11119 14786
rect 9489 14728 9494 14784
rect 9550 14728 11058 14784
rect 11114 14728 11119 14784
rect 9489 14726 11119 14728
rect 11838 14786 11898 14862
rect 12249 14920 12388 14922
rect 12249 14864 12254 14920
rect 12310 14864 12388 14920
rect 12249 14862 12388 14864
rect 12249 14859 12315 14862
rect 12382 14860 12388 14862
rect 12452 14922 12458 14924
rect 16757 14922 16823 14925
rect 12452 14920 16823 14922
rect 12452 14864 16762 14920
rect 16818 14864 16823 14920
rect 12452 14862 16823 14864
rect 12452 14860 12458 14862
rect 16757 14859 16823 14862
rect 18781 14922 18847 14925
rect 24945 14922 25011 14925
rect 18781 14920 25011 14922
rect 18781 14864 18786 14920
rect 18842 14864 24950 14920
rect 25006 14864 25011 14920
rect 18781 14862 25011 14864
rect 18781 14859 18847 14862
rect 24945 14859 25011 14862
rect 12709 14786 12775 14789
rect 13670 14786 13676 14788
rect 11838 14726 12450 14786
rect 9489 14723 9555 14726
rect 11053 14723 11119 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 4705 14650 4771 14653
rect 7189 14650 7255 14653
rect 4705 14648 7255 14650
rect 4705 14592 4710 14648
rect 4766 14592 7194 14648
rect 7250 14592 7255 14648
rect 4705 14590 7255 14592
rect 4705 14587 4771 14590
rect 7189 14587 7255 14590
rect 7925 14650 7991 14653
rect 9489 14652 9555 14653
rect 8518 14650 8524 14652
rect 7925 14648 8524 14650
rect 7925 14592 7930 14648
rect 7986 14592 8524 14648
rect 7925 14590 8524 14592
rect 7925 14587 7991 14590
rect 8518 14588 8524 14590
rect 8588 14588 8594 14652
rect 9438 14588 9444 14652
rect 9508 14650 9555 14652
rect 9857 14650 9923 14653
rect 12249 14650 12315 14653
rect 9508 14648 9600 14650
rect 9550 14592 9600 14648
rect 9508 14590 9600 14592
rect 9857 14648 12315 14650
rect 9857 14592 9862 14648
rect 9918 14592 12254 14648
rect 12310 14592 12315 14648
rect 9857 14590 12315 14592
rect 12390 14650 12450 14726
rect 12709 14784 13676 14786
rect 12709 14728 12714 14784
rect 12770 14728 13676 14784
rect 12709 14726 13676 14728
rect 12709 14723 12775 14726
rect 13670 14724 13676 14726
rect 13740 14724 13746 14788
rect 14273 14786 14339 14789
rect 15285 14786 15351 14789
rect 14273 14784 15351 14786
rect 14273 14728 14278 14784
rect 14334 14728 15290 14784
rect 15346 14728 15351 14784
rect 14273 14726 15351 14728
rect 14273 14723 14339 14726
rect 15285 14723 15351 14726
rect 16757 14786 16823 14789
rect 25589 14786 25655 14789
rect 16757 14784 25655 14786
rect 16757 14728 16762 14784
rect 16818 14728 25594 14784
rect 25650 14728 25655 14784
rect 16757 14726 25655 14728
rect 16757 14723 16823 14726
rect 25589 14723 25655 14726
rect 30833 14786 30899 14789
rect 30966 14786 30972 14788
rect 30833 14784 30972 14786
rect 30833 14728 30838 14784
rect 30894 14728 30972 14784
rect 30833 14726 30972 14728
rect 30833 14723 30899 14726
rect 30966 14724 30972 14726
rect 31036 14724 31042 14788
rect 13813 14650 13879 14653
rect 12390 14648 13879 14650
rect 12390 14592 13818 14648
rect 13874 14592 13879 14648
rect 12390 14590 13879 14592
rect 9508 14588 9555 14590
rect 9489 14587 9555 14588
rect 9857 14587 9923 14590
rect 12249 14587 12315 14590
rect 13813 14587 13879 14590
rect 14273 14650 14339 14653
rect 17677 14650 17743 14653
rect 14273 14648 17743 14650
rect 14273 14592 14278 14648
rect 14334 14592 17682 14648
rect 17738 14592 17743 14648
rect 14273 14590 17743 14592
rect 14273 14587 14339 14590
rect 17677 14587 17743 14590
rect 18597 14650 18663 14653
rect 18781 14650 18847 14653
rect 19149 14650 19215 14653
rect 18597 14648 18706 14650
rect 18597 14592 18602 14648
rect 18658 14592 18706 14648
rect 18597 14587 18706 14592
rect 18781 14648 20730 14650
rect 18781 14592 18786 14648
rect 18842 14592 19154 14648
rect 19210 14592 20730 14648
rect 18781 14590 20730 14592
rect 18781 14587 18847 14590
rect 19149 14587 19215 14590
rect 841 14514 907 14517
rect 798 14512 907 14514
rect 798 14456 846 14512
rect 902 14456 907 14512
rect 798 14451 907 14456
rect 3550 14452 3556 14516
rect 3620 14514 3626 14516
rect 3877 14514 3943 14517
rect 3620 14512 3943 14514
rect 3620 14456 3882 14512
rect 3938 14456 3943 14512
rect 3620 14454 3943 14456
rect 3620 14452 3626 14454
rect 3877 14451 3943 14454
rect 5625 14514 5691 14517
rect 6821 14514 6887 14517
rect 5625 14512 6887 14514
rect 5625 14456 5630 14512
rect 5686 14456 6826 14512
rect 6882 14456 6887 14512
rect 5625 14454 6887 14456
rect 5625 14451 5691 14454
rect 6821 14451 6887 14454
rect 7046 14452 7052 14516
rect 7116 14514 7122 14516
rect 7928 14514 7988 14587
rect 7116 14454 7988 14514
rect 8569 14514 8635 14517
rect 15101 14514 15167 14517
rect 8569 14512 15167 14514
rect 8569 14456 8574 14512
rect 8630 14456 15106 14512
rect 15162 14456 15167 14512
rect 8569 14454 15167 14456
rect 18646 14514 18706 14587
rect 18873 14514 18939 14517
rect 18646 14512 18939 14514
rect 18646 14456 18878 14512
rect 18934 14456 18939 14512
rect 18646 14454 18939 14456
rect 7116 14452 7122 14454
rect 8569 14451 8635 14454
rect 15101 14451 15167 14454
rect 18873 14451 18939 14454
rect 19190 14452 19196 14516
rect 19260 14514 19266 14516
rect 19517 14514 19583 14517
rect 19260 14512 19583 14514
rect 19260 14456 19522 14512
rect 19578 14456 19583 14512
rect 19260 14454 19583 14456
rect 19260 14452 19266 14454
rect 19517 14451 19583 14454
rect 20345 14514 20411 14517
rect 20478 14514 20484 14516
rect 20345 14512 20484 14514
rect 20345 14456 20350 14512
rect 20406 14456 20484 14512
rect 20345 14454 20484 14456
rect 20345 14451 20411 14454
rect 20478 14452 20484 14454
rect 20548 14452 20554 14516
rect 20670 14514 20730 14590
rect 21030 14588 21036 14652
rect 21100 14650 21106 14652
rect 22369 14650 22435 14653
rect 21100 14648 22435 14650
rect 21100 14592 22374 14648
rect 22430 14592 22435 14648
rect 21100 14590 22435 14592
rect 21100 14588 21106 14590
rect 22369 14587 22435 14590
rect 23606 14514 23612 14516
rect 20670 14454 23612 14514
rect 23606 14452 23612 14454
rect 23676 14452 23682 14516
rect 23974 14452 23980 14516
rect 24044 14514 24050 14516
rect 24301 14514 24367 14517
rect 24044 14512 24367 14514
rect 24044 14456 24306 14512
rect 24362 14456 24367 14512
rect 24044 14454 24367 14456
rect 24044 14452 24050 14454
rect 24301 14451 24367 14454
rect 798 14408 858 14451
rect 0 14318 858 14408
rect 0 14288 800 14318
rect 3550 14316 3556 14380
rect 3620 14378 3626 14380
rect 3785 14378 3851 14381
rect 3620 14376 3851 14378
rect 3620 14320 3790 14376
rect 3846 14320 3851 14376
rect 3620 14318 3851 14320
rect 3620 14316 3626 14318
rect 3785 14315 3851 14318
rect 4245 14378 4311 14381
rect 5717 14380 5783 14381
rect 5717 14378 5764 14380
rect 4245 14376 5320 14378
rect 4245 14320 4250 14376
rect 4306 14320 5320 14376
rect 4245 14318 5320 14320
rect 5672 14376 5764 14378
rect 5672 14320 5722 14376
rect 5672 14318 5764 14320
rect 4245 14315 4311 14318
rect 5260 14242 5320 14318
rect 5717 14316 5764 14318
rect 5828 14316 5834 14380
rect 8886 14316 8892 14380
rect 8956 14378 8962 14380
rect 10133 14378 10199 14381
rect 8956 14376 10199 14378
rect 8956 14320 10138 14376
rect 10194 14320 10199 14376
rect 8956 14318 10199 14320
rect 8956 14316 8962 14318
rect 5717 14315 5783 14316
rect 10133 14315 10199 14318
rect 10409 14378 10475 14381
rect 23657 14378 23723 14381
rect 24485 14380 24551 14381
rect 24485 14378 24532 14380
rect 10409 14376 23723 14378
rect 10409 14320 10414 14376
rect 10470 14320 23662 14376
rect 23718 14320 23723 14376
rect 10409 14318 23723 14320
rect 24440 14376 24532 14378
rect 24440 14320 24490 14376
rect 24440 14318 24532 14320
rect 10409 14315 10475 14318
rect 23657 14315 23723 14318
rect 24485 14316 24532 14318
rect 24596 14316 24602 14380
rect 26366 14316 26372 14380
rect 26436 14378 26442 14380
rect 27705 14378 27771 14381
rect 26436 14376 27771 14378
rect 26436 14320 27710 14376
rect 27766 14320 27771 14376
rect 26436 14318 27771 14320
rect 26436 14316 26442 14318
rect 24485 14315 24551 14316
rect 9857 14242 9923 14245
rect 11830 14242 11836 14244
rect 5260 14240 9923 14242
rect 5260 14184 9862 14240
rect 9918 14184 9923 14240
rect 5260 14182 9923 14184
rect 9857 14179 9923 14182
rect 9998 14182 11836 14242
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 657 14106 723 14109
rect 5717 14106 5783 14109
rect 7373 14108 7439 14109
rect 7373 14106 7420 14108
rect 657 14104 2790 14106
rect 657 14048 662 14104
rect 718 14048 2790 14104
rect 657 14046 2790 14048
rect 657 14043 723 14046
rect 2730 13970 2790 14046
rect 5717 14104 7420 14106
rect 5717 14048 5722 14104
rect 5778 14048 7378 14104
rect 5717 14046 7420 14048
rect 5717 14043 5783 14046
rect 7373 14044 7420 14046
rect 7484 14044 7490 14108
rect 7649 14106 7715 14109
rect 9998 14106 10058 14182
rect 11830 14180 11836 14182
rect 11900 14180 11906 14244
rect 12198 14180 12204 14244
rect 12268 14242 12274 14244
rect 12617 14242 12683 14245
rect 12268 14240 12683 14242
rect 12268 14184 12622 14240
rect 12678 14184 12683 14240
rect 12268 14182 12683 14184
rect 12268 14180 12274 14182
rect 12617 14179 12683 14182
rect 13721 14242 13787 14245
rect 20437 14242 20503 14245
rect 13721 14240 20503 14242
rect 13721 14184 13726 14240
rect 13782 14184 20442 14240
rect 20498 14184 20503 14240
rect 13721 14182 20503 14184
rect 13721 14179 13787 14182
rect 20437 14179 20503 14182
rect 21449 14242 21515 14245
rect 22277 14242 22343 14245
rect 21449 14240 22343 14242
rect 21449 14184 21454 14240
rect 21510 14184 22282 14240
rect 22338 14184 22343 14240
rect 21449 14182 22343 14184
rect 21449 14179 21515 14182
rect 22277 14179 22343 14182
rect 7649 14104 10058 14106
rect 7649 14048 7654 14104
rect 7710 14048 10058 14104
rect 7649 14046 10058 14048
rect 7373 14043 7439 14044
rect 7649 14043 7715 14046
rect 10358 14044 10364 14108
rect 10428 14106 10434 14108
rect 10593 14106 10659 14109
rect 10428 14104 10659 14106
rect 10428 14048 10598 14104
rect 10654 14048 10659 14104
rect 10428 14046 10659 14048
rect 10428 14044 10434 14046
rect 10593 14043 10659 14046
rect 10869 14106 10935 14109
rect 11513 14106 11579 14109
rect 10869 14104 11579 14106
rect 10869 14048 10874 14104
rect 10930 14048 11518 14104
rect 11574 14048 11579 14104
rect 10869 14046 11579 14048
rect 10869 14043 10935 14046
rect 11513 14043 11579 14046
rect 11697 14106 11763 14109
rect 12934 14106 12940 14108
rect 11697 14104 12940 14106
rect 11697 14048 11702 14104
rect 11758 14048 12940 14104
rect 11697 14046 12940 14048
rect 11697 14043 11763 14046
rect 12934 14044 12940 14046
rect 13004 14044 13010 14108
rect 17217 14106 17283 14109
rect 13080 14104 17283 14106
rect 13080 14048 17222 14104
rect 17278 14048 17283 14104
rect 13080 14046 17283 14048
rect 7741 13970 7807 13973
rect 11973 13970 12039 13973
rect 12433 13972 12499 13973
rect 12382 13970 12388 13972
rect 2730 13968 12039 13970
rect 2730 13912 7746 13968
rect 7802 13912 11978 13968
rect 12034 13912 12039 13968
rect 2730 13910 12039 13912
rect 12342 13910 12388 13970
rect 12452 13968 12499 13972
rect 12494 13912 12499 13968
rect 7741 13907 7807 13910
rect 11973 13907 12039 13910
rect 12382 13908 12388 13910
rect 12452 13908 12499 13912
rect 12433 13907 12499 13908
rect 12801 13970 12867 13973
rect 13080 13970 13140 14046
rect 17217 14043 17283 14046
rect 17350 14044 17356 14108
rect 17420 14106 17426 14108
rect 20846 14106 20852 14108
rect 17420 14046 20852 14106
rect 17420 14044 17426 14046
rect 20846 14044 20852 14046
rect 20916 14044 20922 14108
rect 21398 14044 21404 14108
rect 21468 14106 21474 14108
rect 26374 14106 26434 14316
rect 27705 14315 27771 14318
rect 21468 14046 26434 14106
rect 21468 14044 21474 14046
rect 12801 13968 13140 13970
rect 12801 13912 12806 13968
rect 12862 13912 13140 13968
rect 12801 13910 13140 13912
rect 13261 13970 13327 13973
rect 14641 13970 14707 13973
rect 13261 13968 14707 13970
rect 13261 13912 13266 13968
rect 13322 13912 14646 13968
rect 14702 13912 14707 13968
rect 13261 13910 14707 13912
rect 12801 13907 12867 13910
rect 13261 13907 13327 13910
rect 14641 13907 14707 13910
rect 14825 13970 14891 13973
rect 17953 13970 18019 13973
rect 18781 13970 18847 13973
rect 14825 13968 18847 13970
rect 14825 13912 14830 13968
rect 14886 13912 17958 13968
rect 18014 13912 18786 13968
rect 18842 13912 18847 13968
rect 14825 13910 18847 13912
rect 14825 13907 14891 13910
rect 17953 13907 18019 13910
rect 18781 13907 18847 13910
rect 19885 13970 19951 13973
rect 20345 13970 20411 13973
rect 19885 13968 20411 13970
rect 19885 13912 19890 13968
rect 19946 13912 20350 13968
rect 20406 13912 20411 13968
rect 19885 13910 20411 13912
rect 19885 13907 19951 13910
rect 20345 13907 20411 13910
rect 22921 13970 22987 13973
rect 28206 13970 28212 13972
rect 22921 13968 28212 13970
rect 22921 13912 22926 13968
rect 22982 13912 28212 13968
rect 22921 13910 28212 13912
rect 22921 13907 22987 13910
rect 28206 13908 28212 13910
rect 28276 13908 28282 13972
rect 3049 13834 3115 13837
rect 4889 13834 4955 13837
rect 5349 13834 5415 13837
rect 7649 13834 7715 13837
rect 3049 13832 4768 13834
rect 3049 13776 3054 13832
rect 3110 13776 4768 13832
rect 3049 13774 4768 13776
rect 3049 13771 3115 13774
rect 4708 13698 4768 13774
rect 4889 13832 7715 13834
rect 4889 13776 4894 13832
rect 4950 13776 5354 13832
rect 5410 13776 7654 13832
rect 7710 13776 7715 13832
rect 4889 13774 7715 13776
rect 4889 13771 4955 13774
rect 5349 13771 5415 13774
rect 7649 13771 7715 13774
rect 8886 13772 8892 13836
rect 8956 13834 8962 13836
rect 9305 13834 9371 13837
rect 9489 13836 9555 13837
rect 8956 13832 9371 13834
rect 8956 13776 9310 13832
rect 9366 13776 9371 13832
rect 8956 13774 9371 13776
rect 8956 13772 8962 13774
rect 9305 13771 9371 13774
rect 9438 13772 9444 13836
rect 9508 13834 9555 13836
rect 9857 13834 9923 13837
rect 10542 13834 10548 13836
rect 9508 13832 9600 13834
rect 9550 13776 9600 13832
rect 9508 13774 9600 13776
rect 9857 13832 10548 13834
rect 9857 13776 9862 13832
rect 9918 13776 10548 13832
rect 9857 13774 10548 13776
rect 9508 13772 9555 13774
rect 9489 13771 9555 13772
rect 9857 13771 9923 13774
rect 10542 13772 10548 13774
rect 10612 13772 10618 13836
rect 10869 13834 10935 13837
rect 11094 13834 11100 13836
rect 10869 13832 11100 13834
rect 10869 13776 10874 13832
rect 10930 13776 11100 13832
rect 10869 13774 11100 13776
rect 10869 13771 10935 13774
rect 11094 13772 11100 13774
rect 11164 13772 11170 13836
rect 11237 13834 11303 13837
rect 11973 13834 12039 13837
rect 12157 13836 12223 13837
rect 12157 13834 12204 13836
rect 11237 13832 12039 13834
rect 11237 13776 11242 13832
rect 11298 13776 11978 13832
rect 12034 13776 12039 13832
rect 11237 13774 12039 13776
rect 12112 13832 12204 13834
rect 12112 13776 12162 13832
rect 12112 13774 12204 13776
rect 11237 13771 11303 13774
rect 11973 13771 12039 13774
rect 12157 13772 12204 13774
rect 12268 13772 12274 13836
rect 21449 13834 21515 13837
rect 12390 13832 21515 13834
rect 12390 13776 21454 13832
rect 21510 13776 21515 13832
rect 12390 13774 21515 13776
rect 12157 13771 12223 13772
rect 9305 13698 9371 13701
rect 4708 13696 9371 13698
rect 4708 13640 9310 13696
rect 9366 13640 9371 13696
rect 4708 13638 9371 13640
rect 9305 13635 9371 13638
rect 9581 13698 9647 13701
rect 12390 13698 12450 13774
rect 21449 13771 21515 13774
rect 23238 13772 23244 13836
rect 23308 13834 23314 13836
rect 23381 13834 23447 13837
rect 23308 13832 23447 13834
rect 23308 13776 23386 13832
rect 23442 13776 23447 13832
rect 23308 13774 23447 13776
rect 23308 13772 23314 13774
rect 23381 13771 23447 13774
rect 23606 13772 23612 13836
rect 23676 13834 23682 13836
rect 23933 13834 23999 13837
rect 26509 13836 26575 13837
rect 26509 13834 26556 13836
rect 23676 13832 23999 13834
rect 23676 13776 23938 13832
rect 23994 13776 23999 13832
rect 23676 13774 23999 13776
rect 26464 13832 26556 13834
rect 26464 13776 26514 13832
rect 26464 13774 26556 13776
rect 23676 13772 23682 13774
rect 23933 13771 23999 13774
rect 26509 13772 26556 13774
rect 26620 13772 26626 13836
rect 26785 13834 26851 13837
rect 27429 13834 27495 13837
rect 26785 13832 27495 13834
rect 26785 13776 26790 13832
rect 26846 13776 27434 13832
rect 27490 13776 27495 13832
rect 26785 13774 27495 13776
rect 26509 13771 26575 13772
rect 26785 13771 26851 13774
rect 27429 13771 27495 13774
rect 9581 13696 12450 13698
rect 9581 13640 9586 13696
rect 9642 13640 12450 13696
rect 9581 13638 12450 13640
rect 9581 13635 9647 13638
rect 14774 13636 14780 13700
rect 14844 13698 14850 13700
rect 16614 13698 16620 13700
rect 14844 13638 16620 13698
rect 14844 13636 14850 13638
rect 16614 13636 16620 13638
rect 16684 13636 16690 13700
rect 17953 13698 18019 13701
rect 18086 13698 18092 13700
rect 17953 13696 18092 13698
rect 17953 13640 17958 13696
rect 18014 13640 18092 13696
rect 17953 13638 18092 13640
rect 17953 13635 18019 13638
rect 18086 13636 18092 13638
rect 18156 13636 18162 13700
rect 19333 13698 19399 13701
rect 20805 13698 20871 13701
rect 19333 13696 20871 13698
rect 19333 13640 19338 13696
rect 19394 13640 20810 13696
rect 20866 13640 20871 13696
rect 19333 13638 20871 13640
rect 19333 13635 19399 13638
rect 20805 13635 20871 13638
rect 21030 13636 21036 13700
rect 21100 13698 21106 13700
rect 21541 13698 21607 13701
rect 21100 13696 21607 13698
rect 21100 13640 21546 13696
rect 21602 13640 21607 13696
rect 21100 13638 21607 13640
rect 21100 13636 21106 13638
rect 21541 13635 21607 13638
rect 22369 13698 22435 13701
rect 22686 13698 22692 13700
rect 22369 13696 22692 13698
rect 22369 13640 22374 13696
rect 22430 13640 22692 13696
rect 22369 13638 22692 13640
rect 22369 13635 22435 13638
rect 22686 13636 22692 13638
rect 22756 13636 22762 13700
rect 23790 13636 23796 13700
rect 23860 13698 23866 13700
rect 23933 13698 23999 13701
rect 23860 13696 23999 13698
rect 23860 13640 23938 13696
rect 23994 13640 23999 13696
rect 23860 13638 23999 13640
rect 23860 13636 23866 13638
rect 23933 13635 23999 13638
rect 24117 13698 24183 13701
rect 27981 13698 28047 13701
rect 24117 13696 28047 13698
rect 24117 13640 24122 13696
rect 24178 13640 27986 13696
rect 28042 13640 28047 13696
rect 24117 13638 28047 13640
rect 24117 13635 24183 13638
rect 27981 13635 28047 13638
rect 32397 13698 32463 13701
rect 33200 13698 34000 13728
rect 32397 13696 34000 13698
rect 32397 13640 32402 13696
rect 32458 13640 34000 13696
rect 32397 13638 34000 13640
rect 32397 13635 32463 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 33200 13608 34000 13638
rect 4210 13567 4526 13568
rect 4797 13562 4863 13565
rect 8334 13562 8340 13564
rect 4797 13560 8340 13562
rect 4797 13504 4802 13560
rect 4858 13504 8340 13560
rect 4797 13502 8340 13504
rect 4797 13499 4863 13502
rect 8334 13500 8340 13502
rect 8404 13562 8410 13564
rect 26233 13562 26299 13565
rect 29310 13562 29316 13564
rect 8404 13560 26299 13562
rect 8404 13504 26238 13560
rect 26294 13504 26299 13560
rect 8404 13502 26299 13504
rect 8404 13500 8410 13502
rect 26233 13499 26299 13502
rect 28950 13502 29316 13562
rect 2313 13426 2379 13429
rect 4429 13426 4495 13429
rect 6862 13426 6868 13428
rect 2313 13424 4495 13426
rect 2313 13368 2318 13424
rect 2374 13368 4434 13424
rect 4490 13368 4495 13424
rect 2313 13366 4495 13368
rect 2313 13363 2379 13366
rect 4429 13363 4495 13366
rect 4662 13366 6868 13426
rect 3141 13290 3207 13293
rect 4337 13290 4403 13293
rect 3141 13288 4403 13290
rect 3141 13232 3146 13288
rect 3202 13232 4342 13288
rect 4398 13232 4403 13288
rect 3141 13230 4403 13232
rect 3141 13227 3207 13230
rect 4337 13227 4403 13230
rect 3141 13154 3207 13157
rect 4662 13154 4722 13366
rect 6862 13364 6868 13366
rect 6932 13364 6938 13428
rect 7281 13426 7347 13429
rect 17350 13426 17356 13428
rect 7281 13424 17356 13426
rect 7281 13368 7286 13424
rect 7342 13368 17356 13424
rect 7281 13366 17356 13368
rect 7281 13363 7347 13366
rect 17350 13364 17356 13366
rect 17420 13364 17426 13428
rect 17585 13426 17651 13429
rect 19793 13426 19859 13429
rect 24485 13426 24551 13429
rect 17585 13424 24551 13426
rect 17585 13368 17590 13424
rect 17646 13368 19798 13424
rect 19854 13368 24490 13424
rect 24546 13368 24551 13424
rect 17585 13366 24551 13368
rect 17585 13363 17651 13366
rect 19793 13363 19859 13366
rect 24485 13363 24551 13366
rect 4889 13290 4955 13293
rect 12985 13290 13051 13293
rect 20110 13290 20116 13292
rect 4889 13288 12450 13290
rect 4889 13232 4894 13288
rect 4950 13232 12450 13288
rect 4889 13230 12450 13232
rect 4889 13227 4955 13230
rect 3141 13152 4722 13154
rect 3141 13096 3146 13152
rect 3202 13096 4722 13152
rect 3141 13094 4722 13096
rect 5533 13154 5599 13157
rect 6126 13154 6132 13156
rect 5533 13152 6132 13154
rect 5533 13096 5538 13152
rect 5594 13096 6132 13152
rect 5533 13094 6132 13096
rect 3141 13091 3207 13094
rect 5533 13091 5599 13094
rect 6126 13092 6132 13094
rect 6196 13092 6202 13156
rect 6310 13092 6316 13156
rect 6380 13154 6386 13156
rect 6729 13154 6795 13157
rect 6380 13152 6795 13154
rect 6380 13096 6734 13152
rect 6790 13096 6795 13152
rect 6380 13094 6795 13096
rect 6380 13092 6386 13094
rect 6729 13091 6795 13094
rect 7189 13156 7255 13157
rect 7189 13152 7236 13156
rect 7300 13154 7306 13156
rect 8937 13154 9003 13157
rect 9070 13154 9076 13156
rect 7189 13096 7194 13152
rect 7189 13092 7236 13096
rect 7300 13094 7346 13154
rect 8937 13152 9076 13154
rect 8937 13096 8942 13152
rect 8998 13096 9076 13152
rect 8937 13094 9076 13096
rect 7300 13092 7306 13094
rect 7189 13091 7255 13092
rect 8937 13091 9003 13094
rect 9070 13092 9076 13094
rect 9140 13092 9146 13156
rect 9305 13154 9371 13157
rect 9489 13154 9555 13157
rect 12390 13154 12450 13230
rect 12985 13288 20116 13290
rect 12985 13232 12990 13288
rect 13046 13232 20116 13288
rect 12985 13230 20116 13232
rect 12985 13227 13051 13230
rect 20110 13228 20116 13230
rect 20180 13228 20186 13292
rect 20294 13228 20300 13292
rect 20364 13290 20370 13292
rect 21725 13290 21791 13293
rect 20364 13288 21791 13290
rect 20364 13232 21730 13288
rect 21786 13232 21791 13288
rect 20364 13230 21791 13232
rect 20364 13228 20370 13230
rect 21725 13227 21791 13230
rect 21950 13228 21956 13292
rect 22020 13290 22026 13292
rect 22093 13290 22159 13293
rect 22645 13292 22711 13293
rect 22645 13290 22692 13292
rect 22020 13288 22159 13290
rect 22020 13232 22098 13288
rect 22154 13232 22159 13288
rect 22020 13230 22159 13232
rect 22600 13288 22692 13290
rect 22600 13232 22650 13288
rect 22600 13230 22692 13232
rect 22020 13228 22026 13230
rect 22093 13227 22159 13230
rect 22645 13228 22692 13230
rect 22756 13228 22762 13292
rect 23054 13228 23060 13292
rect 23124 13290 23130 13292
rect 23289 13290 23355 13293
rect 23124 13288 23355 13290
rect 23124 13232 23294 13288
rect 23350 13232 23355 13288
rect 23124 13230 23355 13232
rect 23124 13228 23130 13230
rect 22645 13227 22711 13228
rect 23289 13227 23355 13230
rect 24117 13290 24183 13293
rect 28950 13290 29010 13502
rect 29310 13500 29316 13502
rect 29380 13500 29386 13564
rect 24117 13288 29010 13290
rect 24117 13232 24122 13288
rect 24178 13232 29010 13288
rect 24117 13230 29010 13232
rect 24117 13227 24183 13230
rect 13813 13154 13879 13157
rect 9305 13152 11898 13154
rect 9305 13096 9310 13152
rect 9366 13096 9494 13152
rect 9550 13096 11898 13152
rect 9305 13094 11898 13096
rect 12390 13152 13879 13154
rect 12390 13096 13818 13152
rect 13874 13096 13879 13152
rect 12390 13094 13879 13096
rect 9305 13091 9371 13094
rect 9489 13091 9555 13094
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 3785 13018 3851 13021
rect 4705 13020 4771 13021
rect 3918 13018 3924 13020
rect 3785 13016 3924 13018
rect 3785 12960 3790 13016
rect 3846 12960 3924 13016
rect 3785 12958 3924 12960
rect 3785 12955 3851 12958
rect 3918 12956 3924 12958
rect 3988 12956 3994 13020
rect 4654 13018 4660 13020
rect 4614 12958 4660 13018
rect 4724 13016 4771 13020
rect 11697 13018 11763 13021
rect 4766 12960 4771 13016
rect 4654 12956 4660 12958
rect 4724 12956 4771 12960
rect 4705 12955 4771 12956
rect 5950 13016 11763 13018
rect 5950 12960 11702 13016
rect 11758 12960 11763 13016
rect 5950 12958 11763 12960
rect 3601 12882 3667 12885
rect 5950 12882 6010 12958
rect 11697 12955 11763 12958
rect 3601 12880 6010 12882
rect 3601 12824 3606 12880
rect 3662 12824 6010 12880
rect 3601 12822 6010 12824
rect 6177 12882 6243 12885
rect 6453 12882 6519 12885
rect 6177 12880 6519 12882
rect 6177 12824 6182 12880
rect 6238 12824 6458 12880
rect 6514 12824 6519 12880
rect 6177 12822 6519 12824
rect 3601 12819 3667 12822
rect 6177 12819 6243 12822
rect 6453 12819 6519 12822
rect 6821 12882 6887 12885
rect 10041 12882 10107 12885
rect 6821 12880 10107 12882
rect 6821 12824 6826 12880
rect 6882 12824 10046 12880
rect 10102 12824 10107 12880
rect 6821 12822 10107 12824
rect 6821 12819 6887 12822
rect 10041 12819 10107 12822
rect 11145 12880 11211 12885
rect 11145 12824 11150 12880
rect 11206 12824 11211 12880
rect 11145 12819 11211 12824
rect 11421 12882 11487 12885
rect 11646 12882 11652 12884
rect 11421 12880 11652 12882
rect 11421 12824 11426 12880
rect 11482 12824 11652 12880
rect 11421 12822 11652 12824
rect 11421 12819 11487 12822
rect 11646 12820 11652 12822
rect 11716 12820 11722 12884
rect 11838 12882 11898 13094
rect 13813 13091 13879 13094
rect 14273 13154 14339 13157
rect 15377 13154 15443 13157
rect 23974 13154 23980 13156
rect 14273 13152 23980 13154
rect 14273 13096 14278 13152
rect 14334 13096 15382 13152
rect 15438 13096 23980 13152
rect 14273 13094 23980 13096
rect 14273 13091 14339 13094
rect 15377 13091 15443 13094
rect 23974 13092 23980 13094
rect 24044 13092 24050 13156
rect 12014 12956 12020 13020
rect 12084 13018 12090 13020
rect 13077 13018 13143 13021
rect 12084 13016 13143 13018
rect 12084 12960 13082 13016
rect 13138 12960 13143 13016
rect 12084 12958 13143 12960
rect 12084 12956 12090 12958
rect 13077 12955 13143 12958
rect 14365 13018 14431 13021
rect 14825 13018 14891 13021
rect 14365 13016 14891 13018
rect 14365 12960 14370 13016
rect 14426 12960 14830 13016
rect 14886 12960 14891 13016
rect 14365 12958 14891 12960
rect 14365 12955 14431 12958
rect 14825 12955 14891 12958
rect 15285 13018 15351 13021
rect 15510 13018 15516 13020
rect 15285 13016 15516 13018
rect 15285 12960 15290 13016
rect 15346 12960 15516 13016
rect 15285 12958 15516 12960
rect 15285 12955 15351 12958
rect 15510 12956 15516 12958
rect 15580 12956 15586 13020
rect 17033 13018 17099 13021
rect 18965 13018 19031 13021
rect 17033 13016 19031 13018
rect 17033 12960 17038 13016
rect 17094 12960 18970 13016
rect 19026 12960 19031 13016
rect 17033 12958 19031 12960
rect 17033 12955 17099 12958
rect 18965 12955 19031 12958
rect 19374 12956 19380 13020
rect 19444 13018 19450 13020
rect 21817 13018 21883 13021
rect 19444 13016 21883 13018
rect 19444 12960 21822 13016
rect 21878 12960 21883 13016
rect 19444 12958 21883 12960
rect 19444 12956 19450 12958
rect 21817 12955 21883 12958
rect 22870 12956 22876 13020
rect 22940 13018 22946 13020
rect 25773 13018 25839 13021
rect 22940 13016 25839 13018
rect 22940 12960 25778 13016
rect 25834 12960 25839 13016
rect 22940 12958 25839 12960
rect 22940 12956 22946 12958
rect 25773 12955 25839 12958
rect 32489 13018 32555 13021
rect 33200 13018 34000 13048
rect 32489 13016 34000 13018
rect 32489 12960 32494 13016
rect 32550 12960 34000 13016
rect 32489 12958 34000 12960
rect 32489 12955 32555 12958
rect 33200 12928 34000 12958
rect 24761 12882 24827 12885
rect 11838 12880 24827 12882
rect 11838 12824 24766 12880
rect 24822 12824 24827 12880
rect 11838 12822 24827 12824
rect 24761 12819 24827 12822
rect 5073 12746 5139 12749
rect 5533 12746 5599 12749
rect 6678 12746 6684 12748
rect 5073 12744 5599 12746
rect 5073 12688 5078 12744
rect 5134 12688 5538 12744
rect 5594 12688 5599 12744
rect 5073 12686 5599 12688
rect 5073 12683 5139 12686
rect 5533 12683 5599 12686
rect 6134 12686 6684 12746
rect 5257 12610 5323 12613
rect 6134 12610 6194 12686
rect 6678 12684 6684 12686
rect 6748 12746 6754 12748
rect 6821 12746 6887 12749
rect 6748 12744 6887 12746
rect 6748 12688 6826 12744
rect 6882 12688 6887 12744
rect 6748 12686 6887 12688
rect 6748 12684 6754 12686
rect 6821 12683 6887 12686
rect 7833 12746 7899 12749
rect 8150 12746 8156 12748
rect 7833 12744 8156 12746
rect 7833 12688 7838 12744
rect 7894 12688 8156 12744
rect 7833 12686 8156 12688
rect 7833 12683 7899 12686
rect 8150 12684 8156 12686
rect 8220 12684 8226 12748
rect 9305 12746 9371 12749
rect 9673 12746 9739 12749
rect 9305 12744 9739 12746
rect 9305 12688 9310 12744
rect 9366 12688 9678 12744
rect 9734 12688 9739 12744
rect 9305 12686 9739 12688
rect 9305 12683 9371 12686
rect 9673 12683 9739 12686
rect 9857 12746 9923 12749
rect 10501 12746 10567 12749
rect 9857 12744 10567 12746
rect 9857 12688 9862 12744
rect 9918 12688 10506 12744
rect 10562 12688 10567 12744
rect 9857 12686 10567 12688
rect 11148 12746 11208 12819
rect 11789 12746 11855 12749
rect 11148 12744 11855 12746
rect 11148 12688 11794 12744
rect 11850 12688 11855 12744
rect 11148 12686 11855 12688
rect 9857 12683 9923 12686
rect 10501 12683 10567 12686
rect 11789 12683 11855 12686
rect 12065 12746 12131 12749
rect 13077 12746 13143 12749
rect 12065 12744 13143 12746
rect 12065 12688 12070 12744
rect 12126 12688 13082 12744
rect 13138 12688 13143 12744
rect 12065 12686 13143 12688
rect 12065 12683 12131 12686
rect 13077 12683 13143 12686
rect 15878 12684 15884 12748
rect 15948 12746 15954 12748
rect 17309 12746 17375 12749
rect 15948 12744 17375 12746
rect 15948 12688 17314 12744
rect 17370 12688 17375 12744
rect 15948 12686 17375 12688
rect 15948 12684 15954 12686
rect 17309 12683 17375 12686
rect 18638 12684 18644 12748
rect 18708 12746 18714 12748
rect 18781 12746 18847 12749
rect 18708 12744 18847 12746
rect 18708 12688 18786 12744
rect 18842 12688 18847 12744
rect 18708 12686 18847 12688
rect 18708 12684 18714 12686
rect 18781 12683 18847 12686
rect 18965 12746 19031 12749
rect 28809 12746 28875 12749
rect 18965 12744 28875 12746
rect 18965 12688 18970 12744
rect 19026 12688 28814 12744
rect 28870 12688 28875 12744
rect 18965 12686 28875 12688
rect 18965 12683 19031 12686
rect 28809 12683 28875 12686
rect 5257 12608 6194 12610
rect 5257 12552 5262 12608
rect 5318 12552 6194 12608
rect 5257 12550 6194 12552
rect 6637 12610 6703 12613
rect 7925 12612 7991 12613
rect 6637 12608 7850 12610
rect 6637 12552 6642 12608
rect 6698 12552 7850 12608
rect 6637 12550 7850 12552
rect 5257 12547 5323 12550
rect 6637 12547 6703 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 5257 12474 5323 12477
rect 6085 12474 6151 12477
rect 7649 12474 7715 12477
rect 5257 12472 5964 12474
rect 5257 12416 5262 12472
rect 5318 12416 5964 12472
rect 5257 12414 5964 12416
rect 5257 12411 5323 12414
rect 3734 12276 3740 12340
rect 3804 12338 3810 12340
rect 5717 12338 5783 12341
rect 3804 12336 5783 12338
rect 3804 12280 5722 12336
rect 5778 12280 5783 12336
rect 3804 12278 5783 12280
rect 5904 12338 5964 12414
rect 6085 12472 7715 12474
rect 6085 12416 6090 12472
rect 6146 12416 7654 12472
rect 7710 12416 7715 12472
rect 6085 12414 7715 12416
rect 7790 12474 7850 12550
rect 7925 12608 7972 12612
rect 8036 12610 8042 12612
rect 9765 12610 9831 12613
rect 10133 12610 10199 12613
rect 7925 12552 7930 12608
rect 7925 12548 7972 12552
rect 8036 12550 8082 12610
rect 9765 12608 10199 12610
rect 9765 12552 9770 12608
rect 9826 12552 10138 12608
rect 10194 12552 10199 12608
rect 9765 12550 10199 12552
rect 8036 12548 8042 12550
rect 7925 12547 7991 12548
rect 9765 12547 9831 12550
rect 10133 12547 10199 12550
rect 11329 12610 11395 12613
rect 22093 12610 22159 12613
rect 11329 12608 22159 12610
rect 11329 12552 11334 12608
rect 11390 12552 22098 12608
rect 22154 12552 22159 12608
rect 11329 12550 22159 12552
rect 11329 12547 11395 12550
rect 22093 12547 22159 12550
rect 22645 12610 22711 12613
rect 22645 12608 23444 12610
rect 22645 12552 22650 12608
rect 22706 12552 23444 12608
rect 22645 12550 23444 12552
rect 22645 12547 22711 12550
rect 14365 12474 14431 12477
rect 7790 12472 14431 12474
rect 7790 12416 14370 12472
rect 14426 12416 14431 12472
rect 7790 12414 14431 12416
rect 6085 12411 6151 12414
rect 7649 12411 7715 12414
rect 14365 12411 14431 12414
rect 14549 12474 14615 12477
rect 16430 12474 16436 12476
rect 14549 12472 16436 12474
rect 14549 12416 14554 12472
rect 14610 12416 16436 12472
rect 14549 12414 16436 12416
rect 14549 12411 14615 12414
rect 16430 12412 16436 12414
rect 16500 12412 16506 12476
rect 17769 12474 17835 12477
rect 18137 12474 18203 12477
rect 23197 12474 23263 12477
rect 17769 12472 18203 12474
rect 17769 12416 17774 12472
rect 17830 12416 18142 12472
rect 18198 12416 18203 12472
rect 17769 12414 18203 12416
rect 17769 12411 17835 12414
rect 18137 12411 18203 12414
rect 19290 12472 23263 12474
rect 19290 12416 23202 12472
rect 23258 12416 23263 12472
rect 19290 12414 23263 12416
rect 23384 12474 23444 12550
rect 24945 12474 25011 12477
rect 23384 12472 25011 12474
rect 23384 12416 24950 12472
rect 25006 12416 25011 12472
rect 23384 12414 25011 12416
rect 6494 12338 6500 12340
rect 5904 12278 6500 12338
rect 3804 12276 3810 12278
rect 5717 12275 5783 12278
rect 6494 12276 6500 12278
rect 6564 12276 6570 12340
rect 6913 12338 6979 12341
rect 12341 12338 12407 12341
rect 14549 12338 14615 12341
rect 15694 12338 15700 12340
rect 6913 12336 12450 12338
rect 6913 12280 6918 12336
rect 6974 12280 12346 12336
rect 12402 12280 12450 12336
rect 6913 12278 12450 12280
rect 6913 12275 6979 12278
rect 12341 12275 12450 12278
rect 14549 12336 15700 12338
rect 14549 12280 14554 12336
rect 14610 12280 15700 12336
rect 14549 12278 15700 12280
rect 14549 12275 14615 12278
rect 15694 12276 15700 12278
rect 15764 12276 15770 12340
rect 15837 12338 15903 12341
rect 19290 12338 19350 12414
rect 23197 12411 23263 12414
rect 24945 12411 25011 12414
rect 25405 12474 25471 12477
rect 25773 12474 25839 12477
rect 28441 12476 28507 12477
rect 25405 12472 25839 12474
rect 25405 12416 25410 12472
rect 25466 12416 25778 12472
rect 25834 12416 25839 12472
rect 25405 12414 25839 12416
rect 25405 12411 25471 12414
rect 25773 12411 25839 12414
rect 28390 12412 28396 12476
rect 28460 12474 28507 12476
rect 28460 12472 28552 12474
rect 28502 12416 28552 12472
rect 28460 12414 28552 12416
rect 28460 12412 28507 12414
rect 28441 12411 28507 12412
rect 15837 12336 19350 12338
rect 15837 12280 15842 12336
rect 15898 12280 19350 12336
rect 15837 12278 19350 12280
rect 19609 12338 19675 12341
rect 20294 12338 20300 12340
rect 19609 12336 20300 12338
rect 19609 12280 19614 12336
rect 19670 12280 20300 12336
rect 19609 12278 20300 12280
rect 15837 12275 15903 12278
rect 19609 12275 19675 12278
rect 20294 12276 20300 12278
rect 20364 12276 20370 12340
rect 21449 12338 21515 12341
rect 23933 12338 23999 12341
rect 21449 12336 23999 12338
rect 21449 12280 21454 12336
rect 21510 12280 23938 12336
rect 23994 12280 23999 12336
rect 21449 12278 23999 12280
rect 21449 12275 21515 12278
rect 23933 12275 23999 12278
rect 24945 12338 25011 12341
rect 25078 12338 25084 12340
rect 24945 12336 25084 12338
rect 24945 12280 24950 12336
rect 25006 12280 25084 12336
rect 24945 12278 25084 12280
rect 24945 12275 25011 12278
rect 25078 12276 25084 12278
rect 25148 12338 25154 12340
rect 25957 12338 26023 12341
rect 25148 12336 26023 12338
rect 25148 12280 25962 12336
rect 26018 12280 26023 12336
rect 25148 12278 26023 12280
rect 25148 12276 25154 12278
rect 25957 12275 26023 12278
rect 29678 12276 29684 12340
rect 29748 12338 29754 12340
rect 29913 12338 29979 12341
rect 29748 12336 29979 12338
rect 29748 12280 29918 12336
rect 29974 12280 29979 12336
rect 29748 12278 29979 12280
rect 29748 12276 29754 12278
rect 29913 12275 29979 12278
rect 2957 12202 3023 12205
rect 5720 12202 5780 12275
rect 7649 12202 7715 12205
rect 2957 12200 5642 12202
rect 2957 12144 2962 12200
rect 3018 12144 5642 12200
rect 2957 12142 5642 12144
rect 5720 12200 7715 12202
rect 5720 12144 7654 12200
rect 7710 12144 7715 12200
rect 5720 12142 7715 12144
rect 2957 12139 3023 12142
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 5582 11933 5642 12142
rect 7649 12139 7715 12142
rect 7782 12140 7788 12204
rect 7852 12202 7858 12204
rect 11421 12202 11487 12205
rect 7852 12142 10932 12202
rect 7852 12140 7858 12142
rect 10872 12069 10932 12142
rect 11056 12200 11487 12202
rect 11056 12144 11426 12200
rect 11482 12144 11487 12200
rect 11056 12142 11487 12144
rect 11056 12069 11116 12142
rect 11421 12139 11487 12142
rect 11697 12202 11763 12205
rect 12390 12202 12450 12275
rect 19425 12202 19491 12205
rect 27245 12202 27311 12205
rect 11697 12200 12036 12202
rect 11697 12144 11702 12200
rect 11758 12144 12036 12200
rect 11697 12142 12036 12144
rect 12390 12200 19491 12202
rect 12390 12144 19430 12200
rect 19486 12144 19491 12200
rect 12390 12142 19491 12144
rect 11697 12139 11763 12142
rect 5717 12066 5783 12069
rect 7557 12066 7623 12069
rect 5717 12064 5964 12066
rect 5717 12008 5722 12064
rect 5778 12008 5964 12064
rect 5717 12006 5964 12008
rect 5717 12003 5783 12006
rect 4337 11930 4403 11933
rect 4654 11930 4660 11932
rect 4337 11928 4660 11930
rect 4337 11872 4342 11928
rect 4398 11872 4660 11928
rect 4337 11870 4660 11872
rect 4337 11867 4403 11870
rect 4654 11868 4660 11870
rect 4724 11868 4730 11932
rect 5582 11928 5691 11933
rect 5582 11872 5630 11928
rect 5686 11872 5691 11928
rect 5582 11870 5691 11872
rect 5625 11867 5691 11870
rect 1158 11732 1164 11796
rect 1228 11794 1234 11796
rect 5625 11794 5691 11797
rect 1228 11792 5691 11794
rect 1228 11736 5630 11792
rect 5686 11736 5691 11792
rect 1228 11734 5691 11736
rect 5904 11794 5964 12006
rect 6870 12064 7623 12066
rect 6870 12008 7562 12064
rect 7618 12008 7623 12064
rect 6870 12006 7623 12008
rect 6545 11932 6611 11933
rect 6494 11930 6500 11932
rect 6454 11870 6500 11930
rect 6564 11928 6611 11932
rect 6606 11872 6611 11928
rect 6494 11868 6500 11870
rect 6564 11868 6611 11872
rect 6545 11867 6611 11868
rect 6729 11930 6795 11933
rect 6870 11930 6930 12006
rect 7557 12003 7623 12006
rect 8109 12066 8175 12069
rect 9581 12066 9647 12069
rect 8109 12064 9647 12066
rect 8109 12008 8114 12064
rect 8170 12008 9586 12064
rect 9642 12008 9647 12064
rect 8109 12006 9647 12008
rect 8109 12003 8175 12006
rect 9581 12003 9647 12006
rect 10869 12064 10935 12069
rect 10869 12008 10874 12064
rect 10930 12008 10935 12064
rect 10869 12003 10935 12008
rect 11053 12064 11119 12069
rect 11053 12008 11058 12064
rect 11114 12008 11119 12064
rect 11053 12003 11119 12008
rect 11237 12068 11303 12069
rect 11237 12064 11284 12068
rect 11348 12066 11354 12068
rect 11237 12008 11242 12064
rect 11237 12004 11284 12008
rect 11348 12006 11394 12066
rect 11348 12004 11354 12006
rect 11462 12004 11468 12068
rect 11532 12066 11538 12068
rect 11789 12066 11855 12069
rect 11532 12064 11855 12066
rect 11532 12008 11794 12064
rect 11850 12008 11855 12064
rect 11532 12006 11855 12008
rect 11976 12066 12036 12142
rect 19425 12139 19491 12142
rect 22050 12200 27311 12202
rect 22050 12144 27250 12200
rect 27306 12144 27311 12200
rect 22050 12142 27311 12144
rect 15837 12066 15903 12069
rect 11976 12064 15903 12066
rect 11976 12008 15842 12064
rect 15898 12008 15903 12064
rect 11976 12006 15903 12008
rect 11532 12004 11538 12006
rect 11237 12003 11303 12004
rect 11789 12003 11855 12006
rect 15837 12003 15903 12006
rect 17217 12066 17283 12069
rect 22050 12066 22110 12142
rect 27245 12139 27311 12142
rect 17217 12064 22110 12066
rect 17217 12008 17222 12064
rect 17278 12008 22110 12064
rect 17217 12006 22110 12008
rect 22185 12066 22251 12069
rect 25589 12066 25655 12069
rect 28625 12068 28691 12069
rect 28574 12066 28580 12068
rect 22185 12064 25655 12066
rect 22185 12008 22190 12064
rect 22246 12008 25594 12064
rect 25650 12008 25655 12064
rect 22185 12006 25655 12008
rect 28534 12006 28580 12066
rect 28644 12064 28691 12068
rect 28686 12008 28691 12064
rect 17217 12003 17283 12006
rect 22185 12003 22251 12006
rect 25589 12003 25655 12006
rect 28574 12004 28580 12006
rect 28644 12004 28691 12008
rect 28625 12003 28691 12004
rect 6729 11928 6930 11930
rect 6729 11872 6734 11928
rect 6790 11872 6930 11928
rect 6729 11870 6930 11872
rect 7005 11930 7071 11933
rect 13813 11930 13879 11933
rect 14457 11930 14523 11933
rect 7005 11928 13879 11930
rect 7005 11872 7010 11928
rect 7066 11872 13818 11928
rect 13874 11872 13879 11928
rect 7005 11870 13879 11872
rect 6729 11867 6795 11870
rect 7005 11867 7071 11870
rect 13813 11867 13879 11870
rect 14230 11928 14523 11930
rect 14230 11872 14462 11928
rect 14518 11872 14523 11928
rect 14230 11870 14523 11872
rect 9121 11794 9187 11797
rect 14230 11794 14290 11870
rect 14457 11867 14523 11870
rect 14958 11868 14964 11932
rect 15028 11930 15034 11932
rect 15469 11930 15535 11933
rect 15028 11928 15535 11930
rect 15028 11872 15474 11928
rect 15530 11872 15535 11928
rect 15028 11870 15535 11872
rect 15028 11868 15034 11870
rect 15469 11867 15535 11870
rect 16246 11868 16252 11932
rect 16316 11930 16322 11932
rect 17861 11930 17927 11933
rect 16316 11928 17927 11930
rect 16316 11872 17866 11928
rect 17922 11872 17927 11928
rect 16316 11870 17927 11872
rect 16316 11868 16322 11870
rect 17861 11867 17927 11870
rect 19425 11930 19491 11933
rect 29269 11930 29335 11933
rect 19425 11928 29335 11930
rect 19425 11872 19430 11928
rect 19486 11872 29274 11928
rect 29330 11872 29335 11928
rect 19425 11870 29335 11872
rect 19425 11867 19491 11870
rect 29269 11867 29335 11870
rect 5904 11792 14290 11794
rect 5904 11736 9126 11792
rect 9182 11736 14290 11792
rect 5904 11734 14290 11736
rect 14457 11794 14523 11797
rect 14590 11794 14596 11796
rect 14457 11792 14596 11794
rect 14457 11736 14462 11792
rect 14518 11736 14596 11792
rect 14457 11734 14596 11736
rect 1228 11732 1234 11734
rect 5625 11731 5691 11734
rect 9121 11731 9187 11734
rect 14457 11731 14523 11734
rect 14590 11732 14596 11734
rect 14660 11732 14666 11796
rect 14733 11794 14799 11797
rect 21398 11794 21404 11796
rect 14733 11792 21404 11794
rect 14733 11736 14738 11792
rect 14794 11736 21404 11792
rect 14733 11734 21404 11736
rect 14733 11731 14799 11734
rect 21398 11732 21404 11734
rect 21468 11732 21474 11796
rect 23933 11794 23999 11797
rect 24710 11794 24716 11796
rect 23933 11792 24716 11794
rect 23933 11736 23938 11792
rect 23994 11736 24716 11792
rect 23933 11734 24716 11736
rect 23933 11731 23999 11734
rect 24710 11732 24716 11734
rect 24780 11732 24786 11796
rect 4153 11658 4219 11661
rect 6453 11658 6519 11661
rect 4153 11656 6519 11658
rect 4153 11600 4158 11656
rect 4214 11600 6458 11656
rect 6514 11600 6519 11656
rect 4153 11598 6519 11600
rect 4153 11595 4219 11598
rect 6453 11595 6519 11598
rect 7005 11658 7071 11661
rect 7649 11660 7715 11661
rect 7414 11658 7420 11660
rect 7005 11656 7420 11658
rect 7005 11600 7010 11656
rect 7066 11600 7420 11656
rect 7005 11598 7420 11600
rect 7005 11595 7071 11598
rect 7414 11596 7420 11598
rect 7484 11596 7490 11660
rect 7598 11596 7604 11660
rect 7668 11658 7715 11660
rect 8661 11658 8727 11661
rect 9489 11658 9555 11661
rect 7668 11656 7760 11658
rect 7710 11600 7760 11656
rect 7668 11598 7760 11600
rect 8661 11656 9555 11658
rect 8661 11600 8666 11656
rect 8722 11600 9494 11656
rect 9550 11600 9555 11656
rect 8661 11598 9555 11600
rect 7668 11596 7715 11598
rect 7649 11595 7715 11596
rect 8661 11595 8727 11598
rect 9489 11595 9555 11598
rect 10041 11658 10107 11661
rect 10409 11660 10475 11661
rect 10174 11658 10180 11660
rect 10041 11656 10180 11658
rect 10041 11600 10046 11656
rect 10102 11600 10180 11656
rect 10041 11598 10180 11600
rect 10041 11595 10107 11598
rect 10174 11596 10180 11598
rect 10244 11596 10250 11660
rect 10358 11658 10364 11660
rect 10318 11598 10364 11658
rect 10428 11656 10475 11660
rect 10470 11600 10475 11656
rect 10358 11596 10364 11598
rect 10428 11596 10475 11600
rect 10409 11595 10475 11596
rect 10869 11658 10935 11661
rect 15009 11658 15075 11661
rect 10869 11656 15075 11658
rect 10869 11600 10874 11656
rect 10930 11600 15014 11656
rect 15070 11600 15075 11656
rect 10869 11598 15075 11600
rect 10869 11595 10935 11598
rect 15009 11595 15075 11598
rect 16430 11596 16436 11660
rect 16500 11658 16506 11660
rect 17125 11658 17191 11661
rect 16500 11656 17191 11658
rect 16500 11600 17130 11656
rect 17186 11600 17191 11656
rect 16500 11598 17191 11600
rect 16500 11596 16506 11598
rect 17125 11595 17191 11598
rect 20345 11658 20411 11661
rect 20662 11658 20668 11660
rect 20345 11656 20668 11658
rect 20345 11600 20350 11656
rect 20406 11600 20668 11656
rect 20345 11598 20668 11600
rect 20345 11595 20411 11598
rect 20662 11596 20668 11598
rect 20732 11596 20738 11660
rect 32397 11658 32463 11661
rect 33200 11658 34000 11688
rect 32397 11656 34000 11658
rect 32397 11600 32402 11656
rect 32458 11600 34000 11656
rect 32397 11598 34000 11600
rect 32397 11595 32463 11598
rect 33200 11568 34000 11598
rect 5165 11522 5231 11525
rect 7005 11522 7071 11525
rect 5165 11520 7071 11522
rect 5165 11464 5170 11520
rect 5226 11464 7010 11520
rect 7066 11464 7071 11520
rect 5165 11462 7071 11464
rect 5165 11459 5231 11462
rect 7005 11459 7071 11462
rect 8569 11522 8635 11525
rect 12065 11522 12131 11525
rect 8569 11520 12131 11522
rect 8569 11464 8574 11520
rect 8630 11464 12070 11520
rect 12126 11464 12131 11520
rect 8569 11462 12131 11464
rect 8569 11459 8635 11462
rect 12065 11459 12131 11462
rect 13813 11522 13879 11525
rect 16573 11522 16639 11525
rect 16982 11522 16988 11524
rect 13813 11520 16988 11522
rect 13813 11464 13818 11520
rect 13874 11464 16578 11520
rect 16634 11464 16988 11520
rect 13813 11462 16988 11464
rect 13813 11459 13879 11462
rect 16573 11459 16639 11462
rect 16982 11460 16988 11462
rect 17052 11460 17058 11524
rect 20846 11522 20852 11524
rect 17128 11462 20852 11522
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 5349 11388 5415 11389
rect 5349 11386 5396 11388
rect 5304 11384 5396 11386
rect 5304 11328 5354 11384
rect 5304 11326 5396 11328
rect 5349 11324 5396 11326
rect 5460 11324 5466 11388
rect 5993 11386 6059 11389
rect 7598 11386 7604 11388
rect 5993 11384 7604 11386
rect 5993 11328 5998 11384
rect 6054 11328 7604 11384
rect 5993 11326 7604 11328
rect 5349 11323 5415 11324
rect 5993 11323 6059 11326
rect 7598 11324 7604 11326
rect 7668 11324 7674 11388
rect 8661 11386 8727 11389
rect 16297 11386 16363 11389
rect 8661 11384 16363 11386
rect 8661 11328 8666 11384
rect 8722 11328 16302 11384
rect 16358 11328 16363 11384
rect 8661 11326 16363 11328
rect 8661 11323 8727 11326
rect 16297 11323 16363 11326
rect 16481 11386 16547 11389
rect 17128 11386 17188 11462
rect 20846 11460 20852 11462
rect 20916 11460 20922 11524
rect 21817 11522 21883 11525
rect 32029 11522 32095 11525
rect 21817 11520 32095 11522
rect 21817 11464 21822 11520
rect 21878 11464 32034 11520
rect 32090 11464 32095 11520
rect 21817 11462 32095 11464
rect 21817 11459 21883 11462
rect 32029 11459 32095 11462
rect 16481 11384 17188 11386
rect 16481 11328 16486 11384
rect 16542 11328 17188 11384
rect 16481 11326 17188 11328
rect 19333 11386 19399 11389
rect 20478 11386 20484 11388
rect 19333 11384 20484 11386
rect 19333 11328 19338 11384
rect 19394 11328 20484 11384
rect 19333 11326 20484 11328
rect 16481 11323 16547 11326
rect 19333 11323 19399 11326
rect 20478 11324 20484 11326
rect 20548 11386 20554 11388
rect 26325 11386 26391 11389
rect 27153 11386 27219 11389
rect 20548 11384 27219 11386
rect 20548 11328 26330 11384
rect 26386 11328 27158 11384
rect 27214 11328 27219 11384
rect 20548 11326 27219 11328
rect 20548 11324 20554 11326
rect 26325 11323 26391 11326
rect 27153 11323 27219 11326
rect 2865 11250 2931 11253
rect 6637 11250 6703 11253
rect 7465 11250 7531 11253
rect 2865 11248 6424 11250
rect 2865 11192 2870 11248
rect 2926 11192 6424 11248
rect 2865 11190 6424 11192
rect 2865 11187 2931 11190
rect 6364 11117 6424 11190
rect 6637 11248 7531 11250
rect 6637 11192 6642 11248
rect 6698 11192 7470 11248
rect 7526 11192 7531 11248
rect 6637 11190 7531 11192
rect 6637 11187 6703 11190
rect 7465 11187 7531 11190
rect 8569 11250 8635 11253
rect 10726 11250 10732 11252
rect 8569 11248 10732 11250
rect 8569 11192 8574 11248
rect 8630 11192 10732 11248
rect 8569 11190 10732 11192
rect 8569 11187 8635 11190
rect 10726 11188 10732 11190
rect 10796 11250 10802 11252
rect 16481 11250 16547 11253
rect 10796 11248 16547 11250
rect 10796 11192 16486 11248
rect 16542 11192 16547 11248
rect 10796 11190 16547 11192
rect 10796 11188 10802 11190
rect 16481 11187 16547 11190
rect 19609 11250 19675 11253
rect 23013 11250 23079 11253
rect 19609 11248 23079 11250
rect 19609 11192 19614 11248
rect 19670 11192 23018 11248
rect 23074 11192 23079 11248
rect 19609 11190 23079 11192
rect 19609 11187 19675 11190
rect 23013 11187 23079 11190
rect 2221 11114 2287 11117
rect 2865 11114 2931 11117
rect 2221 11112 2931 11114
rect 2221 11056 2226 11112
rect 2282 11056 2870 11112
rect 2926 11056 2931 11112
rect 2221 11054 2931 11056
rect 2221 11051 2287 11054
rect 2865 11051 2931 11054
rect 3918 11052 3924 11116
rect 3988 11114 3994 11116
rect 5625 11114 5691 11117
rect 3988 11112 5691 11114
rect 3988 11056 5630 11112
rect 5686 11056 5691 11112
rect 3988 11054 5691 11056
rect 3988 11052 3994 11054
rect 5625 11051 5691 11054
rect 6361 11114 6427 11117
rect 10225 11114 10291 11117
rect 10869 11114 10935 11117
rect 6361 11112 9690 11114
rect 6361 11056 6366 11112
rect 6422 11056 9690 11112
rect 6361 11054 9690 11056
rect 6361 11051 6427 11054
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 5349 10978 5415 10981
rect 5901 10978 5967 10981
rect 5349 10976 5967 10978
rect 5349 10920 5354 10976
rect 5410 10920 5906 10976
rect 5962 10920 5967 10976
rect 5349 10918 5967 10920
rect 5349 10915 5415 10918
rect 5901 10915 5967 10918
rect 6126 10916 6132 10980
rect 6196 10978 6202 10980
rect 6361 10978 6427 10981
rect 6196 10976 6427 10978
rect 6196 10920 6366 10976
rect 6422 10920 6427 10976
rect 6196 10918 6427 10920
rect 6196 10916 6202 10918
rect 6361 10915 6427 10918
rect 6637 10980 6703 10981
rect 6637 10976 6684 10980
rect 6748 10978 6754 10980
rect 7649 10978 7715 10981
rect 6748 10976 7715 10978
rect 6637 10920 6642 10976
rect 6748 10920 7654 10976
rect 7710 10920 7715 10976
rect 6637 10916 6684 10920
rect 6748 10918 7715 10920
rect 9630 10978 9690 11054
rect 10225 11112 10935 11114
rect 10225 11056 10230 11112
rect 10286 11056 10874 11112
rect 10930 11056 10935 11112
rect 10225 11054 10935 11056
rect 10225 11051 10291 11054
rect 10869 11051 10935 11054
rect 12382 11052 12388 11116
rect 12452 11114 12458 11116
rect 16941 11114 17007 11117
rect 12452 11112 17007 11114
rect 12452 11056 16946 11112
rect 17002 11056 17007 11112
rect 12452 11054 17007 11056
rect 12452 11052 12458 11054
rect 16941 11051 17007 11054
rect 17350 11052 17356 11116
rect 17420 11114 17426 11116
rect 17585 11114 17651 11117
rect 17420 11112 17651 11114
rect 17420 11056 17590 11112
rect 17646 11056 17651 11112
rect 17420 11054 17651 11056
rect 17420 11052 17426 11054
rect 17585 11051 17651 11054
rect 18505 11114 18571 11117
rect 19558 11114 19564 11116
rect 18505 11112 19564 11114
rect 18505 11056 18510 11112
rect 18566 11056 19564 11112
rect 18505 11054 19564 11056
rect 18505 11051 18571 11054
rect 19558 11052 19564 11054
rect 19628 11052 19634 11116
rect 19885 11114 19951 11117
rect 20345 11114 20411 11117
rect 20897 11116 20963 11117
rect 20846 11114 20852 11116
rect 19885 11112 20411 11114
rect 19885 11056 19890 11112
rect 19946 11056 20350 11112
rect 20406 11056 20411 11112
rect 19885 11054 20411 11056
rect 20806 11054 20852 11114
rect 20916 11112 20963 11116
rect 20958 11056 20963 11112
rect 19885 11051 19951 11054
rect 20345 11051 20411 11054
rect 20846 11052 20852 11054
rect 20916 11052 20963 11056
rect 21214 11052 21220 11116
rect 21284 11114 21290 11116
rect 22645 11114 22711 11117
rect 21284 11112 22711 11114
rect 21284 11056 22650 11112
rect 22706 11056 22711 11112
rect 21284 11054 22711 11056
rect 21284 11052 21290 11054
rect 20897 11051 20963 11052
rect 22645 11051 22711 11054
rect 24209 11114 24275 11117
rect 27797 11114 27863 11117
rect 24209 11112 27863 11114
rect 24209 11056 24214 11112
rect 24270 11056 27802 11112
rect 27858 11056 27863 11112
rect 24209 11054 27863 11056
rect 24209 11051 24275 11054
rect 27797 11051 27863 11054
rect 15101 10978 15167 10981
rect 9630 10976 15167 10978
rect 9630 10920 15106 10976
rect 15162 10920 15167 10976
rect 9630 10918 15167 10920
rect 6748 10916 6754 10918
rect 6637 10915 6703 10916
rect 7649 10915 7715 10918
rect 15101 10915 15167 10918
rect 15510 10916 15516 10980
rect 15580 10978 15586 10980
rect 18781 10978 18847 10981
rect 15580 10976 18847 10978
rect 15580 10920 18786 10976
rect 18842 10920 18847 10976
rect 15580 10918 18847 10920
rect 15580 10916 15586 10918
rect 18781 10915 18847 10918
rect 19241 10978 19307 10981
rect 20897 10978 20963 10981
rect 19241 10976 20963 10978
rect 19241 10920 19246 10976
rect 19302 10920 20902 10976
rect 20958 10920 20963 10976
rect 19241 10918 20963 10920
rect 19241 10915 19307 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 20348 10845 20408 10918
rect 20897 10915 20963 10918
rect 21081 10978 21147 10981
rect 24301 10978 24367 10981
rect 26918 10978 26924 10980
rect 21081 10976 24226 10978
rect 21081 10920 21086 10976
rect 21142 10920 24226 10976
rect 21081 10918 24226 10920
rect 21081 10915 21147 10918
rect 933 10842 999 10845
rect 4705 10842 4771 10845
rect 933 10840 4771 10842
rect 933 10784 938 10840
rect 994 10784 4710 10840
rect 4766 10784 4771 10840
rect 933 10782 4771 10784
rect 933 10779 999 10782
rect 4705 10779 4771 10782
rect 5533 10842 5599 10845
rect 8661 10842 8727 10845
rect 16757 10842 16823 10845
rect 17493 10842 17559 10845
rect 5533 10840 8586 10842
rect 5533 10784 5538 10840
rect 5594 10784 8586 10840
rect 5533 10782 8586 10784
rect 5533 10779 5599 10782
rect 4429 10706 4495 10709
rect 6862 10706 6868 10708
rect 4429 10704 6868 10706
rect 4429 10648 4434 10704
rect 4490 10648 6868 10704
rect 4429 10646 6868 10648
rect 4429 10643 4495 10646
rect 6862 10644 6868 10646
rect 6932 10644 6938 10708
rect 7373 10706 7439 10709
rect 8334 10706 8340 10708
rect 7373 10704 8340 10706
rect 7373 10648 7378 10704
rect 7434 10648 8340 10704
rect 7373 10646 8340 10648
rect 7373 10643 7439 10646
rect 8334 10644 8340 10646
rect 8404 10644 8410 10708
rect 2262 10508 2268 10572
rect 2332 10570 2338 10572
rect 8526 10570 8586 10782
rect 8661 10840 12450 10842
rect 8661 10784 8666 10840
rect 8722 10784 12450 10840
rect 8661 10782 12450 10784
rect 8661 10779 8727 10782
rect 9070 10644 9076 10708
rect 9140 10706 9146 10708
rect 9397 10706 9463 10709
rect 9140 10704 9463 10706
rect 9140 10648 9402 10704
rect 9458 10648 9463 10704
rect 9140 10646 9463 10648
rect 9140 10644 9146 10646
rect 9397 10643 9463 10646
rect 9622 10644 9628 10708
rect 9692 10706 9698 10708
rect 11697 10706 11763 10709
rect 9692 10704 11763 10706
rect 9692 10648 11702 10704
rect 11758 10648 11763 10704
rect 9692 10646 11763 10648
rect 12390 10706 12450 10782
rect 16757 10840 17559 10842
rect 16757 10784 16762 10840
rect 16818 10784 17498 10840
rect 17554 10784 17559 10840
rect 16757 10782 17559 10784
rect 16757 10779 16823 10782
rect 17493 10779 17559 10782
rect 20345 10840 20411 10845
rect 20345 10784 20350 10840
rect 20406 10784 20411 10840
rect 20345 10779 20411 10784
rect 20529 10842 20595 10845
rect 22737 10844 22803 10845
rect 22318 10842 22324 10844
rect 20529 10840 22324 10842
rect 20529 10784 20534 10840
rect 20590 10784 22324 10840
rect 20529 10782 22324 10784
rect 20529 10779 20595 10782
rect 22318 10780 22324 10782
rect 22388 10780 22394 10844
rect 22686 10842 22692 10844
rect 22646 10782 22692 10842
rect 22756 10840 22803 10844
rect 23933 10844 23999 10845
rect 23933 10842 23980 10844
rect 22798 10784 22803 10840
rect 22686 10780 22692 10782
rect 22756 10780 22803 10784
rect 23888 10840 23980 10842
rect 23888 10784 23938 10840
rect 23888 10782 23980 10784
rect 22737 10779 22803 10780
rect 23933 10780 23980 10782
rect 24044 10780 24050 10844
rect 24166 10842 24226 10918
rect 24301 10976 26924 10978
rect 24301 10920 24306 10976
rect 24362 10920 26924 10976
rect 24301 10918 26924 10920
rect 24301 10915 24367 10918
rect 26918 10916 26924 10918
rect 26988 10916 26994 10980
rect 27981 10842 28047 10845
rect 24166 10840 28047 10842
rect 24166 10784 27986 10840
rect 28042 10784 28047 10840
rect 24166 10782 28047 10784
rect 23933 10779 23999 10780
rect 27981 10779 28047 10782
rect 22001 10706 22067 10709
rect 24117 10708 24183 10709
rect 24117 10706 24164 10708
rect 12390 10704 22067 10706
rect 12390 10648 22006 10704
rect 22062 10648 22067 10704
rect 12390 10646 22067 10648
rect 24072 10704 24164 10706
rect 24072 10648 24122 10704
rect 24072 10646 24164 10648
rect 9692 10644 9698 10646
rect 11697 10643 11763 10646
rect 22001 10643 22067 10646
rect 24117 10644 24164 10646
rect 24228 10644 24234 10708
rect 25681 10706 25747 10709
rect 26785 10706 26851 10709
rect 25681 10704 26851 10706
rect 25681 10648 25686 10704
rect 25742 10648 26790 10704
rect 26846 10648 26851 10704
rect 25681 10646 26851 10648
rect 24117 10643 24183 10644
rect 25681 10643 25747 10646
rect 26785 10643 26851 10646
rect 2332 10510 7666 10570
rect 8526 10510 9690 10570
rect 2332 10508 2338 10510
rect 4797 10434 4863 10437
rect 6729 10434 6795 10437
rect 4797 10432 6795 10434
rect 4797 10376 4802 10432
rect 4858 10376 6734 10432
rect 6790 10376 6795 10432
rect 4797 10374 6795 10376
rect 4797 10371 4863 10374
rect 6729 10371 6795 10374
rect 6862 10372 6868 10436
rect 6932 10434 6938 10436
rect 7097 10434 7163 10437
rect 6932 10432 7163 10434
rect 6932 10376 7102 10432
rect 7158 10376 7163 10432
rect 6932 10374 7163 10376
rect 6932 10372 6938 10374
rect 7097 10371 7163 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 4705 10298 4771 10301
rect 6310 10298 6316 10300
rect 4705 10296 6316 10298
rect 4705 10240 4710 10296
rect 4766 10240 6316 10296
rect 4705 10238 6316 10240
rect 4705 10235 4771 10238
rect 6310 10236 6316 10238
rect 6380 10236 6386 10300
rect 6494 10236 6500 10300
rect 6564 10298 6570 10300
rect 6729 10298 6795 10301
rect 6564 10296 6795 10298
rect 6564 10240 6734 10296
rect 6790 10240 6795 10296
rect 6564 10238 6795 10240
rect 6564 10236 6570 10238
rect 6729 10235 6795 10238
rect 790 10100 796 10164
rect 860 10162 866 10164
rect 4981 10162 5047 10165
rect 860 10160 5047 10162
rect 860 10104 4986 10160
rect 5042 10104 5047 10160
rect 860 10102 5047 10104
rect 860 10100 866 10102
rect 4981 10099 5047 10102
rect 5349 10162 5415 10165
rect 6913 10162 6979 10165
rect 5349 10160 6979 10162
rect 5349 10104 5354 10160
rect 5410 10104 6918 10160
rect 6974 10104 6979 10160
rect 5349 10102 6979 10104
rect 5349 10099 5415 10102
rect 6913 10099 6979 10102
rect 3918 9964 3924 10028
rect 3988 10026 3994 10028
rect 4153 10026 4219 10029
rect 6913 10026 6979 10029
rect 3988 10024 4219 10026
rect 3988 9968 4158 10024
rect 4214 9968 4219 10024
rect 3988 9966 4219 9968
rect 3988 9964 3994 9966
rect 4153 9963 4219 9966
rect 4662 10024 6979 10026
rect 4662 9968 6918 10024
rect 6974 9968 6979 10024
rect 4662 9966 6979 9968
rect 1894 9692 1900 9756
rect 1964 9754 1970 9756
rect 4662 9754 4722 9966
rect 6913 9963 6979 9966
rect 6545 9890 6611 9893
rect 5260 9888 6611 9890
rect 5260 9832 6550 9888
rect 6606 9832 6611 9888
rect 5260 9830 6611 9832
rect 7606 9890 7666 10510
rect 9630 10434 9690 10510
rect 10174 10508 10180 10572
rect 10244 10570 10250 10572
rect 15837 10570 15903 10573
rect 10244 10568 15903 10570
rect 10244 10512 15842 10568
rect 15898 10512 15903 10568
rect 10244 10510 15903 10512
rect 10244 10508 10250 10510
rect 15837 10507 15903 10510
rect 16021 10570 16087 10573
rect 18781 10570 18847 10573
rect 16021 10568 18847 10570
rect 16021 10512 16026 10568
rect 16082 10512 18786 10568
rect 18842 10512 18847 10568
rect 16021 10510 18847 10512
rect 16021 10507 16087 10510
rect 18781 10507 18847 10510
rect 19793 10570 19859 10573
rect 21173 10570 21239 10573
rect 19793 10568 21239 10570
rect 19793 10512 19798 10568
rect 19854 10512 21178 10568
rect 21234 10512 21239 10568
rect 19793 10510 21239 10512
rect 19793 10507 19859 10510
rect 21173 10507 21239 10510
rect 21357 10570 21423 10573
rect 30782 10570 30788 10572
rect 21357 10568 30788 10570
rect 21357 10512 21362 10568
rect 21418 10512 30788 10568
rect 21357 10510 30788 10512
rect 21357 10507 21423 10510
rect 30782 10508 30788 10510
rect 30852 10508 30858 10572
rect 10501 10434 10567 10437
rect 12525 10436 12591 10437
rect 9630 10432 12450 10434
rect 9630 10376 10506 10432
rect 10562 10376 12450 10432
rect 9630 10374 12450 10376
rect 10501 10371 10567 10374
rect 8569 10298 8635 10301
rect 12065 10298 12131 10301
rect 8569 10296 12131 10298
rect 8569 10240 8574 10296
rect 8630 10240 12070 10296
rect 12126 10240 12131 10296
rect 8569 10238 12131 10240
rect 12390 10298 12450 10374
rect 12525 10432 12572 10436
rect 12636 10434 12642 10436
rect 16297 10434 16363 10437
rect 25405 10434 25471 10437
rect 32581 10434 32647 10437
rect 12525 10376 12530 10432
rect 12525 10372 12572 10376
rect 12636 10374 12682 10434
rect 16297 10432 25471 10434
rect 16297 10376 16302 10432
rect 16358 10376 25410 10432
rect 25466 10376 25471 10432
rect 16297 10374 25471 10376
rect 12636 10372 12642 10374
rect 12525 10371 12591 10372
rect 16297 10371 16363 10374
rect 25405 10371 25471 10374
rect 31710 10432 32647 10434
rect 31710 10376 32586 10432
rect 32642 10376 32647 10432
rect 31710 10374 32647 10376
rect 12709 10298 12775 10301
rect 12390 10296 12775 10298
rect 12390 10240 12714 10296
rect 12770 10240 12775 10296
rect 12390 10238 12775 10240
rect 8569 10235 8635 10238
rect 12065 10235 12131 10238
rect 12709 10235 12775 10238
rect 14457 10298 14523 10301
rect 19374 10298 19380 10300
rect 14457 10296 19380 10298
rect 14457 10240 14462 10296
rect 14518 10240 19380 10296
rect 14457 10238 19380 10240
rect 14457 10235 14523 10238
rect 19374 10236 19380 10238
rect 19444 10236 19450 10300
rect 20621 10298 20687 10301
rect 20846 10298 20852 10300
rect 20621 10296 20852 10298
rect 20621 10240 20626 10296
rect 20682 10240 20852 10296
rect 20621 10238 20852 10240
rect 20621 10235 20687 10238
rect 20846 10236 20852 10238
rect 20916 10236 20922 10300
rect 22645 10298 22711 10301
rect 23013 10298 23079 10301
rect 22645 10296 23079 10298
rect 22645 10240 22650 10296
rect 22706 10240 23018 10296
rect 23074 10240 23079 10296
rect 22645 10238 23079 10240
rect 22645 10235 22711 10238
rect 23013 10235 23079 10238
rect 23422 10236 23428 10300
rect 23492 10298 23498 10300
rect 23565 10298 23631 10301
rect 23492 10296 23631 10298
rect 23492 10240 23570 10296
rect 23626 10240 23631 10296
rect 23492 10238 23631 10240
rect 23492 10236 23498 10238
rect 23565 10235 23631 10238
rect 24117 10298 24183 10301
rect 29862 10298 29868 10300
rect 24117 10296 29868 10298
rect 24117 10240 24122 10296
rect 24178 10240 29868 10296
rect 24117 10238 29868 10240
rect 24117 10235 24183 10238
rect 29862 10236 29868 10238
rect 29932 10236 29938 10300
rect 7966 10100 7972 10164
rect 8036 10162 8042 10164
rect 16757 10162 16823 10165
rect 8036 10160 16823 10162
rect 8036 10104 16762 10160
rect 16818 10104 16823 10160
rect 8036 10102 16823 10104
rect 8036 10100 8042 10102
rect 16757 10099 16823 10102
rect 17401 10162 17467 10165
rect 31710 10162 31770 10374
rect 32581 10371 32647 10374
rect 32397 10298 32463 10301
rect 33200 10298 34000 10328
rect 32397 10296 34000 10298
rect 32397 10240 32402 10296
rect 32458 10240 34000 10296
rect 32397 10238 34000 10240
rect 32397 10235 32463 10238
rect 33200 10208 34000 10238
rect 17401 10160 31770 10162
rect 17401 10104 17406 10160
rect 17462 10104 31770 10160
rect 17401 10102 31770 10104
rect 17401 10099 17467 10102
rect 8886 9964 8892 10028
rect 8956 10026 8962 10028
rect 9489 10026 9555 10029
rect 8956 10024 9555 10026
rect 8956 9968 9494 10024
rect 9550 9968 9555 10024
rect 8956 9966 9555 9968
rect 8956 9964 8962 9966
rect 9489 9963 9555 9966
rect 10225 10026 10291 10029
rect 10358 10026 10364 10028
rect 10225 10024 10364 10026
rect 10225 9968 10230 10024
rect 10286 9968 10364 10024
rect 10225 9966 10364 9968
rect 10225 9963 10291 9966
rect 10358 9964 10364 9966
rect 10428 9964 10434 10028
rect 11237 10026 11303 10029
rect 27153 10026 27219 10029
rect 11237 10024 27219 10026
rect 11237 9968 11242 10024
rect 11298 9968 27158 10024
rect 27214 9968 27219 10024
rect 11237 9966 27219 9968
rect 11237 9963 11303 9966
rect 27153 9963 27219 9966
rect 16389 9890 16455 9893
rect 7606 9888 16455 9890
rect 7606 9832 16394 9888
rect 16450 9832 16455 9888
rect 7606 9830 16455 9832
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 1964 9694 4722 9754
rect 1964 9692 1970 9694
rect 4429 9618 4495 9621
rect 5260 9618 5320 9830
rect 6545 9827 6611 9830
rect 16389 9827 16455 9830
rect 19241 9890 19307 9893
rect 24117 9890 24183 9893
rect 19241 9888 24183 9890
rect 19241 9832 19246 9888
rect 19302 9832 24122 9888
rect 24178 9832 24183 9888
rect 19241 9830 24183 9832
rect 19241 9827 19307 9830
rect 24117 9827 24183 9830
rect 25446 9828 25452 9892
rect 25516 9890 25522 9892
rect 25589 9890 25655 9893
rect 25516 9888 25655 9890
rect 25516 9832 25594 9888
rect 25650 9832 25655 9888
rect 25516 9830 25655 9832
rect 25516 9828 25522 9830
rect 25589 9827 25655 9830
rect 5809 9754 5875 9757
rect 6269 9754 6335 9757
rect 5809 9752 6335 9754
rect 5809 9696 5814 9752
rect 5870 9696 6274 9752
rect 6330 9696 6335 9752
rect 5809 9694 6335 9696
rect 5809 9691 5875 9694
rect 6269 9691 6335 9694
rect 6453 9754 6519 9757
rect 6453 9752 9690 9754
rect 6453 9696 6458 9752
rect 6514 9696 9690 9752
rect 6453 9694 9690 9696
rect 6453 9691 6519 9694
rect 4429 9616 5320 9618
rect 4429 9560 4434 9616
rect 4490 9560 5320 9616
rect 4429 9558 5320 9560
rect 4429 9555 4495 9558
rect 5574 9556 5580 9620
rect 5644 9618 5650 9620
rect 7465 9618 7531 9621
rect 8569 9618 8635 9621
rect 8937 9618 9003 9621
rect 5644 9616 7531 9618
rect 5644 9560 7470 9616
rect 7526 9560 7531 9616
rect 5644 9558 7531 9560
rect 5644 9556 5650 9558
rect 7465 9555 7531 9558
rect 7606 9616 9003 9618
rect 7606 9560 8574 9616
rect 8630 9560 8942 9616
rect 8998 9560 9003 9616
rect 7606 9558 9003 9560
rect 3877 9482 3943 9485
rect 7606 9482 7666 9558
rect 8569 9555 8635 9558
rect 8937 9555 9003 9558
rect 9121 9618 9187 9621
rect 9254 9618 9260 9620
rect 9121 9616 9260 9618
rect 9121 9560 9126 9616
rect 9182 9560 9260 9616
rect 9121 9558 9260 9560
rect 9121 9555 9187 9558
rect 9254 9556 9260 9558
rect 9324 9556 9330 9620
rect 9630 9618 9690 9694
rect 10542 9692 10548 9756
rect 10612 9754 10618 9756
rect 11237 9754 11303 9757
rect 10612 9752 11303 9754
rect 10612 9696 11242 9752
rect 11298 9696 11303 9752
rect 10612 9694 11303 9696
rect 10612 9692 10618 9694
rect 11237 9691 11303 9694
rect 12617 9754 12683 9757
rect 19425 9754 19491 9757
rect 19609 9756 19675 9757
rect 12617 9752 19491 9754
rect 12617 9696 12622 9752
rect 12678 9696 19430 9752
rect 19486 9696 19491 9752
rect 12617 9694 19491 9696
rect 12617 9691 12683 9694
rect 19425 9691 19491 9694
rect 19558 9692 19564 9756
rect 19628 9754 19675 9756
rect 24301 9754 24367 9757
rect 27654 9754 27660 9756
rect 19628 9752 19720 9754
rect 19670 9696 19720 9752
rect 19628 9694 19720 9696
rect 24301 9752 27660 9754
rect 24301 9696 24306 9752
rect 24362 9696 27660 9752
rect 24301 9694 27660 9696
rect 19628 9692 19675 9694
rect 19609 9691 19675 9692
rect 24301 9691 24367 9694
rect 27654 9692 27660 9694
rect 27724 9692 27730 9756
rect 15101 9618 15167 9621
rect 9630 9616 15167 9618
rect 9630 9560 15106 9616
rect 15162 9560 15167 9616
rect 9630 9558 15167 9560
rect 15101 9555 15167 9558
rect 15561 9618 15627 9621
rect 16665 9618 16731 9621
rect 15561 9616 16731 9618
rect 15561 9560 15566 9616
rect 15622 9560 16670 9616
rect 16726 9560 16731 9616
rect 15561 9558 16731 9560
rect 15561 9555 15627 9558
rect 16665 9555 16731 9558
rect 19333 9618 19399 9621
rect 20345 9618 20411 9621
rect 19333 9616 20411 9618
rect 19333 9560 19338 9616
rect 19394 9560 20350 9616
rect 20406 9560 20411 9616
rect 19333 9558 20411 9560
rect 19333 9555 19399 9558
rect 20345 9555 20411 9558
rect 20662 9556 20668 9620
rect 20732 9618 20738 9620
rect 32121 9618 32187 9621
rect 20732 9616 32187 9618
rect 20732 9560 32126 9616
rect 32182 9560 32187 9616
rect 20732 9558 32187 9560
rect 20732 9556 20738 9558
rect 32121 9555 32187 9558
rect 32305 9618 32371 9621
rect 33200 9618 34000 9648
rect 32305 9616 34000 9618
rect 32305 9560 32310 9616
rect 32366 9560 34000 9616
rect 32305 9558 34000 9560
rect 32305 9555 32371 9558
rect 33200 9528 34000 9558
rect 3877 9480 7666 9482
rect 3877 9424 3882 9480
rect 3938 9424 7666 9480
rect 3877 9422 7666 9424
rect 8753 9482 8819 9485
rect 8886 9482 8892 9484
rect 8753 9480 8892 9482
rect 8753 9424 8758 9480
rect 8814 9424 8892 9480
rect 8753 9422 8892 9424
rect 3877 9419 3943 9422
rect 8753 9419 8819 9422
rect 8886 9420 8892 9422
rect 8956 9420 8962 9484
rect 11973 9482 12039 9485
rect 9262 9480 12039 9482
rect 9262 9424 11978 9480
rect 12034 9424 12039 9480
rect 9262 9422 12039 9424
rect 4889 9346 4955 9349
rect 8477 9346 8543 9349
rect 4889 9344 8543 9346
rect 4889 9288 4894 9344
rect 4950 9288 8482 9344
rect 8538 9288 8543 9344
rect 4889 9286 8543 9288
rect 4889 9283 4955 9286
rect 8477 9283 8543 9286
rect 8845 9346 8911 9349
rect 9262 9346 9322 9422
rect 11973 9419 12039 9422
rect 12249 9482 12315 9485
rect 14273 9482 14339 9485
rect 12249 9480 14339 9482
rect 12249 9424 12254 9480
rect 12310 9424 14278 9480
rect 14334 9424 14339 9480
rect 12249 9422 14339 9424
rect 12249 9419 12315 9422
rect 14273 9419 14339 9422
rect 15469 9482 15535 9485
rect 16297 9482 16363 9485
rect 15469 9480 16363 9482
rect 15469 9424 15474 9480
rect 15530 9424 16302 9480
rect 16358 9424 16363 9480
rect 15469 9422 16363 9424
rect 15469 9419 15535 9422
rect 16297 9419 16363 9422
rect 18454 9420 18460 9484
rect 18524 9482 18530 9484
rect 18597 9482 18663 9485
rect 18524 9480 18663 9482
rect 18524 9424 18602 9480
rect 18658 9424 18663 9480
rect 18524 9422 18663 9424
rect 18524 9420 18530 9422
rect 18597 9419 18663 9422
rect 19190 9420 19196 9484
rect 19260 9482 19266 9484
rect 19517 9482 19583 9485
rect 19260 9480 19583 9482
rect 19260 9424 19522 9480
rect 19578 9424 19583 9480
rect 19260 9422 19583 9424
rect 19260 9420 19266 9422
rect 19517 9419 19583 9422
rect 21541 9482 21607 9485
rect 22277 9482 22343 9485
rect 21541 9480 22343 9482
rect 21541 9424 21546 9480
rect 21602 9424 22282 9480
rect 22338 9424 22343 9480
rect 21541 9422 22343 9424
rect 21541 9419 21607 9422
rect 22277 9419 22343 9422
rect 25262 9420 25268 9484
rect 25332 9482 25338 9484
rect 26785 9482 26851 9485
rect 25332 9480 26851 9482
rect 25332 9424 26790 9480
rect 26846 9424 26851 9480
rect 25332 9422 26851 9424
rect 25332 9420 25338 9422
rect 26785 9419 26851 9422
rect 8845 9344 9322 9346
rect 8845 9288 8850 9344
rect 8906 9288 9322 9344
rect 8845 9286 9322 9288
rect 9397 9346 9463 9349
rect 22553 9346 22619 9349
rect 9397 9344 22619 9346
rect 9397 9288 9402 9344
rect 9458 9288 22558 9344
rect 22614 9288 22619 9344
rect 9397 9286 22619 9288
rect 8845 9283 8911 9286
rect 9397 9283 9463 9286
rect 22553 9283 22619 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 6085 9210 6151 9213
rect 6637 9210 6703 9213
rect 6085 9208 6703 9210
rect 6085 9152 6090 9208
rect 6146 9152 6642 9208
rect 6698 9152 6703 9208
rect 6085 9150 6703 9152
rect 6085 9147 6151 9150
rect 6637 9147 6703 9150
rect 7465 9210 7531 9213
rect 11145 9210 11211 9213
rect 7465 9208 11211 9210
rect 7465 9152 7470 9208
rect 7526 9152 11150 9208
rect 11206 9152 11211 9208
rect 7465 9150 11211 9152
rect 7465 9147 7531 9150
rect 11145 9147 11211 9150
rect 11697 9210 11763 9213
rect 14273 9210 14339 9213
rect 11697 9208 14339 9210
rect 11697 9152 11702 9208
rect 11758 9152 14278 9208
rect 14334 9152 14339 9208
rect 11697 9150 14339 9152
rect 11697 9147 11763 9150
rect 14273 9147 14339 9150
rect 14549 9210 14615 9213
rect 14774 9210 14780 9212
rect 14549 9208 14780 9210
rect 14549 9152 14554 9208
rect 14610 9152 14780 9208
rect 14549 9150 14780 9152
rect 14549 9147 14615 9150
rect 14774 9148 14780 9150
rect 14844 9148 14850 9212
rect 14958 9148 14964 9212
rect 15028 9210 15034 9212
rect 20345 9210 20411 9213
rect 15028 9208 20411 9210
rect 15028 9152 20350 9208
rect 20406 9152 20411 9208
rect 15028 9150 20411 9152
rect 15028 9148 15034 9150
rect 20345 9147 20411 9150
rect 22277 9210 22343 9213
rect 25497 9210 25563 9213
rect 22277 9208 25563 9210
rect 22277 9152 22282 9208
rect 22338 9152 25502 9208
rect 25558 9152 25563 9208
rect 22277 9150 25563 9152
rect 22277 9147 22343 9150
rect 25497 9147 25563 9150
rect 2497 9074 2563 9077
rect 7414 9074 7420 9076
rect 2497 9072 7420 9074
rect 2497 9016 2502 9072
rect 2558 9016 7420 9072
rect 2497 9014 7420 9016
rect 2497 9011 2563 9014
rect 7414 9012 7420 9014
rect 7484 9012 7490 9076
rect 7598 9012 7604 9076
rect 7668 9074 7674 9076
rect 8753 9074 8819 9077
rect 7668 9072 8819 9074
rect 7668 9016 8758 9072
rect 8814 9016 8819 9072
rect 7668 9014 8819 9016
rect 7668 9012 7674 9014
rect 8753 9011 8819 9014
rect 9254 9012 9260 9076
rect 9324 9074 9330 9076
rect 16021 9074 16087 9077
rect 9324 9072 16087 9074
rect 9324 9016 16026 9072
rect 16082 9016 16087 9072
rect 9324 9014 16087 9016
rect 9324 9012 9330 9014
rect 16021 9011 16087 9014
rect 16297 9074 16363 9077
rect 25773 9074 25839 9077
rect 16297 9072 25839 9074
rect 16297 9016 16302 9072
rect 16358 9016 25778 9072
rect 25834 9016 25839 9072
rect 16297 9014 25839 9016
rect 16297 9011 16363 9014
rect 25773 9011 25839 9014
rect 26141 9074 26207 9077
rect 26601 9074 26667 9077
rect 26141 9072 26667 9074
rect 26141 9016 26146 9072
rect 26202 9016 26606 9072
rect 26662 9016 26667 9072
rect 26141 9014 26667 9016
rect 26141 9011 26207 9014
rect 26601 9011 26667 9014
rect 5073 8938 5139 8941
rect 7230 8938 7236 8940
rect 5073 8936 7236 8938
rect 5073 8880 5078 8936
rect 5134 8880 7236 8936
rect 5073 8878 7236 8880
rect 5073 8875 5139 8878
rect 7230 8876 7236 8878
rect 7300 8876 7306 8940
rect 8385 8938 8451 8941
rect 9397 8938 9463 8941
rect 13169 8938 13235 8941
rect 8385 8936 13235 8938
rect 8385 8880 8390 8936
rect 8446 8880 9402 8936
rect 9458 8880 13174 8936
rect 13230 8880 13235 8936
rect 8385 8878 13235 8880
rect 8385 8875 8451 8878
rect 9397 8875 9463 8878
rect 13169 8875 13235 8878
rect 14273 8938 14339 8941
rect 17125 8938 17191 8941
rect 17585 8938 17651 8941
rect 14273 8936 17651 8938
rect 14273 8880 14278 8936
rect 14334 8880 17130 8936
rect 17186 8880 17590 8936
rect 17646 8880 17651 8936
rect 14273 8878 17651 8880
rect 14273 8875 14339 8878
rect 17125 8875 17191 8878
rect 17585 8875 17651 8878
rect 17769 8938 17835 8941
rect 18689 8938 18755 8941
rect 17769 8936 18755 8938
rect 17769 8880 17774 8936
rect 17830 8880 18694 8936
rect 18750 8880 18755 8936
rect 17769 8878 18755 8880
rect 17769 8875 17835 8878
rect 18689 8875 18755 8878
rect 21582 8876 21588 8940
rect 21652 8938 21658 8940
rect 22001 8938 22067 8941
rect 21652 8936 22067 8938
rect 21652 8880 22006 8936
rect 22062 8880 22067 8936
rect 21652 8878 22067 8880
rect 21652 8876 21658 8878
rect 22001 8875 22067 8878
rect 5257 8802 5323 8805
rect 6637 8802 6703 8805
rect 5257 8800 6703 8802
rect 5257 8744 5262 8800
rect 5318 8744 6642 8800
rect 6698 8744 6703 8800
rect 5257 8742 6703 8744
rect 5257 8739 5323 8742
rect 6637 8739 6703 8742
rect 6862 8740 6868 8804
rect 6932 8802 6938 8804
rect 10041 8802 10107 8805
rect 6932 8800 10107 8802
rect 6932 8744 10046 8800
rect 10102 8744 10107 8800
rect 6932 8742 10107 8744
rect 6932 8740 6938 8742
rect 10041 8739 10107 8742
rect 11053 8802 11119 8805
rect 21449 8802 21515 8805
rect 11053 8800 21515 8802
rect 11053 8744 11058 8800
rect 11114 8744 21454 8800
rect 21510 8744 21515 8800
rect 11053 8742 21515 8744
rect 11053 8739 11119 8742
rect 21449 8739 21515 8742
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 6361 8666 6427 8669
rect 11697 8666 11763 8669
rect 6361 8664 11763 8666
rect 6361 8608 6366 8664
rect 6422 8608 11702 8664
rect 11758 8608 11763 8664
rect 6361 8606 11763 8608
rect 6361 8603 6427 8606
rect 11697 8603 11763 8606
rect 11973 8666 12039 8669
rect 12893 8666 12959 8669
rect 14089 8666 14155 8669
rect 11973 8664 12634 8666
rect 11973 8608 11978 8664
rect 12034 8608 12634 8664
rect 11973 8606 12634 8608
rect 11973 8603 12039 8606
rect 4654 8468 4660 8532
rect 4724 8530 4730 8532
rect 4797 8530 4863 8533
rect 4724 8528 4863 8530
rect 4724 8472 4802 8528
rect 4858 8472 4863 8528
rect 4724 8470 4863 8472
rect 4724 8468 4730 8470
rect 4797 8467 4863 8470
rect 4981 8530 5047 8533
rect 8753 8530 8819 8533
rect 9581 8530 9647 8533
rect 4981 8528 9647 8530
rect 4981 8472 4986 8528
rect 5042 8472 8758 8528
rect 8814 8472 9586 8528
rect 9642 8472 9647 8528
rect 4981 8470 9647 8472
rect 4981 8467 5047 8470
rect 8753 8467 8819 8470
rect 9581 8467 9647 8470
rect 9949 8530 10015 8533
rect 11053 8530 11119 8533
rect 9949 8528 11119 8530
rect 9949 8472 9954 8528
rect 10010 8472 11058 8528
rect 11114 8472 11119 8528
rect 9949 8470 11119 8472
rect 9949 8467 10015 8470
rect 11053 8467 11119 8470
rect 12014 8468 12020 8532
rect 12084 8530 12090 8532
rect 12249 8530 12315 8533
rect 12433 8530 12499 8533
rect 12084 8528 12499 8530
rect 12084 8472 12254 8528
rect 12310 8472 12438 8528
rect 12494 8472 12499 8528
rect 12084 8470 12499 8472
rect 12574 8530 12634 8606
rect 12893 8664 14155 8666
rect 12893 8608 12898 8664
rect 12954 8608 14094 8664
rect 14150 8608 14155 8664
rect 12893 8606 14155 8608
rect 12893 8603 12959 8606
rect 14089 8603 14155 8606
rect 15009 8666 15075 8669
rect 19885 8666 19951 8669
rect 15009 8664 19951 8666
rect 15009 8608 15014 8664
rect 15070 8608 19890 8664
rect 19946 8608 19951 8664
rect 15009 8606 19951 8608
rect 15009 8603 15075 8606
rect 19885 8603 19951 8606
rect 20345 8666 20411 8669
rect 23473 8666 23539 8669
rect 24761 8666 24827 8669
rect 20345 8664 24827 8666
rect 20345 8608 20350 8664
rect 20406 8608 23478 8664
rect 23534 8608 24766 8664
rect 24822 8608 24827 8664
rect 20345 8606 24827 8608
rect 20345 8603 20411 8606
rect 23473 8603 23539 8606
rect 24761 8603 24827 8606
rect 15009 8530 15075 8533
rect 12574 8528 15075 8530
rect 12574 8472 15014 8528
rect 15070 8472 15075 8528
rect 12574 8470 15075 8472
rect 12084 8468 12090 8470
rect 12249 8467 12315 8470
rect 12433 8467 12499 8470
rect 15009 8467 15075 8470
rect 15193 8530 15259 8533
rect 15326 8530 15332 8532
rect 15193 8528 15332 8530
rect 15193 8472 15198 8528
rect 15254 8472 15332 8528
rect 15193 8470 15332 8472
rect 15193 8467 15259 8470
rect 15326 8468 15332 8470
rect 15396 8468 15402 8532
rect 18045 8530 18111 8533
rect 18822 8530 18828 8532
rect 18045 8528 18828 8530
rect 18045 8472 18050 8528
rect 18106 8472 18828 8528
rect 18045 8470 18828 8472
rect 18045 8467 18111 8470
rect 18822 8468 18828 8470
rect 18892 8468 18898 8532
rect 19425 8530 19491 8533
rect 25773 8530 25839 8533
rect 19425 8528 25839 8530
rect 19425 8472 19430 8528
rect 19486 8472 25778 8528
rect 25834 8472 25839 8528
rect 19425 8470 25839 8472
rect 19425 8467 19491 8470
rect 25773 8467 25839 8470
rect 5441 8396 5507 8397
rect 5390 8394 5396 8396
rect 5350 8334 5396 8394
rect 5460 8392 5507 8396
rect 5502 8336 5507 8392
rect 5390 8332 5396 8334
rect 5460 8332 5507 8336
rect 5441 8331 5507 8332
rect 5809 8394 5875 8397
rect 5942 8394 5948 8396
rect 5809 8392 5948 8394
rect 5809 8336 5814 8392
rect 5870 8336 5948 8392
rect 5809 8334 5948 8336
rect 5809 8331 5875 8334
rect 5942 8332 5948 8334
rect 6012 8332 6018 8396
rect 6729 8394 6795 8397
rect 6862 8394 6868 8396
rect 6729 8392 6868 8394
rect 6729 8336 6734 8392
rect 6790 8336 6868 8392
rect 6729 8334 6868 8336
rect 6729 8331 6795 8334
rect 6862 8332 6868 8334
rect 6932 8332 6938 8396
rect 8109 8394 8175 8397
rect 9029 8394 9095 8397
rect 8109 8392 9095 8394
rect 8109 8336 8114 8392
rect 8170 8336 9034 8392
rect 9090 8336 9095 8392
rect 8109 8334 9095 8336
rect 8109 8331 8175 8334
rect 9029 8331 9095 8334
rect 11421 8394 11487 8397
rect 14549 8394 14615 8397
rect 15009 8394 15075 8397
rect 11421 8392 15075 8394
rect 11421 8336 11426 8392
rect 11482 8336 14554 8392
rect 14610 8336 15014 8392
rect 15070 8336 15075 8392
rect 11421 8334 15075 8336
rect 11421 8331 11487 8334
rect 14549 8331 14615 8334
rect 15009 8331 15075 8334
rect 15377 8394 15443 8397
rect 24577 8394 24643 8397
rect 15377 8392 24643 8394
rect 15377 8336 15382 8392
rect 15438 8336 24582 8392
rect 24638 8336 24643 8392
rect 15377 8334 24643 8336
rect 15377 8331 15443 8334
rect 24577 8331 24643 8334
rect 4613 8258 4679 8261
rect 6085 8258 6151 8261
rect 8201 8258 8267 8261
rect 4613 8256 8267 8258
rect 4613 8200 4618 8256
rect 4674 8200 6090 8256
rect 6146 8200 8206 8256
rect 8262 8200 8267 8256
rect 4613 8198 8267 8200
rect 4613 8195 4679 8198
rect 6085 8195 6151 8198
rect 8201 8195 8267 8198
rect 8385 8258 8451 8261
rect 9213 8258 9279 8261
rect 8385 8256 9279 8258
rect 8385 8200 8390 8256
rect 8446 8200 9218 8256
rect 9274 8200 9279 8256
rect 8385 8198 9279 8200
rect 8385 8195 8451 8198
rect 9213 8195 9279 8198
rect 12801 8258 12867 8261
rect 15377 8258 15443 8261
rect 12801 8256 15443 8258
rect 12801 8200 12806 8256
rect 12862 8200 15382 8256
rect 15438 8200 15443 8256
rect 12801 8198 15443 8200
rect 12801 8195 12867 8198
rect 15377 8195 15443 8198
rect 15929 8258 15995 8261
rect 23606 8258 23612 8260
rect 15929 8256 23612 8258
rect 15929 8200 15934 8256
rect 15990 8200 23612 8256
rect 15929 8198 23612 8200
rect 15929 8195 15995 8198
rect 23606 8196 23612 8198
rect 23676 8258 23682 8260
rect 23749 8258 23815 8261
rect 23676 8256 23815 8258
rect 23676 8200 23754 8256
rect 23810 8200 23815 8256
rect 23676 8198 23815 8200
rect 23676 8196 23682 8198
rect 23749 8195 23815 8198
rect 32397 8258 32463 8261
rect 33200 8258 34000 8288
rect 32397 8256 34000 8258
rect 32397 8200 32402 8256
rect 32458 8200 34000 8256
rect 32397 8198 34000 8200
rect 32397 8195 32463 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 33200 8168 34000 8198
rect 4210 8127 4526 8128
rect 11973 8122 12039 8125
rect 22829 8122 22895 8125
rect 11973 8120 22895 8122
rect 11973 8064 11978 8120
rect 12034 8064 22834 8120
rect 22890 8064 22895 8120
rect 11973 8062 22895 8064
rect 11973 8059 12039 8062
rect 22829 8059 22895 8062
rect 23105 8122 23171 8125
rect 31150 8122 31156 8124
rect 23105 8120 31156 8122
rect 23105 8064 23110 8120
rect 23166 8064 31156 8120
rect 23105 8062 31156 8064
rect 23105 8059 23171 8062
rect 31150 8060 31156 8062
rect 31220 8060 31226 8124
rect 381 7986 447 7989
rect 14549 7986 14615 7989
rect 381 7984 14615 7986
rect 381 7928 386 7984
rect 442 7928 14554 7984
rect 14610 7928 14615 7984
rect 381 7926 14615 7928
rect 381 7923 447 7926
rect 14549 7923 14615 7926
rect 15653 7986 15719 7989
rect 28809 7986 28875 7989
rect 15653 7984 28875 7986
rect 15653 7928 15658 7984
rect 15714 7928 28814 7984
rect 28870 7928 28875 7984
rect 15653 7926 28875 7928
rect 15653 7923 15719 7926
rect 28809 7923 28875 7926
rect 9070 7788 9076 7852
rect 9140 7850 9146 7852
rect 18781 7850 18847 7853
rect 9140 7848 18847 7850
rect 9140 7792 18786 7848
rect 18842 7792 18847 7848
rect 9140 7790 18847 7792
rect 9140 7788 9146 7790
rect 18781 7787 18847 7790
rect 12750 7652 12756 7716
rect 12820 7714 12826 7716
rect 20989 7714 21055 7717
rect 12820 7712 21055 7714
rect 12820 7656 20994 7712
rect 21050 7656 21055 7712
rect 12820 7654 21055 7656
rect 12820 7652 12826 7654
rect 20989 7651 21055 7654
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 8201 7578 8267 7581
rect 9489 7578 9555 7581
rect 8201 7576 9555 7578
rect 8201 7520 8206 7576
rect 8262 7520 9494 7576
rect 9550 7520 9555 7576
rect 8201 7518 9555 7520
rect 8201 7515 8267 7518
rect 9489 7515 9555 7518
rect 13353 7578 13419 7581
rect 13486 7578 13492 7580
rect 13353 7576 13492 7578
rect 13353 7520 13358 7576
rect 13414 7520 13492 7576
rect 13353 7518 13492 7520
rect 13353 7515 13419 7518
rect 13486 7516 13492 7518
rect 13556 7516 13562 7580
rect 13629 7578 13695 7581
rect 16665 7578 16731 7581
rect 30281 7578 30347 7581
rect 13629 7576 16731 7578
rect 13629 7520 13634 7576
rect 13690 7520 16670 7576
rect 16726 7520 16731 7576
rect 13629 7518 16731 7520
rect 13629 7515 13695 7518
rect 16665 7515 16731 7518
rect 22050 7576 30347 7578
rect 22050 7520 30286 7576
rect 30342 7520 30347 7576
rect 22050 7518 30347 7520
rect 3785 7442 3851 7445
rect 4245 7442 4311 7445
rect 4981 7442 5047 7445
rect 3785 7440 5047 7442
rect 3785 7384 3790 7440
rect 3846 7384 4250 7440
rect 4306 7384 4986 7440
rect 5042 7384 5047 7440
rect 3785 7382 5047 7384
rect 3785 7379 3851 7382
rect 4245 7379 4311 7382
rect 4981 7379 5047 7382
rect 12617 7442 12683 7445
rect 15510 7442 15516 7444
rect 12617 7440 15516 7442
rect 12617 7384 12622 7440
rect 12678 7384 15516 7440
rect 12617 7382 15516 7384
rect 12617 7379 12683 7382
rect 15510 7380 15516 7382
rect 15580 7380 15586 7444
rect 19333 7442 19399 7445
rect 22050 7442 22110 7518
rect 30281 7515 30347 7518
rect 31661 7578 31727 7581
rect 33200 7578 34000 7608
rect 31661 7576 34000 7578
rect 31661 7520 31666 7576
rect 31722 7520 34000 7576
rect 31661 7518 34000 7520
rect 31661 7515 31727 7518
rect 33200 7488 34000 7518
rect 19333 7440 22110 7442
rect 19333 7384 19338 7440
rect 19394 7384 22110 7440
rect 19333 7382 22110 7384
rect 19333 7379 19399 7382
rect 23238 7380 23244 7444
rect 23308 7442 23314 7444
rect 23381 7442 23447 7445
rect 23308 7440 23447 7442
rect 23308 7384 23386 7440
rect 23442 7384 23447 7440
rect 23308 7382 23447 7384
rect 23308 7380 23314 7382
rect 23381 7379 23447 7382
rect 24117 7442 24183 7445
rect 24526 7442 24532 7444
rect 24117 7440 24532 7442
rect 24117 7384 24122 7440
rect 24178 7384 24532 7440
rect 24117 7382 24532 7384
rect 24117 7379 24183 7382
rect 24526 7380 24532 7382
rect 24596 7380 24602 7444
rect 7230 7244 7236 7308
rect 7300 7306 7306 7308
rect 16849 7306 16915 7309
rect 7300 7304 16915 7306
rect 7300 7248 16854 7304
rect 16910 7248 16915 7304
rect 7300 7246 16915 7248
rect 7300 7244 7306 7246
rect 16849 7243 16915 7246
rect 17217 7306 17283 7309
rect 27797 7306 27863 7309
rect 17217 7304 27863 7306
rect 17217 7248 17222 7304
rect 17278 7248 27802 7304
rect 27858 7248 27863 7304
rect 17217 7246 27863 7248
rect 17217 7243 17283 7246
rect 27797 7243 27863 7246
rect 11094 7108 11100 7172
rect 11164 7170 11170 7172
rect 11513 7170 11579 7173
rect 11164 7168 11579 7170
rect 11164 7112 11518 7168
rect 11574 7112 11579 7168
rect 11164 7110 11579 7112
rect 11164 7108 11170 7110
rect 11513 7107 11579 7110
rect 12617 7170 12683 7173
rect 14089 7170 14155 7173
rect 12617 7168 14155 7170
rect 12617 7112 12622 7168
rect 12678 7112 14094 7168
rect 14150 7112 14155 7168
rect 12617 7110 14155 7112
rect 12617 7107 12683 7110
rect 14089 7107 14155 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 8150 6972 8156 7036
rect 8220 7034 8226 7036
rect 18638 7034 18644 7036
rect 8220 6974 18644 7034
rect 8220 6972 8226 6974
rect 18638 6972 18644 6974
rect 18708 6972 18714 7036
rect 8702 6836 8708 6900
rect 8772 6898 8778 6900
rect 9305 6898 9371 6901
rect 8772 6896 9371 6898
rect 8772 6840 9310 6896
rect 9366 6840 9371 6896
rect 8772 6838 9371 6840
rect 8772 6836 8778 6838
rect 9305 6835 9371 6838
rect 9489 6898 9555 6901
rect 9806 6898 9812 6900
rect 9489 6896 9812 6898
rect 9489 6840 9494 6896
rect 9550 6840 9812 6896
rect 9489 6838 9812 6840
rect 9489 6835 9555 6838
rect 9806 6836 9812 6838
rect 9876 6836 9882 6900
rect 12709 6898 12775 6901
rect 15193 6898 15259 6901
rect 12709 6896 15259 6898
rect 12709 6840 12714 6896
rect 12770 6840 15198 6896
rect 15254 6840 15259 6896
rect 12709 6838 15259 6840
rect 12709 6835 12775 6838
rect 15193 6835 15259 6838
rect 17769 6898 17835 6901
rect 20253 6898 20319 6901
rect 29085 6898 29151 6901
rect 17769 6896 29151 6898
rect 17769 6840 17774 6896
rect 17830 6840 20258 6896
rect 20314 6840 29090 6896
rect 29146 6840 29151 6896
rect 17769 6838 29151 6840
rect 17769 6835 17835 6838
rect 20253 6835 20319 6838
rect 29085 6835 29151 6838
rect 32305 6898 32371 6901
rect 33200 6898 34000 6928
rect 32305 6896 34000 6898
rect 32305 6840 32310 6896
rect 32366 6840 34000 6896
rect 32305 6838 34000 6840
rect 32305 6835 32371 6838
rect 33200 6808 34000 6838
rect 3550 6700 3556 6764
rect 3620 6762 3626 6764
rect 8201 6762 8267 6765
rect 13629 6762 13695 6765
rect 14038 6762 14044 6764
rect 3620 6702 5320 6762
rect 3620 6700 3626 6702
rect 5260 6626 5320 6702
rect 8201 6760 14044 6762
rect 8201 6704 8206 6760
rect 8262 6704 13634 6760
rect 13690 6704 14044 6760
rect 8201 6702 14044 6704
rect 8201 6699 8267 6702
rect 13629 6699 13695 6702
rect 14038 6700 14044 6702
rect 14108 6700 14114 6764
rect 20529 6762 20595 6765
rect 22921 6762 22987 6765
rect 20529 6760 22987 6762
rect 20529 6704 20534 6760
rect 20590 6704 22926 6760
rect 22982 6704 22987 6760
rect 20529 6702 22987 6704
rect 20529 6699 20595 6702
rect 22921 6699 22987 6702
rect 10777 6626 10843 6629
rect 5260 6624 10843 6626
rect 5260 6568 10782 6624
rect 10838 6568 10843 6624
rect 5260 6566 10843 6568
rect 10777 6563 10843 6566
rect 11145 6626 11211 6629
rect 11789 6626 11855 6629
rect 17217 6626 17283 6629
rect 21214 6626 21220 6628
rect 11145 6624 17283 6626
rect 11145 6568 11150 6624
rect 11206 6568 11794 6624
rect 11850 6568 17222 6624
rect 17278 6568 17283 6624
rect 11145 6566 17283 6568
rect 11145 6563 11211 6566
rect 11789 6563 11855 6566
rect 17217 6563 17283 6566
rect 17358 6566 21220 6626
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 7414 6428 7420 6492
rect 7484 6490 7490 6492
rect 17358 6490 17418 6566
rect 21214 6564 21220 6566
rect 21284 6564 21290 6628
rect 7484 6430 17418 6490
rect 17585 6490 17651 6493
rect 20529 6490 20595 6493
rect 20662 6490 20668 6492
rect 17585 6488 20668 6490
rect 17585 6432 17590 6488
rect 17646 6432 20534 6488
rect 20590 6432 20668 6488
rect 17585 6430 20668 6432
rect 7484 6428 7490 6430
rect 17585 6427 17651 6430
rect 20529 6427 20595 6430
rect 20662 6428 20668 6430
rect 20732 6428 20738 6492
rect 6913 6354 6979 6357
rect 7373 6354 7439 6357
rect 15878 6354 15884 6356
rect 6913 6352 15884 6354
rect 6913 6296 6918 6352
rect 6974 6296 7378 6352
rect 7434 6296 15884 6352
rect 6913 6294 15884 6296
rect 6913 6291 6979 6294
rect 7373 6291 7439 6294
rect 15878 6292 15884 6294
rect 15948 6292 15954 6356
rect 18413 6354 18479 6357
rect 25957 6354 26023 6357
rect 18413 6352 26023 6354
rect 18413 6296 18418 6352
rect 18474 6296 25962 6352
rect 26018 6296 26023 6352
rect 18413 6294 26023 6296
rect 18413 6291 18479 6294
rect 25957 6291 26023 6294
rect 2078 6156 2084 6220
rect 2148 6218 2154 6220
rect 11053 6218 11119 6221
rect 12198 6218 12204 6220
rect 2148 6158 10978 6218
rect 2148 6156 2154 6158
rect 7097 6082 7163 6085
rect 8886 6082 8892 6084
rect 7097 6080 8892 6082
rect 7097 6024 7102 6080
rect 7158 6024 8892 6080
rect 7097 6022 8892 6024
rect 7097 6019 7163 6022
rect 8886 6020 8892 6022
rect 8956 6082 8962 6084
rect 9305 6082 9371 6085
rect 8956 6080 9371 6082
rect 8956 6024 9310 6080
rect 9366 6024 9371 6080
rect 8956 6022 9371 6024
rect 10918 6082 10978 6158
rect 11053 6216 12204 6218
rect 11053 6160 11058 6216
rect 11114 6160 12204 6216
rect 11053 6158 12204 6160
rect 11053 6155 11119 6158
rect 12198 6156 12204 6158
rect 12268 6218 12274 6220
rect 23197 6218 23263 6221
rect 25681 6220 25747 6221
rect 12268 6216 23263 6218
rect 12268 6160 23202 6216
rect 23258 6160 23263 6216
rect 12268 6158 23263 6160
rect 12268 6156 12274 6158
rect 23197 6155 23263 6158
rect 25630 6156 25636 6220
rect 25700 6218 25747 6220
rect 25700 6216 25792 6218
rect 25742 6160 25792 6216
rect 25700 6158 25792 6160
rect 25700 6156 25747 6158
rect 25681 6155 25747 6156
rect 11973 6082 12039 6085
rect 10918 6080 12039 6082
rect 10918 6024 11978 6080
rect 12034 6024 12039 6080
rect 10918 6022 12039 6024
rect 8956 6020 8962 6022
rect 9305 6019 9371 6022
rect 11973 6019 12039 6022
rect 17769 6082 17835 6085
rect 22870 6082 22876 6084
rect 17769 6080 22876 6082
rect 17769 6024 17774 6080
rect 17830 6024 22876 6080
rect 17769 6022 22876 6024
rect 17769 6019 17835 6022
rect 22870 6020 22876 6022
rect 22940 6020 22946 6084
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 11237 5946 11303 5949
rect 18413 5946 18479 5949
rect 11237 5944 18479 5946
rect 11237 5888 11242 5944
rect 11298 5888 18418 5944
rect 18474 5888 18479 5944
rect 11237 5886 18479 5888
rect 11237 5883 11303 5886
rect 18413 5883 18479 5886
rect 11329 5810 11395 5813
rect 17953 5810 18019 5813
rect 11329 5808 18019 5810
rect 11329 5752 11334 5808
rect 11390 5752 17958 5808
rect 18014 5752 18019 5808
rect 11329 5750 18019 5752
rect 11329 5747 11395 5750
rect 17953 5747 18019 5750
rect 2313 5674 2379 5677
rect 11145 5674 11211 5677
rect 2313 5672 11211 5674
rect 2313 5616 2318 5672
rect 2374 5616 11150 5672
rect 11206 5616 11211 5672
rect 2313 5614 11211 5616
rect 2313 5611 2379 5614
rect 11145 5611 11211 5614
rect 17033 5674 17099 5677
rect 19517 5674 19583 5677
rect 17033 5672 19583 5674
rect 17033 5616 17038 5672
rect 17094 5616 19522 5672
rect 19578 5616 19583 5672
rect 17033 5614 19583 5616
rect 17033 5611 17099 5614
rect 19517 5611 19583 5614
rect 20713 5674 20779 5677
rect 21357 5674 21423 5677
rect 23473 5674 23539 5677
rect 20713 5672 23539 5674
rect 20713 5616 20718 5672
rect 20774 5616 21362 5672
rect 21418 5616 23478 5672
rect 23534 5616 23539 5672
rect 20713 5614 23539 5616
rect 20713 5611 20779 5614
rect 21357 5611 21423 5614
rect 23473 5611 23539 5614
rect 12157 5538 12223 5541
rect 32673 5538 32739 5541
rect 12157 5536 32739 5538
rect 12157 5480 12162 5536
rect 12218 5480 32678 5536
rect 32734 5480 32739 5536
rect 12157 5478 32739 5480
rect 12157 5475 12223 5478
rect 32673 5475 32739 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 13721 5402 13787 5405
rect 22737 5402 22803 5405
rect 13721 5400 22803 5402
rect 13721 5344 13726 5400
rect 13782 5344 22742 5400
rect 22798 5344 22803 5400
rect 13721 5342 22803 5344
rect 13721 5339 13787 5342
rect 22737 5339 22803 5342
rect 24577 5402 24643 5405
rect 30966 5402 30972 5404
rect 24577 5400 30972 5402
rect 24577 5344 24582 5400
rect 24638 5344 30972 5400
rect 24577 5342 30972 5344
rect 24577 5339 24643 5342
rect 30966 5340 30972 5342
rect 31036 5340 31042 5404
rect 9990 5204 9996 5268
rect 10060 5266 10066 5268
rect 14365 5266 14431 5269
rect 23197 5266 23263 5269
rect 26550 5266 26556 5268
rect 10060 5264 14431 5266
rect 10060 5208 14370 5264
rect 14426 5208 14431 5264
rect 10060 5206 14431 5208
rect 10060 5204 10066 5206
rect 14365 5203 14431 5206
rect 22050 5264 26556 5266
rect 22050 5208 23202 5264
rect 23258 5208 26556 5264
rect 22050 5206 26556 5208
rect 2037 5130 2103 5133
rect 22050 5130 22110 5206
rect 23197 5203 23263 5206
rect 26550 5204 26556 5206
rect 26620 5204 26626 5268
rect 2037 5128 22110 5130
rect 2037 5072 2042 5128
rect 2098 5072 22110 5128
rect 2037 5070 22110 5072
rect 2037 5067 2103 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 12617 4722 12683 4725
rect 23238 4722 23244 4724
rect 12617 4720 23244 4722
rect 12617 4664 12622 4720
rect 12678 4664 23244 4720
rect 12617 4662 23244 4664
rect 12617 4659 12683 4662
rect 23238 4660 23244 4662
rect 23308 4660 23314 4724
rect 9949 4586 10015 4589
rect 20713 4586 20779 4589
rect 9949 4584 20779 4586
rect 9949 4528 9954 4584
rect 10010 4528 20718 4584
rect 20774 4528 20779 4584
rect 9949 4526 20779 4528
rect 9949 4523 10015 4526
rect 20713 4523 20779 4526
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 15837 4042 15903 4045
rect 29126 4042 29132 4044
rect 15837 4040 29132 4042
rect 15837 3984 15842 4040
rect 15898 3984 29132 4040
rect 15837 3982 29132 3984
rect 15837 3979 15903 3982
rect 29126 3980 29132 3982
rect 29196 3980 29202 4044
rect 13670 3844 13676 3908
rect 13740 3906 13746 3908
rect 22829 3906 22895 3909
rect 13740 3904 22895 3906
rect 13740 3848 22834 3904
rect 22890 3848 22895 3904
rect 13740 3846 22895 3848
rect 13740 3844 13746 3846
rect 22829 3843 22895 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 12893 3770 12959 3773
rect 26182 3770 26188 3772
rect 12893 3768 26188 3770
rect 12893 3712 12898 3768
rect 12954 3712 26188 3768
rect 12893 3710 26188 3712
rect 12893 3707 12959 3710
rect 26182 3708 26188 3710
rect 26252 3708 26258 3772
rect 15101 3634 15167 3637
rect 25814 3634 25820 3636
rect 15101 3632 25820 3634
rect 15101 3576 15106 3632
rect 15162 3576 25820 3632
rect 15101 3574 25820 3576
rect 15101 3571 15167 3574
rect 25814 3572 25820 3574
rect 25884 3572 25890 3636
rect 5758 3436 5764 3500
rect 5828 3498 5834 3500
rect 24025 3498 24091 3501
rect 5828 3496 24091 3498
rect 5828 3440 24030 3496
rect 24086 3440 24091 3496
rect 5828 3438 24091 3440
rect 5828 3436 5834 3438
rect 24025 3435 24091 3438
rect 13537 3362 13603 3365
rect 30414 3362 30420 3364
rect 13537 3360 30420 3362
rect 13537 3304 13542 3360
rect 13598 3304 30420 3360
rect 13537 3302 30420 3304
rect 13537 3299 13603 3302
rect 30414 3300 30420 3302
rect 30484 3300 30490 3364
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 9438 3164 9444 3228
rect 9508 3226 9514 3228
rect 17401 3226 17467 3229
rect 9508 3224 17467 3226
rect 9508 3168 17406 3224
rect 17462 3168 17467 3224
rect 9508 3166 17467 3168
rect 9508 3164 9514 3166
rect 17401 3163 17467 3166
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 10869 2682 10935 2685
rect 21030 2682 21036 2684
rect 10869 2680 21036 2682
rect 10869 2624 10874 2680
rect 10930 2624 21036 2680
rect 10869 2622 21036 2624
rect 10869 2619 10935 2622
rect 21030 2620 21036 2622
rect 21100 2620 21106 2684
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 980 31316 1044 31380
rect 20668 31316 20732 31380
rect 2084 31180 2148 31244
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 14412 30908 14476 30972
rect 30420 30772 30484 30836
rect 30604 30500 30668 30564
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 17908 30364 17972 30428
rect 612 30092 676 30156
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 2636 29684 2700 29748
rect 1164 29548 1228 29612
rect 5396 29412 5460 29476
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 29316 29276 29380 29340
rect 2452 29140 2516 29204
rect 8156 29004 8220 29068
rect 18276 29004 18340 29068
rect 6316 28868 6380 28932
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 12940 28732 13004 28796
rect 7420 28596 7484 28660
rect 3372 28384 3436 28388
rect 3372 28328 3386 28384
rect 3386 28328 3436 28384
rect 3372 28324 3436 28328
rect 6500 28324 6564 28388
rect 10180 28384 10244 28388
rect 10180 28328 10194 28384
rect 10194 28328 10244 28384
rect 10180 28324 10244 28328
rect 21036 28324 21100 28388
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 11100 28188 11164 28252
rect 13492 28188 13556 28252
rect 4660 28112 4724 28116
rect 4660 28056 4674 28112
rect 4674 28056 4724 28112
rect 4660 28052 4724 28056
rect 6868 27916 6932 27980
rect 9444 27780 9508 27844
rect 11284 27780 11348 27844
rect 12756 27780 12820 27844
rect 27844 27780 27908 27844
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 12572 27644 12636 27708
rect 15148 27704 15212 27708
rect 15148 27648 15198 27704
rect 15198 27648 15212 27704
rect 15148 27644 15212 27648
rect 16068 27704 16132 27708
rect 16068 27648 16082 27704
rect 16082 27648 16132 27704
rect 16068 27644 16132 27648
rect 20484 27644 20548 27708
rect 19380 27508 19444 27572
rect 22508 27508 22572 27572
rect 23428 27644 23492 27708
rect 24532 27508 24596 27572
rect 7236 27432 7300 27436
rect 7236 27376 7250 27432
rect 7250 27376 7300 27432
rect 7236 27372 7300 27376
rect 19932 27372 19996 27436
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 7052 27296 7116 27300
rect 7052 27240 7066 27296
rect 7066 27240 7116 27296
rect 7052 27236 7116 27240
rect 7972 27296 8036 27300
rect 7972 27240 7986 27296
rect 7986 27240 8036 27296
rect 7972 27236 8036 27240
rect 18828 27236 18892 27300
rect 6132 26964 6196 27028
rect 9260 26828 9324 26892
rect 19012 26964 19076 27028
rect 12756 26828 12820 26892
rect 18828 26828 18892 26892
rect 21404 26828 21468 26892
rect 19564 26692 19628 26756
rect 29868 26964 29932 27028
rect 30788 26692 30852 26756
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 13308 26556 13372 26620
rect 5580 26480 5644 26484
rect 5580 26424 5594 26480
rect 5594 26424 5644 26480
rect 5580 26420 5644 26424
rect 5948 26420 6012 26484
rect 26924 26480 26988 26484
rect 26924 26424 26974 26480
rect 26974 26424 26988 26480
rect 26924 26420 26988 26424
rect 17724 26344 17788 26348
rect 17724 26288 17774 26344
rect 17774 26288 17788 26344
rect 17724 26284 17788 26288
rect 8708 26148 8772 26212
rect 10180 26148 10244 26212
rect 21220 26344 21284 26348
rect 21220 26288 21234 26344
rect 21234 26288 21284 26344
rect 21220 26284 21284 26288
rect 24900 26284 24964 26348
rect 26188 26148 26252 26212
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 19380 25876 19444 25940
rect 19748 25876 19812 25940
rect 25820 25876 25884 25940
rect 21772 25740 21836 25804
rect 5764 25604 5828 25668
rect 7236 25604 7300 25668
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 19380 25604 19444 25668
rect 12388 25468 12452 25532
rect 28948 25468 29012 25532
rect 13676 25392 13740 25396
rect 13676 25336 13726 25392
rect 13726 25336 13740 25392
rect 13676 25332 13740 25336
rect 16988 25332 17052 25396
rect 10548 25196 10612 25260
rect 26372 25196 26436 25260
rect 16620 25060 16684 25124
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 9444 24924 9508 24988
rect 11100 24924 11164 24988
rect 15884 24924 15948 24988
rect 3740 24788 3804 24852
rect 9812 24788 9876 24852
rect 20668 24924 20732 24988
rect 20852 24924 20916 24988
rect 28580 24924 28644 24988
rect 19564 24652 19628 24716
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 20668 24516 20732 24580
rect 7420 24244 7484 24308
rect 13124 24244 13188 24308
rect 20852 24244 20916 24308
rect 6316 23972 6380 24036
rect 10916 23972 10980 24036
rect 13308 23972 13372 24036
rect 16804 23972 16868 24036
rect 20852 24108 20916 24172
rect 28396 23972 28460 24036
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 11468 23564 11532 23628
rect 4660 23428 4724 23492
rect 6500 23428 6564 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 11100 23292 11164 23356
rect 12388 23292 12452 23356
rect 14596 23488 14660 23492
rect 14596 23432 14610 23488
rect 14610 23432 14660 23488
rect 14596 23428 14660 23432
rect 17908 23488 17972 23492
rect 17908 23432 17958 23488
rect 17958 23432 17972 23488
rect 17908 23428 17972 23432
rect 21956 23428 22020 23492
rect 22140 23428 22204 23492
rect 23980 23428 24044 23492
rect 28212 23488 28276 23492
rect 28212 23432 28226 23488
rect 28226 23432 28276 23488
rect 28212 23428 28276 23432
rect 4660 23020 4724 23084
rect 7420 23156 7484 23220
rect 5396 23020 5460 23084
rect 5764 23020 5828 23084
rect 11284 23156 11348 23220
rect 22876 23156 22940 23220
rect 8524 22884 8588 22948
rect 19564 23020 19628 23084
rect 19380 22944 19444 22948
rect 19380 22888 19394 22944
rect 19394 22888 19444 22944
rect 19380 22884 19444 22888
rect 20116 22944 20180 22948
rect 20116 22888 20166 22944
rect 20166 22888 20180 22944
rect 20116 22884 20180 22888
rect 25268 22884 25332 22948
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 20300 22748 20364 22812
rect 20668 22748 20732 22812
rect 18460 22612 18524 22676
rect 25084 22340 25148 22404
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 6500 22264 6564 22268
rect 6500 22208 6550 22264
rect 6550 22208 6564 22264
rect 6500 22204 6564 22208
rect 12020 22204 12084 22268
rect 12204 22204 12268 22268
rect 20300 22204 20364 22268
rect 24716 22204 24780 22268
rect 5580 22068 5644 22132
rect 6132 22068 6196 22132
rect 6868 22068 6932 22132
rect 19748 22068 19812 22132
rect 21404 22068 21468 22132
rect 3556 21796 3620 21860
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 2268 21660 2332 21724
rect 5580 21992 5644 21996
rect 5580 21936 5594 21992
rect 5594 21936 5644 21992
rect 5580 21932 5644 21936
rect 12388 21932 12452 21996
rect 13492 21932 13556 21996
rect 25820 21932 25884 21996
rect 14228 21796 14292 21860
rect 22692 21796 22756 21860
rect 10732 21524 10796 21588
rect 13308 21660 13372 21724
rect 13492 21660 13556 21724
rect 14044 21660 14108 21724
rect 22876 21660 22940 21724
rect 23428 21660 23492 21724
rect 24348 21660 24412 21724
rect 18092 21524 18156 21588
rect 20300 21524 20364 21588
rect 20484 21524 20548 21588
rect 23428 21524 23492 21588
rect 5396 21448 5460 21452
rect 5396 21392 5410 21448
rect 5410 21392 5460 21448
rect 5396 21388 5460 21392
rect 9996 21388 10060 21452
rect 12388 21448 12452 21452
rect 12388 21392 12438 21448
rect 12438 21392 12452 21448
rect 5764 21252 5828 21316
rect 7420 21252 7484 21316
rect 12388 21388 12452 21392
rect 12756 21388 12820 21452
rect 12940 21448 13004 21452
rect 12940 21392 12954 21448
rect 12954 21392 13004 21448
rect 12940 21388 13004 21392
rect 13492 21252 13556 21316
rect 19932 21448 19996 21452
rect 19932 21392 19982 21448
rect 19982 21392 19996 21448
rect 19932 21388 19996 21392
rect 20852 21388 20916 21452
rect 22140 21252 22204 21316
rect 31156 21252 31220 21316
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 14780 21116 14844 21180
rect 23060 21116 23124 21180
rect 17908 20980 17972 21044
rect 19564 21040 19628 21044
rect 19564 20984 19578 21040
rect 19578 20984 19628 21040
rect 19564 20980 19628 20984
rect 21588 21040 21652 21044
rect 21588 20984 21638 21040
rect 21638 20984 21652 21040
rect 21588 20980 21652 20984
rect 796 20708 860 20772
rect 3924 20708 3988 20772
rect 7052 20708 7116 20772
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 13676 20844 13740 20908
rect 14044 20904 14108 20908
rect 14044 20848 14058 20904
rect 14058 20848 14108 20904
rect 14044 20844 14108 20848
rect 15516 20844 15580 20908
rect 8708 20572 8772 20636
rect 12940 20708 13004 20772
rect 18092 20708 18156 20772
rect 20668 20708 20732 20772
rect 25452 20708 25516 20772
rect 26556 20708 26620 20772
rect 30420 20436 30484 20500
rect 3188 20300 3252 20364
rect 12204 20300 12268 20364
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 1900 19892 1964 19956
rect 5948 19756 6012 19820
rect 2268 19620 2332 19684
rect 3372 19620 3436 19684
rect 11836 20224 11900 20228
rect 11836 20168 11850 20224
rect 11850 20168 11900 20224
rect 11836 20164 11900 20168
rect 12204 20164 12268 20228
rect 18092 20028 18156 20092
rect 19380 20028 19444 20092
rect 24900 20028 24964 20092
rect 11652 19952 11716 19956
rect 11652 19896 11666 19952
rect 11666 19896 11716 19952
rect 11652 19892 11716 19896
rect 13676 19892 13740 19956
rect 21772 19892 21836 19956
rect 26004 19952 26068 19956
rect 26004 19896 26054 19952
rect 26054 19896 26068 19952
rect 26004 19892 26068 19896
rect 25268 19756 25332 19820
rect 25820 19816 25884 19820
rect 25820 19760 25834 19816
rect 25834 19760 25884 19816
rect 25820 19756 25884 19760
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 2268 19484 2332 19548
rect 2084 19348 2148 19412
rect 9812 19484 9876 19548
rect 9444 19348 9508 19412
rect 10548 19348 10612 19412
rect 13676 19620 13740 19684
rect 21036 19620 21100 19684
rect 14780 19348 14844 19412
rect 10916 19272 10980 19276
rect 10916 19216 10930 19272
rect 10930 19216 10980 19272
rect 10916 19212 10980 19216
rect 13124 19212 13188 19276
rect 13676 19212 13740 19276
rect 7972 19076 8036 19140
rect 13492 19076 13556 19140
rect 16252 19076 16316 19140
rect 20116 19348 20180 19412
rect 21220 19348 21284 19412
rect 22324 19348 22388 19412
rect 20852 19076 20916 19140
rect 28396 19212 28460 19276
rect 24716 19076 24780 19140
rect 29684 19076 29748 19140
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 6316 18940 6380 19004
rect 22140 18940 22204 19004
rect 22508 19000 22572 19004
rect 22508 18944 22522 19000
rect 22522 18944 22572 19000
rect 22508 18940 22572 18944
rect 30420 18940 30484 19004
rect 30972 18864 31036 18868
rect 30972 18808 30986 18864
rect 30986 18808 31036 18864
rect 30972 18804 31036 18808
rect 22140 18668 22204 18732
rect 6684 18532 6748 18596
rect 7604 18592 7668 18596
rect 7604 18536 7654 18592
rect 7654 18536 7668 18592
rect 7604 18532 7668 18536
rect 10364 18532 10428 18596
rect 11100 18532 11164 18596
rect 14228 18532 14292 18596
rect 18276 18532 18340 18596
rect 21036 18532 21100 18596
rect 30604 18668 30668 18732
rect 25636 18532 25700 18596
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 5764 18396 5828 18460
rect 12020 18396 12084 18460
rect 12940 18396 13004 18460
rect 612 18260 676 18324
rect 9076 18320 9140 18324
rect 9076 18264 9090 18320
rect 9090 18264 9140 18320
rect 9076 18260 9140 18264
rect 11652 18124 11716 18188
rect 23428 18124 23492 18188
rect 10548 18048 10612 18052
rect 10548 17992 10562 18048
rect 10562 17992 10612 18048
rect 10548 17988 10612 17992
rect 11468 17988 11532 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 2084 17852 2148 17916
rect 2452 17852 2516 17916
rect 6500 17912 6564 17916
rect 6500 17856 6514 17912
rect 6514 17856 6564 17912
rect 6500 17852 6564 17856
rect 8156 17852 8220 17916
rect 8892 17852 8956 17916
rect 12204 17852 12268 17916
rect 14964 17988 15028 18052
rect 18828 17988 18892 18052
rect 27660 17988 27724 18052
rect 28948 18048 29012 18052
rect 28948 17992 28998 18048
rect 28998 17992 29012 18048
rect 28948 17988 29012 17992
rect 23244 17852 23308 17916
rect 2636 17716 2700 17780
rect 9996 17716 10060 17780
rect 7788 17580 7852 17644
rect 14412 17580 14476 17644
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 15148 17308 15212 17372
rect 15884 17308 15948 17372
rect 23980 17308 24044 17372
rect 24716 17308 24780 17372
rect 21772 17172 21836 17236
rect 23060 17172 23124 17236
rect 25084 17172 25148 17236
rect 26004 17172 26068 17236
rect 9812 16900 9876 16964
rect 14412 16900 14476 16964
rect 17908 16900 17972 16964
rect 24164 16900 24228 16964
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 4660 16492 4724 16556
rect 5764 16628 5828 16692
rect 15332 16764 15396 16828
rect 15700 16764 15764 16828
rect 12572 16628 12636 16692
rect 12940 16628 13004 16692
rect 19748 16628 19812 16692
rect 9628 16492 9692 16556
rect 10364 16492 10428 16556
rect 11284 16492 11348 16556
rect 12572 16552 12636 16556
rect 12572 16496 12586 16552
rect 12586 16496 12636 16552
rect 12572 16492 12636 16496
rect 12020 16356 12084 16420
rect 16068 16492 16132 16556
rect 25268 16492 25332 16556
rect 26556 16492 26620 16556
rect 19564 16356 19628 16420
rect 24348 16416 24412 16420
rect 24348 16360 24362 16416
rect 24362 16360 24412 16416
rect 24348 16356 24412 16360
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 7236 16220 7300 16284
rect 13124 15948 13188 16012
rect 5396 15812 5460 15876
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 4660 15676 4724 15740
rect 3924 15600 3988 15604
rect 3924 15544 3938 15600
rect 3938 15544 3988 15600
rect 3924 15540 3988 15544
rect 10916 15812 10980 15876
rect 6868 15676 6932 15740
rect 13492 15676 13556 15740
rect 16804 15736 16868 15740
rect 16804 15680 16818 15736
rect 16818 15680 16868 15736
rect 16804 15676 16868 15680
rect 21956 15736 22020 15740
rect 21956 15680 22006 15736
rect 22006 15680 22020 15736
rect 21956 15676 22020 15680
rect 27844 15676 27908 15740
rect 13124 15540 13188 15604
rect 3556 15404 3620 15468
rect 18092 15404 18156 15468
rect 28396 15404 28460 15468
rect 5948 15268 6012 15332
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 3188 15132 3252 15196
rect 9996 15132 10060 15196
rect 23428 15268 23492 15332
rect 11836 15132 11900 15196
rect 19564 15192 19628 15196
rect 19564 15136 19578 15192
rect 19578 15136 19628 15192
rect 19564 15132 19628 15136
rect 29132 15132 29196 15196
rect 980 14996 1044 15060
rect 12204 14996 12268 15060
rect 17724 14996 17788 15060
rect 21220 14996 21284 15060
rect 30972 15056 31036 15060
rect 30972 15000 31022 15056
rect 31022 15000 31036 15056
rect 30972 14996 31036 15000
rect 5580 14860 5644 14924
rect 8708 14860 8772 14924
rect 9260 14724 9324 14788
rect 12388 14860 12452 14924
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 8524 14588 8588 14652
rect 9444 14648 9508 14652
rect 9444 14592 9494 14648
rect 9494 14592 9508 14648
rect 9444 14588 9508 14592
rect 13676 14724 13740 14788
rect 30972 14724 31036 14788
rect 3556 14452 3620 14516
rect 7052 14452 7116 14516
rect 19196 14452 19260 14516
rect 20484 14452 20548 14516
rect 21036 14588 21100 14652
rect 23612 14452 23676 14516
rect 23980 14452 24044 14516
rect 3556 14316 3620 14380
rect 5764 14376 5828 14380
rect 5764 14320 5778 14376
rect 5778 14320 5828 14376
rect 5764 14316 5828 14320
rect 8892 14316 8956 14380
rect 24532 14376 24596 14380
rect 24532 14320 24546 14376
rect 24546 14320 24596 14376
rect 24532 14316 24596 14320
rect 26372 14316 26436 14380
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 7420 14104 7484 14108
rect 7420 14048 7434 14104
rect 7434 14048 7484 14104
rect 7420 14044 7484 14048
rect 11836 14180 11900 14244
rect 12204 14180 12268 14244
rect 10364 14044 10428 14108
rect 12940 14044 13004 14108
rect 12388 13968 12452 13972
rect 12388 13912 12438 13968
rect 12438 13912 12452 13968
rect 12388 13908 12452 13912
rect 17356 14044 17420 14108
rect 20852 14044 20916 14108
rect 21404 14044 21468 14108
rect 28212 13908 28276 13972
rect 8892 13772 8956 13836
rect 9444 13832 9508 13836
rect 9444 13776 9494 13832
rect 9494 13776 9508 13832
rect 9444 13772 9508 13776
rect 10548 13772 10612 13836
rect 11100 13772 11164 13836
rect 12204 13832 12268 13836
rect 12204 13776 12218 13832
rect 12218 13776 12268 13832
rect 12204 13772 12268 13776
rect 23244 13772 23308 13836
rect 23612 13772 23676 13836
rect 26556 13832 26620 13836
rect 26556 13776 26570 13832
rect 26570 13776 26620 13832
rect 26556 13772 26620 13776
rect 14780 13636 14844 13700
rect 16620 13636 16684 13700
rect 18092 13636 18156 13700
rect 21036 13636 21100 13700
rect 22692 13636 22756 13700
rect 23796 13636 23860 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 8340 13500 8404 13564
rect 6868 13364 6932 13428
rect 17356 13364 17420 13428
rect 6132 13092 6196 13156
rect 6316 13092 6380 13156
rect 7236 13152 7300 13156
rect 7236 13096 7250 13152
rect 7250 13096 7300 13152
rect 7236 13092 7300 13096
rect 9076 13092 9140 13156
rect 20116 13228 20180 13292
rect 20300 13228 20364 13292
rect 21956 13228 22020 13292
rect 22692 13288 22756 13292
rect 22692 13232 22706 13288
rect 22706 13232 22756 13288
rect 22692 13228 22756 13232
rect 23060 13228 23124 13292
rect 29316 13500 29380 13564
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 3924 12956 3988 13020
rect 4660 13016 4724 13020
rect 4660 12960 4710 13016
rect 4710 12960 4724 13016
rect 4660 12956 4724 12960
rect 11652 12820 11716 12884
rect 23980 13092 24044 13156
rect 12020 12956 12084 13020
rect 15516 12956 15580 13020
rect 19380 12956 19444 13020
rect 22876 12956 22940 13020
rect 6684 12684 6748 12748
rect 8156 12684 8220 12748
rect 15884 12684 15948 12748
rect 18644 12684 18708 12748
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 3740 12276 3804 12340
rect 7972 12608 8036 12612
rect 7972 12552 7986 12608
rect 7986 12552 8036 12608
rect 7972 12548 8036 12552
rect 16436 12412 16500 12476
rect 6500 12276 6564 12340
rect 15700 12276 15764 12340
rect 28396 12472 28460 12476
rect 28396 12416 28446 12472
rect 28446 12416 28460 12472
rect 28396 12412 28460 12416
rect 20300 12276 20364 12340
rect 25084 12276 25148 12340
rect 29684 12276 29748 12340
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 7788 12140 7852 12204
rect 4660 11868 4724 11932
rect 1164 11732 1228 11796
rect 6500 11928 6564 11932
rect 6500 11872 6550 11928
rect 6550 11872 6564 11928
rect 6500 11868 6564 11872
rect 11284 12064 11348 12068
rect 11284 12008 11298 12064
rect 11298 12008 11348 12064
rect 11284 12004 11348 12008
rect 11468 12004 11532 12068
rect 28580 12064 28644 12068
rect 28580 12008 28630 12064
rect 28630 12008 28644 12064
rect 28580 12004 28644 12008
rect 14964 11868 15028 11932
rect 16252 11868 16316 11932
rect 14596 11732 14660 11796
rect 21404 11732 21468 11796
rect 24716 11732 24780 11796
rect 7420 11596 7484 11660
rect 7604 11656 7668 11660
rect 7604 11600 7654 11656
rect 7654 11600 7668 11656
rect 7604 11596 7668 11600
rect 10180 11596 10244 11660
rect 10364 11656 10428 11660
rect 10364 11600 10414 11656
rect 10414 11600 10428 11656
rect 10364 11596 10428 11600
rect 16436 11596 16500 11660
rect 20668 11596 20732 11660
rect 16988 11460 17052 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 5396 11384 5460 11388
rect 5396 11328 5410 11384
rect 5410 11328 5460 11384
rect 5396 11324 5460 11328
rect 7604 11324 7668 11388
rect 20852 11460 20916 11524
rect 20484 11324 20548 11388
rect 10732 11188 10796 11252
rect 3924 11052 3988 11116
rect 6132 10916 6196 10980
rect 6684 10976 6748 10980
rect 6684 10920 6698 10976
rect 6698 10920 6748 10976
rect 6684 10916 6748 10920
rect 12388 11052 12452 11116
rect 17356 11052 17420 11116
rect 19564 11052 19628 11116
rect 20852 11112 20916 11116
rect 20852 11056 20902 11112
rect 20902 11056 20916 11112
rect 20852 11052 20916 11056
rect 21220 11052 21284 11116
rect 15516 10916 15580 10980
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 6868 10644 6932 10708
rect 8340 10644 8404 10708
rect 2268 10508 2332 10572
rect 9076 10644 9140 10708
rect 9628 10644 9692 10708
rect 22324 10780 22388 10844
rect 22692 10840 22756 10844
rect 22692 10784 22742 10840
rect 22742 10784 22756 10840
rect 22692 10780 22756 10784
rect 23980 10840 24044 10844
rect 23980 10784 23994 10840
rect 23994 10784 24044 10840
rect 23980 10780 24044 10784
rect 26924 10916 26988 10980
rect 24164 10704 24228 10708
rect 24164 10648 24178 10704
rect 24178 10648 24228 10704
rect 24164 10644 24228 10648
rect 6868 10372 6932 10436
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 6316 10236 6380 10300
rect 6500 10236 6564 10300
rect 796 10100 860 10164
rect 3924 9964 3988 10028
rect 1900 9692 1964 9756
rect 10180 10508 10244 10572
rect 30788 10508 30852 10572
rect 12572 10432 12636 10436
rect 12572 10376 12586 10432
rect 12586 10376 12636 10432
rect 12572 10372 12636 10376
rect 19380 10236 19444 10300
rect 20852 10236 20916 10300
rect 23428 10236 23492 10300
rect 29868 10236 29932 10300
rect 7972 10100 8036 10164
rect 8892 9964 8956 10028
rect 10364 9964 10428 10028
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 25452 9828 25516 9892
rect 5580 9556 5644 9620
rect 9260 9556 9324 9620
rect 10548 9692 10612 9756
rect 19564 9752 19628 9756
rect 19564 9696 19614 9752
rect 19614 9696 19628 9752
rect 19564 9692 19628 9696
rect 27660 9692 27724 9756
rect 20668 9556 20732 9620
rect 8892 9420 8956 9484
rect 18460 9420 18524 9484
rect 19196 9420 19260 9484
rect 25268 9420 25332 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 14780 9148 14844 9212
rect 14964 9148 15028 9212
rect 7420 9012 7484 9076
rect 7604 9012 7668 9076
rect 9260 9012 9324 9076
rect 7236 8876 7300 8940
rect 21588 8876 21652 8940
rect 6868 8740 6932 8804
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4660 8468 4724 8532
rect 12020 8468 12084 8532
rect 15332 8468 15396 8532
rect 18828 8468 18892 8532
rect 5396 8392 5460 8396
rect 5396 8336 5446 8392
rect 5446 8336 5460 8392
rect 5396 8332 5460 8336
rect 5948 8332 6012 8396
rect 6868 8332 6932 8396
rect 23612 8196 23676 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 31156 8060 31220 8124
rect 9076 7788 9140 7852
rect 12756 7652 12820 7716
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 13492 7516 13556 7580
rect 15516 7380 15580 7444
rect 23244 7380 23308 7444
rect 24532 7380 24596 7444
rect 7236 7244 7300 7308
rect 11100 7108 11164 7172
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 8156 6972 8220 7036
rect 18644 6972 18708 7036
rect 8708 6836 8772 6900
rect 9812 6836 9876 6900
rect 3556 6700 3620 6764
rect 14044 6700 14108 6764
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 7420 6428 7484 6492
rect 21220 6564 21284 6628
rect 20668 6428 20732 6492
rect 15884 6292 15948 6356
rect 2084 6156 2148 6220
rect 8892 6020 8956 6084
rect 12204 6156 12268 6220
rect 25636 6216 25700 6220
rect 25636 6160 25686 6216
rect 25686 6160 25700 6216
rect 25636 6156 25700 6160
rect 22876 6020 22940 6084
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 30972 5340 31036 5404
rect 9996 5204 10060 5268
rect 26556 5204 26620 5268
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 23244 4660 23308 4724
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 29132 3980 29196 4044
rect 13676 3844 13740 3908
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 26188 3708 26252 3772
rect 25820 3572 25884 3636
rect 5764 3436 5828 3500
rect 30420 3300 30484 3364
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 9444 3164 9508 3228
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 21036 2620 21100 2684
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 979 31380 1045 31381
rect 979 31316 980 31380
rect 1044 31316 1045 31380
rect 979 31315 1045 31316
rect 611 30156 677 30157
rect 611 30092 612 30156
rect 676 30092 677 30156
rect 611 30091 677 30092
rect 614 18325 674 30091
rect 795 20772 861 20773
rect 795 20708 796 20772
rect 860 20708 861 20772
rect 795 20707 861 20708
rect 611 18324 677 18325
rect 611 18260 612 18324
rect 676 18260 677 18324
rect 611 18259 677 18260
rect 798 10165 858 20707
rect 982 15061 1042 31315
rect 2083 31244 2149 31245
rect 2083 31180 2084 31244
rect 2148 31180 2149 31244
rect 2083 31179 2149 31180
rect 1163 29612 1229 29613
rect 1163 29548 1164 29612
rect 1228 29548 1229 29612
rect 1163 29547 1229 29548
rect 979 15060 1045 15061
rect 979 14996 980 15060
rect 1044 14996 1045 15060
rect 979 14995 1045 14996
rect 1166 11797 1226 29547
rect 1899 19956 1965 19957
rect 1899 19892 1900 19956
rect 1964 19892 1965 19956
rect 1899 19891 1965 19892
rect 1163 11796 1229 11797
rect 1163 11732 1164 11796
rect 1228 11732 1229 11796
rect 1163 11731 1229 11732
rect 795 10164 861 10165
rect 795 10100 796 10164
rect 860 10100 861 10164
rect 795 10099 861 10100
rect 1902 9757 1962 19891
rect 2086 19413 2146 31179
rect 4208 31040 4528 31600
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 2635 29748 2701 29749
rect 2635 29684 2636 29748
rect 2700 29684 2701 29748
rect 2635 29683 2701 29684
rect 2451 29204 2517 29205
rect 2451 29140 2452 29204
rect 2516 29140 2517 29204
rect 2451 29139 2517 29140
rect 2267 21724 2333 21725
rect 2267 21660 2268 21724
rect 2332 21660 2333 21724
rect 2267 21659 2333 21660
rect 2270 19685 2330 21659
rect 2267 19684 2333 19685
rect 2267 19620 2268 19684
rect 2332 19620 2333 19684
rect 2267 19619 2333 19620
rect 2267 19548 2333 19549
rect 2267 19484 2268 19548
rect 2332 19484 2333 19548
rect 2267 19483 2333 19484
rect 2083 19412 2149 19413
rect 2083 19348 2084 19412
rect 2148 19348 2149 19412
rect 2083 19347 2149 19348
rect 2083 17916 2149 17917
rect 2083 17852 2084 17916
rect 2148 17852 2149 17916
rect 2083 17851 2149 17852
rect 1899 9756 1965 9757
rect 1899 9692 1900 9756
rect 1964 9692 1965 9756
rect 1899 9691 1965 9692
rect 2086 6221 2146 17851
rect 2270 10573 2330 19483
rect 2454 17917 2514 29139
rect 2451 17916 2517 17917
rect 2451 17852 2452 17916
rect 2516 17852 2517 17916
rect 2451 17851 2517 17852
rect 2638 17781 2698 29683
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 3371 28388 3437 28389
rect 3371 28324 3372 28388
rect 3436 28324 3437 28388
rect 3371 28323 3437 28324
rect 3187 20364 3253 20365
rect 3187 20300 3188 20364
rect 3252 20300 3253 20364
rect 3187 20299 3253 20300
rect 2635 17780 2701 17781
rect 2635 17716 2636 17780
rect 2700 17716 2701 17780
rect 2635 17715 2701 17716
rect 3190 15197 3250 20299
rect 3374 19685 3434 28323
rect 4208 27776 4528 28800
rect 4868 31584 5188 31600
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 20667 31380 20733 31381
rect 20667 31316 20668 31380
rect 20732 31316 20733 31380
rect 20667 31315 20733 31316
rect 14411 30972 14477 30973
rect 14411 30908 14412 30972
rect 14476 30908 14477 30972
rect 14411 30907 14477 30908
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 5395 29476 5461 29477
rect 5395 29412 5396 29476
rect 5460 29412 5461 29476
rect 5395 29411 5461 29412
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4659 28116 4725 28117
rect 4659 28052 4660 28116
rect 4724 28052 4725 28116
rect 4659 28051 4725 28052
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 3739 24852 3805 24853
rect 3739 24788 3740 24852
rect 3804 24788 3805 24852
rect 3739 24787 3805 24788
rect 3555 21860 3621 21861
rect 3555 21796 3556 21860
rect 3620 21796 3621 21860
rect 3555 21795 3621 21796
rect 3371 19684 3437 19685
rect 3371 19620 3372 19684
rect 3436 19620 3437 19684
rect 3371 19619 3437 19620
rect 3558 15469 3618 21795
rect 3555 15468 3621 15469
rect 3555 15404 3556 15468
rect 3620 15404 3621 15468
rect 3555 15403 3621 15404
rect 3187 15196 3253 15197
rect 3187 15132 3188 15196
rect 3252 15132 3253 15196
rect 3187 15131 3253 15132
rect 3558 14517 3618 15403
rect 3555 14516 3621 14517
rect 3555 14452 3556 14516
rect 3620 14452 3621 14516
rect 3555 14451 3621 14452
rect 3555 14380 3621 14381
rect 3555 14316 3556 14380
rect 3620 14316 3621 14380
rect 3555 14315 3621 14316
rect 2267 10572 2333 10573
rect 2267 10508 2268 10572
rect 2332 10508 2333 10572
rect 2267 10507 2333 10508
rect 3558 6765 3618 14315
rect 3742 12341 3802 24787
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4662 23493 4722 28051
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4659 23492 4725 23493
rect 4659 23428 4660 23492
rect 4724 23428 4725 23492
rect 4659 23427 4725 23428
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4659 23084 4725 23085
rect 4659 23020 4660 23084
rect 4724 23020 4725 23084
rect 4659 23019 4725 23020
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 3923 20772 3989 20773
rect 3923 20708 3924 20772
rect 3988 20708 3989 20772
rect 3923 20707 3989 20708
rect 3926 15605 3986 20707
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4662 16557 4722 23019
rect 4868 22880 5188 23904
rect 5398 23085 5458 29411
rect 8155 29068 8221 29069
rect 8155 29004 8156 29068
rect 8220 29004 8221 29068
rect 8155 29003 8221 29004
rect 6315 28932 6381 28933
rect 6315 28868 6316 28932
rect 6380 28868 6381 28932
rect 6315 28867 6381 28868
rect 6131 27028 6197 27029
rect 6131 26964 6132 27028
rect 6196 26964 6197 27028
rect 6131 26963 6197 26964
rect 5579 26484 5645 26485
rect 5579 26420 5580 26484
rect 5644 26420 5645 26484
rect 5579 26419 5645 26420
rect 5947 26484 6013 26485
rect 5947 26420 5948 26484
rect 6012 26420 6013 26484
rect 5947 26419 6013 26420
rect 5395 23084 5461 23085
rect 5395 23020 5396 23084
rect 5460 23020 5461 23084
rect 5395 23019 5461 23020
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 5582 22133 5642 26419
rect 5763 25668 5829 25669
rect 5763 25604 5764 25668
rect 5828 25604 5829 25668
rect 5763 25603 5829 25604
rect 5766 23085 5826 25603
rect 5763 23084 5829 23085
rect 5763 23020 5764 23084
rect 5828 23020 5829 23084
rect 5763 23019 5829 23020
rect 5579 22132 5645 22133
rect 5579 22068 5580 22132
rect 5644 22068 5645 22132
rect 5579 22067 5645 22068
rect 5579 21996 5645 21997
rect 5579 21932 5580 21996
rect 5644 21932 5645 21996
rect 5579 21931 5645 21932
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 5395 21452 5461 21453
rect 5395 21388 5396 21452
rect 5460 21388 5461 21452
rect 5395 21387 5461 21388
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4659 16556 4725 16557
rect 4659 16492 4660 16556
rect 4724 16492 4725 16556
rect 4659 16491 4725 16492
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 3923 15604 3989 15605
rect 3923 15540 3924 15604
rect 3988 15540 3989 15604
rect 3923 15539 3989 15540
rect 4208 14720 4528 15744
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4659 15740 4725 15741
rect 4659 15676 4660 15740
rect 4724 15676 4725 15740
rect 4659 15675 4725 15676
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 3923 13020 3989 13021
rect 3923 12956 3924 13020
rect 3988 12956 3989 13020
rect 3923 12955 3989 12956
rect 3739 12340 3805 12341
rect 3739 12276 3740 12340
rect 3804 12276 3805 12340
rect 3739 12275 3805 12276
rect 3926 11117 3986 12955
rect 4208 12544 4528 13568
rect 4662 13021 4722 15675
rect 4868 15264 5188 16288
rect 5398 15877 5458 21387
rect 5395 15876 5461 15877
rect 5395 15812 5396 15876
rect 5460 15812 5461 15876
rect 5395 15811 5461 15812
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 5582 14925 5642 21931
rect 5763 21316 5829 21317
rect 5763 21252 5764 21316
rect 5828 21252 5829 21316
rect 5763 21251 5829 21252
rect 5766 18461 5826 21251
rect 5950 19821 6010 26419
rect 6134 22133 6194 26963
rect 6318 24037 6378 28867
rect 7419 28660 7485 28661
rect 7419 28596 7420 28660
rect 7484 28596 7485 28660
rect 7419 28595 7485 28596
rect 6499 28388 6565 28389
rect 6499 28324 6500 28388
rect 6564 28324 6565 28388
rect 6499 28323 6565 28324
rect 6315 24036 6381 24037
rect 6315 23972 6316 24036
rect 6380 23972 6381 24036
rect 6315 23971 6381 23972
rect 6502 23493 6562 28323
rect 6867 27980 6933 27981
rect 6867 27916 6868 27980
rect 6932 27916 6933 27980
rect 6867 27915 6933 27916
rect 6870 26210 6930 27915
rect 7235 27436 7301 27437
rect 7235 27372 7236 27436
rect 7300 27372 7301 27436
rect 7235 27371 7301 27372
rect 7051 27300 7117 27301
rect 7051 27236 7052 27300
rect 7116 27236 7117 27300
rect 7051 27235 7117 27236
rect 6686 26150 6930 26210
rect 6499 23492 6565 23493
rect 6499 23428 6500 23492
rect 6564 23428 6565 23492
rect 6499 23427 6565 23428
rect 6502 22269 6562 23427
rect 6499 22268 6565 22269
rect 6499 22204 6500 22268
rect 6564 22204 6565 22268
rect 6499 22203 6565 22204
rect 6131 22132 6197 22133
rect 6131 22068 6132 22132
rect 6196 22068 6197 22132
rect 6686 22110 6746 26150
rect 6131 22067 6197 22068
rect 6502 22050 6746 22110
rect 6867 22132 6933 22133
rect 6867 22068 6868 22132
rect 6932 22068 6933 22132
rect 6867 22067 6933 22068
rect 5947 19820 6013 19821
rect 5947 19756 5948 19820
rect 6012 19756 6013 19820
rect 5947 19755 6013 19756
rect 6315 19004 6381 19005
rect 6315 18940 6316 19004
rect 6380 18940 6381 19004
rect 6315 18939 6381 18940
rect 5763 18460 5829 18461
rect 5763 18396 5764 18460
rect 5828 18396 5829 18460
rect 5763 18395 5829 18396
rect 6318 17370 6378 18939
rect 6502 17917 6562 22050
rect 6683 18596 6749 18597
rect 6683 18532 6684 18596
rect 6748 18532 6749 18596
rect 6683 18531 6749 18532
rect 6499 17916 6565 17917
rect 6499 17852 6500 17916
rect 6564 17852 6565 17916
rect 6499 17851 6565 17852
rect 6318 17310 6562 17370
rect 5763 16692 5829 16693
rect 5763 16628 5764 16692
rect 5828 16628 5829 16692
rect 5763 16627 5829 16628
rect 5579 14924 5645 14925
rect 5579 14860 5580 14924
rect 5644 14860 5645 14924
rect 5579 14859 5645 14860
rect 5766 14650 5826 16627
rect 5947 15332 6013 15333
rect 5947 15268 5948 15332
rect 6012 15268 6013 15332
rect 5947 15267 6013 15268
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4659 13020 4725 13021
rect 4659 12956 4660 13020
rect 4724 12956 4725 13020
rect 4659 12955 4725 12956
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4659 11932 4725 11933
rect 4659 11868 4660 11932
rect 4724 11868 4725 11932
rect 4659 11867 4725 11868
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 3923 11116 3989 11117
rect 3923 11052 3924 11116
rect 3988 11052 3989 11116
rect 3923 11051 3989 11052
rect 3926 10029 3986 11051
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 3923 10028 3989 10029
rect 3923 9964 3924 10028
rect 3988 9964 3989 10028
rect 3923 9963 3989 9964
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4662 8533 4722 11867
rect 4868 10912 5188 11936
rect 5398 14590 5826 14650
rect 5398 11930 5458 14590
rect 5763 14380 5829 14381
rect 5763 14316 5764 14380
rect 5828 14316 5829 14380
rect 5763 14315 5829 14316
rect 5398 11870 5642 11930
rect 5395 11388 5461 11389
rect 5395 11324 5396 11388
rect 5460 11324 5461 11388
rect 5395 11323 5461 11324
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4659 8532 4725 8533
rect 4659 8468 4660 8532
rect 4724 8468 4725 8532
rect 4659 8467 4725 8468
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 3555 6764 3621 6765
rect 3555 6700 3556 6764
rect 3620 6700 3621 6764
rect 3555 6699 3621 6700
rect 2083 6220 2149 6221
rect 2083 6156 2084 6220
rect 2148 6156 2149 6220
rect 2083 6155 2149 6156
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 7648 5188 8672
rect 5398 8397 5458 11323
rect 5582 9621 5642 11870
rect 5579 9620 5645 9621
rect 5579 9556 5580 9620
rect 5644 9556 5645 9620
rect 5579 9555 5645 9556
rect 5395 8396 5461 8397
rect 5395 8332 5396 8396
rect 5460 8332 5461 8396
rect 5395 8331 5461 8332
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 5766 3501 5826 14315
rect 5950 8397 6010 15267
rect 6131 13156 6197 13157
rect 6131 13092 6132 13156
rect 6196 13092 6197 13156
rect 6131 13091 6197 13092
rect 6315 13156 6381 13157
rect 6315 13092 6316 13156
rect 6380 13092 6381 13156
rect 6315 13091 6381 13092
rect 6134 10981 6194 13091
rect 6131 10980 6197 10981
rect 6131 10916 6132 10980
rect 6196 10916 6197 10980
rect 6131 10915 6197 10916
rect 6318 10301 6378 13091
rect 6502 12341 6562 17310
rect 6686 12749 6746 18531
rect 6870 15741 6930 22067
rect 7054 20773 7114 27235
rect 7238 25669 7298 27371
rect 7235 25668 7301 25669
rect 7235 25604 7236 25668
rect 7300 25604 7301 25668
rect 7235 25603 7301 25604
rect 7422 24309 7482 28595
rect 7971 27300 8037 27301
rect 7971 27236 7972 27300
rect 8036 27236 8037 27300
rect 7971 27235 8037 27236
rect 7419 24308 7485 24309
rect 7419 24244 7420 24308
rect 7484 24244 7485 24308
rect 7419 24243 7485 24244
rect 7422 23221 7482 24243
rect 7419 23220 7485 23221
rect 7419 23156 7420 23220
rect 7484 23156 7485 23220
rect 7419 23155 7485 23156
rect 7419 21316 7485 21317
rect 7419 21252 7420 21316
rect 7484 21252 7485 21316
rect 7419 21251 7485 21252
rect 7051 20772 7117 20773
rect 7051 20708 7052 20772
rect 7116 20708 7117 20772
rect 7051 20707 7117 20708
rect 7235 16284 7301 16285
rect 7235 16220 7236 16284
rect 7300 16220 7301 16284
rect 7235 16219 7301 16220
rect 6867 15740 6933 15741
rect 6867 15676 6868 15740
rect 6932 15676 6933 15740
rect 6867 15675 6933 15676
rect 7238 14650 7298 16219
rect 6870 14590 7298 14650
rect 6870 13429 6930 14590
rect 7051 14516 7117 14517
rect 7051 14452 7052 14516
rect 7116 14452 7117 14516
rect 7051 14451 7117 14452
rect 6867 13428 6933 13429
rect 6867 13364 6868 13428
rect 6932 13364 6933 13428
rect 6867 13363 6933 13364
rect 6683 12748 6749 12749
rect 6683 12684 6684 12748
rect 6748 12684 6749 12748
rect 6683 12683 6749 12684
rect 6499 12340 6565 12341
rect 6499 12276 6500 12340
rect 6564 12276 6565 12340
rect 6499 12275 6565 12276
rect 6499 11932 6565 11933
rect 6499 11868 6500 11932
rect 6564 11868 6565 11932
rect 6499 11867 6565 11868
rect 6502 10301 6562 11867
rect 6683 10980 6749 10981
rect 6683 10916 6684 10980
rect 6748 10916 6749 10980
rect 6683 10915 6749 10916
rect 6686 10570 6746 10915
rect 6867 10708 6933 10709
rect 6867 10644 6868 10708
rect 6932 10706 6933 10708
rect 7054 10706 7114 14451
rect 7422 14109 7482 21251
rect 7974 19141 8034 27235
rect 7971 19140 8037 19141
rect 7971 19076 7972 19140
rect 8036 19076 8037 19140
rect 7971 19075 8037 19076
rect 7603 18596 7669 18597
rect 7603 18532 7604 18596
rect 7668 18532 7669 18596
rect 7603 18531 7669 18532
rect 7419 14108 7485 14109
rect 7419 14044 7420 14108
rect 7484 14044 7485 14108
rect 7419 14043 7485 14044
rect 7235 13156 7301 13157
rect 7235 13092 7236 13156
rect 7300 13092 7301 13156
rect 7235 13091 7301 13092
rect 6932 10646 7114 10706
rect 6932 10644 6933 10646
rect 6867 10643 6933 10644
rect 6686 10510 6930 10570
rect 6870 10437 6930 10510
rect 6867 10436 6933 10437
rect 6867 10372 6868 10436
rect 6932 10372 6933 10436
rect 6867 10371 6933 10372
rect 6315 10300 6381 10301
rect 6315 10236 6316 10300
rect 6380 10236 6381 10300
rect 6315 10235 6381 10236
rect 6499 10300 6565 10301
rect 6499 10236 6500 10300
rect 6564 10236 6565 10300
rect 6499 10235 6565 10236
rect 7238 8941 7298 13091
rect 7606 11661 7666 18531
rect 8158 17917 8218 29003
rect 12939 28796 13005 28797
rect 12939 28732 12940 28796
rect 13004 28732 13005 28796
rect 12939 28731 13005 28732
rect 10179 28388 10245 28389
rect 10179 28324 10180 28388
rect 10244 28324 10245 28388
rect 10179 28323 10245 28324
rect 9443 27844 9509 27845
rect 9443 27780 9444 27844
rect 9508 27780 9509 27844
rect 9443 27779 9509 27780
rect 9259 26892 9325 26893
rect 9259 26828 9260 26892
rect 9324 26828 9325 26892
rect 9259 26827 9325 26828
rect 8707 26212 8773 26213
rect 8707 26148 8708 26212
rect 8772 26148 8773 26212
rect 8707 26147 8773 26148
rect 8523 22948 8589 22949
rect 8523 22884 8524 22948
rect 8588 22884 8589 22948
rect 8523 22883 8589 22884
rect 8155 17916 8221 17917
rect 8155 17852 8156 17916
rect 8220 17852 8221 17916
rect 8155 17851 8221 17852
rect 7787 17644 7853 17645
rect 7787 17580 7788 17644
rect 7852 17580 7853 17644
rect 7787 17579 7853 17580
rect 7790 12205 7850 17579
rect 8526 14653 8586 22883
rect 8710 20637 8770 26147
rect 8707 20636 8773 20637
rect 8707 20572 8708 20636
rect 8772 20572 8773 20636
rect 8707 20571 8773 20572
rect 9075 18324 9141 18325
rect 9075 18260 9076 18324
rect 9140 18260 9141 18324
rect 9075 18259 9141 18260
rect 8891 17916 8957 17917
rect 8891 17852 8892 17916
rect 8956 17852 8957 17916
rect 8891 17851 8957 17852
rect 8707 14924 8773 14925
rect 8707 14860 8708 14924
rect 8772 14860 8773 14924
rect 8707 14859 8773 14860
rect 8523 14652 8589 14653
rect 8523 14588 8524 14652
rect 8588 14588 8589 14652
rect 8523 14587 8589 14588
rect 8339 13564 8405 13565
rect 8339 13500 8340 13564
rect 8404 13500 8405 13564
rect 8339 13499 8405 13500
rect 8155 12748 8221 12749
rect 8155 12684 8156 12748
rect 8220 12684 8221 12748
rect 8155 12683 8221 12684
rect 7971 12612 8037 12613
rect 7971 12548 7972 12612
rect 8036 12548 8037 12612
rect 7971 12547 8037 12548
rect 7787 12204 7853 12205
rect 7787 12140 7788 12204
rect 7852 12140 7853 12204
rect 7787 12139 7853 12140
rect 7419 11660 7485 11661
rect 7419 11596 7420 11660
rect 7484 11596 7485 11660
rect 7419 11595 7485 11596
rect 7603 11660 7669 11661
rect 7603 11596 7604 11660
rect 7668 11596 7669 11660
rect 7603 11595 7669 11596
rect 7422 9077 7482 11595
rect 7603 11388 7669 11389
rect 7603 11324 7604 11388
rect 7668 11324 7669 11388
rect 7603 11323 7669 11324
rect 7606 9077 7666 11323
rect 7974 10165 8034 12547
rect 7971 10164 8037 10165
rect 7971 10100 7972 10164
rect 8036 10100 8037 10164
rect 7971 10099 8037 10100
rect 7419 9076 7485 9077
rect 7419 9012 7420 9076
rect 7484 9012 7485 9076
rect 7419 9011 7485 9012
rect 7603 9076 7669 9077
rect 7603 9012 7604 9076
rect 7668 9012 7669 9076
rect 7603 9011 7669 9012
rect 7235 8940 7301 8941
rect 7235 8876 7236 8940
rect 7300 8876 7301 8940
rect 7235 8875 7301 8876
rect 6867 8804 6933 8805
rect 6867 8740 6868 8804
rect 6932 8740 6933 8804
rect 6867 8739 6933 8740
rect 6870 8397 6930 8739
rect 5947 8396 6013 8397
rect 5947 8332 5948 8396
rect 6012 8332 6013 8396
rect 5947 8331 6013 8332
rect 6867 8396 6933 8397
rect 6867 8332 6868 8396
rect 6932 8332 6933 8396
rect 6867 8331 6933 8332
rect 7238 7309 7298 8875
rect 7235 7308 7301 7309
rect 7235 7244 7236 7308
rect 7300 7244 7301 7308
rect 7235 7243 7301 7244
rect 7422 6493 7482 9011
rect 8158 7037 8218 12683
rect 8342 10709 8402 13499
rect 8339 10708 8405 10709
rect 8339 10644 8340 10708
rect 8404 10644 8405 10708
rect 8339 10643 8405 10644
rect 8155 7036 8221 7037
rect 8155 6972 8156 7036
rect 8220 6972 8221 7036
rect 8155 6971 8221 6972
rect 8710 6901 8770 14859
rect 8894 14381 8954 17851
rect 8891 14380 8957 14381
rect 8891 14316 8892 14380
rect 8956 14316 8957 14380
rect 8891 14315 8957 14316
rect 8891 13836 8957 13837
rect 8891 13772 8892 13836
rect 8956 13772 8957 13836
rect 8891 13771 8957 13772
rect 8894 10029 8954 13771
rect 9078 13157 9138 18259
rect 9262 14789 9322 26827
rect 9446 24989 9506 27779
rect 10182 26213 10242 28323
rect 11099 28252 11165 28253
rect 11099 28188 11100 28252
rect 11164 28188 11165 28252
rect 11099 28187 11165 28188
rect 11102 26890 11162 28187
rect 11283 27844 11349 27845
rect 11283 27780 11284 27844
rect 11348 27780 11349 27844
rect 11283 27779 11349 27780
rect 12755 27844 12821 27845
rect 12755 27780 12756 27844
rect 12820 27780 12821 27844
rect 12755 27779 12821 27780
rect 10734 26830 11162 26890
rect 10179 26212 10245 26213
rect 10179 26148 10180 26212
rect 10244 26148 10245 26212
rect 10179 26147 10245 26148
rect 10547 25260 10613 25261
rect 10547 25196 10548 25260
rect 10612 25196 10613 25260
rect 10547 25195 10613 25196
rect 9443 24988 9509 24989
rect 9443 24924 9444 24988
rect 9508 24924 9509 24988
rect 9443 24923 9509 24924
rect 9811 24852 9877 24853
rect 9811 24788 9812 24852
rect 9876 24788 9877 24852
rect 9811 24787 9877 24788
rect 9814 19549 9874 24787
rect 9995 21452 10061 21453
rect 9995 21388 9996 21452
rect 10060 21388 10061 21452
rect 9995 21387 10061 21388
rect 9811 19548 9877 19549
rect 9811 19484 9812 19548
rect 9876 19484 9877 19548
rect 9811 19483 9877 19484
rect 9443 19412 9509 19413
rect 9443 19348 9444 19412
rect 9508 19348 9509 19412
rect 9443 19347 9509 19348
rect 9259 14788 9325 14789
rect 9259 14724 9260 14788
rect 9324 14724 9325 14788
rect 9259 14723 9325 14724
rect 9446 14653 9506 19347
rect 9998 17781 10058 21387
rect 10550 19413 10610 25195
rect 10734 21589 10794 26830
rect 11099 24988 11165 24989
rect 11099 24924 11100 24988
rect 11164 24924 11165 24988
rect 11099 24923 11165 24924
rect 10915 24036 10981 24037
rect 10915 23972 10916 24036
rect 10980 23972 10981 24036
rect 10915 23971 10981 23972
rect 10731 21588 10797 21589
rect 10731 21524 10732 21588
rect 10796 21524 10797 21588
rect 10731 21523 10797 21524
rect 10547 19412 10613 19413
rect 10547 19348 10548 19412
rect 10612 19348 10613 19412
rect 10547 19347 10613 19348
rect 10363 18596 10429 18597
rect 10363 18532 10364 18596
rect 10428 18532 10429 18596
rect 10363 18531 10429 18532
rect 9995 17780 10061 17781
rect 9995 17716 9996 17780
rect 10060 17716 10061 17780
rect 9995 17715 10061 17716
rect 9811 16964 9877 16965
rect 9811 16900 9812 16964
rect 9876 16900 9877 16964
rect 9811 16899 9877 16900
rect 9627 16556 9693 16557
rect 9627 16492 9628 16556
rect 9692 16492 9693 16556
rect 9627 16491 9693 16492
rect 9443 14652 9509 14653
rect 9443 14588 9444 14652
rect 9508 14588 9509 14652
rect 9443 14587 9509 14588
rect 9443 13836 9509 13837
rect 9443 13772 9444 13836
rect 9508 13772 9509 13836
rect 9443 13771 9509 13772
rect 9075 13156 9141 13157
rect 9075 13092 9076 13156
rect 9140 13092 9141 13156
rect 9075 13091 9141 13092
rect 9075 10708 9141 10709
rect 9075 10644 9076 10708
rect 9140 10644 9141 10708
rect 9075 10643 9141 10644
rect 8891 10028 8957 10029
rect 8891 9964 8892 10028
rect 8956 9964 8957 10028
rect 8891 9963 8957 9964
rect 8891 9484 8957 9485
rect 8891 9420 8892 9484
rect 8956 9420 8957 9484
rect 8891 9419 8957 9420
rect 8707 6900 8773 6901
rect 8707 6836 8708 6900
rect 8772 6836 8773 6900
rect 8707 6835 8773 6836
rect 7419 6492 7485 6493
rect 7419 6428 7420 6492
rect 7484 6428 7485 6492
rect 7419 6427 7485 6428
rect 8894 6085 8954 9419
rect 9078 7853 9138 10643
rect 9259 9620 9325 9621
rect 9259 9556 9260 9620
rect 9324 9556 9325 9620
rect 9259 9555 9325 9556
rect 9262 9077 9322 9555
rect 9259 9076 9325 9077
rect 9259 9012 9260 9076
rect 9324 9012 9325 9076
rect 9259 9011 9325 9012
rect 9075 7852 9141 7853
rect 9075 7788 9076 7852
rect 9140 7788 9141 7852
rect 9075 7787 9141 7788
rect 8891 6084 8957 6085
rect 8891 6020 8892 6084
rect 8956 6020 8957 6084
rect 8891 6019 8957 6020
rect 5763 3500 5829 3501
rect 5763 3436 5764 3500
rect 5828 3436 5829 3500
rect 5763 3435 5829 3436
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 9446 3229 9506 13771
rect 9630 10709 9690 16491
rect 9627 10708 9693 10709
rect 9627 10644 9628 10708
rect 9692 10644 9693 10708
rect 9627 10643 9693 10644
rect 9814 6901 9874 16899
rect 10366 16557 10426 18531
rect 10547 18052 10613 18053
rect 10547 17988 10548 18052
rect 10612 17988 10613 18052
rect 10547 17987 10613 17988
rect 10363 16556 10429 16557
rect 10363 16492 10364 16556
rect 10428 16492 10429 16556
rect 10363 16491 10429 16492
rect 9995 15196 10061 15197
rect 9995 15132 9996 15196
rect 10060 15132 10061 15196
rect 9995 15131 10061 15132
rect 9811 6900 9877 6901
rect 9811 6836 9812 6900
rect 9876 6836 9877 6900
rect 9811 6835 9877 6836
rect 9998 5269 10058 15131
rect 10363 14108 10429 14109
rect 10363 14044 10364 14108
rect 10428 14044 10429 14108
rect 10363 14043 10429 14044
rect 10366 13698 10426 14043
rect 10550 13837 10610 17987
rect 10547 13836 10613 13837
rect 10547 13772 10548 13836
rect 10612 13772 10613 13836
rect 10547 13771 10613 13772
rect 10366 13638 10610 13698
rect 10179 11660 10245 11661
rect 10179 11596 10180 11660
rect 10244 11596 10245 11660
rect 10179 11595 10245 11596
rect 10363 11660 10429 11661
rect 10363 11596 10364 11660
rect 10428 11596 10429 11660
rect 10363 11595 10429 11596
rect 10182 10573 10242 11595
rect 10179 10572 10245 10573
rect 10179 10508 10180 10572
rect 10244 10508 10245 10572
rect 10179 10507 10245 10508
rect 10366 10029 10426 11595
rect 10363 10028 10429 10029
rect 10363 9964 10364 10028
rect 10428 9964 10429 10028
rect 10363 9963 10429 9964
rect 10550 9757 10610 13638
rect 10734 11253 10794 21523
rect 10918 19277 10978 23971
rect 11102 23357 11162 24923
rect 11099 23356 11165 23357
rect 11099 23292 11100 23356
rect 11164 23292 11165 23356
rect 11099 23291 11165 23292
rect 11286 23221 11346 27779
rect 12571 27708 12637 27709
rect 12571 27644 12572 27708
rect 12636 27644 12637 27708
rect 12571 27643 12637 27644
rect 12387 25532 12453 25533
rect 12387 25468 12388 25532
rect 12452 25468 12453 25532
rect 12387 25467 12453 25468
rect 11467 23628 11533 23629
rect 11467 23564 11468 23628
rect 11532 23564 11533 23628
rect 11467 23563 11533 23564
rect 11283 23220 11349 23221
rect 11283 23156 11284 23220
rect 11348 23156 11349 23220
rect 11283 23155 11349 23156
rect 10915 19276 10981 19277
rect 10915 19212 10916 19276
rect 10980 19212 10981 19276
rect 10915 19211 10981 19212
rect 11099 18596 11165 18597
rect 11099 18532 11100 18596
rect 11164 18532 11165 18596
rect 11099 18531 11165 18532
rect 10915 15876 10981 15877
rect 10915 15812 10916 15876
rect 10980 15874 10981 15876
rect 11102 15874 11162 18531
rect 11470 18053 11530 23563
rect 12390 23357 12450 25467
rect 12387 23356 12453 23357
rect 12387 23292 12388 23356
rect 12452 23292 12453 23356
rect 12387 23291 12453 23292
rect 12019 22268 12085 22269
rect 12019 22204 12020 22268
rect 12084 22204 12085 22268
rect 12019 22203 12085 22204
rect 12203 22268 12269 22269
rect 12203 22204 12204 22268
rect 12268 22204 12269 22268
rect 12574 22266 12634 27643
rect 12758 26893 12818 27779
rect 12755 26892 12821 26893
rect 12755 26828 12756 26892
rect 12820 26828 12821 26892
rect 12755 26827 12821 26828
rect 12203 22203 12269 22204
rect 12390 22206 12634 22266
rect 11835 20228 11901 20229
rect 11835 20164 11836 20228
rect 11900 20164 11901 20228
rect 11835 20163 11901 20164
rect 11651 19956 11717 19957
rect 11651 19892 11652 19956
rect 11716 19892 11717 19956
rect 11651 19891 11717 19892
rect 11654 18189 11714 19891
rect 11651 18188 11717 18189
rect 11651 18124 11652 18188
rect 11716 18124 11717 18188
rect 11651 18123 11717 18124
rect 11467 18052 11533 18053
rect 11467 17988 11468 18052
rect 11532 17988 11533 18052
rect 11467 17987 11533 17988
rect 11283 16556 11349 16557
rect 11283 16492 11284 16556
rect 11348 16492 11349 16556
rect 11283 16491 11349 16492
rect 10980 15814 11162 15874
rect 10980 15812 10981 15814
rect 10915 15811 10981 15812
rect 11099 13836 11165 13837
rect 11099 13772 11100 13836
rect 11164 13772 11165 13836
rect 11099 13771 11165 13772
rect 10731 11252 10797 11253
rect 10731 11188 10732 11252
rect 10796 11188 10797 11252
rect 10731 11187 10797 11188
rect 10547 9756 10613 9757
rect 10547 9692 10548 9756
rect 10612 9692 10613 9756
rect 10547 9691 10613 9692
rect 11102 7173 11162 13771
rect 11286 12069 11346 16491
rect 11470 12069 11530 17987
rect 11838 15197 11898 20163
rect 12022 18461 12082 22203
rect 12206 20365 12266 22203
rect 12390 21997 12450 22206
rect 12758 22130 12818 26827
rect 12574 22070 12818 22130
rect 12387 21996 12453 21997
rect 12387 21932 12388 21996
rect 12452 21932 12453 21996
rect 12387 21931 12453 21932
rect 12387 21452 12453 21453
rect 12387 21388 12388 21452
rect 12452 21388 12453 21452
rect 12387 21387 12453 21388
rect 12203 20364 12269 20365
rect 12203 20300 12204 20364
rect 12268 20300 12269 20364
rect 12203 20299 12269 20300
rect 12203 20228 12269 20229
rect 12203 20164 12204 20228
rect 12268 20164 12269 20228
rect 12203 20163 12269 20164
rect 12019 18460 12085 18461
rect 12019 18396 12020 18460
rect 12084 18396 12085 18460
rect 12019 18395 12085 18396
rect 12206 18322 12266 20163
rect 12022 18262 12266 18322
rect 12022 16421 12082 18262
rect 12203 17916 12269 17917
rect 12203 17852 12204 17916
rect 12268 17852 12269 17916
rect 12203 17851 12269 17852
rect 12019 16420 12085 16421
rect 12019 16356 12020 16420
rect 12084 16356 12085 16420
rect 12019 16355 12085 16356
rect 11835 15196 11901 15197
rect 11835 15132 11836 15196
rect 11900 15132 11901 15196
rect 11835 15131 11901 15132
rect 11838 14245 11898 15131
rect 12206 15061 12266 17851
rect 12203 15060 12269 15061
rect 12203 14996 12204 15060
rect 12268 14996 12269 15060
rect 12203 14995 12269 14996
rect 12206 14245 12266 14995
rect 12390 14925 12450 21387
rect 12574 16693 12634 22070
rect 12942 21453 13002 28731
rect 13491 28252 13557 28253
rect 13491 28188 13492 28252
rect 13556 28188 13557 28252
rect 13491 28187 13557 28188
rect 13307 26620 13373 26621
rect 13307 26556 13308 26620
rect 13372 26556 13373 26620
rect 13307 26555 13373 26556
rect 13123 24308 13189 24309
rect 13123 24244 13124 24308
rect 13188 24244 13189 24308
rect 13123 24243 13189 24244
rect 12755 21452 12821 21453
rect 12755 21388 12756 21452
rect 12820 21388 12821 21452
rect 12755 21387 12821 21388
rect 12939 21452 13005 21453
rect 12939 21388 12940 21452
rect 13004 21388 13005 21452
rect 12939 21387 13005 21388
rect 12571 16692 12637 16693
rect 12571 16628 12572 16692
rect 12636 16628 12637 16692
rect 12571 16627 12637 16628
rect 12571 16556 12637 16557
rect 12571 16492 12572 16556
rect 12636 16492 12637 16556
rect 12571 16491 12637 16492
rect 12387 14924 12453 14925
rect 12387 14860 12388 14924
rect 12452 14860 12453 14924
rect 12387 14859 12453 14860
rect 11835 14244 11901 14245
rect 11835 14180 11836 14244
rect 11900 14180 11901 14244
rect 11835 14179 11901 14180
rect 12203 14244 12269 14245
rect 12203 14180 12204 14244
rect 12268 14180 12269 14244
rect 12203 14179 12269 14180
rect 12387 13972 12453 13973
rect 12387 13908 12388 13972
rect 12452 13908 12453 13972
rect 12387 13907 12453 13908
rect 12203 13836 12269 13837
rect 12203 13772 12204 13836
rect 12268 13772 12269 13836
rect 12203 13771 12269 13772
rect 12019 13020 12085 13021
rect 12019 13018 12020 13020
rect 11654 12958 12020 13018
rect 11654 12885 11714 12958
rect 12019 12956 12020 12958
rect 12084 12956 12085 13020
rect 12019 12955 12085 12956
rect 11651 12884 11717 12885
rect 11651 12820 11652 12884
rect 11716 12820 11717 12884
rect 11651 12819 11717 12820
rect 12206 12450 12266 13771
rect 12022 12390 12266 12450
rect 11283 12068 11349 12069
rect 11283 12004 11284 12068
rect 11348 12004 11349 12068
rect 11283 12003 11349 12004
rect 11467 12068 11533 12069
rect 11467 12004 11468 12068
rect 11532 12004 11533 12068
rect 11467 12003 11533 12004
rect 12022 8533 12082 12390
rect 12390 11117 12450 13907
rect 12387 11116 12453 11117
rect 12387 11052 12388 11116
rect 12452 11052 12453 11116
rect 12387 11051 12453 11052
rect 12390 9690 12450 11051
rect 12574 10437 12634 16491
rect 12571 10436 12637 10437
rect 12571 10372 12572 10436
rect 12636 10372 12637 10436
rect 12571 10371 12637 10372
rect 12390 9630 12634 9690
rect 12019 8532 12085 8533
rect 12019 8468 12020 8532
rect 12084 8468 12085 8532
rect 12019 8467 12085 8468
rect 11099 7172 11165 7173
rect 11099 7108 11100 7172
rect 11164 7108 11165 7172
rect 11099 7107 11165 7108
rect 12574 6930 12634 9630
rect 12758 7717 12818 21387
rect 12939 20772 13005 20773
rect 12939 20708 12940 20772
rect 13004 20708 13005 20772
rect 12939 20707 13005 20708
rect 12942 18461 13002 20707
rect 13126 19277 13186 24243
rect 13310 24037 13370 26555
rect 13307 24036 13373 24037
rect 13307 23972 13308 24036
rect 13372 23972 13373 24036
rect 13307 23971 13373 23972
rect 13494 23490 13554 28187
rect 14414 27630 14474 30907
rect 17907 30428 17973 30429
rect 17907 30364 17908 30428
rect 17972 30364 17973 30428
rect 17907 30363 17973 30364
rect 15147 27708 15213 27709
rect 15147 27644 15148 27708
rect 15212 27644 15213 27708
rect 15147 27643 15213 27644
rect 16067 27708 16133 27709
rect 16067 27644 16068 27708
rect 16132 27644 16133 27708
rect 16067 27643 16133 27644
rect 14046 27570 14474 27630
rect 13675 25396 13741 25397
rect 13675 25332 13676 25396
rect 13740 25332 13741 25396
rect 13675 25331 13741 25332
rect 13310 23430 13554 23490
rect 13310 21725 13370 23430
rect 13491 21996 13557 21997
rect 13491 21932 13492 21996
rect 13556 21932 13557 21996
rect 13491 21931 13557 21932
rect 13494 21725 13554 21931
rect 13307 21724 13373 21725
rect 13307 21660 13308 21724
rect 13372 21660 13373 21724
rect 13307 21659 13373 21660
rect 13491 21724 13557 21725
rect 13491 21660 13492 21724
rect 13556 21660 13557 21724
rect 13491 21659 13557 21660
rect 13491 21316 13557 21317
rect 13491 21252 13492 21316
rect 13556 21252 13557 21316
rect 13491 21251 13557 21252
rect 13123 19276 13189 19277
rect 13123 19212 13124 19276
rect 13188 19212 13189 19276
rect 13123 19211 13189 19212
rect 13494 19141 13554 21251
rect 13678 20909 13738 25331
rect 14046 21725 14106 27570
rect 14595 23492 14661 23493
rect 14595 23428 14596 23492
rect 14660 23428 14661 23492
rect 14595 23427 14661 23428
rect 14227 21860 14293 21861
rect 14227 21796 14228 21860
rect 14292 21796 14293 21860
rect 14227 21795 14293 21796
rect 14043 21724 14109 21725
rect 14043 21660 14044 21724
rect 14108 21660 14109 21724
rect 14043 21659 14109 21660
rect 13675 20908 13741 20909
rect 13675 20844 13676 20908
rect 13740 20844 13741 20908
rect 13675 20843 13741 20844
rect 14043 20908 14109 20909
rect 14043 20844 14044 20908
rect 14108 20844 14109 20908
rect 14043 20843 14109 20844
rect 13675 19956 13741 19957
rect 13675 19892 13676 19956
rect 13740 19892 13741 19956
rect 13675 19891 13741 19892
rect 13678 19685 13738 19891
rect 13675 19684 13741 19685
rect 13675 19620 13676 19684
rect 13740 19620 13741 19684
rect 13675 19619 13741 19620
rect 13675 19276 13741 19277
rect 13675 19212 13676 19276
rect 13740 19212 13741 19276
rect 13675 19211 13741 19212
rect 13491 19140 13557 19141
rect 13491 19076 13492 19140
rect 13556 19076 13557 19140
rect 13491 19075 13557 19076
rect 13678 19002 13738 19211
rect 13494 18942 13738 19002
rect 12939 18460 13005 18461
rect 12939 18396 12940 18460
rect 13004 18396 13005 18460
rect 12939 18395 13005 18396
rect 12939 16692 13005 16693
rect 12939 16628 12940 16692
rect 13004 16628 13005 16692
rect 12939 16627 13005 16628
rect 12942 14109 13002 16627
rect 13123 16012 13189 16013
rect 13123 15948 13124 16012
rect 13188 15948 13189 16012
rect 13123 15947 13189 15948
rect 13126 15605 13186 15947
rect 13494 15741 13554 18942
rect 13491 15740 13557 15741
rect 13491 15676 13492 15740
rect 13556 15676 13557 15740
rect 13491 15675 13557 15676
rect 13123 15604 13189 15605
rect 13123 15540 13124 15604
rect 13188 15540 13189 15604
rect 13123 15539 13189 15540
rect 12939 14108 13005 14109
rect 12939 14044 12940 14108
rect 13004 14044 13005 14108
rect 12939 14043 13005 14044
rect 12755 7716 12821 7717
rect 12755 7652 12756 7716
rect 12820 7652 12821 7716
rect 12755 7651 12821 7652
rect 13494 7581 13554 15675
rect 13675 14788 13741 14789
rect 13675 14724 13676 14788
rect 13740 14724 13741 14788
rect 13675 14723 13741 14724
rect 13491 7580 13557 7581
rect 13491 7516 13492 7580
rect 13556 7516 13557 7580
rect 13491 7515 13557 7516
rect 12206 6870 12634 6930
rect 12206 6221 12266 6870
rect 12203 6220 12269 6221
rect 12203 6156 12204 6220
rect 12268 6156 12269 6220
rect 12203 6155 12269 6156
rect 9995 5268 10061 5269
rect 9995 5204 9996 5268
rect 10060 5204 10061 5268
rect 9995 5203 10061 5204
rect 13678 3909 13738 14723
rect 14046 6765 14106 20843
rect 14230 18597 14290 21795
rect 14227 18596 14293 18597
rect 14227 18532 14228 18596
rect 14292 18532 14293 18596
rect 14227 18531 14293 18532
rect 14411 17644 14477 17645
rect 14411 17580 14412 17644
rect 14476 17580 14477 17644
rect 14411 17579 14477 17580
rect 14414 16965 14474 17579
rect 14411 16964 14477 16965
rect 14411 16900 14412 16964
rect 14476 16900 14477 16964
rect 14411 16899 14477 16900
rect 14598 11797 14658 23427
rect 14779 21180 14845 21181
rect 14779 21116 14780 21180
rect 14844 21116 14845 21180
rect 14779 21115 14845 21116
rect 14782 19413 14842 21115
rect 14779 19412 14845 19413
rect 14779 19348 14780 19412
rect 14844 19348 14845 19412
rect 14779 19347 14845 19348
rect 14963 18052 15029 18053
rect 14963 17988 14964 18052
rect 15028 17988 15029 18052
rect 14963 17987 15029 17988
rect 14779 13700 14845 13701
rect 14779 13636 14780 13700
rect 14844 13636 14845 13700
rect 14779 13635 14845 13636
rect 14595 11796 14661 11797
rect 14595 11732 14596 11796
rect 14660 11732 14661 11796
rect 14595 11731 14661 11732
rect 14782 9213 14842 13635
rect 14966 11933 15026 17987
rect 15150 17373 15210 27643
rect 15883 24988 15949 24989
rect 15883 24924 15884 24988
rect 15948 24924 15949 24988
rect 15883 24923 15949 24924
rect 15515 20908 15581 20909
rect 15515 20844 15516 20908
rect 15580 20844 15581 20908
rect 15515 20843 15581 20844
rect 15147 17372 15213 17373
rect 15147 17308 15148 17372
rect 15212 17308 15213 17372
rect 15147 17307 15213 17308
rect 15331 16828 15397 16829
rect 15331 16764 15332 16828
rect 15396 16764 15397 16828
rect 15331 16763 15397 16764
rect 14963 11932 15029 11933
rect 14963 11868 14964 11932
rect 15028 11868 15029 11932
rect 14963 11867 15029 11868
rect 14966 9213 15026 11867
rect 14779 9212 14845 9213
rect 14779 9148 14780 9212
rect 14844 9148 14845 9212
rect 14779 9147 14845 9148
rect 14963 9212 15029 9213
rect 14963 9148 14964 9212
rect 15028 9148 15029 9212
rect 14963 9147 15029 9148
rect 15334 8533 15394 16763
rect 15518 13021 15578 20843
rect 15886 17373 15946 24923
rect 15883 17372 15949 17373
rect 15883 17308 15884 17372
rect 15948 17308 15949 17372
rect 15883 17307 15949 17308
rect 15699 16828 15765 16829
rect 15699 16764 15700 16828
rect 15764 16764 15765 16828
rect 15699 16763 15765 16764
rect 15515 13020 15581 13021
rect 15515 12956 15516 13020
rect 15580 12956 15581 13020
rect 15515 12955 15581 12956
rect 15702 12341 15762 16763
rect 16070 16557 16130 27643
rect 17723 26348 17789 26349
rect 17723 26284 17724 26348
rect 17788 26284 17789 26348
rect 17723 26283 17789 26284
rect 16987 25396 17053 25397
rect 16987 25332 16988 25396
rect 17052 25332 17053 25396
rect 16987 25331 17053 25332
rect 16619 25124 16685 25125
rect 16619 25060 16620 25124
rect 16684 25060 16685 25124
rect 16619 25059 16685 25060
rect 16251 19140 16317 19141
rect 16251 19076 16252 19140
rect 16316 19076 16317 19140
rect 16251 19075 16317 19076
rect 16067 16556 16133 16557
rect 16067 16492 16068 16556
rect 16132 16492 16133 16556
rect 16067 16491 16133 16492
rect 15883 12748 15949 12749
rect 15883 12684 15884 12748
rect 15948 12684 15949 12748
rect 15883 12683 15949 12684
rect 15699 12340 15765 12341
rect 15699 12276 15700 12340
rect 15764 12276 15765 12340
rect 15699 12275 15765 12276
rect 15515 10980 15581 10981
rect 15515 10916 15516 10980
rect 15580 10916 15581 10980
rect 15515 10915 15581 10916
rect 15331 8532 15397 8533
rect 15331 8468 15332 8532
rect 15396 8468 15397 8532
rect 15331 8467 15397 8468
rect 15518 7445 15578 10915
rect 15515 7444 15581 7445
rect 15515 7380 15516 7444
rect 15580 7380 15581 7444
rect 15515 7379 15581 7380
rect 14043 6764 14109 6765
rect 14043 6700 14044 6764
rect 14108 6700 14109 6764
rect 14043 6699 14109 6700
rect 15886 6357 15946 12683
rect 16254 11933 16314 19075
rect 16622 13701 16682 25059
rect 16803 24036 16869 24037
rect 16803 23972 16804 24036
rect 16868 23972 16869 24036
rect 16803 23971 16869 23972
rect 16806 15741 16866 23971
rect 16803 15740 16869 15741
rect 16803 15676 16804 15740
rect 16868 15676 16869 15740
rect 16803 15675 16869 15676
rect 16619 13700 16685 13701
rect 16619 13636 16620 13700
rect 16684 13636 16685 13700
rect 16619 13635 16685 13636
rect 16435 12476 16501 12477
rect 16435 12412 16436 12476
rect 16500 12412 16501 12476
rect 16435 12411 16501 12412
rect 16251 11932 16317 11933
rect 16251 11868 16252 11932
rect 16316 11868 16317 11932
rect 16251 11867 16317 11868
rect 16438 11661 16498 12411
rect 16435 11660 16501 11661
rect 16435 11596 16436 11660
rect 16500 11596 16501 11660
rect 16435 11595 16501 11596
rect 16990 11525 17050 25331
rect 17726 15061 17786 26283
rect 17910 23493 17970 30363
rect 18275 29068 18341 29069
rect 18275 29004 18276 29068
rect 18340 29004 18341 29068
rect 18275 29003 18341 29004
rect 17907 23492 17973 23493
rect 17907 23428 17908 23492
rect 17972 23428 17973 23492
rect 17907 23427 17973 23428
rect 18091 21588 18157 21589
rect 18091 21524 18092 21588
rect 18156 21524 18157 21588
rect 18091 21523 18157 21524
rect 17907 21044 17973 21045
rect 17907 20980 17908 21044
rect 17972 20980 17973 21044
rect 17907 20979 17973 20980
rect 17910 16965 17970 20979
rect 18094 20773 18154 21523
rect 18091 20772 18157 20773
rect 18091 20708 18092 20772
rect 18156 20708 18157 20772
rect 18091 20707 18157 20708
rect 18094 20093 18154 20707
rect 18091 20092 18157 20093
rect 18091 20028 18092 20092
rect 18156 20028 18157 20092
rect 18091 20027 18157 20028
rect 18278 18597 18338 29003
rect 20483 27708 20549 27709
rect 20483 27644 20484 27708
rect 20548 27644 20549 27708
rect 20483 27643 20549 27644
rect 19379 27572 19445 27573
rect 19379 27570 19380 27572
rect 19014 27510 19380 27570
rect 18827 27300 18893 27301
rect 18827 27236 18828 27300
rect 18892 27236 18893 27300
rect 18827 27235 18893 27236
rect 18830 26893 18890 27235
rect 19014 27029 19074 27510
rect 19379 27508 19380 27510
rect 19444 27508 19445 27572
rect 19379 27507 19445 27508
rect 19931 27436 19997 27437
rect 19931 27372 19932 27436
rect 19996 27372 19997 27436
rect 19931 27371 19997 27372
rect 19011 27028 19077 27029
rect 19011 26964 19012 27028
rect 19076 26964 19077 27028
rect 19011 26963 19077 26964
rect 18827 26892 18893 26893
rect 18827 26828 18828 26892
rect 18892 26828 18893 26892
rect 18827 26827 18893 26828
rect 19563 26756 19629 26757
rect 19563 26692 19564 26756
rect 19628 26692 19629 26756
rect 19563 26691 19629 26692
rect 19379 25940 19445 25941
rect 19379 25876 19380 25940
rect 19444 25876 19445 25940
rect 19379 25875 19445 25876
rect 19382 25669 19442 25875
rect 19379 25668 19445 25669
rect 19379 25604 19380 25668
rect 19444 25604 19445 25668
rect 19379 25603 19445 25604
rect 19566 24717 19626 26691
rect 19747 25940 19813 25941
rect 19747 25876 19748 25940
rect 19812 25876 19813 25940
rect 19747 25875 19813 25876
rect 19563 24716 19629 24717
rect 19563 24652 19564 24716
rect 19628 24652 19629 24716
rect 19563 24651 19629 24652
rect 19563 23084 19629 23085
rect 19563 23020 19564 23084
rect 19628 23020 19629 23084
rect 19563 23019 19629 23020
rect 19379 22948 19445 22949
rect 19379 22884 19380 22948
rect 19444 22884 19445 22948
rect 19379 22883 19445 22884
rect 18459 22676 18525 22677
rect 18459 22612 18460 22676
rect 18524 22612 18525 22676
rect 18459 22611 18525 22612
rect 18275 18596 18341 18597
rect 18275 18532 18276 18596
rect 18340 18532 18341 18596
rect 18275 18531 18341 18532
rect 17907 16964 17973 16965
rect 17907 16900 17908 16964
rect 17972 16900 17973 16964
rect 17907 16899 17973 16900
rect 18091 15468 18157 15469
rect 18091 15404 18092 15468
rect 18156 15404 18157 15468
rect 18091 15403 18157 15404
rect 17723 15060 17789 15061
rect 17723 14996 17724 15060
rect 17788 14996 17789 15060
rect 17723 14995 17789 14996
rect 17355 14108 17421 14109
rect 17355 14044 17356 14108
rect 17420 14044 17421 14108
rect 17355 14043 17421 14044
rect 17358 13429 17418 14043
rect 18094 13701 18154 15403
rect 18091 13700 18157 13701
rect 18091 13636 18092 13700
rect 18156 13636 18157 13700
rect 18091 13635 18157 13636
rect 17355 13428 17421 13429
rect 17355 13364 17356 13428
rect 17420 13364 17421 13428
rect 17355 13363 17421 13364
rect 16987 11524 17053 11525
rect 16987 11460 16988 11524
rect 17052 11460 17053 11524
rect 16987 11459 17053 11460
rect 17358 11117 17418 13363
rect 17355 11116 17421 11117
rect 17355 11052 17356 11116
rect 17420 11052 17421 11116
rect 17355 11051 17421 11052
rect 18462 9485 18522 22611
rect 19382 20093 19442 22883
rect 19566 21045 19626 23019
rect 19750 22133 19810 25875
rect 19747 22132 19813 22133
rect 19747 22068 19748 22132
rect 19812 22068 19813 22132
rect 19747 22067 19813 22068
rect 19934 21453 19994 27371
rect 20115 22948 20181 22949
rect 20115 22884 20116 22948
rect 20180 22884 20181 22948
rect 20115 22883 20181 22884
rect 19931 21452 19997 21453
rect 19931 21388 19932 21452
rect 19996 21388 19997 21452
rect 19931 21387 19997 21388
rect 19563 21044 19629 21045
rect 19563 20980 19564 21044
rect 19628 20980 19629 21044
rect 19563 20979 19629 20980
rect 19379 20092 19445 20093
rect 19379 20028 19380 20092
rect 19444 20028 19445 20092
rect 19379 20027 19445 20028
rect 18827 18052 18893 18053
rect 18827 17988 18828 18052
rect 18892 17988 18893 18052
rect 18827 17987 18893 17988
rect 18643 12748 18709 12749
rect 18643 12684 18644 12748
rect 18708 12684 18709 12748
rect 18643 12683 18709 12684
rect 18459 9484 18525 9485
rect 18459 9420 18460 9484
rect 18524 9420 18525 9484
rect 18459 9419 18525 9420
rect 18646 7037 18706 12683
rect 18830 8533 18890 17987
rect 19566 16421 19626 20979
rect 20118 19413 20178 22883
rect 20299 22812 20365 22813
rect 20299 22748 20300 22812
rect 20364 22748 20365 22812
rect 20299 22747 20365 22748
rect 20302 22269 20362 22747
rect 20299 22268 20365 22269
rect 20299 22204 20300 22268
rect 20364 22204 20365 22268
rect 20299 22203 20365 22204
rect 20486 21589 20546 27643
rect 20670 24989 20730 31315
rect 30419 30836 30485 30837
rect 30419 30772 30420 30836
rect 30484 30772 30485 30836
rect 30419 30771 30485 30772
rect 29315 29340 29381 29341
rect 29315 29276 29316 29340
rect 29380 29276 29381 29340
rect 29315 29275 29381 29276
rect 21035 28388 21101 28389
rect 21035 28324 21036 28388
rect 21100 28324 21101 28388
rect 21035 28323 21101 28324
rect 20667 24988 20733 24989
rect 20667 24924 20668 24988
rect 20732 24924 20733 24988
rect 20667 24923 20733 24924
rect 20851 24988 20917 24989
rect 20851 24924 20852 24988
rect 20916 24924 20917 24988
rect 20851 24923 20917 24924
rect 20667 24580 20733 24581
rect 20667 24516 20668 24580
rect 20732 24516 20733 24580
rect 20667 24515 20733 24516
rect 20670 22813 20730 24515
rect 20854 24309 20914 24923
rect 20851 24308 20917 24309
rect 20851 24244 20852 24308
rect 20916 24244 20917 24308
rect 20851 24243 20917 24244
rect 20851 24172 20917 24173
rect 20851 24108 20852 24172
rect 20916 24108 20917 24172
rect 20851 24107 20917 24108
rect 20667 22812 20733 22813
rect 20667 22748 20668 22812
rect 20732 22748 20733 22812
rect 20667 22747 20733 22748
rect 20299 21588 20365 21589
rect 20299 21524 20300 21588
rect 20364 21524 20365 21588
rect 20299 21523 20365 21524
rect 20483 21588 20549 21589
rect 20483 21524 20484 21588
rect 20548 21524 20549 21588
rect 20483 21523 20549 21524
rect 20115 19412 20181 19413
rect 20115 19348 20116 19412
rect 20180 19348 20181 19412
rect 20115 19347 20181 19348
rect 19747 16692 19813 16693
rect 19747 16628 19748 16692
rect 19812 16628 19813 16692
rect 19747 16627 19813 16628
rect 19563 16420 19629 16421
rect 19563 16356 19564 16420
rect 19628 16356 19629 16420
rect 19563 16355 19629 16356
rect 19563 15196 19629 15197
rect 19563 15132 19564 15196
rect 19628 15132 19629 15196
rect 19563 15131 19629 15132
rect 19195 14516 19261 14517
rect 19195 14452 19196 14516
rect 19260 14452 19261 14516
rect 19195 14451 19261 14452
rect 19198 9485 19258 14451
rect 19379 13020 19445 13021
rect 19379 12956 19380 13020
rect 19444 12956 19445 13020
rect 19379 12955 19445 12956
rect 19382 10301 19442 12955
rect 19566 11117 19626 15131
rect 19563 11116 19629 11117
rect 19563 11052 19564 11116
rect 19628 11052 19629 11116
rect 19563 11051 19629 11052
rect 19379 10300 19445 10301
rect 19379 10236 19380 10300
rect 19444 10236 19445 10300
rect 19379 10235 19445 10236
rect 19563 9756 19629 9757
rect 19563 9692 19564 9756
rect 19628 9754 19629 9756
rect 19750 9754 19810 16627
rect 20118 13293 20178 19347
rect 20302 13293 20362 21523
rect 20854 21453 20914 24107
rect 20851 21452 20917 21453
rect 20851 21388 20852 21452
rect 20916 21388 20917 21452
rect 20851 21387 20917 21388
rect 20667 20772 20733 20773
rect 20667 20708 20668 20772
rect 20732 20708 20733 20772
rect 20667 20707 20733 20708
rect 20483 14516 20549 14517
rect 20483 14452 20484 14516
rect 20548 14452 20549 14516
rect 20483 14451 20549 14452
rect 20115 13292 20181 13293
rect 20115 13228 20116 13292
rect 20180 13228 20181 13292
rect 20115 13227 20181 13228
rect 20299 13292 20365 13293
rect 20299 13228 20300 13292
rect 20364 13228 20365 13292
rect 20299 13227 20365 13228
rect 20302 12341 20362 13227
rect 20299 12340 20365 12341
rect 20299 12276 20300 12340
rect 20364 12276 20365 12340
rect 20299 12275 20365 12276
rect 20486 11389 20546 14451
rect 20670 12450 20730 20707
rect 21038 19685 21098 28323
rect 27843 27844 27909 27845
rect 27843 27780 27844 27844
rect 27908 27780 27909 27844
rect 27843 27779 27909 27780
rect 23427 27708 23493 27709
rect 23427 27644 23428 27708
rect 23492 27644 23493 27708
rect 23427 27643 23493 27644
rect 22507 27572 22573 27573
rect 22507 27508 22508 27572
rect 22572 27508 22573 27572
rect 22507 27507 22573 27508
rect 21403 26892 21469 26893
rect 21403 26828 21404 26892
rect 21468 26828 21469 26892
rect 21403 26827 21469 26828
rect 21219 26348 21285 26349
rect 21219 26284 21220 26348
rect 21284 26284 21285 26348
rect 21219 26283 21285 26284
rect 21035 19684 21101 19685
rect 21035 19620 21036 19684
rect 21100 19620 21101 19684
rect 21035 19619 21101 19620
rect 21222 19413 21282 26283
rect 21406 22133 21466 26827
rect 21771 25804 21837 25805
rect 21771 25740 21772 25804
rect 21836 25740 21837 25804
rect 21771 25739 21837 25740
rect 21403 22132 21469 22133
rect 21403 22068 21404 22132
rect 21468 22068 21469 22132
rect 21403 22067 21469 22068
rect 21587 21044 21653 21045
rect 21587 20980 21588 21044
rect 21652 20980 21653 21044
rect 21587 20979 21653 20980
rect 21219 19412 21285 19413
rect 21219 19348 21220 19412
rect 21284 19348 21285 19412
rect 21219 19347 21285 19348
rect 20851 19140 20917 19141
rect 20851 19076 20852 19140
rect 20916 19076 20917 19140
rect 20851 19075 20917 19076
rect 20854 14109 20914 19075
rect 21035 18596 21101 18597
rect 21035 18532 21036 18596
rect 21100 18532 21101 18596
rect 21035 18531 21101 18532
rect 21038 14653 21098 18531
rect 21222 15061 21282 19347
rect 21219 15060 21285 15061
rect 21219 14996 21220 15060
rect 21284 14996 21285 15060
rect 21219 14995 21285 14996
rect 21035 14652 21101 14653
rect 21035 14588 21036 14652
rect 21100 14588 21101 14652
rect 21035 14587 21101 14588
rect 20851 14108 20917 14109
rect 20851 14044 20852 14108
rect 20916 14044 20917 14108
rect 20851 14043 20917 14044
rect 21403 14108 21469 14109
rect 21403 14044 21404 14108
rect 21468 14044 21469 14108
rect 21403 14043 21469 14044
rect 21035 13700 21101 13701
rect 21035 13636 21036 13700
rect 21100 13636 21101 13700
rect 21035 13635 21101 13636
rect 20670 12390 20914 12450
rect 20667 11660 20733 11661
rect 20667 11596 20668 11660
rect 20732 11596 20733 11660
rect 20667 11595 20733 11596
rect 20483 11388 20549 11389
rect 20483 11324 20484 11388
rect 20548 11324 20549 11388
rect 20483 11323 20549 11324
rect 19628 9694 19810 9754
rect 19628 9692 19629 9694
rect 19563 9691 19629 9692
rect 20670 9621 20730 11595
rect 20854 11525 20914 12390
rect 20851 11524 20917 11525
rect 20851 11460 20852 11524
rect 20916 11460 20917 11524
rect 20851 11459 20917 11460
rect 20851 11116 20917 11117
rect 20851 11052 20852 11116
rect 20916 11052 20917 11116
rect 20851 11051 20917 11052
rect 20854 10301 20914 11051
rect 20851 10300 20917 10301
rect 20851 10236 20852 10300
rect 20916 10236 20917 10300
rect 20851 10235 20917 10236
rect 20667 9620 20733 9621
rect 20667 9556 20668 9620
rect 20732 9556 20733 9620
rect 20667 9555 20733 9556
rect 19195 9484 19261 9485
rect 19195 9420 19196 9484
rect 19260 9420 19261 9484
rect 19195 9419 19261 9420
rect 18827 8532 18893 8533
rect 18827 8468 18828 8532
rect 18892 8468 18893 8532
rect 18827 8467 18893 8468
rect 18643 7036 18709 7037
rect 18643 6972 18644 7036
rect 18708 6972 18709 7036
rect 18643 6971 18709 6972
rect 20670 6493 20730 9555
rect 20667 6492 20733 6493
rect 20667 6428 20668 6492
rect 20732 6428 20733 6492
rect 20667 6427 20733 6428
rect 15883 6356 15949 6357
rect 15883 6292 15884 6356
rect 15948 6292 15949 6356
rect 15883 6291 15949 6292
rect 13675 3908 13741 3909
rect 13675 3844 13676 3908
rect 13740 3844 13741 3908
rect 13675 3843 13741 3844
rect 9443 3228 9509 3229
rect 9443 3164 9444 3228
rect 9508 3164 9509 3228
rect 9443 3163 9509 3164
rect 21038 2685 21098 13635
rect 21406 11797 21466 14043
rect 21403 11796 21469 11797
rect 21403 11732 21404 11796
rect 21468 11732 21469 11796
rect 21403 11731 21469 11732
rect 21219 11116 21285 11117
rect 21219 11052 21220 11116
rect 21284 11052 21285 11116
rect 21219 11051 21285 11052
rect 21222 6629 21282 11051
rect 21590 8941 21650 20979
rect 21774 19957 21834 25739
rect 21955 23492 22021 23493
rect 21955 23428 21956 23492
rect 22020 23428 22021 23492
rect 21955 23427 22021 23428
rect 22139 23492 22205 23493
rect 22139 23428 22140 23492
rect 22204 23428 22205 23492
rect 22139 23427 22205 23428
rect 21771 19956 21837 19957
rect 21771 19892 21772 19956
rect 21836 19892 21837 19956
rect 21771 19891 21837 19892
rect 21771 17236 21837 17237
rect 21771 17172 21772 17236
rect 21836 17172 21837 17236
rect 21771 17171 21837 17172
rect 21774 13290 21834 17171
rect 21958 15741 22018 23427
rect 22142 21317 22202 23427
rect 22139 21316 22205 21317
rect 22139 21252 22140 21316
rect 22204 21252 22205 21316
rect 22139 21251 22205 21252
rect 22323 19412 22389 19413
rect 22323 19348 22324 19412
rect 22388 19348 22389 19412
rect 22323 19347 22389 19348
rect 22139 19004 22205 19005
rect 22139 18940 22140 19004
rect 22204 18940 22205 19004
rect 22139 18939 22205 18940
rect 22142 18733 22202 18939
rect 22139 18732 22205 18733
rect 22139 18668 22140 18732
rect 22204 18668 22205 18732
rect 22139 18667 22205 18668
rect 21955 15740 22021 15741
rect 21955 15676 21956 15740
rect 22020 15676 22021 15740
rect 21955 15675 22021 15676
rect 21955 13292 22021 13293
rect 21955 13290 21956 13292
rect 21774 13230 21956 13290
rect 21955 13228 21956 13230
rect 22020 13228 22021 13292
rect 21955 13227 22021 13228
rect 22326 10845 22386 19347
rect 22510 19005 22570 27507
rect 22875 23220 22941 23221
rect 22875 23156 22876 23220
rect 22940 23156 22941 23220
rect 22875 23155 22941 23156
rect 22691 21860 22757 21861
rect 22691 21796 22692 21860
rect 22756 21796 22757 21860
rect 22691 21795 22757 21796
rect 22507 19004 22573 19005
rect 22507 18940 22508 19004
rect 22572 18940 22573 19004
rect 22507 18939 22573 18940
rect 22694 13701 22754 21795
rect 22878 21725 22938 23155
rect 23430 21725 23490 27643
rect 24531 27572 24597 27573
rect 24531 27508 24532 27572
rect 24596 27508 24597 27572
rect 24531 27507 24597 27508
rect 23979 23492 24045 23493
rect 23979 23428 23980 23492
rect 24044 23428 24045 23492
rect 23979 23427 24045 23428
rect 22875 21724 22941 21725
rect 22875 21660 22876 21724
rect 22940 21660 22941 21724
rect 22875 21659 22941 21660
rect 23427 21724 23493 21725
rect 23427 21660 23428 21724
rect 23492 21660 23493 21724
rect 23427 21659 23493 21660
rect 23427 21588 23493 21589
rect 23427 21524 23428 21588
rect 23492 21524 23493 21588
rect 23427 21523 23493 21524
rect 23059 21180 23125 21181
rect 23059 21116 23060 21180
rect 23124 21116 23125 21180
rect 23059 21115 23125 21116
rect 23062 17237 23122 21115
rect 23430 18189 23490 21523
rect 23427 18188 23493 18189
rect 23427 18124 23428 18188
rect 23492 18124 23493 18188
rect 23427 18123 23493 18124
rect 23243 17916 23309 17917
rect 23243 17852 23244 17916
rect 23308 17852 23309 17916
rect 23243 17851 23309 17852
rect 23246 17370 23306 17851
rect 23982 17373 24042 23427
rect 24347 21724 24413 21725
rect 24347 21660 24348 21724
rect 24412 21660 24413 21724
rect 24347 21659 24413 21660
rect 23979 17372 24045 17373
rect 23246 17310 23858 17370
rect 23059 17236 23125 17237
rect 23059 17172 23060 17236
rect 23124 17172 23125 17236
rect 23059 17171 23125 17172
rect 22691 13700 22757 13701
rect 22691 13636 22692 13700
rect 22756 13636 22757 13700
rect 22691 13635 22757 13636
rect 23062 13293 23122 17171
rect 23427 15332 23493 15333
rect 23427 15268 23428 15332
rect 23492 15268 23493 15332
rect 23427 15267 23493 15268
rect 23243 13836 23309 13837
rect 23243 13772 23244 13836
rect 23308 13772 23309 13836
rect 23243 13771 23309 13772
rect 22691 13292 22757 13293
rect 22691 13228 22692 13292
rect 22756 13228 22757 13292
rect 22691 13227 22757 13228
rect 23059 13292 23125 13293
rect 23059 13228 23060 13292
rect 23124 13228 23125 13292
rect 23059 13227 23125 13228
rect 22694 10845 22754 13227
rect 22875 13020 22941 13021
rect 22875 12956 22876 13020
rect 22940 12956 22941 13020
rect 22875 12955 22941 12956
rect 22323 10844 22389 10845
rect 22323 10780 22324 10844
rect 22388 10780 22389 10844
rect 22323 10779 22389 10780
rect 22691 10844 22757 10845
rect 22691 10780 22692 10844
rect 22756 10780 22757 10844
rect 22691 10779 22757 10780
rect 21587 8940 21653 8941
rect 21587 8876 21588 8940
rect 21652 8876 21653 8940
rect 21587 8875 21653 8876
rect 21219 6628 21285 6629
rect 21219 6564 21220 6628
rect 21284 6564 21285 6628
rect 21219 6563 21285 6564
rect 22878 6085 22938 12955
rect 23246 7445 23306 13771
rect 23430 10301 23490 15267
rect 23611 14516 23677 14517
rect 23611 14452 23612 14516
rect 23676 14452 23677 14516
rect 23611 14451 23677 14452
rect 23614 13837 23674 14451
rect 23611 13836 23677 13837
rect 23611 13772 23612 13836
rect 23676 13772 23677 13836
rect 23611 13771 23677 13772
rect 23427 10300 23493 10301
rect 23427 10236 23428 10300
rect 23492 10236 23493 10300
rect 23427 10235 23493 10236
rect 23614 8261 23674 13771
rect 23798 13701 23858 17310
rect 23979 17308 23980 17372
rect 24044 17308 24045 17372
rect 23979 17307 24045 17308
rect 24163 16964 24229 16965
rect 24163 16900 24164 16964
rect 24228 16900 24229 16964
rect 24163 16899 24229 16900
rect 23979 14516 24045 14517
rect 23979 14452 23980 14516
rect 24044 14452 24045 14516
rect 23979 14451 24045 14452
rect 23795 13700 23861 13701
rect 23795 13636 23796 13700
rect 23860 13636 23861 13700
rect 23795 13635 23861 13636
rect 23982 13157 24042 14451
rect 23979 13156 24045 13157
rect 23979 13092 23980 13156
rect 24044 13092 24045 13156
rect 23979 13091 24045 13092
rect 23982 10845 24042 13091
rect 23979 10844 24045 10845
rect 23979 10780 23980 10844
rect 24044 10780 24045 10844
rect 23979 10779 24045 10780
rect 24166 10709 24226 16899
rect 24350 16421 24410 21659
rect 24347 16420 24413 16421
rect 24347 16356 24348 16420
rect 24412 16356 24413 16420
rect 24347 16355 24413 16356
rect 24534 14381 24594 27507
rect 26923 26484 26989 26485
rect 26923 26420 26924 26484
rect 26988 26420 26989 26484
rect 26923 26419 26989 26420
rect 24899 26348 24965 26349
rect 24899 26284 24900 26348
rect 24964 26284 24965 26348
rect 24899 26283 24965 26284
rect 24715 22268 24781 22269
rect 24715 22204 24716 22268
rect 24780 22204 24781 22268
rect 24715 22203 24781 22204
rect 24718 19141 24778 22203
rect 24902 20093 24962 26283
rect 26187 26212 26253 26213
rect 26187 26148 26188 26212
rect 26252 26148 26253 26212
rect 26187 26147 26253 26148
rect 25819 25940 25885 25941
rect 25819 25876 25820 25940
rect 25884 25876 25885 25940
rect 25819 25875 25885 25876
rect 25267 22948 25333 22949
rect 25267 22884 25268 22948
rect 25332 22884 25333 22948
rect 25267 22883 25333 22884
rect 25083 22404 25149 22405
rect 25083 22340 25084 22404
rect 25148 22340 25149 22404
rect 25083 22339 25149 22340
rect 24899 20092 24965 20093
rect 24899 20028 24900 20092
rect 24964 20028 24965 20092
rect 24899 20027 24965 20028
rect 24715 19140 24781 19141
rect 24715 19076 24716 19140
rect 24780 19076 24781 19140
rect 24715 19075 24781 19076
rect 24715 17372 24781 17373
rect 24715 17308 24716 17372
rect 24780 17308 24781 17372
rect 24715 17307 24781 17308
rect 24531 14380 24597 14381
rect 24531 14316 24532 14380
rect 24596 14316 24597 14380
rect 24531 14315 24597 14316
rect 24163 10708 24229 10709
rect 24163 10644 24164 10708
rect 24228 10644 24229 10708
rect 24163 10643 24229 10644
rect 23611 8260 23677 8261
rect 23611 8196 23612 8260
rect 23676 8196 23677 8260
rect 23611 8195 23677 8196
rect 24534 7445 24594 14315
rect 24718 11797 24778 17307
rect 25086 17237 25146 22339
rect 25270 19821 25330 22883
rect 25822 21997 25882 25875
rect 25819 21996 25885 21997
rect 25819 21932 25820 21996
rect 25884 21932 25885 21996
rect 25819 21931 25885 21932
rect 25451 20772 25517 20773
rect 25451 20708 25452 20772
rect 25516 20708 25517 20772
rect 25451 20707 25517 20708
rect 25267 19820 25333 19821
rect 25267 19756 25268 19820
rect 25332 19756 25333 19820
rect 25267 19755 25333 19756
rect 25083 17236 25149 17237
rect 25083 17172 25084 17236
rect 25148 17172 25149 17236
rect 25083 17171 25149 17172
rect 25086 12341 25146 17171
rect 25267 16556 25333 16557
rect 25267 16492 25268 16556
rect 25332 16492 25333 16556
rect 25267 16491 25333 16492
rect 25083 12340 25149 12341
rect 25083 12276 25084 12340
rect 25148 12276 25149 12340
rect 25083 12275 25149 12276
rect 24715 11796 24781 11797
rect 24715 11732 24716 11796
rect 24780 11732 24781 11796
rect 24715 11731 24781 11732
rect 25270 9485 25330 16491
rect 25454 9893 25514 20707
rect 26003 19956 26069 19957
rect 26003 19892 26004 19956
rect 26068 19892 26069 19956
rect 26003 19891 26069 19892
rect 25819 19820 25885 19821
rect 25819 19756 25820 19820
rect 25884 19756 25885 19820
rect 25819 19755 25885 19756
rect 25635 18596 25701 18597
rect 25635 18532 25636 18596
rect 25700 18532 25701 18596
rect 25635 18531 25701 18532
rect 25451 9892 25517 9893
rect 25451 9828 25452 9892
rect 25516 9828 25517 9892
rect 25451 9827 25517 9828
rect 25267 9484 25333 9485
rect 25267 9420 25268 9484
rect 25332 9420 25333 9484
rect 25267 9419 25333 9420
rect 23243 7444 23309 7445
rect 23243 7380 23244 7444
rect 23308 7380 23309 7444
rect 23243 7379 23309 7380
rect 24531 7444 24597 7445
rect 24531 7380 24532 7444
rect 24596 7380 24597 7444
rect 24531 7379 24597 7380
rect 22875 6084 22941 6085
rect 22875 6020 22876 6084
rect 22940 6020 22941 6084
rect 22875 6019 22941 6020
rect 23246 4725 23306 7379
rect 25638 6221 25698 18531
rect 25635 6220 25701 6221
rect 25635 6156 25636 6220
rect 25700 6156 25701 6220
rect 25635 6155 25701 6156
rect 23243 4724 23309 4725
rect 23243 4660 23244 4724
rect 23308 4660 23309 4724
rect 23243 4659 23309 4660
rect 25822 3637 25882 19755
rect 26006 17237 26066 19891
rect 26003 17236 26069 17237
rect 26003 17172 26004 17236
rect 26068 17172 26069 17236
rect 26003 17171 26069 17172
rect 26190 3773 26250 26147
rect 26371 25260 26437 25261
rect 26371 25196 26372 25260
rect 26436 25196 26437 25260
rect 26371 25195 26437 25196
rect 26374 14381 26434 25195
rect 26555 20772 26621 20773
rect 26555 20708 26556 20772
rect 26620 20708 26621 20772
rect 26555 20707 26621 20708
rect 26558 16557 26618 20707
rect 26555 16556 26621 16557
rect 26555 16492 26556 16556
rect 26620 16492 26621 16556
rect 26555 16491 26621 16492
rect 26371 14380 26437 14381
rect 26371 14316 26372 14380
rect 26436 14316 26437 14380
rect 26371 14315 26437 14316
rect 26555 13836 26621 13837
rect 26555 13772 26556 13836
rect 26620 13772 26621 13836
rect 26555 13771 26621 13772
rect 26558 5269 26618 13771
rect 26926 10981 26986 26419
rect 27659 18052 27725 18053
rect 27659 17988 27660 18052
rect 27724 17988 27725 18052
rect 27659 17987 27725 17988
rect 26923 10980 26989 10981
rect 26923 10916 26924 10980
rect 26988 10916 26989 10980
rect 26923 10915 26989 10916
rect 27662 9757 27722 17987
rect 27846 15741 27906 27779
rect 28947 25532 29013 25533
rect 28947 25468 28948 25532
rect 29012 25468 29013 25532
rect 28947 25467 29013 25468
rect 28579 24988 28645 24989
rect 28579 24924 28580 24988
rect 28644 24924 28645 24988
rect 28579 24923 28645 24924
rect 28395 24036 28461 24037
rect 28395 23972 28396 24036
rect 28460 23972 28461 24036
rect 28395 23971 28461 23972
rect 28211 23492 28277 23493
rect 28211 23428 28212 23492
rect 28276 23428 28277 23492
rect 28211 23427 28277 23428
rect 27843 15740 27909 15741
rect 27843 15676 27844 15740
rect 27908 15676 27909 15740
rect 27843 15675 27909 15676
rect 28214 13973 28274 23427
rect 28398 19277 28458 23971
rect 28395 19276 28461 19277
rect 28395 19212 28396 19276
rect 28460 19212 28461 19276
rect 28395 19211 28461 19212
rect 28395 15468 28461 15469
rect 28395 15404 28396 15468
rect 28460 15404 28461 15468
rect 28395 15403 28461 15404
rect 28211 13972 28277 13973
rect 28211 13908 28212 13972
rect 28276 13908 28277 13972
rect 28211 13907 28277 13908
rect 28398 12477 28458 15403
rect 28395 12476 28461 12477
rect 28395 12412 28396 12476
rect 28460 12412 28461 12476
rect 28395 12411 28461 12412
rect 28582 12069 28642 24923
rect 28950 18053 29010 25467
rect 28947 18052 29013 18053
rect 28947 17988 28948 18052
rect 29012 17988 29013 18052
rect 28947 17987 29013 17988
rect 29131 15196 29197 15197
rect 29131 15132 29132 15196
rect 29196 15132 29197 15196
rect 29131 15131 29197 15132
rect 28579 12068 28645 12069
rect 28579 12004 28580 12068
rect 28644 12004 28645 12068
rect 28579 12003 28645 12004
rect 27659 9756 27725 9757
rect 27659 9692 27660 9756
rect 27724 9692 27725 9756
rect 27659 9691 27725 9692
rect 26555 5268 26621 5269
rect 26555 5204 26556 5268
rect 26620 5204 26621 5268
rect 26555 5203 26621 5204
rect 29134 4045 29194 15131
rect 29318 13565 29378 29275
rect 29867 27028 29933 27029
rect 29867 26964 29868 27028
rect 29932 26964 29933 27028
rect 29867 26963 29933 26964
rect 29683 19140 29749 19141
rect 29683 19076 29684 19140
rect 29748 19076 29749 19140
rect 29683 19075 29749 19076
rect 29315 13564 29381 13565
rect 29315 13500 29316 13564
rect 29380 13500 29381 13564
rect 29315 13499 29381 13500
rect 29686 12341 29746 19075
rect 29683 12340 29749 12341
rect 29683 12276 29684 12340
rect 29748 12276 29749 12340
rect 29683 12275 29749 12276
rect 29870 10301 29930 26963
rect 30422 20501 30482 30771
rect 30603 30564 30669 30565
rect 30603 30500 30604 30564
rect 30668 30500 30669 30564
rect 30603 30499 30669 30500
rect 30419 20500 30485 20501
rect 30419 20436 30420 20500
rect 30484 20436 30485 20500
rect 30419 20435 30485 20436
rect 30419 19004 30485 19005
rect 30419 18940 30420 19004
rect 30484 18940 30485 19004
rect 30419 18939 30485 18940
rect 29867 10300 29933 10301
rect 29867 10236 29868 10300
rect 29932 10236 29933 10300
rect 29867 10235 29933 10236
rect 29131 4044 29197 4045
rect 29131 3980 29132 4044
rect 29196 3980 29197 4044
rect 29131 3979 29197 3980
rect 26187 3772 26253 3773
rect 26187 3708 26188 3772
rect 26252 3708 26253 3772
rect 26187 3707 26253 3708
rect 25819 3636 25885 3637
rect 25819 3572 25820 3636
rect 25884 3572 25885 3636
rect 25819 3571 25885 3572
rect 30422 3365 30482 18939
rect 30606 18733 30666 30499
rect 30787 26756 30853 26757
rect 30787 26692 30788 26756
rect 30852 26692 30853 26756
rect 30787 26691 30853 26692
rect 30603 18732 30669 18733
rect 30603 18668 30604 18732
rect 30668 18668 30669 18732
rect 30603 18667 30669 18668
rect 30790 10573 30850 26691
rect 31155 21316 31221 21317
rect 31155 21252 31156 21316
rect 31220 21252 31221 21316
rect 31155 21251 31221 21252
rect 30971 18868 31037 18869
rect 30971 18804 30972 18868
rect 31036 18804 31037 18868
rect 30971 18803 31037 18804
rect 30974 15061 31034 18803
rect 30971 15060 31037 15061
rect 30971 14996 30972 15060
rect 31036 14996 31037 15060
rect 30971 14995 31037 14996
rect 30971 14788 31037 14789
rect 30971 14724 30972 14788
rect 31036 14724 31037 14788
rect 30971 14723 31037 14724
rect 30787 10572 30853 10573
rect 30787 10508 30788 10572
rect 30852 10508 30853 10572
rect 30787 10507 30853 10508
rect 30974 5405 31034 14723
rect 31158 8125 31218 21251
rect 31155 8124 31221 8125
rect 31155 8060 31156 8124
rect 31220 8060 31221 8124
rect 31155 8059 31221 8060
rect 30971 5404 31037 5405
rect 30971 5340 30972 5404
rect 31036 5340 31037 5404
rect 30971 5339 31037 5340
rect 30419 3364 30485 3365
rect 30419 3300 30420 3364
rect 30484 3300 30485 3364
rect 30419 3299 30485 3300
rect 21035 2684 21101 2685
rect 21035 2620 21036 2684
rect 21100 2620 21101 2684
rect 21035 2619 21101 2620
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1
transform 1 0 30268 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _0717_
timestamp 1
transform 1 0 2760 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0718_
timestamp 1
transform 1 0 3864 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0719_
timestamp 1
transform 1 0 3772 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _0720_
timestamp 1
transform 1 0 3036 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0721_
timestamp 1
transform 1 0 11500 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0722_
timestamp 1
transform 1 0 3864 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0723_
timestamp 1
transform -1 0 5520 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0724_
timestamp 1
transform 1 0 11500 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0725_
timestamp 1
transform 1 0 14996 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0726_
timestamp 1
transform 1 0 3772 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0727_
timestamp 1
transform 1 0 2668 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _0728_
timestamp 1
transform -1 0 9016 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _0729_
timestamp 1
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0730_
timestamp 1
transform 1 0 3772 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0731_
timestamp 1
transform 1 0 6992 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0732_
timestamp 1
transform 1 0 23828 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0733_
timestamp 1
transform 1 0 2852 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0734_
timestamp 1
transform 1 0 2576 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0735_
timestamp 1
transform 1 0 5336 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0736_
timestamp 1
transform -1 0 23368 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0737_
timestamp 1
transform 1 0 2852 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_1  _0738_
timestamp 1
transform 1 0 2208 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0739_
timestamp 1
transform 1 0 9568 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0740_
timestamp 1
transform 1 0 4692 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0741_
timestamp 1
transform 1 0 4784 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0742_
timestamp 1
transform 1 0 8740 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0743_
timestamp 1
transform 1 0 4784 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nor4b_1  _0744_
timestamp 1
transform -1 0 6164 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0745_
timestamp 1
transform 1 0 10396 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0746_
timestamp 1
transform 1 0 11316 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0747_
timestamp 1
transform 1 0 23368 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0748_
timestamp 1
transform 1 0 22908 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0749_
timestamp 1
transform 1 0 23460 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0750_
timestamp 1
transform 1 0 22724 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0751_
timestamp 1
transform 1 0 21896 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0752_
timestamp 1
transform 1 0 2116 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0753_
timestamp 1
transform 1 0 4692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0754_
timestamp 1
transform -1 0 11776 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0755_
timestamp 1
transform 1 0 11776 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0756_
timestamp 1
transform 1 0 10396 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0757_
timestamp 1
transform -1 0 15088 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0758_
timestamp 1
transform 1 0 9936 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0759_
timestamp 1
transform 1 0 12512 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0760_
timestamp 1
transform 1 0 21252 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0761_
timestamp 1
transform 1 0 22448 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0762_
timestamp 1
transform 1 0 20148 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0763_
timestamp 1
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0764_
timestamp 1
transform -1 0 10856 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0765_
timestamp 1
transform 1 0 11592 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0766_
timestamp 1
transform 1 0 12604 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0767_
timestamp 1
transform 1 0 18124 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0768_
timestamp 1
transform 1 0 18308 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0769_
timestamp 1
transform 1 0 18216 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0770_
timestamp 1
transform 1 0 12052 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0771_
timestamp 1
transform 1 0 10304 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0772_
timestamp 1
transform -1 0 12236 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0773_
timestamp 1
transform 1 0 11408 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0774_
timestamp 1
transform 1 0 9660 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0775_
timestamp 1
transform -1 0 24380 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0776_
timestamp 1
transform 1 0 5704 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0777_
timestamp 1
transform 1 0 10212 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0778_
timestamp 1
transform -1 0 14076 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0779_
timestamp 1
transform 1 0 8924 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0780_
timestamp 1
transform 1 0 6900 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0781_
timestamp 1
transform -1 0 21712 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0782_
timestamp 1
transform -1 0 28152 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0783_
timestamp 1
transform -1 0 9292 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0784_
timestamp 1
transform 1 0 5520 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0785_
timestamp 1
transform 1 0 7268 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0786_
timestamp 1
transform -1 0 9660 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0787_
timestamp 1
transform 1 0 7912 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0788_
timestamp 1
transform 1 0 27968 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0789_
timestamp 1
transform -1 0 9844 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0790_
timestamp 1
transform 1 0 28244 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0791_
timestamp 1
transform 1 0 2760 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0792_
timestamp 1
transform 1 0 2576 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0793_
timestamp 1
transform 1 0 5336 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0794_
timestamp 1
transform 1 0 2668 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0795_
timestamp 1
transform 1 0 7268 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_1  _0796_
timestamp 1
transform -1 0 4876 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0797_
timestamp 1
transform 1 0 2392 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0798_
timestamp 1
transform -1 0 23552 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0799_
timestamp 1
transform 1 0 26956 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0800_
timestamp 1
transform 1 0 4324 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0801_
timestamp 1
transform 1 0 4968 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0802_
timestamp 1
transform 1 0 6256 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0803_
timestamp 1
transform -1 0 17848 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0804_
timestamp 1
transform 1 0 4048 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0805_
timestamp 1
transform -1 0 25760 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0806_
timestamp 1
transform 1 0 26128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0807_
timestamp 1
transform -1 0 2944 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0808_
timestamp 1
transform 1 0 5244 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0809_
timestamp 1
transform 1 0 4968 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0810_
timestamp 1
transform 1 0 4048 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0811_
timestamp 1
transform 1 0 23460 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0812_
timestamp 1
transform 1 0 14076 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0813_
timestamp 1
transform 1 0 23828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0814_
timestamp 1
transform 1 0 5612 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0815_
timestamp 1
transform 1 0 2576 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0816_
timestamp 1
transform 1 0 2668 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0817_
timestamp 1
transform 1 0 3312 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0818_
timestamp 1
transform -1 0 23460 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0819_
timestamp 1
transform -1 0 6900 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0820_
timestamp 1
transform 1 0 17204 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0821_
timestamp 1
transform 1 0 26312 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0822_
timestamp 1
transform 1 0 10580 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0823_
timestamp 1
transform 1 0 5796 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0824_
timestamp 1
transform 1 0 6992 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0825_
timestamp 1
transform 1 0 15916 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0826_
timestamp 1
transform 1 0 25300 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0827_
timestamp 1
transform 1 0 8740 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0828_
timestamp 1
transform 1 0 9108 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0829_
timestamp 1
transform -1 0 22264 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0830_
timestamp 1
transform 1 0 25024 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0831_
timestamp 1
transform -1 0 4416 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0832_
timestamp 1
transform 1 0 2852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0833_
timestamp 1
transform 1 0 6532 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0834_
timestamp 1
transform -1 0 3496 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0835_
timestamp 1
transform -1 0 6624 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0836_
timestamp 1
transform -1 0 9476 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0837_
timestamp 1
transform -1 0 5060 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0838_
timestamp 1
transform 1 0 6808 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0839_
timestamp 1
transform 1 0 17296 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0840_
timestamp 1
transform 1 0 16928 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0841_
timestamp 1
transform 1 0 5244 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0842_
timestamp 1
transform 1 0 5428 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0843_
timestamp 1
transform 1 0 14996 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0844_
timestamp 1
transform 1 0 6532 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0845_
timestamp 1
transform 1 0 3956 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0846_
timestamp 1
transform 1 0 17112 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0847_
timestamp 1
transform 1 0 6992 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0848_
timestamp 1
transform 1 0 7176 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0849_
timestamp 1
transform 1 0 5336 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0850_
timestamp 1
transform 1 0 4232 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0851_
timestamp 1
transform -1 0 14628 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0852_
timestamp 1
transform -1 0 9568 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0853_
timestamp 1
transform 1 0 18032 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0854_
timestamp 1
transform 1 0 3588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_1  _0855_
timestamp 1
transform -1 0 4416 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0856_
timestamp 1
transform 1 0 6900 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0857_
timestamp 1
transform 1 0 4324 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0858_
timestamp 1
transform 1 0 13064 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0859_
timestamp 1
transform 1 0 6532 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0860_
timestamp 1
transform 1 0 8556 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0861_
timestamp 1
transform 1 0 11500 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0862_
timestamp 1
transform 1 0 16928 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0863_
timestamp 1
transform 1 0 12236 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0864_
timestamp 1
transform -1 0 9660 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0865_
timestamp 1
transform 1 0 8556 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0866_
timestamp 1
transform 1 0 14996 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0867_
timestamp 1
transform 1 0 7912 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0868_
timestamp 1
transform 1 0 7912 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0869_
timestamp 1
transform -1 0 8924 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0870_
timestamp 1
transform 1 0 14260 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0871_
timestamp 1
transform 1 0 28060 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _0872_
timestamp 1
transform 1 0 3588 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0873_
timestamp 1
transform 1 0 2944 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0874_
timestamp 1
transform 1 0 9476 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0875_
timestamp 1
transform 1 0 7176 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0876_
timestamp 1
transform 1 0 16008 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0877_
timestamp 1
transform 1 0 10120 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0878_
timestamp 1
transform 1 0 8188 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0879_
timestamp 1
transform 1 0 15088 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0880_
timestamp 1
transform 1 0 15364 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0881_
timestamp 1
transform 1 0 9384 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0882_
timestamp 1
transform -1 0 9936 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0883_
timestamp 1
transform 1 0 13524 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0884_
timestamp 1
transform 1 0 9016 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0885_
timestamp 1
transform 1 0 10120 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0886_
timestamp 1
transform 1 0 21436 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _0887_
timestamp 1
transform -1 0 22356 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0888_
timestamp 1
transform 1 0 9200 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0889_
timestamp 1
transform -1 0 9568 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0890_
timestamp 1
transform 1 0 7268 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0891_
timestamp 1
transform 1 0 8556 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0892_
timestamp 1
transform 1 0 24840 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0893_
timestamp 1
transform 1 0 15364 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0894_
timestamp 1
transform 1 0 26128 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0895_
timestamp 1
transform 1 0 2024 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0896_
timestamp 1
transform 1 0 5612 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0897_
timestamp 1
transform 1 0 6164 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0898_
timestamp 1
transform 1 0 4692 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0899_
timestamp 1
transform -1 0 6072 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0900_
timestamp 1
transform 1 0 19228 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0901_
timestamp 1
transform 1 0 2484 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0902_
timestamp 1
transform 1 0 5704 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0903_
timestamp 1
transform -1 0 24104 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0904_
timestamp 1
transform 1 0 25760 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0905_
timestamp 1
transform 1 0 2576 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0906_
timestamp 1
transform 1 0 1932 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0907_
timestamp 1
transform 1 0 7820 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0908_
timestamp 1
transform 1 0 6348 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0909_
timestamp 1
transform 1 0 3956 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0910_
timestamp 1
transform 1 0 16928 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0911_
timestamp 1
transform 1 0 19872 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0912_
timestamp 1
transform 1 0 7084 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0913_
timestamp 1
transform 1 0 4784 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0914_
timestamp 1
transform 1 0 6348 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0915_
timestamp 1
transform 1 0 10580 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0916_
timestamp 1
transform 1 0 3864 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0917_
timestamp 1
transform -1 0 3680 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0918_
timestamp 1
transform -1 0 10396 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0919_
timestamp 1
transform 1 0 10212 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0920_
timestamp 1
transform -1 0 26496 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0921_
timestamp 1
transform 1 0 7820 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0922_
timestamp 1
transform 1 0 5152 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0923_
timestamp 1
transform 1 0 7176 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0924_
timestamp 1
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0925_
timestamp 1
transform 1 0 11132 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0926_
timestamp 1
transform 1 0 15180 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0927_
timestamp 1
transform 1 0 16008 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0928_
timestamp 1
transform 1 0 11500 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0929_
timestamp 1
transform 1 0 3312 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0930_
timestamp 1
transform 1 0 6348 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0931_
timestamp 1
transform 1 0 11960 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0932_
timestamp 1
transform 1 0 5060 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0933_
timestamp 1
transform 1 0 8924 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0934_
timestamp 1
transform -1 0 10396 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0935_
timestamp 1
transform 1 0 19688 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0936_
timestamp 1
transform 1 0 12420 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0937_
timestamp 1
transform 1 0 9752 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0938_
timestamp 1
transform -1 0 20884 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0939_
timestamp 1
transform 1 0 6624 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0940_
timestamp 1
transform 1 0 4416 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0941_
timestamp 1
transform 1 0 15824 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0942_
timestamp 1
transform 1 0 19504 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0943_
timestamp 1
transform 1 0 14168 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0944_
timestamp 1
transform 1 0 23276 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0945_
timestamp 1
transform 1 0 8556 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0946_
timestamp 1
transform 1 0 11316 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0947_
timestamp 1
transform 1 0 10488 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0948_
timestamp 1
transform -1 0 7728 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0949_
timestamp 1
transform 1 0 24840 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0950_
timestamp 1
transform 1 0 9292 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0951_
timestamp 1
transform 1 0 11776 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0952_
timestamp 1
transform -1 0 18860 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0953_
timestamp 1
transform 1 0 6348 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0954_
timestamp 1
transform 1 0 7912 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0955_
timestamp 1
transform 1 0 17572 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0956_
timestamp 1
transform 1 0 22264 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0957_
timestamp 1
transform 1 0 25576 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0958_
timestamp 1
transform 1 0 8188 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0959_
timestamp 1
transform 1 0 10764 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0960_
timestamp 1
transform 1 0 15456 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0961_
timestamp 1
transform 1 0 5060 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0962_
timestamp 1
transform 1 0 4784 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0963_
timestamp 1
transform 1 0 16100 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0964_
timestamp 1
transform 1 0 6348 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0965_
timestamp 1
transform 1 0 8188 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0966_
timestamp 1
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0967_
timestamp 1
transform 1 0 4140 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0968_
timestamp 1
transform 1 0 7544 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0969_
timestamp 1
transform 1 0 4508 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0970_
timestamp 1
transform 1 0 6072 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0971_
timestamp 1
transform 1 0 20056 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0972_
timestamp 1
transform 1 0 19872 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0973_
timestamp 1
transform -1 0 4416 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0974_
timestamp 1
transform -1 0 7912 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0975_
timestamp 1
transform 1 0 16652 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0976_
timestamp 1
transform 1 0 3772 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0977_
timestamp 1
transform 1 0 3772 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0978_
timestamp 1
transform -1 0 2760 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0979_
timestamp 1
transform 1 0 14076 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0980_
timestamp 1
transform 1 0 10948 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0981_
timestamp 1
transform 1 0 15916 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0982_
timestamp 1
transform 1 0 27600 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0983_
timestamp 1
transform -1 0 28980 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0984_
timestamp 1
transform -1 0 11684 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0985_
timestamp 1
transform 1 0 14812 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0986_
timestamp 1
transform 1 0 24932 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0987_
timestamp 1
transform -1 0 28888 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0988_
timestamp 1
transform 1 0 26956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _0989_
timestamp 1
transform 1 0 27692 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0990_
timestamp 1
transform 1 0 25484 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0991_
timestamp 1
transform 1 0 16744 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0992_
timestamp 1
transform 1 0 26680 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0993_
timestamp 1
transform 1 0 27140 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _0994_
timestamp 1
transform -1 0 29348 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0995_
timestamp 1
transform -1 0 11132 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0996_
timestamp 1
transform 1 0 11592 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0997_
timestamp 1
transform -1 0 18032 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0998_
timestamp 1
transform 1 0 17296 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0999_
timestamp 1
transform 1 0 17756 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1000_
timestamp 1
transform 1 0 12880 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1001_
timestamp 1
transform 1 0 10028 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1002_
timestamp 1
transform 1 0 13708 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1003_
timestamp 1
transform 1 0 24380 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1004_
timestamp 1
transform 1 0 12052 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1005_
timestamp 1
transform 1 0 12972 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1006_
timestamp 1
transform 1 0 12696 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1007_
timestamp 1
transform 1 0 12788 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1008_
timestamp 1
transform -1 0 19044 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1009_
timestamp 1
transform 1 0 12788 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1010_
timestamp 1
transform 1 0 12696 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1011_
timestamp 1
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1012_
timestamp 1
transform 1 0 13524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1013_
timestamp 1
transform -1 0 13616 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1014_
timestamp 1
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1015_
timestamp 1
transform 1 0 18400 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1016_
timestamp 1
transform 1 0 18216 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _1017_
timestamp 1
transform 1 0 16376 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1018_
timestamp 1
transform 1 0 25668 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1019_
timestamp 1
transform 1 0 16928 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1020_
timestamp 1
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1021_
timestamp 1
transform 1 0 18400 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1022_
timestamp 1
transform 1 0 26404 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1023_
timestamp 1
transform 1 0 16376 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1024_
timestamp 1
transform 1 0 13340 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1025_
timestamp 1
transform 1 0 13340 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1026_
timestamp 1
transform 1 0 25300 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1027_
timestamp 1
transform 1 0 18676 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1028_
timestamp 1
transform -1 0 19688 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1029_
timestamp 1
transform 1 0 23552 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1030_
timestamp 1
transform 1 0 28428 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1031_
timestamp 1
transform 1 0 20240 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1032_
timestamp 1
transform 1 0 29072 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1033_
timestamp 1
transform 1 0 28888 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1034_
timestamp 1
transform 1 0 29532 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1035_
timestamp 1
transform -1 0 25484 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1036_
timestamp 1
transform 1 0 18216 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1037_
timestamp 1
transform 1 0 22540 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1038_
timestamp 1
transform 1 0 22632 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1039_
timestamp 1
transform 1 0 23920 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1040_
timestamp 1
transform 1 0 23644 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1041_
timestamp 1
transform 1 0 18400 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1042_
timestamp 1
transform 1 0 24380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1043_
timestamp 1
transform 1 0 25576 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1044_
timestamp 1
transform 1 0 25668 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1045_
timestamp 1
transform 1 0 26128 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1046_
timestamp 1
transform 1 0 30176 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1047_
timestamp 1
transform 1 0 29900 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1048_
timestamp 1
transform 1 0 20332 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1049_
timestamp 1
transform 1 0 14352 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1050_
timestamp 1
transform -1 0 14076 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1051_
timestamp 1
transform 1 0 20976 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1052_
timestamp 1
transform 1 0 14444 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1053_
timestamp 1
transform 1 0 16008 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1054_
timestamp 1
transform -1 0 7176 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1055_
timestamp 1
transform -1 0 7820 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1056_
timestamp 1
transform 1 0 9844 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1057_
timestamp 1
transform -1 0 10304 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1058_
timestamp 1
transform 1 0 9292 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1059_
timestamp 1
transform -1 0 10120 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1060_
timestamp 1
transform -1 0 17204 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1061_
timestamp 1
transform -1 0 9476 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1062_
timestamp 1
transform -1 0 17480 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1063_
timestamp 1
transform -1 0 10304 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1064_
timestamp 1
transform 1 0 8188 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1065_
timestamp 1
transform 1 0 7912 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1066_
timestamp 1
transform -1 0 9660 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1067_
timestamp 1
transform 1 0 9200 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1068_
timestamp 1
transform 1 0 16560 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1069_
timestamp 1
transform 1 0 18124 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1070_
timestamp 1
transform -1 0 17940 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1071_
timestamp 1
transform 1 0 18676 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1072_
timestamp 1
transform -1 0 20424 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1073_
timestamp 1
transform 1 0 26404 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1074_
timestamp 1
transform 1 0 18584 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1075_
timestamp 1
transform 1 0 27692 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1076_
timestamp 1
transform 1 0 27876 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1077_
timestamp 1
transform 1 0 26404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1078_
timestamp 1
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1079_
timestamp 1
transform 1 0 16928 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1080_
timestamp 1
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1081_
timestamp 1
transform 1 0 28612 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1082_
timestamp 1
transform 1 0 17940 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1083_
timestamp 1
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1084_
timestamp 1
transform 1 0 18400 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1085_
timestamp 1
transform 1 0 29532 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1086_
timestamp 1
transform 1 0 29716 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1087_
timestamp 1
transform -1 0 21160 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1088_
timestamp 1
transform 1 0 21804 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1089_
timestamp 1
transform -1 0 13708 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1090_
timestamp 1
transform 1 0 25024 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1091_
timestamp 1
transform 1 0 17296 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1092_
timestamp 1
transform 1 0 26036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1093_
timestamp 1
transform 1 0 19596 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1094_
timestamp 1
transform 1 0 14352 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1095_
timestamp 1
transform 1 0 20056 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1096_
timestamp 1
transform 1 0 26588 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1097_
timestamp 1
transform 1 0 19228 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1098_
timestamp 1
transform 1 0 19780 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1099_
timestamp 1
transform 1 0 18676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1100_
timestamp 1
transform 1 0 20608 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1101_
timestamp 1
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1102_
timestamp 1
transform 1 0 25484 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1103_
timestamp 1
transform 1 0 28796 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1104_
timestamp 1
transform 1 0 14720 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1105_
timestamp 1
transform -1 0 13984 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1106_
timestamp 1
transform 1 0 14996 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1107_
timestamp 1
transform 1 0 21068 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1108_
timestamp 1
transform -1 0 22908 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1109_
timestamp 1
transform -1 0 22540 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1110_
timestamp 1
transform -1 0 24288 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1111_
timestamp 1
transform -1 0 22448 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1112_
timestamp 1
transform 1 0 21804 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1113_
timestamp 1
transform -1 0 19688 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1114_
timestamp 1
transform 1 0 20240 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1115_
timestamp 1
transform 1 0 20240 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1116_
timestamp 1
transform -1 0 7820 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1117_
timestamp 1
transform 1 0 7360 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1118_
timestamp 1
transform -1 0 12144 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1119_
timestamp 1
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1120_
timestamp 1
transform 1 0 6624 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1121_
timestamp 1
transform -1 0 15180 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1122_
timestamp 1
transform -1 0 8648 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1123_
timestamp 1
transform 1 0 20700 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1124_
timestamp 1
transform -1 0 21344 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1125_
timestamp 1
transform 1 0 23736 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1126_
timestamp 1
transform 1 0 26588 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1127_
timestamp 1
transform -1 0 6900 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1128_
timestamp 1
transform 1 0 7544 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1129_
timestamp 1
transform 1 0 10764 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1
transform -1 0 6164 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1131_
timestamp 1
transform 1 0 19780 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1132_
timestamp 1
transform 1 0 19964 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1133_
timestamp 1
transform 1 0 15824 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1134_
timestamp 1
transform 1 0 24932 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1135_
timestamp 1
transform -1 0 27692 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1136_
timestamp 1
transform 1 0 25668 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1137_
timestamp 1
transform 1 0 20424 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1138_
timestamp 1
transform 1 0 26220 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1139_
timestamp 1
transform 1 0 23552 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1140_
timestamp 1
transform 1 0 23644 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1141_
timestamp 1
transform 1 0 20240 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1142_
timestamp 1
transform 1 0 24196 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1143_
timestamp 1
transform -1 0 27876 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1144_
timestamp 1
transform -1 0 25300 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1145_
timestamp 1
transform 1 0 24472 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1146_
timestamp 1
transform 1 0 28152 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1147_
timestamp 1
transform -1 0 10580 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1148_
timestamp 1
transform -1 0 17020 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1149_
timestamp 1
transform -1 0 11960 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1150_
timestamp 1
transform -1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1151_
timestamp 1
transform -1 0 21620 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1152_
timestamp 1
transform 1 0 17204 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1153_
timestamp 1
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1154_
timestamp 1
transform 1 0 17204 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1155_
timestamp 1
transform -1 0 19228 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1156_
timestamp 1
transform 1 0 16008 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1157_
timestamp 1
transform -1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1158_
timestamp 1
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1159_
timestamp 1
transform 1 0 21528 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1160_
timestamp 1
transform 1 0 22080 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1161_
timestamp 1
transform 1 0 21896 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1162_
timestamp 1
transform 1 0 9016 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1163_
timestamp 1
transform 1 0 9384 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1164_
timestamp 1
transform 1 0 9200 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1165_
timestamp 1
transform 1 0 8740 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1166_
timestamp 1
transform 1 0 9936 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1167_
timestamp 1
transform 1 0 23184 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1168_
timestamp 1
transform 1 0 23552 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1169_
timestamp 1
transform -1 0 23736 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1170_
timestamp 1
transform -1 0 23368 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1171_
timestamp 1
transform 1 0 22816 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1172_
timestamp 1
transform 1 0 26680 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1173_
timestamp 1
transform 1 0 12144 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1174_
timestamp 1
transform 1 0 22172 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1175_
timestamp 1
transform 1 0 22632 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1176_
timestamp 1
transform 1 0 23368 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1177_
timestamp 1
transform 1 0 23736 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1178_
timestamp 1
transform 1 0 23920 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1179_
timestamp 1
transform -1 0 4048 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1180_
timestamp 1
transform -1 0 5060 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1181_
timestamp 1
transform 1 0 25852 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1182_
timestamp 1
transform 1 0 27876 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1183_
timestamp 1
transform 1 0 29716 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1184_
timestamp 1
transform -1 0 3588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1185_
timestamp 1
transform 1 0 14996 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1186_
timestamp 1
transform 1 0 14720 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1187_
timestamp 1
transform 1 0 15272 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1188_
timestamp 1
transform 1 0 15732 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1189_
timestamp 1
transform 1 0 27140 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1190_
timestamp 1
transform 1 0 29716 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1191_
timestamp 1
transform 1 0 29992 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1192_
timestamp 1
transform 1 0 30728 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1193_
timestamp 1
transform 1 0 22540 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1194_
timestamp 1
transform 1 0 28152 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1195_
timestamp 1
transform 1 0 18860 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1196_
timestamp 1
transform 1 0 27600 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1197_
timestamp 1
transform 1 0 24472 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1198_
timestamp 1
transform 1 0 28704 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1199_
timestamp 1
transform 1 0 11684 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1200_
timestamp 1
transform 1 0 13156 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1201_
timestamp 1
transform 1 0 16744 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1202_
timestamp 1
transform 1 0 19688 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1203_
timestamp 1
transform 1 0 13064 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1204_
timestamp 1
transform 1 0 23092 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1205_
timestamp 1
transform 1 0 23552 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1206_
timestamp 1
transform 1 0 29532 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1207_
timestamp 1
transform 1 0 29624 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1208_
timestamp 1
transform -1 0 16468 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1209_
timestamp 1
transform 1 0 11592 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1210_
timestamp 1
transform 1 0 15732 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1211_
timestamp 1
transform 1 0 15272 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1212_
timestamp 1
transform -1 0 9660 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1213_
timestamp 1
transform 1 0 9752 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1214_
timestamp 1
transform 1 0 12144 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1215_
timestamp 1
transform 1 0 11592 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1216_
timestamp 1
transform -1 0 11960 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1217_
timestamp 1
transform 1 0 11960 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1218_
timestamp 1
transform -1 0 17020 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1219_
timestamp 1
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1220_
timestamp 1
transform 1 0 30636 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1221_
timestamp 1
transform 1 0 10764 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1222_
timestamp 1
transform 1 0 20884 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1223_
timestamp 1
transform 1 0 20884 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1224_
timestamp 1
transform 1 0 15272 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1225_
timestamp 1
transform 1 0 21252 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1226_
timestamp 1
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1227_
timestamp 1
transform 1 0 16008 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1228_
timestamp 1
transform -1 0 22632 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1229_
timestamp 1
transform 1 0 22356 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1230_
timestamp 1
transform -1 0 23092 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1231_
timestamp 1
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1232_
timestamp 1
transform 1 0 12236 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1233_
timestamp 1
transform 1 0 21712 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1234_
timestamp 1
transform -1 0 22448 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1235_
timestamp 1
transform 1 0 21896 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1236_
timestamp 1
transform 1 0 22264 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1237_
timestamp 1
transform 1 0 27508 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1238_
timestamp 1
transform -1 0 25024 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1239_
timestamp 1
transform -1 0 12604 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1240_
timestamp 1
transform 1 0 17756 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1241_
timestamp 1
transform -1 0 24196 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1242_
timestamp 1
transform 1 0 19228 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1243_
timestamp 1
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1244_
timestamp 1
transform 1 0 20056 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1245_
timestamp 1
transform 1 0 12512 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1246_
timestamp 1
transform 1 0 25760 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1247_
timestamp 1
transform 1 0 21988 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1248_
timestamp 1
transform 1 0 13432 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1249_
timestamp 1
transform 1 0 23828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1250_
timestamp 1
transform 1 0 25852 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1251_
timestamp 1
transform 1 0 30636 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1252_
timestamp 1
transform 1 0 19412 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1253_
timestamp 1
transform 1 0 24196 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1254_
timestamp 1
transform -1 0 10120 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1255_
timestamp 1
transform 1 0 7820 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1256_
timestamp 1
transform -1 0 8464 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1257_
timestamp 1
transform -1 0 11132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1258_
timestamp 1
transform -1 0 11040 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1259_
timestamp 1
transform 1 0 10120 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1260_
timestamp 1
transform 1 0 20516 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1261_
timestamp 1
transform 1 0 22724 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1262_
timestamp 1
transform 1 0 23736 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1263_
timestamp 1
transform 1 0 24380 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1264_
timestamp 1
transform 1 0 30912 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1265_
timestamp 1
transform 1 0 12144 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1266_
timestamp 1
transform 1 0 14720 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1267_
timestamp 1
transform 1 0 14444 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1268_
timestamp 1
transform 1 0 15088 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1269_
timestamp 1
transform 1 0 13800 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1270_
timestamp 1
transform 1 0 14904 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1271_
timestamp 1
transform 1 0 15456 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1272_
timestamp 1
transform 1 0 20148 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1273_
timestamp 1
transform -1 0 24288 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1274_
timestamp 1
transform -1 0 24288 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1275_
timestamp 1
transform 1 0 15916 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1276_
timestamp 1
transform 1 0 16652 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1277_
timestamp 1
transform 1 0 13984 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1278_
timestamp 1
transform -1 0 20884 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1279_
timestamp 1
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1280_
timestamp 1
transform -1 0 14904 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1281_
timestamp 1
transform 1 0 13432 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1282_
timestamp 1
transform 1 0 14352 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1283_
timestamp 1
transform 1 0 21804 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1284_
timestamp 1
transform 1 0 19688 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1285_
timestamp 1
transform 1 0 26036 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1286_
timestamp 1
transform 1 0 21988 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1287_
timestamp 1
transform -1 0 28152 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1288_
timestamp 1
transform 1 0 8648 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1289_
timestamp 1
transform 1 0 9108 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1290_
timestamp 1
transform 1 0 22080 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1291_
timestamp 1
transform 1 0 22264 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1292_
timestamp 1
transform 1 0 23552 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1293_
timestamp 1
transform 1 0 6992 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1294_
timestamp 1
transform 1 0 20976 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1295_
timestamp 1
transform 1 0 25300 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1296_
timestamp 1
transform 1 0 27692 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1297_
timestamp 1
transform 1 0 26312 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1298_
timestamp 1
transform 1 0 27692 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1299_
timestamp 1
transform 1 0 28428 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1300_
timestamp 1
transform 1 0 14168 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1301_
timestamp 1
transform 1 0 7452 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1302_
timestamp 1
transform 1 0 14444 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1303_
timestamp 1
transform -1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1304_
timestamp 1
transform 1 0 14904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1305_
timestamp 1
transform 1 0 28888 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1306_
timestamp 1
transform 1 0 29532 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1307_
timestamp 1
transform 1 0 28152 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1308_
timestamp 1
transform 1 0 18308 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1309_
timestamp 1
transform -1 0 20056 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1310_
timestamp 1
transform -1 0 30452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1311_
timestamp 1
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1312_
timestamp 1
transform 1 0 18124 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1313_
timestamp 1
transform 1 0 18952 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1314_
timestamp 1
transform 1 0 18216 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1315_
timestamp 1
transform 1 0 12604 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1316_
timestamp 1
transform 1 0 17664 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1317_
timestamp 1
transform 1 0 18952 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1318_
timestamp 1
transform 1 0 29624 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1319_
timestamp 1
transform 1 0 30912 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1320_
timestamp 1
transform 1 0 22908 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1321_
timestamp 1
transform 1 0 13800 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1322_
timestamp 1
transform 1 0 16744 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1323_
timestamp 1
transform 1 0 17296 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1324_
timestamp 1
transform 1 0 17848 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1325_
timestamp 1
transform -1 0 18768 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1326_
timestamp 1
transform 1 0 18124 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1327_
timestamp 1
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1328_
timestamp 1
transform 1 0 19780 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1329_
timestamp 1
transform 1 0 22356 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1330_
timestamp 1
transform 1 0 30176 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1331_
timestamp 1
transform -1 0 11408 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1332_
timestamp 1
transform 1 0 11592 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1333_
timestamp 1
transform 1 0 10580 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1334_
timestamp 1
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1335_
timestamp 1
transform 1 0 12144 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1336_
timestamp 1
transform 1 0 19780 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1337_
timestamp 1
transform 1 0 20424 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1338_
timestamp 1
transform 1 0 25760 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1339_
timestamp 1
transform 1 0 21528 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1340_
timestamp 1
transform 1 0 21528 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1341_
timestamp 1
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1342_
timestamp 1
transform -1 0 22448 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1343_
timestamp 1
transform -1 0 21436 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1344_
timestamp 1
transform 1 0 20792 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1345_
timestamp 1
transform 1 0 23460 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1346_
timestamp 1
transform 1 0 21988 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1347_
timestamp 1
transform 1 0 23368 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1348_
timestamp 1
transform 1 0 23000 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1349_
timestamp 1
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1350_
timestamp 1
transform 1 0 23920 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1351_
timestamp 1
transform 1 0 24656 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1352_
timestamp 1
transform 1 0 25484 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1353_
timestamp 1
transform 1 0 26772 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1354_
timestamp 1
transform 1 0 30176 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1355_
timestamp 1
transform -1 0 17480 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1356_
timestamp 1
transform 1 0 15824 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1357_
timestamp 1
transform 1 0 17204 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1358_
timestamp 1
transform 1 0 17020 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1359_
timestamp 1
transform 1 0 15824 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1360_
timestamp 1
transform 1 0 16652 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1361_
timestamp 1
transform 1 0 17480 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1362_
timestamp 1
transform 1 0 27600 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1363_
timestamp 1
transform 1 0 29532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1364_
timestamp 1
transform 1 0 22356 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1365_
timestamp 1
transform 1 0 30084 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1366_
timestamp 1
transform -1 0 22356 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1367_
timestamp 1
transform 1 0 21804 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1368_
timestamp 1
transform 1 0 28980 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1369_
timestamp 1
transform 1 0 29532 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1370_
timestamp 1
transform 1 0 29716 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1371_
timestamp 1
transform 1 0 30452 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1372_
timestamp 1
transform 1 0 20608 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1373_
timestamp 1
transform -1 0 21160 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1374_
timestamp 1
transform 1 0 19964 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1375_
timestamp 1
transform -1 0 5520 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1376_
timestamp 1
transform 1 0 5520 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1377_
timestamp 1
transform 1 0 5520 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1378_
timestamp 1
transform 1 0 6072 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1379_
timestamp 1
transform 1 0 17848 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1380_
timestamp 1
transform 1 0 14352 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1381_
timestamp 1
transform 1 0 17940 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1382_
timestamp 1
transform 1 0 20792 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1383_
timestamp 1
transform 1 0 30636 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1384_
timestamp 1
transform 1 0 11684 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1385_
timestamp 1
transform 1 0 11960 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1386_
timestamp 1
transform 1 0 12512 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1387_
timestamp 1
transform 1 0 12788 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1388_
timestamp 1
transform -1 0 14812 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1389_
timestamp 1
transform 1 0 13248 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1390_
timestamp 1
transform 1 0 14076 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1391_
timestamp 1
transform 1 0 14444 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1392_
timestamp 1
transform -1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1393_
timestamp 1
transform 1 0 15272 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1394_
timestamp 1
transform 1 0 28796 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1395_
timestamp 1
transform 1 0 29624 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1396_
timestamp 1
transform 1 0 17940 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1397_
timestamp 1
transform -1 0 20240 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1398_
timestamp 1
transform -1 0 4692 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1399_
timestamp 1
transform 1 0 3772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1400_
timestamp 1
transform -1 0 20424 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1401_
timestamp 1
transform 1 0 19964 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1402_
timestamp 1
transform 1 0 27048 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1403_
timestamp 1
transform 1 0 23552 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1404_
timestamp 1
transform 1 0 16744 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1405_
timestamp 1
transform 1 0 26956 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1406_
timestamp 1
transform 1 0 30176 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1407_
timestamp 1
transform 1 0 30636 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1408_
timestamp 1
transform 1 0 24932 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1409_
timestamp 1
transform -1 0 27140 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1410_
timestamp 1
transform 1 0 25576 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1411_
timestamp 1
transform 1 0 28152 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1412_
timestamp 1
transform 1 0 26772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1413_
timestamp 1
transform 1 0 26036 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1414_
timestamp 1
transform -1 0 28152 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1415_
timestamp 1
transform 1 0 27600 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1416_
timestamp 1
transform 1 0 30912 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1417_
timestamp 1
transform 1 0 27876 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1418_
timestamp 1
transform 1 0 25208 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1419_
timestamp 1
transform 1 0 24196 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1420_
timestamp 1
transform 1 0 25576 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1421_
timestamp 1
transform 1 0 25484 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1422_
timestamp 1
transform 1 0 26956 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1423_
timestamp 1
transform 1 0 28152 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1424_
timestamp 1
transform 1 0 30912 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1425_
timestamp 1
transform 1 0 26220 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1426_
timestamp 1
transform 1 0 27876 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1427_
timestamp 1
transform 1 0 28704 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1428_
timestamp 1
transform 1 0 31004 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1429_
timestamp 1
transform 1 0 28152 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1430_
timestamp 1
transform 1 0 30912 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1431_
timestamp 1
transform 1 0 16192 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1432_
timestamp 1
transform 1 0 1380 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1433_
timestamp 1
transform 1 0 1380 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1434_
timestamp 1
transform 1 0 1380 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1435_
timestamp 1
transform 1 0 1380 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1436_
timestamp 1
transform 1 0 1380 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1437_
timestamp 1
transform 1 0 1380 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1438_
timestamp 1
transform 1 0 1380 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1439_
timestamp 1
transform 1 0 1380 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1440_
timestamp 1
transform -1 0 32016 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1441_
timestamp 1
transform -1 0 20332 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1442_
timestamp 1
transform 1 0 30084 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1443_
timestamp 1
transform 1 0 17388 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1444_
timestamp 1
transform 1 0 30360 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1445_
timestamp 1
transform 1 0 30544 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1446_
timestamp 1
transform 1 0 20240 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1447_
timestamp 1
transform 1 0 24840 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1448_
timestamp 1
transform 1 0 21988 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1449_
timestamp 1
transform -1 0 25852 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1450_
timestamp 1
transform 1 0 30544 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1451_
timestamp 1
transform 1 0 30268 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1452_
timestamp 1
transform 1 0 31096 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1453_
timestamp 1
transform 1 0 22172 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1454_
timestamp 1
transform 1 0 31096 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1455_
timestamp 1
transform 1 0 31096 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1456_
timestamp 1
transform -1 0 17388 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1457_
timestamp 1
transform 1 0 23828 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1458_
timestamp 1
transform 1 0 30176 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1459_
timestamp 1
transform 1 0 30544 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1460_
timestamp 1
transform 1 0 30820 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1461_
timestamp 1
transform -1 0 21988 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1462_
timestamp 1
transform 1 0 31096 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1463_
timestamp 1
transform 1 0 31096 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1464_
timestamp 1
transform 1 0 31096 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1465_
timestamp 1
transform 1 0 29532 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1466_
timestamp 1
transform 1 0 31096 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1467_
timestamp 1
transform 1 0 31096 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1468_
timestamp 1
transform 1 0 30544 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1469_
timestamp 1
transform 1 0 30544 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1470_
timestamp 1
transform 1 0 30544 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1471_
timestamp 1
transform 1 0 16652 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform 1 0 23368 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1
transform 1 0 12144 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1
transform -1 0 19412 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1
transform -1 0 25116 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1
transform 1 0 24012 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1
transform 1 0 28244 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1
transform -1 0 17756 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1
transform -1 0 27692 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1
transform 1 0 19228 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1
transform -1 0 23092 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1
transform -1 0 12788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1
transform 1 0 22540 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1
transform -1 0 24932 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1
transform -1 0 14352 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1
transform -1 0 30176 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1
transform -1 0 15732 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1
transform -1 0 16560 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1
transform 1 0 24564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1
transform 1 0 22448 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1
transform 1 0 20056 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1
transform -1 0 17204 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1
transform 1 0 28612 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1
transform 1 0 23736 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1
transform -1 0 16468 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1
transform 1 0 23552 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1
transform -1 0 22264 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1
transform -1 0 22080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1
transform 1 0 29440 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1
transform -1 0 18124 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1
transform -1 0 17940 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1
transform 1 0 19780 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1
transform -1 0 22724 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1
transform -1 0 12512 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1
transform 1 0 15916 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1
transform 1 0 14628 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1
transform -1 0 18860 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1
transform -1 0 16928 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1
transform 1 0 25944 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1
transform 1 0 18584 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1
transform -1 0 23184 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1
transform -1 0 26404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1
transform 1 0 29900 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1
transform 1 0 26956 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1
transform 1 0 27784 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_47
timestamp 1
transform 1 0 20332 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_48
timestamp 1
transform 1 0 16928 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_49
timestamp 1
transform -1 0 23644 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_50
timestamp 1
transform -1 0 27324 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_51
timestamp 1
transform -1 0 23736 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_52
timestamp 1
transform -1 0 22908 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_53
timestamp 1
transform -1 0 18308 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk0
timestamp 1
transform 1 0 16652 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk0
timestamp 1
transform -1 0 12144 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk0
timestamp 1
transform -1 0 21068 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk0
timestamp 1
transform 1 0 24380 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk0
timestamp 1
transform 1 0 24380 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinv_4  clkload0
timestamp 1
transform 1 0 10304 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload1
timestamp 1
transform 1 0 18492 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__bufinv_16  clkload2
timestamp 1
transform -1 0 26496 0 -1 18496
box -38 -48 2246 592
use sky130_fd_sc_hd__conb_1  cust_rom0_630
timestamp 1
transform -1 0 29992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout41
timestamp 1
transform -1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout42
timestamp 1
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout43
timestamp 1
transform -1 0 30452 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout44
timestamp 1
transform -1 0 30728 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout45
timestamp 1
transform -1 0 31004 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout46
timestamp 1
transform -1 0 30636 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout47
timestamp 1
transform 1 0 31188 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout48
timestamp 1
transform -1 0 30820 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout49
timestamp 1
transform -1 0 31096 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout50
timestamp 1
transform 1 0 30268 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout51
timestamp 1
transform 1 0 32292 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout52
timestamp 1
transform -1 0 30820 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout53
timestamp 1
transform 1 0 30176 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout54
timestamp 1
transform -1 0 31096 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout55
timestamp 1
transform -1 0 21988 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout56
timestamp 1
transform 1 0 31096 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout58
timestamp 1
transform 1 0 9016 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout59
timestamp 1
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout60
timestamp 1
transform -1 0 17756 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout61
timestamp 1
transform -1 0 11408 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout62
timestamp 1
transform -1 0 8648 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout63
timestamp 1
transform 1 0 24840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout64
timestamp 1
transform -1 0 20056 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout65
timestamp 1
transform -1 0 15456 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout66
timestamp 1
transform 1 0 12696 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout67
timestamp 1
transform -1 0 13064 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout68
timestamp 1
transform 1 0 12328 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout69
timestamp 1
transform -1 0 8648 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout70
timestamp 1
transform 1 0 16284 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout71
timestamp 1
transform 1 0 8004 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout72
timestamp 1
transform -1 0 2760 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout73
timestamp 1
transform -1 0 16468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout74
timestamp 1
transform -1 0 12328 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout75
timestamp 1
transform 1 0 11960 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout76
timestamp 1
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout77
timestamp 1
transform -1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout78
timestamp 1
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout79
timestamp 1
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout80
timestamp 1
transform -1 0 9844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout81
timestamp 1
transform 1 0 19688 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout82
timestamp 1
transform 1 0 11132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout83
timestamp 1
transform -1 0 11408 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout84
timestamp 1
transform -1 0 20608 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout85
timestamp 1
transform -1 0 20148 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout86
timestamp 1
transform -1 0 9844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout87
timestamp 1
transform 1 0 9108 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout88
timestamp 1
transform 1 0 6532 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout89
timestamp 1
transform -1 0 20332 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout90
timestamp 1
transform 1 0 5888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout91
timestamp 1
transform -1 0 16928 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout92
timestamp 1
transform 1 0 6808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout93
timestamp 1
transform 1 0 4692 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout94
timestamp 1
transform 1 0 15548 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout95
timestamp 1
transform -1 0 7268 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout96
timestamp 1
transform -1 0 12420 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout97
timestamp 1
transform 1 0 6348 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout98
timestamp 1
transform -1 0 11500 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout99
timestamp 1
transform 1 0 11316 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout100
timestamp 1
transform 1 0 11500 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout101
timestamp 1
transform -1 0 14352 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout102
timestamp 1
transform -1 0 15180 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout103
timestamp 1
transform -1 0 14812 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout104
timestamp 1
transform 1 0 15180 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout105
timestamp 1
transform 1 0 12788 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout106
timestamp 1
transform 1 0 18768 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout107
timestamp 1
transform 1 0 16468 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout108
timestamp 1
transform 1 0 21620 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout109
timestamp 1
transform 1 0 16836 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout110
timestamp 1
transform 1 0 16928 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout111
timestamp 1
transform -1 0 22632 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout112
timestamp 1
transform 1 0 11684 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout113
timestamp 1
transform 1 0 19688 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout114
timestamp 1
transform -1 0 25760 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout115
timestamp 1
transform -1 0 15088 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout116
timestamp 1
transform 1 0 13340 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout117
timestamp 1
transform -1 0 4416 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout118
timestamp 1
transform 1 0 16284 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout119
timestamp 1
transform -1 0 23736 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout120
timestamp 1
transform 1 0 16100 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout121
timestamp 1
transform 1 0 7820 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout122
timestamp 1
transform 1 0 19688 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout123
timestamp 1
transform -1 0 12972 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout124
timestamp 1
transform 1 0 20148 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout125
timestamp 1
transform -1 0 18032 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout126
timestamp 1
transform -1 0 18492 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout127
timestamp 1
transform 1 0 17848 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout128
timestamp 1
transform -1 0 17848 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout129
timestamp 1
transform 1 0 17848 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout130
timestamp 1
transform 1 0 7452 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout131
timestamp 1
transform 1 0 20148 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout132
timestamp 1
transform 1 0 20148 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout133
timestamp 1
transform 1 0 20240 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout134
timestamp 1
transform -1 0 13064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout135
timestamp 1
transform 1 0 4324 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout136
timestamp 1
transform 1 0 15272 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout137
timestamp 1
transform -1 0 10580 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout138
timestamp 1
transform 1 0 8372 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout139
timestamp 1
transform 1 0 9752 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout140
timestamp 1
transform 1 0 10488 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout141
timestamp 1
transform -1 0 10304 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout142
timestamp 1
transform -1 0 11500 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout143
timestamp 1
transform 1 0 12328 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout144
timestamp 1
transform 1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout145
timestamp 1
transform -1 0 3956 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout146
timestamp 1
transform 1 0 8096 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout147
timestamp 1
transform -1 0 5612 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout148
timestamp 1
transform 1 0 10396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout149
timestamp 1
transform -1 0 5336 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout150
timestamp 1
transform 1 0 5244 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout151
timestamp 1
transform 1 0 6900 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout152
timestamp 1
transform 1 0 7912 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout153
timestamp 1
transform -1 0 17664 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout154
timestamp 1
transform 1 0 7084 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout155
timestamp 1
transform 1 0 7268 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout156
timestamp 1
transform 1 0 22448 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout157
timestamp 1
transform 1 0 24288 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout158
timestamp 1
transform -1 0 20424 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout159
timestamp 1
transform 1 0 11960 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout160
timestamp 1
transform -1 0 9568 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout161
timestamp 1
transform 1 0 24564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout162
timestamp 1
transform -1 0 12420 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout163
timestamp 1
transform 1 0 17848 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout164
timestamp 1
transform 1 0 11408 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout165
timestamp 1
transform 1 0 17572 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout166
timestamp 1
transform -1 0 7452 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout167
timestamp 1
transform 1 0 17296 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout168
timestamp 1
transform 1 0 25760 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout169
timestamp 1
transform 1 0 22540 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout170
timestamp 1
transform -1 0 19320 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout171
timestamp 1
transform 1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout172
timestamp 1
transform 1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout173
timestamp 1
transform 1 0 8924 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout174
timestamp 1
transform -1 0 15916 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout175
timestamp 1
transform 1 0 19412 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout176
timestamp 1
transform 1 0 11132 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout177
timestamp 1
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout178
timestamp 1
transform 1 0 8648 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout179
timestamp 1
transform -1 0 21712 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout180
timestamp 1
transform 1 0 8924 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout181
timestamp 1
transform -1 0 14904 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout182
timestamp 1
transform 1 0 12788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout183
timestamp 1
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout184
timestamp 1
transform -1 0 14904 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout185
timestamp 1
transform -1 0 8004 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout186
timestamp 1
transform 1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout187
timestamp 1
transform -1 0 16560 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout188
timestamp 1
transform -1 0 13524 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout189
timestamp 1
transform -1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout190
timestamp 1
transform -1 0 12972 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout191
timestamp 1
transform 1 0 12972 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout192
timestamp 1
transform 1 0 12788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout193
timestamp 1
transform -1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout194
timestamp 1
transform 1 0 13064 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout195
timestamp 1
transform -1 0 10120 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout196
timestamp 1
transform -1 0 9752 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout197
timestamp 1
transform -1 0 16928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout198
timestamp 1
transform 1 0 11960 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout199
timestamp 1
transform 1 0 11960 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout200
timestamp 1
transform 1 0 13432 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout201
timestamp 1
transform 1 0 4876 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout202
timestamp 1
transform 1 0 15824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout203
timestamp 1
transform 1 0 12236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout204
timestamp 1
transform 1 0 9476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout205
timestamp 1
transform -1 0 18584 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout206
timestamp 1
transform -1 0 6164 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout207
timestamp 1
transform -1 0 9936 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout208
timestamp 1
transform 1 0 10856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout209
timestamp 1
transform 1 0 16376 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout210
timestamp 1
transform -1 0 10580 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout211
timestamp 1
transform 1 0 13892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout212
timestamp 1
transform 1 0 13524 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout213
timestamp 1
transform 1 0 5152 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout214
timestamp 1
transform -1 0 15456 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout215
timestamp 1
transform -1 0 17204 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout216
timestamp 1
transform -1 0 11960 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout217
timestamp 1
transform 1 0 14720 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout218
timestamp 1
transform 1 0 14536 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout219
timestamp 1
transform -1 0 7820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout220
timestamp 1
transform -1 0 10304 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout221
timestamp 1
transform -1 0 17020 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout222
timestamp 1
transform -1 0 17848 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout223
timestamp 1
transform 1 0 4508 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout224
timestamp 1
transform -1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout225
timestamp 1
transform -1 0 10580 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout226
timestamp 1
transform 1 0 17756 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout227
timestamp 1
transform -1 0 10856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout228
timestamp 1
transform 1 0 13064 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout229
timestamp 1
transform -1 0 10672 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout230
timestamp 1
transform 1 0 22724 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout231
timestamp 1
transform 1 0 18032 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout232
timestamp 1
transform -1 0 14628 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout233
timestamp 1
transform 1 0 22540 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout234
timestamp 1
transform -1 0 19136 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout235
timestamp 1
transform -1 0 16468 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout236
timestamp 1
transform 1 0 19136 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout237
timestamp 1
transform -1 0 14536 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout238
timestamp 1
transform -1 0 22172 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout239
timestamp 1
transform 1 0 12788 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout240
timestamp 1
transform -1 0 24288 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout241
timestamp 1
transform 1 0 11224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout242
timestamp 1
transform 1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout243
timestamp 1
transform 1 0 23184 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout244
timestamp 1
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout245
timestamp 1
transform 1 0 6900 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout246
timestamp 1
transform -1 0 6532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout247
timestamp 1
transform 1 0 17480 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout248
timestamp 1
transform -1 0 28428 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout249
timestamp 1
transform 1 0 17940 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout250
timestamp 1
transform 1 0 7176 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout251
timestamp 1
transform 1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout252
timestamp 1
transform 1 0 7912 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout253
timestamp 1
transform -1 0 19412 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout254
timestamp 1
transform -1 0 21068 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout255
timestamp 1
transform 1 0 19412 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout256
timestamp 1
transform -1 0 6624 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout257
timestamp 1
transform -1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout258
timestamp 1
transform 1 0 14720 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout259
timestamp 1
transform 1 0 25760 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout260
timestamp 1
transform 1 0 11684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout261
timestamp 1
transform -1 0 10120 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout262
timestamp 1
transform -1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout263
timestamp 1
transform 1 0 17112 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout264
timestamp 1
transform -1 0 18492 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout265
timestamp 1
transform -1 0 7268 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout266
timestamp 1
transform -1 0 17756 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout267
timestamp 1
transform 1 0 17940 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout268
timestamp 1
transform 1 0 6164 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout269
timestamp 1
transform 1 0 17756 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout270
timestamp 1
transform 1 0 6900 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout271
timestamp 1
transform 1 0 6900 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout272
timestamp 1
transform -1 0 14720 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout273
timestamp 1
transform -1 0 23828 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout275
timestamp 1
transform 1 0 6900 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout276
timestamp 1
transform 1 0 6624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout277
timestamp 1
transform 1 0 6624 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout278
timestamp 1
transform 1 0 18768 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout279
timestamp 1
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout280
timestamp 1
transform 1 0 6440 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout281
timestamp 1
transform 1 0 27692 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout282
timestamp 1
transform -1 0 13248 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout283
timestamp 1
transform 1 0 7636 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout284
timestamp 1
transform -1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout285
timestamp 1
transform -1 0 14168 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout286
timestamp 1
transform -1 0 27508 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout287
timestamp 1
transform -1 0 8740 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout288
timestamp 1
transform 1 0 28428 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout289
timestamp 1
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout290
timestamp 1
transform 1 0 26956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout291
timestamp 1
transform -1 0 14352 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout292
timestamp 1
transform 1 0 21712 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout293
timestamp 1
transform 1 0 20792 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout294
timestamp 1
transform 1 0 27784 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout295
timestamp 1
transform -1 0 27784 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout296
timestamp 1
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout297
timestamp 1
transform -1 0 12880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout298
timestamp 1
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout299
timestamp 1
transform -1 0 11224 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout300
timestamp 1
transform 1 0 24380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout301
timestamp 1
transform 1 0 14168 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout302
timestamp 1
transform -1 0 18308 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout303
timestamp 1
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout304
timestamp 1
transform -1 0 23184 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout305
timestamp 1
transform -1 0 13248 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout306
timestamp 1
transform -1 0 22264 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout307
timestamp 1
transform -1 0 13524 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout308
timestamp 1
transform -1 0 14352 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout309
timestamp 1
transform 1 0 12328 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout310
timestamp 1
transform 1 0 11960 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout311
timestamp 1
transform 1 0 19228 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout312
timestamp 1
transform 1 0 19872 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout313
timestamp 1
transform -1 0 21528 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout314
timestamp 1
transform 1 0 17296 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout315
timestamp 1
transform 1 0 10212 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout316
timestamp 1
transform 1 0 10764 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout317
timestamp 1
transform -1 0 21252 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout318
timestamp 1
transform -1 0 13248 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout319
timestamp 1
transform -1 0 21344 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout320
timestamp 1
transform -1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout321
timestamp 1
transform 1 0 22264 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout322
timestamp 1
transform 1 0 11040 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout323
timestamp 1
transform -1 0 12696 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout324
timestamp 1
transform 1 0 22816 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout325
timestamp 1
transform -1 0 18032 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout326
timestamp 1
transform 1 0 10304 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout327
timestamp 1
transform 1 0 22816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout328
timestamp 1
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout329
timestamp 1
transform -1 0 23460 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout330
timestamp 1
transform -1 0 23460 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout331
timestamp 1
transform 1 0 10580 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout332
timestamp 1
transform -1 0 11408 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout333
timestamp 1
transform 1 0 22908 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout334
timestamp 1
transform -1 0 15732 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout335
timestamp 1
transform 1 0 17756 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout336
timestamp 1
transform -1 0 13340 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout337
timestamp 1
transform 1 0 5704 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout338
timestamp 1
transform -1 0 6348 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout339
timestamp 1
transform 1 0 10212 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout340
timestamp 1
transform 1 0 11500 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout341
timestamp 1
transform -1 0 10120 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout342
timestamp 1
transform -1 0 10120 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout343
timestamp 1
transform 1 0 5428 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout344
timestamp 1
transform -1 0 4968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout345
timestamp 1
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout346
timestamp 1
transform 1 0 2760 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout347
timestamp 1
transform -1 0 4784 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout348
timestamp 1
transform 1 0 4600 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout349
timestamp 1
transform -1 0 7820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout350
timestamp 1
transform 1 0 11040 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout351
timestamp 1
transform 1 0 8740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout352
timestamp 1
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout353
timestamp 1
transform 1 0 3404 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout354
timestamp 1
transform 1 0 7912 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout355
timestamp 1
transform 1 0 3956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout356
timestamp 1
transform -1 0 8096 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout357
timestamp 1
transform 1 0 10764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout358
timestamp 1
transform 1 0 9844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout359
timestamp 1
transform 1 0 4048 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout360
timestamp 1
transform 1 0 4048 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout361
timestamp 1
transform 1 0 4692 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout362
timestamp 1
transform 1 0 8004 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout363
timestamp 1
transform 1 0 6992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout364
timestamp 1
transform 1 0 7268 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout365
timestamp 1
transform -1 0 5244 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout366
timestamp 1
transform 1 0 4600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout367
timestamp 1
transform 1 0 8280 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout368
timestamp 1
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout369
timestamp 1
transform 1 0 8280 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout370
timestamp 1
transform 1 0 7636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout371
timestamp 1
transform 1 0 7544 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout372
timestamp 1
transform 1 0 4692 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout373
timestamp 1
transform 1 0 4784 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout374
timestamp 1
transform 1 0 5152 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout375
timestamp 1
transform -1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout376
timestamp 1
transform -1 0 6256 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout377
timestamp 1
transform -1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout378
timestamp 1
transform 1 0 3036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout379
timestamp 1
transform -1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout380
timestamp 1
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout381
timestamp 1
transform -1 0 5704 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout382
timestamp 1
transform 1 0 5428 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout383
timestamp 1
transform -1 0 4416 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout384
timestamp 1
transform -1 0 4784 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout385
timestamp 1
transform 1 0 6992 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout386
timestamp 1
transform -1 0 5704 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout387
timestamp 1
transform 1 0 5704 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout388
timestamp 1
transform -1 0 4876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout389
timestamp 1
transform -1 0 4508 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout390
timestamp 1
transform 1 0 7268 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout391
timestamp 1
transform -1 0 7820 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout392
timestamp 1
transform -1 0 5428 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout393
timestamp 1
transform 1 0 5152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout394
timestamp 1
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout395
timestamp 1
transform 1 0 5980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout396
timestamp 1
transform -1 0 3680 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout397
timestamp 1
transform -1 0 3864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout398
timestamp 1
transform -1 0 2668 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout399
timestamp 1
transform -1 0 5336 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout400
timestamp 1
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout401
timestamp 1
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout402
timestamp 1
transform 1 0 4416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout403
timestamp 1
transform 1 0 5244 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout404
timestamp 1
transform -1 0 3588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout405
timestamp 1
transform -1 0 3312 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout406
timestamp 1
transform 1 0 3312 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout407
timestamp 1
transform -1 0 5888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout408
timestamp 1
transform -1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout409
timestamp 1
transform -1 0 4140 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout410
timestamp 1
transform 1 0 7176 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout411
timestamp 1
transform -1 0 6992 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout412
timestamp 1
transform -1 0 8740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout413
timestamp 1
transform -1 0 6256 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout414
timestamp 1
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout415
timestamp 1
transform -1 0 11316 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout416
timestamp 1
transform 1 0 9660 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout417
timestamp 1
transform -1 0 8280 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout418
timestamp 1
transform 1 0 6348 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout419
timestamp 1
transform -1 0 6716 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout420
timestamp 1
transform 1 0 6992 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout421
timestamp 1
transform -1 0 9844 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout422
timestamp 1
transform -1 0 12788 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout423
timestamp 1
transform -1 0 9660 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout424
timestamp 1
transform -1 0 10212 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout425
timestamp 1
transform 1 0 7268 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout426
timestamp 1
transform 1 0 6256 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout427
timestamp 1
transform 1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout428
timestamp 1
transform -1 0 6256 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout429
timestamp 1
transform 1 0 10856 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout430
timestamp 1
transform -1 0 6900 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout431
timestamp 1
transform -1 0 7268 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout432
timestamp 1
transform -1 0 8096 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout433
timestamp 1
transform -1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout434
timestamp 1
transform 1 0 9200 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout435
timestamp 1
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout436
timestamp 1
transform 1 0 10580 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout437
timestamp 1
transform 1 0 6900 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout438
timestamp 1
transform -1 0 7544 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout439
timestamp 1
transform -1 0 7820 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout440
timestamp 1
transform 1 0 4692 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout441
timestamp 1
transform -1 0 5336 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout442
timestamp 1
transform -1 0 10396 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout443
timestamp 1
transform 1 0 9752 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout444
timestamp 1
transform -1 0 8556 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout445
timestamp 1
transform -1 0 10764 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout446
timestamp 1
transform -1 0 9936 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout447
timestamp 1
transform -1 0 10580 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout448
timestamp 1
transform 1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout449
timestamp 1
transform 1 0 5336 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout450
timestamp 1
transform -1 0 8740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout451
timestamp 1
transform -1 0 9568 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout452
timestamp 1
transform 1 0 10120 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout453
timestamp 1
transform -1 0 10488 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout454
timestamp 1
transform -1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout455
timestamp 1
transform 1 0 10028 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout456
timestamp 1
transform -1 0 2484 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout457
timestamp 1
transform -1 0 4600 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout458
timestamp 1
transform 1 0 3496 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout459
timestamp 1
transform -1 0 3496 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout460
timestamp 1
transform 1 0 9200 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout461
timestamp 1
transform -1 0 8832 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout462
timestamp 1
transform 1 0 9200 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout463
timestamp 1
transform -1 0 9752 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout464
timestamp 1
transform 1 0 8924 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout466
timestamp 1
transform -1 0 3680 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout467
timestamp 1
transform -1 0 4692 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout468
timestamp 1
transform 1 0 3772 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout469
timestamp 1
transform -1 0 3220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout470
timestamp 1
transform 1 0 8924 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout471
timestamp 1
transform -1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout472
timestamp 1
transform -1 0 8280 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout473
timestamp 1
transform -1 0 8924 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout474
timestamp 1
transform -1 0 9384 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout475
timestamp 1
transform -1 0 2944 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout476
timestamp 1
transform -1 0 5428 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout477
timestamp 1
transform -1 0 3404 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout478
timestamp 1
transform 1 0 4508 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout479
timestamp 1
transform -1 0 5244 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout480
timestamp 1
transform 1 0 5796 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout481
timestamp 1
transform -1 0 6348 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout482
timestamp 1
transform -1 0 6624 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout483
timestamp 1
transform -1 0 5152 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout484
timestamp 1
transform -1 0 3864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout485
timestamp 1
transform -1 0 4692 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout486
timestamp 1
transform -1 0 5796 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout487
timestamp 1
transform 1 0 6624 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout488
timestamp 1
transform -1 0 5520 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout489
timestamp 1
transform -1 0 6072 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout490
timestamp 1
transform 1 0 5244 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout491
timestamp 1
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout492
timestamp 1
transform 1 0 6624 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout493
timestamp 1
transform -1 0 5244 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout494
timestamp 1
transform -1 0 5888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout495
timestamp 1
transform 1 0 7912 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout496
timestamp 1
transform -1 0 7084 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout497
timestamp 1
transform 1 0 8188 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout498
timestamp 1
transform 1 0 7728 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout499
timestamp 1
transform 1 0 7636 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout500
timestamp 1
transform -1 0 6348 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout501
timestamp 1
transform -1 0 5980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout502
timestamp 1
transform -1 0 5612 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout503
timestamp 1
transform 1 0 7636 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout504
timestamp 1
transform -1 0 7360 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout505
timestamp 1
transform 1 0 7360 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout506
timestamp 1
transform -1 0 7912 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout507
timestamp 1
transform -1 0 8188 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout508
timestamp 1
transform 1 0 4784 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout509
timestamp 1
transform 1 0 6348 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout510
timestamp 1
transform -1 0 13340 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout511
timestamp 1
transform -1 0 10856 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout512
timestamp 1
transform -1 0 11040 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout513
timestamp 1
transform 1 0 11224 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout514
timestamp 1
transform 1 0 5520 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout515
timestamp 1
transform 1 0 8188 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout516
timestamp 1
transform -1 0 4140 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout517
timestamp 1
transform 1 0 4048 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout518
timestamp 1
transform -1 0 5152 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout519
timestamp 1
transform -1 0 5428 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout520
timestamp 1
transform -1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout521
timestamp 1
transform 1 0 5428 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout522
timestamp 1
transform -1 0 12512 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout523
timestamp 1
transform 1 0 12788 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout524
timestamp 1
transform 1 0 5704 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout525
timestamp 1
transform 1 0 5796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout526
timestamp 1
transform -1 0 5152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout527
timestamp 1
transform -1 0 5244 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout528
timestamp 1
transform 1 0 4324 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout529
timestamp 1
transform 1 0 11500 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout530
timestamp 1
transform -1 0 11408 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout531
timestamp 1
transform 1 0 5980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout532
timestamp 1
transform -1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout533
timestamp 1
transform -1 0 5520 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout534
timestamp 1
transform 1 0 3864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout535
timestamp 1
transform -1 0 12236 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout536
timestamp 1
transform -1 0 12512 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout537
timestamp 1
transform 1 0 12788 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout538
timestamp 1
transform 1 0 2944 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout539
timestamp 1
transform -1 0 6624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout540
timestamp 1
transform -1 0 9292 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout541
timestamp 1
transform 1 0 10856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout542
timestamp 1
transform 1 0 12144 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout543
timestamp 1
transform 1 0 9568 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout544
timestamp 1
transform -1 0 6256 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout545
timestamp 1
transform -1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout546
timestamp 1
transform -1 0 4232 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout547
timestamp 1
transform -1 0 4508 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout548
timestamp 1
transform -1 0 13524 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout549
timestamp 1
transform 1 0 12512 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout550
timestamp 1
transform 1 0 13524 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout551
timestamp 1
transform -1 0 5152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout552
timestamp 1
transform -1 0 5704 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout553
timestamp 1
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout554
timestamp 1
transform 1 0 11132 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout555
timestamp 1
transform 1 0 11040 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout556
timestamp 1
transform 1 0 9292 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout557
timestamp 1
transform -1 0 6624 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout558
timestamp 1
transform -1 0 24288 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout559
timestamp 1
transform 1 0 24196 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout560
timestamp 1
transform -1 0 32016 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout561
timestamp 1
transform -1 0 31832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout562
timestamp 1
transform 1 0 31004 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout563
timestamp 1
transform 1 0 30084 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout564
timestamp 1
transform 1 0 30636 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout565
timestamp 1
transform -1 0 31188 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout566
timestamp 1
transform -1 0 30636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout567
timestamp 1
transform 1 0 30636 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout568
timestamp 1
transform -1 0 30912 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout569
timestamp 1
transform -1 0 30360 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout570
timestamp 1
transform -1 0 30084 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout571
timestamp 1
transform -1 0 30636 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout572
timestamp 1
transform -1 0 22816 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout573
timestamp 1
transform 1 0 31648 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout574
timestamp 1
transform 1 0 1472 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout575
timestamp 1
transform 1 0 4508 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout576
timestamp 1
transform -1 0 2944 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout577
timestamp 1
transform 1 0 1840 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout578
timestamp 1
transform -1 0 4048 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout579
timestamp 1
transform 1 0 2392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout580
timestamp 1
transform -1 0 2392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout581
timestamp 1
transform -1 0 3956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout582
timestamp 1
transform -1 0 2852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout583
timestamp 1
transform 1 0 4232 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout584
timestamp 1
transform -1 0 2576 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout585
timestamp 1
transform -1 0 2116 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout586
timestamp 1
transform -1 0 4416 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout587
timestamp 1
transform -1 0 2668 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout588
timestamp 1
transform 1 0 2760 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout589
timestamp 1
transform -1 0 2300 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout590
timestamp 1
transform -1 0 2024 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout591
timestamp 1
transform 1 0 1748 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout592
timestamp 1
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout593
timestamp 1
transform 1 0 4968 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout594
timestamp 1
transform -1 0 3128 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout595
timestamp 1
transform -1 0 3312 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout596
timestamp 1
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout597
timestamp 1
transform -1 0 2576 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout598
timestamp 1
transform -1 0 3128 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout599
timestamp 1
transform 1 0 3220 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout600
timestamp 1
transform 1 0 4416 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout601
timestamp 1
transform -1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout602
timestamp 1
transform 1 0 2116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout603
timestamp 1
transform -1 0 2760 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout604
timestamp 1
transform -1 0 2300 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout605
timestamp 1
transform 1 0 2024 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout606
timestamp 1
transform -1 0 3036 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout607
timestamp 1
transform 1 0 5704 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout608
timestamp 1
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout609
timestamp 1
transform -1 0 4968 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout610
timestamp 1
transform 1 0 4048 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout611
timestamp 1
transform -1 0 3772 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout612
timestamp 1
transform -1 0 4048 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout613
timestamp 1
transform 1 0 2944 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout614
timestamp 1
transform 1 0 4048 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout615
timestamp 1
transform 1 0 5244 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout616
timestamp 1
transform 1 0 3220 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout617
timestamp 1
transform 1 0 2300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout618
timestamp 1
transform -1 0 3404 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout619
timestamp 1
transform 1 0 4968 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout620
timestamp 1
transform -1 0 4692 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout621
timestamp 1
transform -1 0 4048 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout622
timestamp 1
transform -1 0 4324 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout623
timestamp 1
transform -1 0 3496 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout624
timestamp 1
transform 1 0 3496 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout625
timestamp 1
transform -1 0 2760 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout626
timestamp 1
transform -1 0 4600 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout627
timestamp 1
transform -1 0 4968 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout628
timestamp 1
transform -1 0 4692 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout629
timestamp 1
transform 1 0 3772 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1636968456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1636968456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_169
timestamp 1
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_177
timestamp 1
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_182
timestamp 1636968456
transform 1 0 17848 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_194
timestamp 1
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_197
timestamp 1
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_203
timestamp 1636968456
transform 1 0 19780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_215
timestamp 1
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_219
timestamp 1
transform 1 0 21252 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_225
timestamp 1
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_233
timestamp 1
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_238
timestamp 1636968456
transform 1 0 23000 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_250
timestamp 1
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_253
timestamp 1
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_259
timestamp 1
transform 1 0 24932 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_267
timestamp 1
transform 1 0 25668 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_273
timestamp 1
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 1
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1636968456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1636968456
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_309
timestamp 1
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_314
timestamp 1636968456
transform 1 0 29992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_326
timestamp 1
transform 1 0 31096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_334
timestamp 1
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_337
timestamp 1
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_341
timestamp 1
transform 1 0 32476 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1636968456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1636968456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1636968456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1636968456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1636968456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1636968456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1636968456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1636968456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1636968456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1636968456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1636968456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1636968456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1636968456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1636968456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1636968456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1636968456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_337
timestamp 1
transform 1 0 32108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_341
timestamp 1
transform 1 0 32476 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1636968456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1636968456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1636968456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1636968456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1636968456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_153
timestamp 1
transform 1 0 15180 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_161
timestamp 1
transform 1 0 15916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_179
timestamp 1
transform 1 0 17572 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_185
timestamp 1
transform 1 0 18124 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_193
timestamp 1
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1636968456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_209
timestamp 1
transform 1 0 20332 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_227
timestamp 1636968456
transform 1 0 21988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_239
timestamp 1636968456
transform 1 0 23092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1636968456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1636968456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1636968456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1636968456
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1636968456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1636968456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_333
timestamp 1
transform 1 0 31740 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_341
timestamp 1
transform 1 0 32476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1636968456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1636968456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1636968456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1636968456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1636968456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_187
timestamp 1
transform 1 0 18308 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_209
timestamp 1
transform 1 0 20332 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_225
timestamp 1
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_245
timestamp 1
transform 1 0 23644 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_271
timestamp 1
transform 1 0 26036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1636968456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1636968456
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1636968456
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1636968456
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_337
timestamp 1
transform 1 0 32108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_341
timestamp 1
transform 1 0 32476 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1636968456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1636968456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_85
timestamp 1
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_93
timestamp 1
transform 1 0 9660 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_101
timestamp 1636968456
transform 1 0 10396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_113
timestamp 1
transform 1 0 11500 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_119
timestamp 1
transform 1 0 12052 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_130
timestamp 1
transform 1 0 13064 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp 1
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_141
timestamp 1
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_150
timestamp 1
transform 1 0 14904 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_158
timestamp 1
transform 1 0 15640 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_166
timestamp 1636968456
transform 1 0 16376 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_178
timestamp 1636968456
transform 1 0 17480 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_190
timestamp 1
transform 1 0 18584 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_205
timestamp 1
transform 1 0 19964 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_213
timestamp 1
transform 1 0 20700 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_221
timestamp 1
transform 1 0 21436 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_229
timestamp 1
transform 1 0 22172 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_237
timestamp 1
transform 1 0 22908 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_256
timestamp 1
transform 1 0 24656 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_274
timestamp 1636968456
transform 1 0 26312 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_286
timestamp 1636968456
transform 1 0 27416 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_298
timestamp 1
transform 1 0 28520 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_306
timestamp 1
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1636968456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1636968456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_333
timestamp 1
transform 1 0 31740 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_341
timestamp 1
transform 1 0 32476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636968456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1636968456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1636968456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1636968456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636968456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_69
timestamp 1
transform 1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_83
timestamp 1636968456
transform 1 0 8740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_95
timestamp 1636968456
transform 1 0 9844 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_107
timestamp 1
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_113
timestamp 1
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_120
timestamp 1636968456
transform 1 0 12144 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_132
timestamp 1
transform 1 0 13248 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_140
timestamp 1
transform 1 0 13984 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_150
timestamp 1636968456
transform 1 0 14904 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_162
timestamp 1
transform 1 0 16008 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1636968456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_181
timestamp 1
transform 1 0 17756 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_191
timestamp 1636968456
transform 1 0 18676 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_203
timestamp 1636968456
transform 1 0 19780 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_215
timestamp 1
transform 1 0 20884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1636968456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_237
timestamp 1
transform 1 0 22908 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_240
timestamp 1
transform 1 0 23184 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_269
timestamp 1
transform 1 0 25852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_277
timestamp 1
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1636968456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1636968456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1636968456
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1636968456
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_337
timestamp 1
transform 1 0 32108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_341
timestamp 1
transform 1 0 32476 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1636968456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1636968456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1636968456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_53
timestamp 1
transform 1 0 5980 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_69
timestamp 1
transform 1 0 7452 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_75
timestamp 1
transform 1 0 8004 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_89
timestamp 1636968456
transform 1 0 9292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_101
timestamp 1636968456
transform 1 0 10396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_113
timestamp 1636968456
transform 1 0 11500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_125
timestamp 1
transform 1 0 12604 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_136
timestamp 1
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1636968456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1636968456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_165
timestamp 1
transform 1 0 16284 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_171
timestamp 1
transform 1 0 16836 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_177
timestamp 1
transform 1 0 17388 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_185
timestamp 1
transform 1 0 18124 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_192
timestamp 1
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1636968456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1636968456
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1636968456
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_233
timestamp 1
transform 1 0 22540 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_237
timestamp 1
transform 1 0 22908 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_249
timestamp 1
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1636968456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1636968456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1636968456
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1636968456
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1636968456
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1636968456
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_333
timestamp 1
transform 1 0 31740 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_341
timestamp 1
transform 1 0 32476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1636968456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1636968456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1636968456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1636968456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1636968456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1636968456
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1636968456
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_93
timestamp 1
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_101
timestamp 1
transform 1 0 10396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_108
timestamp 1
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_119
timestamp 1636968456
transform 1 0 12052 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_131
timestamp 1
transform 1 0 13156 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_139
timestamp 1
transform 1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_147
timestamp 1
transform 1 0 14628 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_160
timestamp 1
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_169
timestamp 1
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_185
timestamp 1
transform 1 0 18124 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_189
timestamp 1
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_198
timestamp 1
transform 1 0 19320 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_210
timestamp 1
transform 1 0 20424 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_214
timestamp 1
transform 1 0 20792 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_220
timestamp 1
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_236
timestamp 1
transform 1 0 22816 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_246
timestamp 1636968456
transform 1 0 23736 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_269
timestamp 1
transform 1 0 25852 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_278
timestamp 1
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1636968456
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1636968456
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1636968456
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1636968456
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_337
timestamp 1
transform 1 0 32108 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_29
timestamp 1
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_37
timestamp 1
transform 1 0 4508 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_42
timestamp 1636968456
transform 1 0 4968 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_54
timestamp 1636968456
transform 1 0 6072 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_66
timestamp 1
transform 1 0 7176 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_70
timestamp 1
transform 1 0 7544 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_74
timestamp 1
transform 1 0 7912 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 1
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_93
timestamp 1
transform 1 0 9660 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_122
timestamp 1
transform 1 0 12328 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_126
timestamp 1
transform 1 0 12696 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_130
timestamp 1
transform 1 0 13064 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1636968456
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_161
timestamp 1
transform 1 0 15916 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_167
timestamp 1636968456
transform 1 0 16468 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_197
timestamp 1
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_205
timestamp 1
transform 1 0 19964 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_212
timestamp 1636968456
transform 1 0 20608 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_224
timestamp 1
transform 1 0 21712 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_236
timestamp 1636968456
transform 1 0 22816 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_248
timestamp 1
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_258
timestamp 1636968456
transform 1 0 24840 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_270
timestamp 1
transform 1 0 25944 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_274
timestamp 1
transform 1 0 26312 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_280
timestamp 1636968456
transform 1 0 26864 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_292
timestamp 1636968456
transform 1 0 27968 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_304
timestamp 1
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_309
timestamp 1
transform 1 0 29532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_317
timestamp 1
transform 1 0 30268 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1636968456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1636968456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_27
timestamp 1
transform 1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_47
timestamp 1
transform 1 0 5428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_98
timestamp 1
transform 1 0 10120 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_104
timestamp 1
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_113
timestamp 1
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_121
timestamp 1
transform 1 0 12236 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1636968456
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1636968456
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_161
timestamp 1
transform 1 0 15916 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1636968456
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1636968456
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_193
timestamp 1
transform 1 0 18860 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_199
timestamp 1636968456
transform 1 0 19412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_211
timestamp 1636968456
transform 1 0 20516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_225
timestamp 1
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_234
timestamp 1636968456
transform 1 0 22632 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_246
timestamp 1
transform 1 0 23736 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_253
timestamp 1636968456
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_265
timestamp 1
transform 1 0 25484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_274
timestamp 1
transform 1 0 26312 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_281
timestamp 1
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_287
timestamp 1
transform 1 0 27508 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_294
timestamp 1636968456
transform 1 0 28152 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_306
timestamp 1
transform 1 0 29256 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_314
timestamp 1
transform 1 0 29992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_323
timestamp 1
transform 1 0 30820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_327
timestamp 1
transform 1 0 31188 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_341
timestamp 1
transform 1 0 32476 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1636968456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1636968456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1636968456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1636968456
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_53
timestamp 1
transform 1 0 5980 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_62
timestamp 1636968456
transform 1 0 6808 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_74
timestamp 1
transform 1 0 7912 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_78
timestamp 1
transform 1 0 8280 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_92
timestamp 1636968456
transform 1 0 9568 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_104
timestamp 1
transform 1 0 10672 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_116
timestamp 1
transform 1 0 11776 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_124
timestamp 1
transform 1 0 12512 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_132
timestamp 1
transform 1 0 13248 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_141
timestamp 1
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_150
timestamp 1636968456
transform 1 0 14904 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_167
timestamp 1
transform 1 0 16468 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_180
timestamp 1636968456
transform 1 0 17664 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_192
timestamp 1
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1636968456
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_221
timestamp 1
transform 1 0 21436 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_239
timestamp 1636968456
transform 1 0 23092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1636968456
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_265
timestamp 1
transform 1 0 25484 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_274
timestamp 1636968456
transform 1 0 26312 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_286
timestamp 1636968456
transform 1 0 27416 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_298
timestamp 1
transform 1 0 28520 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_325
timestamp 1
transform 1 0 31004 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1636968456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1636968456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_27
timestamp 1
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_31
timestamp 1
transform 1 0 3956 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_35
timestamp 1
transform 1 0 4324 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_39
timestamp 1
transform 1 0 4692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_57
timestamp 1
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_65
timestamp 1
transform 1 0 7084 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_73
timestamp 1
transform 1 0 7820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_130
timestamp 1
transform 1 0 13064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_134
timestamp 1
transform 1 0 13432 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_141
timestamp 1
transform 1 0 14076 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_149
timestamp 1
transform 1 0 14812 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_162
timestamp 1
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_177
timestamp 1
transform 1 0 17388 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_183
timestamp 1636968456
transform 1 0 17940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_195
timestamp 1
transform 1 0 19044 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_203
timestamp 1
transform 1 0 19780 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_214
timestamp 1
transform 1 0 20792 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_222
timestamp 1
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1636968456
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_237
timestamp 1
transform 1 0 22908 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_257
timestamp 1636968456
transform 1 0 24748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_269
timestamp 1
transform 1 0 25852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_277
timestamp 1
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1636968456
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1636968456
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_305
timestamp 1
transform 1 0 29164 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_316
timestamp 1
transform 1 0 30176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_320
timestamp 1
transform 1 0 30544 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_337
timestamp 1
transform 1 0 32108 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1636968456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_15
timestamp 1
transform 1 0 2484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_23
timestamp 1
transform 1 0 3220 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_63
timestamp 1
transform 1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_76
timestamp 1
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_91
timestamp 1636968456
transform 1 0 9476 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_103
timestamp 1
transform 1 0 10580 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_128
timestamp 1636968456
transform 1 0 12880 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_149
timestamp 1636968456
transform 1 0 14812 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_161
timestamp 1
transform 1 0 15916 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_169
timestamp 1
transform 1 0 16652 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_182
timestamp 1
transform 1 0 17848 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_194
timestamp 1
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1636968456
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1636968456
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_221
timestamp 1
transform 1 0 21436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_225
timestamp 1
transform 1 0 21804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_232
timestamp 1636968456
transform 1 0 22448 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_244
timestamp 1
transform 1 0 23552 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_253
timestamp 1
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_261
timestamp 1
transform 1 0 25116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_271
timestamp 1
transform 1 0 26036 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_284
timestamp 1
transform 1 0 27232 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_297
timestamp 1
transform 1 0 28428 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_301
timestamp 1
transform 1 0 28796 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1636968456
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_321
timestamp 1
transform 1 0 30636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_325
timestamp 1
transform 1 0 31004 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_15
timestamp 1
transform 1 0 2484 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_38
timestamp 1
transform 1 0 4600 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_42
timestamp 1
transform 1 0 4968 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_84
timestamp 1
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_113
timestamp 1
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_117
timestamp 1
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_124
timestamp 1
transform 1 0 12512 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_136
timestamp 1
transform 1 0 13616 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_143
timestamp 1636968456
transform 1 0 14260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_155
timestamp 1
transform 1 0 15364 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_161
timestamp 1
transform 1 0 15916 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1636968456
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_191
timestamp 1
transform 1 0 18676 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_207
timestamp 1
transform 1 0 20148 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_220
timestamp 1
transform 1 0 21344 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_225
timestamp 1
transform 1 0 21804 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_239
timestamp 1636968456
transform 1 0 23092 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_251
timestamp 1
transform 1 0 24196 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_263
timestamp 1
transform 1 0 25300 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_271
timestamp 1
transform 1 0 26036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_277
timestamp 1
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1636968456
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1636968456
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_305
timestamp 1
transform 1 0 29164 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_332
timestamp 1
transform 1 0 31648 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_337
timestamp 1
transform 1 0 32108 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1636968456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_15
timestamp 1
transform 1 0 2484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_23
timestamp 1
transform 1 0 3220 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_36
timestamp 1
transform 1 0 4416 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_44
timestamp 1
transform 1 0 5152 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_49
timestamp 1
transform 1 0 5612 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_59
timestamp 1
transform 1 0 6532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_66
timestamp 1
transform 1 0 7176 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_73
timestamp 1
transform 1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_85
timestamp 1
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_96
timestamp 1
transform 1 0 9936 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_104
timestamp 1
transform 1 0 10672 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_111
timestamp 1636968456
transform 1 0 11316 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_123
timestamp 1636968456
transform 1 0 12420 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_135
timestamp 1
transform 1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1636968456
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_153
timestamp 1
transform 1 0 15180 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_163
timestamp 1
transform 1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_179
timestamp 1
transform 1 0 17572 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_190
timestamp 1
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_202
timestamp 1
transform 1 0 19688 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_208
timestamp 1636968456
transform 1 0 20240 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_220
timestamp 1
transform 1 0 21344 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_234
timestamp 1636968456
transform 1 0 22632 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_246
timestamp 1
transform 1 0 23736 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_259
timestamp 1636968456
transform 1 0 24932 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_271
timestamp 1636968456
transform 1 0 26036 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_291
timestamp 1636968456
transform 1 0 27876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_303
timestamp 1
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_315
timestamp 1
transform 1 0 30084 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1636968456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1636968456
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_27
timestamp 1
transform 1 0 3588 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_31
timestamp 1
transform 1 0 3956 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_48
timestamp 1
transform 1 0 5520 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_75
timestamp 1
transform 1 0 8004 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_83
timestamp 1
transform 1 0 8740 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_94
timestamp 1636968456
transform 1 0 9752 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_106
timestamp 1
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_121
timestamp 1
transform 1 0 12236 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_131
timestamp 1636968456
transform 1 0 13156 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_150
timestamp 1
transform 1 0 14904 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_158
timestamp 1
transform 1 0 15640 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_166
timestamp 1
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_169
timestamp 1
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_185
timestamp 1
transform 1 0 18124 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_193
timestamp 1
transform 1 0 18860 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_218
timestamp 1
transform 1 0 21160 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_230
timestamp 1
transform 1 0 22264 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_242
timestamp 1
transform 1 0 23368 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_254
timestamp 1
transform 1 0 24472 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_262
timestamp 1
transform 1 0 25208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_276
timestamp 1
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_281
timestamp 1
transform 1 0 26956 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_298
timestamp 1636968456
transform 1 0 28520 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_310
timestamp 1
transform 1 0 29624 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_337
timestamp 1
transform 1 0 32108 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_6
timestamp 1
transform 1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_23
timestamp 1
transform 1 0 3220 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_29
timestamp 1
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_50
timestamp 1
transform 1 0 5704 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1636968456
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_109
timestamp 1
transform 1 0 11132 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_119
timestamp 1636968456
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_131
timestamp 1
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_141
timestamp 1
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_151
timestamp 1
transform 1 0 14996 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_159
timestamp 1
transform 1 0 15732 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_168
timestamp 1
transform 1 0 16560 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_174
timestamp 1
transform 1 0 17112 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_180
timestamp 1636968456
transform 1 0 17664 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_192
timestamp 1
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1636968456
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_209
timestamp 1
transform 1 0 20332 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_221
timestamp 1
transform 1 0 21436 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_235
timestamp 1
transform 1 0 22724 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_243
timestamp 1
transform 1 0 23460 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 1
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1636968456
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_265
timestamp 1
transform 1 0 25484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_272
timestamp 1
transform 1 0 26128 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_284
timestamp 1
transform 1 0 27232 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_288
timestamp 1
transform 1 0 27600 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_294
timestamp 1636968456
transform 1 0 28152 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_306
timestamp 1
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_309
timestamp 1
transform 1 0 29532 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_315
timestamp 1
transform 1 0 30084 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_339
timestamp 1
transform 1 0 32292 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1636968456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_15
timestamp 1
transform 1 0 2484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_30
timestamp 1
transform 1 0 3864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_37
timestamp 1
transform 1 0 4508 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_41
timestamp 1
transform 1 0 4876 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_48
timestamp 1
transform 1 0 5520 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_52
timestamp 1
transform 1 0 5888 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_57
timestamp 1
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_66
timestamp 1
transform 1 0 7176 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_70
timestamp 1
transform 1 0 7544 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_76
timestamp 1
transform 1 0 8096 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_89
timestamp 1636968456
transform 1 0 9292 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_110
timestamp 1
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_119
timestamp 1
transform 1 0 12052 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_125
timestamp 1
transform 1 0 12604 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_134
timestamp 1
transform 1 0 13432 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_142
timestamp 1
transform 1 0 14168 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_154
timestamp 1636968456
transform 1 0 15272 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_175
timestamp 1
transform 1 0 17204 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_181
timestamp 1
transform 1 0 17756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_196
timestamp 1
transform 1 0 19136 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_207
timestamp 1
transform 1 0 20148 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1636968456
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_237
timestamp 1
transform 1 0 22908 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_245
timestamp 1
transform 1 0 23644 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_251
timestamp 1636968456
transform 1 0 24196 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_263
timestamp 1636968456
transform 1 0 25300 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_275
timestamp 1
transform 1 0 26404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1636968456
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_293
timestamp 1
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_303
timestamp 1
transform 1 0 28980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_315
timestamp 1
transform 1 0 30084 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_319
timestamp 1
transform 1 0 30452 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_337
timestamp 1
transform 1 0 32108 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_3
timestamp 1
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_11
timestamp 1
transform 1 0 2116 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_29
timestamp 1
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_37
timestamp 1
transform 1 0 4508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_57
timestamp 1
transform 1 0 6348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_62
timestamp 1
transform 1 0 6808 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_78
timestamp 1
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_85
timestamp 1
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_93
timestamp 1636968456
transform 1 0 9660 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_105
timestamp 1
transform 1 0 10764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_112
timestamp 1
transform 1 0 11408 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_120
timestamp 1636968456
transform 1 0 12144 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_132
timestamp 1
transform 1 0 13248 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1636968456
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_153
timestamp 1
transform 1 0 15180 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_161
timestamp 1
transform 1 0 15916 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_167
timestamp 1
transform 1 0 16468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_176
timestamp 1
transform 1 0 17296 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_182
timestamp 1
transform 1 0 17848 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_193
timestamp 1
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_202
timestamp 1636968456
transform 1 0 19688 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_214
timestamp 1
transform 1 0 20792 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_222
timestamp 1
transform 1 0 21528 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_237
timestamp 1
transform 1 0 22908 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_271
timestamp 1
transform 1 0 26036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_277
timestamp 1
transform 1 0 26588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_283
timestamp 1
transform 1 0 27140 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_295
timestamp 1636968456
transform 1 0 28244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_309
timestamp 1
transform 1 0 29532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_320
timestamp 1
transform 1 0 30544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_331
timestamp 1
transform 1 0 31556 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_340
timestamp 1
transform 1 0 32384 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1636968456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_15
timestamp 1
transform 1 0 2484 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_32
timestamp 1
transform 1 0 4048 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_49
timestamp 1
transform 1 0 5612 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_63
timestamp 1
transform 1 0 6900 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_75
timestamp 1
transform 1 0 8004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_88
timestamp 1
transform 1 0 9200 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_95
timestamp 1
transform 1 0 9844 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_103
timestamp 1
transform 1 0 10580 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_123
timestamp 1636968456
transform 1 0 12420 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_135
timestamp 1636968456
transform 1 0 13524 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_147
timestamp 1
transform 1 0 14628 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_169
timestamp 1
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_179
timestamp 1
transform 1 0 17572 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_187
timestamp 1
transform 1 0 18308 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_195
timestamp 1
transform 1 0 19044 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_203
timestamp 1
transform 1 0 19780 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_209
timestamp 1636968456
transform 1 0 20332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_221
timestamp 1
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_225
timestamp 1
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_232
timestamp 1
transform 1 0 22448 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_240
timestamp 1
transform 1 0 23184 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_261
timestamp 1
transform 1 0 25116 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_267
timestamp 1
transform 1 0 25668 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_274
timestamp 1
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_281
timestamp 1
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_289
timestamp 1
transform 1 0 27692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_293
timestamp 1
transform 1 0 28060 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_300
timestamp 1636968456
transform 1 0 28704 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_312
timestamp 1
transform 1 0 29808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_316
timestamp 1
transform 1 0 30176 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_337
timestamp 1
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_3
timestamp 1
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_11
timestamp 1
transform 1 0 2116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_18
timestamp 1
transform 1 0 2760 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_24
timestamp 1
transform 1 0 3312 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_39
timestamp 1
transform 1 0 4692 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_78
timestamp 1
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_85
timestamp 1
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_93
timestamp 1636968456
transform 1 0 9660 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_105
timestamp 1
transform 1 0 10764 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_109
timestamp 1
transform 1 0 11132 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_113
timestamp 1636968456
transform 1 0 11500 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_125
timestamp 1
transform 1 0 12604 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_135
timestamp 1
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_146
timestamp 1
transform 1 0 14536 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_157
timestamp 1636968456
transform 1 0 15548 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_169
timestamp 1636968456
transform 1 0 16652 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_181
timestamp 1
transform 1 0 17756 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_188
timestamp 1
transform 1 0 18400 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_197
timestamp 1
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_205
timestamp 1
transform 1 0 19964 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1636968456
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 1636968456
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 1
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_276
timestamp 1
transform 1 0 26496 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_284
timestamp 1
transform 1 0 27232 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1636968456
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_321
timestamp 1
transform 1 0 30636 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_331
timestamp 1
transform 1 0 31556 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_340
timestamp 1
transform 1 0 32384 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1636968456
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_18
timestamp 1
transform 1 0 2760 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_38
timestamp 1
transform 1 0 4600 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_46
timestamp 1
transform 1 0 5336 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 1
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_73
timestamp 1
transform 1 0 7820 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_79
timestamp 1
transform 1 0 8372 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_101
timestamp 1
transform 1 0 10396 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_113
timestamp 1
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_124
timestamp 1
transform 1 0 12512 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_138
timestamp 1
transform 1 0 13800 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_146
timestamp 1
transform 1 0 14536 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_156
timestamp 1636968456
transform 1 0 15456 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1636968456
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_181
timestamp 1
transform 1 0 17756 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_196
timestamp 1636968456
transform 1 0 19136 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_208
timestamp 1
transform 1 0 20240 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_238
timestamp 1
transform 1 0 23000 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_246
timestamp 1
transform 1 0 23736 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_253
timestamp 1636968456
transform 1 0 24380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_265
timestamp 1
transform 1 0 25484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_273
timestamp 1
transform 1 0 26220 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_292
timestamp 1636968456
transform 1 0 27968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_304
timestamp 1
transform 1 0 29072 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_319
timestamp 1
transform 1 0 30452 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_337
timestamp 1
transform 1 0 32108 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_6
timestamp 1636968456
transform 1 0 1656 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_18
timestamp 1
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_26
timestamp 1
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_35
timestamp 1
transform 1 0 4324 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_67
timestamp 1
transform 1 0 7268 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_102
timestamp 1
transform 1 0 10488 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_123
timestamp 1
transform 1 0 12420 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_131
timestamp 1
transform 1 0 13156 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_138
timestamp 1
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1636968456
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_153
timestamp 1
transform 1 0 15180 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_171
timestamp 1
transform 1 0 16836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_181
timestamp 1
transform 1 0 17756 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_193
timestamp 1
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_197
timestamp 1
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_211
timestamp 1
transform 1 0 20516 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_219
timestamp 1
transform 1 0 21252 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_231
timestamp 1636968456
transform 1 0 22356 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_243
timestamp 1
transform 1 0 23460 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp 1
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_268
timestamp 1636968456
transform 1 0 25760 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_280
timestamp 1636968456
transform 1 0 26864 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_292
timestamp 1
transform 1 0 27968 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_309
timestamp 1
transform 1 0 29532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_330
timestamp 1
transform 1 0 31464 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_3
timestamp 1
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_11
timestamp 1
transform 1 0 2116 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_31
timestamp 1
transform 1 0 3956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_39
timestamp 1
transform 1 0 4692 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_67
timestamp 1
transform 1 0 7268 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_71
timestamp 1
transform 1 0 7636 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_96
timestamp 1
transform 1 0 9936 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_109
timestamp 1
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_113
timestamp 1
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_120
timestamp 1636968456
transform 1 0 12144 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_132
timestamp 1
transform 1 0 13248 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1636968456
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_169
timestamp 1
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_184
timestamp 1
transform 1 0 18032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_199
timestamp 1
transform 1 0 19412 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_205
timestamp 1
transform 1 0 19964 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_213
timestamp 1
transform 1 0 20700 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_221
timestamp 1
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1636968456
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_237
timestamp 1
transform 1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_241
timestamp 1
transform 1 0 23276 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_248
timestamp 1636968456
transform 1 0 23920 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_260
timestamp 1
transform 1 0 25024 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_266
timestamp 1
transform 1 0 25576 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_272
timestamp 1
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_281
timestamp 1
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_289
timestamp 1
transform 1 0 27692 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_296
timestamp 1636968456
transform 1 0 28336 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_308
timestamp 1636968456
transform 1 0 29440 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_337
timestamp 1
transform 1 0 32108 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1636968456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_15
timestamp 1
transform 1 0 2484 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_23
timestamp 1
transform 1 0 3220 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_33
timestamp 1
transform 1 0 4140 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_48
timestamp 1
transform 1 0 5520 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_66
timestamp 1636968456
transform 1 0 7176 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_78
timestamp 1
transform 1 0 8280 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_85
timestamp 1
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_91
timestamp 1
transform 1 0 9476 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_98
timestamp 1
transform 1 0 10120 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1636968456
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1636968456
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_141
timestamp 1
transform 1 0 14076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_147
timestamp 1
transform 1 0 14628 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_160
timestamp 1
transform 1 0 15824 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_172
timestamp 1636968456
transform 1 0 16928 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_184
timestamp 1636968456
transform 1 0 18032 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_197
timestamp 1
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_210
timestamp 1636968456
transform 1 0 20424 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_222
timestamp 1
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_237
timestamp 1
transform 1 0 22908 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_244
timestamp 1
transform 1 0 23552 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_253
timestamp 1
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_261
timestamp 1
transform 1 0 25116 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_268
timestamp 1636968456
transform 1 0 25760 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_280
timestamp 1
transform 1 0 26864 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_287
timestamp 1
transform 1 0 27508 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_296
timestamp 1636968456
transform 1 0 28336 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_309
timestamp 1
transform 1 0 29532 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_321
timestamp 1
transform 1 0 30636 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_325
timestamp 1
transform 1 0 31004 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1636968456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_15
timestamp 1
transform 1 0 2484 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_23
timestamp 1
transform 1 0 3220 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_31
timestamp 1
transform 1 0 3956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_36
timestamp 1
transform 1 0 4416 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_40
timestamp 1636968456
transform 1 0 4784 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_57
timestamp 1
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_67
timestamp 1636968456
transform 1 0 7268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_79
timestamp 1
transform 1 0 8372 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_85
timestamp 1636968456
transform 1 0 8924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_97
timestamp 1
transform 1 0 10028 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_101
timestamp 1
transform 1 0 10396 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_113
timestamp 1
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_121
timestamp 1
transform 1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_130
timestamp 1636968456
transform 1 0 13064 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_142
timestamp 1636968456
transform 1 0 14168 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_160
timestamp 1
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1636968456
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1636968456
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_193
timestamp 1
transform 1 0 18860 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_201
timestamp 1
transform 1 0 19596 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_225
timestamp 1
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_233
timestamp 1
transform 1 0 22540 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1636968456
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_261
timestamp 1
transform 1 0 25116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_270
timestamp 1
transform 1 0 25944 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1636968456
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1636968456
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_305
timestamp 1
transform 1 0 29164 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_317
timestamp 1
transform 1 0 30268 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_337
timestamp 1
transform 1 0 32108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_6
timestamp 1
transform 1 0 1656 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_14
timestamp 1
transform 1 0 2392 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_24
timestamp 1
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_29
timestamp 1
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_42
timestamp 1
transform 1 0 4968 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1636968456
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_65
timestamp 1
transform 1 0 7084 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_73
timestamp 1
transform 1 0 7820 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_80
timestamp 1
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_85
timestamp 1
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_94
timestamp 1
transform 1 0 9752 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_101
timestamp 1636968456
transform 1 0 10396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_113
timestamp 1636968456
transform 1 0 11500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_125
timestamp 1
transform 1 0 12604 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_137
timestamp 1
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_141
timestamp 1
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_147
timestamp 1
transform 1 0 14628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_173
timestamp 1
transform 1 0 17020 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_180
timestamp 1
transform 1 0 17664 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_194
timestamp 1
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_197
timestamp 1
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_203
timestamp 1
transform 1 0 19780 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_210
timestamp 1636968456
transform 1 0 20424 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_222
timestamp 1636968456
transform 1 0 21528 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_234
timestamp 1636968456
transform 1 0 22632 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_246
timestamp 1
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_253
timestamp 1
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_261
timestamp 1
transform 1 0 25116 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_268
timestamp 1636968456
transform 1 0 25760 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_280
timestamp 1
transform 1 0 26864 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_288
timestamp 1
transform 1 0 27600 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_302
timestamp 1
transform 1 0 28888 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1636968456
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_321
timestamp 1
transform 1 0 30636 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_332
timestamp 1
transform 1 0 31648 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_341
timestamp 1
transform 1 0 32476 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_3
timestamp 1
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_11
timestamp 1
transform 1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_21
timestamp 1636968456
transform 1 0 3036 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_33
timestamp 1
transform 1 0 4140 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_41
timestamp 1
transform 1 0 4876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_52
timestamp 1
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_79
timestamp 1
transform 1 0 8372 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_104
timestamp 1
transform 1 0 10672 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_113
timestamp 1
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_127
timestamp 1636968456
transform 1 0 12788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_142
timestamp 1
transform 1 0 14168 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_153
timestamp 1636968456
transform 1 0 15180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_165
timestamp 1
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_189
timestamp 1636968456
transform 1 0 18492 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_201
timestamp 1636968456
transform 1 0 19596 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_213
timestamp 1
transform 1 0 20700 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_221
timestamp 1
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_225
timestamp 1
transform 1 0 21804 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_240
timestamp 1
transform 1 0 23184 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_248
timestamp 1
transform 1 0 23920 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_257
timestamp 1
transform 1 0 24748 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_265
timestamp 1
transform 1 0 25484 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_271
timestamp 1
transform 1 0 26036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_287
timestamp 1
transform 1 0 27508 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1636968456
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_317
timestamp 1
transform 1 0 30268 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_337
timestamp 1
transform 1 0 32108 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1636968456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_15
timestamp 1
transform 1 0 2484 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_26
timestamp 1
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_29
timestamp 1
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_44
timestamp 1
transform 1 0 5152 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_52
timestamp 1636968456
transform 1 0 5888 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_64
timestamp 1
transform 1 0 6992 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_73
timestamp 1
transform 1 0 7820 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_81
timestamp 1
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_85
timestamp 1
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_93
timestamp 1
transform 1 0 9660 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_103
timestamp 1636968456
transform 1 0 10580 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_115
timestamp 1
transform 1 0 11684 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_119
timestamp 1
transform 1 0 12052 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_129
timestamp 1
transform 1 0 12972 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_150
timestamp 1
transform 1 0 14904 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_156
timestamp 1636968456
transform 1 0 15456 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_168
timestamp 1
transform 1 0 16560 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_182
timestamp 1636968456
transform 1 0 17848 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_194
timestamp 1
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_197
timestamp 1
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_208
timestamp 1
transform 1 0 20240 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_215
timestamp 1
transform 1 0 20884 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_223
timestamp 1
transform 1 0 21620 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_231
timestamp 1
transform 1 0 22356 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_243
timestamp 1
transform 1 0 23460 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_285
timestamp 1636968456
transform 1 0 27324 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_297
timestamp 1
transform 1 0 28428 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_303
timestamp 1
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1636968456
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_331
timestamp 1
transform 1 0 31556 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_340
timestamp 1
transform 1 0 32384 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_3
timestamp 1
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_11
timestamp 1
transform 1 0 2116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_30
timestamp 1
transform 1 0 3864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_36
timestamp 1
transform 1 0 4416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_47
timestamp 1
transform 1 0 5428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_57
timestamp 1
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_65
timestamp 1
transform 1 0 7084 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_76
timestamp 1636968456
transform 1 0 8096 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_88
timestamp 1
transform 1 0 9200 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_95
timestamp 1636968456
transform 1 0 9844 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_107
timestamp 1
transform 1 0 10948 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_113
timestamp 1
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_119
timestamp 1
transform 1 0 12052 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_125
timestamp 1
transform 1 0 12604 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_133
timestamp 1
transform 1 0 13340 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_137
timestamp 1
transform 1 0 13708 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_141
timestamp 1
transform 1 0 14076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_150
timestamp 1
transform 1 0 14904 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_156
timestamp 1636968456
transform 1 0 15456 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_169
timestamp 1
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_178
timestamp 1636968456
transform 1 0 17480 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_190
timestamp 1
transform 1 0 18584 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_197
timestamp 1636968456
transform 1 0 19228 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_209
timestamp 1636968456
transform 1 0 20332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_221
timestamp 1
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1636968456
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_237
timestamp 1
transform 1 0 22908 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_248
timestamp 1
transform 1 0 23920 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_276
timestamp 1
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_281
timestamp 1
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_289
timestamp 1
transform 1 0 27692 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_297
timestamp 1636968456
transform 1 0 28428 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_309
timestamp 1
transform 1 0 29532 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_316
timestamp 1
transform 1 0 30176 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_337
timestamp 1
transform 1 0 32108 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_19
timestamp 1
transform 1 0 2852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_37
timestamp 1
transform 1 0 4508 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_43
timestamp 1
transform 1 0 5060 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_47
timestamp 1
transform 1 0 5428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_51
timestamp 1
transform 1 0 5796 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_72
timestamp 1
transform 1 0 7728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_79
timestamp 1
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_85
timestamp 1
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_106
timestamp 1
transform 1 0 10856 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_128
timestamp 1636968456
transform 1 0 12880 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_141
timestamp 1
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_149
timestamp 1636968456
transform 1 0 14812 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_161
timestamp 1
transform 1 0 15916 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_169
timestamp 1
transform 1 0 16652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_184
timestamp 1636968456
transform 1 0 18032 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_203
timestamp 1636968456
transform 1 0 19780 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_215
timestamp 1
transform 1 0 20884 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_253
timestamp 1
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_264
timestamp 1636968456
transform 1 0 25392 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_276
timestamp 1636968456
transform 1 0 26496 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_288
timestamp 1636968456
transform 1 0 27600 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_300
timestamp 1
transform 1 0 28704 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_309
timestamp 1
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_317
timestamp 1
transform 1 0 30268 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_6
timestamp 1636968456
transform 1 0 1656 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_18
timestamp 1636968456
transform 1 0 2760 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_33
timestamp 1
transform 1 0 4140 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_40
timestamp 1
transform 1 0 4784 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_46
timestamp 1
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_54
timestamp 1
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1636968456
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_73
timestamp 1636968456
transform 1 0 7820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_85
timestamp 1636968456
transform 1 0 8924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_97
timestamp 1636968456
transform 1 0 10028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_109
timestamp 1
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_124
timestamp 1
transform 1 0 12512 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_132
timestamp 1
transform 1 0 13248 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1636968456
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1636968456
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_193
timestamp 1
transform 1 0 18860 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_201
timestamp 1
transform 1 0 19596 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_213
timestamp 1
transform 1 0 20700 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_221
timestamp 1
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_225
timestamp 1
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_233
timestamp 1
transform 1 0 22540 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_238
timestamp 1
transform 1 0 23000 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_244
timestamp 1
transform 1 0 23552 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_251
timestamp 1
transform 1 0 24196 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_259
timestamp 1
transform 1 0 24932 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_265
timestamp 1
transform 1 0 25484 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_278
timestamp 1
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_281
timestamp 1
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_294
timestamp 1
transform 1 0 28152 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_308
timestamp 1
transform 1 0 29440 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_314
timestamp 1
transform 1 0 29992 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_337
timestamp 1
transform 1 0 32108 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_26
timestamp 1
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_32
timestamp 1
transform 1 0 4048 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_52
timestamp 1
transform 1 0 5888 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_61
timestamp 1
transform 1 0 6716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_93
timestamp 1
transform 1 0 9660 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_103
timestamp 1636968456
transform 1 0 10580 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_115
timestamp 1
transform 1 0 11684 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_128
timestamp 1
transform 1 0 12880 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_150
timestamp 1636968456
transform 1 0 14904 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_162
timestamp 1
transform 1 0 16008 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_166
timestamp 1
transform 1 0 16376 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_173
timestamp 1636968456
transform 1 0 17020 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_185
timestamp 1
transform 1 0 18124 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_193
timestamp 1
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1636968456
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_209
timestamp 1
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_218
timestamp 1636968456
transform 1 0 21160 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_230
timestamp 1636968456
transform 1 0 22264 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_242
timestamp 1
transform 1 0 23368 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_250
timestamp 1
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_258
timestamp 1
transform 1 0 24840 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_266
timestamp 1
transform 1 0 25576 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_283
timestamp 1
transform 1 0 27140 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_289
timestamp 1
transform 1 0 27692 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_302
timestamp 1
transform 1 0 28888 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_324
timestamp 1
transform 1 0 30912 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_3
timestamp 1
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_40
timestamp 1
transform 1 0 4784 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_54
timestamp 1
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1636968456
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_69
timestamp 1
transform 1 0 7452 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_73
timestamp 1
transform 1 0 7820 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1636968456
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_93
timestamp 1
transform 1 0 9660 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_101
timestamp 1
transform 1 0 10396 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_110
timestamp 1
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1636968456
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_137
timestamp 1
transform 1 0 13708 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_148
timestamp 1
transform 1 0 14720 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_164
timestamp 1
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_175
timestamp 1
transform 1 0 17204 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_189
timestamp 1
transform 1 0 18492 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_198
timestamp 1
transform 1 0 19320 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_204
timestamp 1
transform 1 0 19872 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_211
timestamp 1
transform 1 0 20516 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_220
timestamp 1
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_225
timestamp 1
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_238
timestamp 1636968456
transform 1 0 23000 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_250
timestamp 1
transform 1 0 24104 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_257
timestamp 1636968456
transform 1 0 24748 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_269
timestamp 1
transform 1 0 25852 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_277
timestamp 1
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1636968456
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1636968456
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_305
timestamp 1
transform 1 0 29164 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_313
timestamp 1
transform 1 0 29900 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_319
timestamp 1
transform 1 0 30452 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_337
timestamp 1
transform 1 0 32108 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_3
timestamp 1
transform 1 0 1380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_26
timestamp 1
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_36
timestamp 1
transform 1 0 4416 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_57
timestamp 1636968456
transform 1 0 6348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_69
timestamp 1
transform 1 0 7452 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_85
timestamp 1
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_89
timestamp 1
transform 1 0 9292 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_141
timestamp 1
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_151
timestamp 1636968456
transform 1 0 14996 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_163
timestamp 1636968456
transform 1 0 16100 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_175
timestamp 1636968456
transform 1 0 17204 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_187
timestamp 1
transform 1 0 18308 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_197
timestamp 1
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_205
timestamp 1
transform 1 0 19964 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_210
timestamp 1636968456
transform 1 0 20424 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_228
timestamp 1636968456
transform 1 0 22080 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_240
timestamp 1636968456
transform 1 0 23184 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1636968456
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_265
timestamp 1
transform 1 0 25484 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_274
timestamp 1
transform 1 0 26312 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_280
timestamp 1
transform 1 0 26864 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_289
timestamp 1636968456
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_301
timestamp 1
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1636968456
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_321
timestamp 1
transform 1 0 30636 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_329
timestamp 1
transform 1 0 31372 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_19
timestamp 1
transform 1 0 2852 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_57
timestamp 1
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_77
timestamp 1
transform 1 0 8188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_85
timestamp 1
transform 1 0 8924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_113
timestamp 1
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_136
timestamp 1
transform 1 0 13616 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_144
timestamp 1
transform 1 0 14352 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_150
timestamp 1636968456
transform 1 0 14904 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_162
timestamp 1
transform 1 0 16008 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_169
timestamp 1
transform 1 0 16652 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_176
timestamp 1
transform 1 0 17296 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_189
timestamp 1
transform 1 0 18492 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_218
timestamp 1
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1636968456
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_237
timestamp 1
transform 1 0 22908 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_245
timestamp 1
transform 1 0 23644 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_260
timestamp 1636968456
transform 1 0 25024 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_272
timestamp 1
transform 1 0 26128 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_306
timestamp 1636968456
transform 1 0 29256 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_318
timestamp 1
transform 1 0 30360 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_337
timestamp 1
transform 1 0 32108 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_3
timestamp 1
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_9
timestamp 1
transform 1 0 1932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_45
timestamp 1
transform 1 0 5244 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_56
timestamp 1
transform 1 0 6256 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_69
timestamp 1
transform 1 0 7452 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_77
timestamp 1
transform 1 0 8188 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_93
timestamp 1
transform 1 0 9660 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_128
timestamp 1
transform 1 0 12880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_132
timestamp 1
transform 1 0 13248 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_141
timestamp 1
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_149
timestamp 1
transform 1 0 14812 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_156
timestamp 1636968456
transform 1 0 15456 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_168
timestamp 1
transform 1 0 16560 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_175
timestamp 1
transform 1 0 17204 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_184
timestamp 1
transform 1 0 18032 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_188
timestamp 1
transform 1 0 18400 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_220
timestamp 1
transform 1 0 21344 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_232
timestamp 1
transform 1 0 22448 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_240
timestamp 1
transform 1 0 23184 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1636968456
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_265
timestamp 1
transform 1 0 25484 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_274
timestamp 1636968456
transform 1 0 26312 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_286
timestamp 1636968456
transform 1 0 27416 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_298
timestamp 1
transform 1 0 28520 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_306
timestamp 1
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1636968456
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_321
timestamp 1
transform 1 0 30636 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_331
timestamp 1
transform 1 0 31556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_35
timestamp 1
transform 1 0 4324 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_43
timestamp 1
transform 1 0 5060 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_73
timestamp 1
transform 1 0 7820 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_88
timestamp 1
transform 1 0 9200 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_92
timestamp 1
transform 1 0 9568 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_98
timestamp 1
transform 1 0 10120 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_125
timestamp 1
transform 1 0 12604 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_132
timestamp 1636968456
transform 1 0 13248 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_144
timestamp 1636968456
transform 1 0 14352 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_156
timestamp 1
transform 1 0 15456 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_169
timestamp 1
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_177
timestamp 1
transform 1 0 17388 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_182
timestamp 1
transform 1 0 17848 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_190
timestamp 1
transform 1 0 18584 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_202
timestamp 1
transform 1 0 19688 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 1
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_231
timestamp 1
transform 1 0 22356 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_235
timestamp 1
transform 1 0 22724 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_239
timestamp 1636968456
transform 1 0 23092 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_251
timestamp 1
transform 1 0 24196 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_259
timestamp 1
transform 1 0 24932 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_265
timestamp 1636968456
transform 1 0 25484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_277
timestamp 1
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_281
timestamp 1
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_287
timestamp 1
transform 1 0 27508 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1636968456
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_305
timestamp 1
transform 1 0 29164 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_334
timestamp 1
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_337
timestamp 1
transform 1 0 32108 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_3
timestamp 1
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_26
timestamp 1
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_57
timestamp 1
transform 1 0 6348 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_80
timestamp 1
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1636968456
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_97
timestamp 1
transform 1 0 10028 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_126
timestamp 1636968456
transform 1 0 12696 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_138
timestamp 1
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_147
timestamp 1636968456
transform 1 0 14628 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_159
timestamp 1
transform 1 0 15732 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_167
timestamp 1636968456
transform 1 0 16468 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_187
timestamp 1
transform 1 0 18308 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 1
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_197
timestamp 1
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_203
timestamp 1
transform 1 0 19780 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_215
timestamp 1
transform 1 0 20884 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_221
timestamp 1
transform 1 0 21436 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_242
timestamp 1
transform 1 0 23368 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_250
timestamp 1
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_261
timestamp 1
transform 1 0 25116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_271
timestamp 1
transform 1 0 26036 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_281
timestamp 1636968456
transform 1 0 26956 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_293
timestamp 1
transform 1 0 28060 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_305
timestamp 1
transform 1 0 29164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_314
timestamp 1
transform 1 0 29992 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1636968456
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_60
timestamp 1636968456
transform 1 0 6624 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_72
timestamp 1
transform 1 0 7728 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_80
timestamp 1
transform 1 0 8464 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_90
timestamp 1
transform 1 0 9384 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_98
timestamp 1
transform 1 0 10120 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_108
timestamp 1
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_123
timestamp 1
transform 1 0 12420 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_132
timestamp 1
transform 1 0 13248 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_144
timestamp 1
transform 1 0 14352 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_150
timestamp 1
transform 1 0 14904 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_159
timestamp 1
transform 1 0 15732 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_174
timestamp 1
transform 1 0 17112 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_182
timestamp 1
transform 1 0 17848 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_189
timestamp 1636968456
transform 1 0 18492 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_201
timestamp 1
transform 1 0 19596 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 1636968456
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_225
timestamp 1
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_230
timestamp 1
transform 1 0 22264 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_236
timestamp 1
transform 1 0 22816 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_240
timestamp 1
transform 1 0 23184 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_256
timestamp 1636968456
transform 1 0 24656 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_268
timestamp 1
transform 1 0 25760 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_276
timestamp 1
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1636968456
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1636968456
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_305
timestamp 1
transform 1 0 29164 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_337
timestamp 1
transform 1 0 32108 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_6
timestamp 1
transform 1 0 1656 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_60
timestamp 1
transform 1 0 6624 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_70
timestamp 1
transform 1 0 7544 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_78
timestamp 1
transform 1 0 8280 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_112
timestamp 1
transform 1 0 11408 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1636968456
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1636968456
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1636968456
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 1636968456
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 1636968456
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 1
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1636968456
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_209
timestamp 1
transform 1 0 20332 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_218
timestamp 1
transform 1 0 21160 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_227
timestamp 1
transform 1 0 21988 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_235
timestamp 1
transform 1 0 22724 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_239
timestamp 1
transform 1 0 23092 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_243
timestamp 1
transform 1 0 23460 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_249
timestamp 1
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_253
timestamp 1
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_261
timestamp 1
transform 1 0 25116 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_268
timestamp 1636968456
transform 1 0 25760 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_280
timestamp 1
transform 1 0 26864 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_299
timestamp 1
transform 1 0 28612 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_309
timestamp 1
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_339
timestamp 1
transform 1 0 32292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_3
timestamp 1
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_7
timestamp 1
transform 1 0 1748 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_27
timestamp 1
transform 1 0 3588 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_45
timestamp 1
transform 1 0 5244 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_57
timestamp 1
transform 1 0 6348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_63
timestamp 1
transform 1 0 6900 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_71
timestamp 1
transform 1 0 7636 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_77
timestamp 1
transform 1 0 8188 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_95
timestamp 1636968456
transform 1 0 9844 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_107
timestamp 1
transform 1 0 10948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_120
timestamp 1
transform 1 0 12144 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_126
timestamp 1
transform 1 0 12696 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_133
timestamp 1
transform 1 0 13340 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_137
timestamp 1
transform 1 0 13708 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_152
timestamp 1636968456
transform 1 0 15088 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_164
timestamp 1
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_175
timestamp 1
transform 1 0 17204 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_184
timestamp 1
transform 1 0 18032 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_191
timestamp 1
transform 1 0 18676 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_200
timestamp 1
transform 1 0 19504 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_252
timestamp 1636968456
transform 1 0 24288 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_264
timestamp 1636968456
transform 1 0 25392 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_276
timestamp 1
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_281
timestamp 1
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_293
timestamp 1
transform 1 0 28060 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_300
timestamp 1636968456
transform 1 0 28704 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_312
timestamp 1
transform 1 0 29808 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_326
timestamp 1
transform 1 0 31096 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_337
timestamp 1
transform 1 0 32108 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_29
timestamp 1
transform 1 0 3772 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_39
timestamp 1
transform 1 0 4692 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_64
timestamp 1636968456
transform 1 0 6992 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_76
timestamp 1
transform 1 0 8096 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_111
timestamp 1
transform 1 0 11316 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_126
timestamp 1
transform 1 0 12696 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_141
timestamp 1
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_146
timestamp 1636968456
transform 1 0 14536 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_158
timestamp 1
transform 1 0 15640 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_187
timestamp 1
transform 1 0 18308 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_202
timestamp 1
transform 1 0 19688 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_217
timestamp 1
transform 1 0 21068 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_224
timestamp 1
transform 1 0 21712 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_229
timestamp 1
transform 1 0 22172 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_243
timestamp 1
transform 1 0 23460 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_253
timestamp 1
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_259
timestamp 1
transform 1 0 24932 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_273
timestamp 1
transform 1 0 26220 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_280
timestamp 1636968456
transform 1 0 26864 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_292
timestamp 1636968456
transform 1 0 27968 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_304
timestamp 1
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_314
timestamp 1
transform 1 0 29992 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_6
timestamp 1636968456
transform 1 0 1656 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_18
timestamp 1
transform 1 0 2760 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_35
timestamp 1
transform 1 0 4324 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_70
timestamp 1
transform 1 0 7544 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_76
timestamp 1
transform 1 0 8096 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_96
timestamp 1
transform 1 0 9936 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_100
timestamp 1
transform 1 0 10304 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_108
timestamp 1
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1636968456
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_125
timestamp 1
transform 1 0 12604 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_135
timestamp 1636968456
transform 1 0 13524 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_147
timestamp 1636968456
transform 1 0 14628 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_159
timestamp 1
transform 1 0 15732 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_173
timestamp 1
transform 1 0 17020 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_181
timestamp 1
transform 1 0 17756 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_188
timestamp 1
transform 1 0 18400 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_196
timestamp 1
transform 1 0 19136 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_213
timestamp 1
transform 1 0 20700 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_222
timestamp 1
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_231
timestamp 1
transform 1 0 22356 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_239
timestamp 1
transform 1 0 23092 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_243
timestamp 1
transform 1 0 23460 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_252
timestamp 1636968456
transform 1 0 24288 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_264
timestamp 1636968456
transform 1 0 25392 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_276
timestamp 1
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1636968456
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1636968456
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_305
timestamp 1
transform 1 0 29164 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_309
timestamp 1
transform 1 0 29532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_333
timestamp 1
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_337
timestamp 1
transform 1 0 32108 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_19
timestamp 1
transform 1 0 2852 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_55
timestamp 1
transform 1 0 6164 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_63
timestamp 1
transform 1 0 6900 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_91
timestamp 1
transform 1 0 9476 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_101
timestamp 1
transform 1 0 10396 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_123
timestamp 1
transform 1 0 12420 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_131
timestamp 1
transform 1 0 13156 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_141
timestamp 1
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_147
timestamp 1
transform 1 0 14628 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_154
timestamp 1
transform 1 0 15272 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_168
timestamp 1636968456
transform 1 0 16560 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_180
timestamp 1
transform 1 0 17664 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_193
timestamp 1
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1636968456
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_209
timestamp 1
transform 1 0 20332 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_217
timestamp 1
transform 1 0 21068 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_226
timestamp 1
transform 1 0 21896 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_234
timestamp 1
transform 1 0 22632 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 1
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1636968456
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1636968456
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_292
timestamp 1
transform 1 0 27968 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 1
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1636968456
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_321
timestamp 1
transform 1 0 30636 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_332
timestamp 1
transform 1 0 31648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_3
timestamp 1
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_9
timestamp 1
transform 1 0 1932 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_35
timestamp 1
transform 1 0 4324 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_47
timestamp 1
transform 1 0 5428 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_54
timestamp 1
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_81
timestamp 1
transform 1 0 8556 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_109
timestamp 1
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1636968456
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_125
timestamp 1
transform 1 0 12604 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_151
timestamp 1636968456
transform 1 0 14996 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_163
timestamp 1
transform 1 0 16100 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_169
timestamp 1
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_174
timestamp 1
transform 1 0 17112 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_182
timestamp 1
transform 1 0 17848 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_186
timestamp 1
transform 1 0 18216 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_195
timestamp 1
transform 1 0 19044 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 1636968456
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 1
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_225
timestamp 1
transform 1 0 21804 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_231
timestamp 1
transform 1 0 22356 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_237
timestamp 1
transform 1 0 22908 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_247
timestamp 1636968456
transform 1 0 23828 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_265
timestamp 1
transform 1 0 25484 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_272
timestamp 1
transform 1 0 26128 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_287
timestamp 1
transform 1 0 27508 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_300
timestamp 1636968456
transform 1 0 28704 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_312
timestamp 1636968456
transform 1 0 29808 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_331
timestamp 1
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_337
timestamp 1
transform 1 0 32108 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_6
timestamp 1
transform 1 0 1656 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_29
timestamp 1
transform 1 0 3772 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_50
timestamp 1
transform 1 0 5704 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_60
timestamp 1
transform 1 0 6624 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_80
timestamp 1
transform 1 0 8464 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_85
timestamp 1
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_101
timestamp 1
transform 1 0 10396 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_158
timestamp 1
transform 1 0 15640 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_166
timestamp 1
transform 1 0 16376 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_182
timestamp 1
transform 1 0 17848 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_190
timestamp 1
transform 1 0 18584 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_213
timestamp 1636968456
transform 1 0 20700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_225
timestamp 1
transform 1 0 21804 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_229
timestamp 1
transform 1 0 22172 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_236
timestamp 1
transform 1 0 22816 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1636968456
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_265
timestamp 1
transform 1 0 25484 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_273
timestamp 1
transform 1 0 26220 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_282
timestamp 1636968456
transform 1 0 27048 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_294
timestamp 1636968456
transform 1 0 28152 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_306
timestamp 1
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1636968456
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1636968456
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_333
timestamp 1
transform 1 0 31740 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_341
timestamp 1
transform 1 0 32476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_19
timestamp 1
transform 1 0 2852 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_29
timestamp 1
transform 1 0 3772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_88
timestamp 1
transform 1 0 9200 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_113
timestamp 1
transform 1 0 11500 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_130
timestamp 1
transform 1 0 13064 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_136
timestamp 1
transform 1 0 13616 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_143
timestamp 1
transform 1 0 14260 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_156
timestamp 1636968456
transform 1 0 15456 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_169
timestamp 1
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_185
timestamp 1
transform 1 0 18124 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_191
timestamp 1
transform 1 0 18676 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_199
timestamp 1
transform 1 0 19412 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 1
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_234
timestamp 1
transform 1 0 22632 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_240
timestamp 1
transform 1 0 23184 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_247
timestamp 1
transform 1 0 23828 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_255
timestamp 1
transform 1 0 24564 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_268
timestamp 1636968456
transform 1 0 25760 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1636968456
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1636968456
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1636968456
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 1636968456
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 1
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 1
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_337
timestamp 1
transform 1 0 32108 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_341
timestamp 1
transform 1 0 32476 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_55
timestamp 1
transform 1 0 6164 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_59
timestamp 1
transform 1 0 6532 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_69
timestamp 1
transform 1 0 7452 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_74
timestamp 1
transform 1 0 7912 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_92
timestamp 1
transform 1 0 9568 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_97
timestamp 1
transform 1 0 10028 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_109
timestamp 1
transform 1 0 11132 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_138
timestamp 1
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_147
timestamp 1636968456
transform 1 0 14628 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_159
timestamp 1
transform 1 0 15732 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_168
timestamp 1
transform 1 0 16560 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_184
timestamp 1
transform 1 0 18032 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_190
timestamp 1
transform 1 0 18584 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_197
timestamp 1
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_201
timestamp 1
transform 1 0 19596 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_218
timestamp 1636968456
transform 1 0 21160 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_230
timestamp 1
transform 1 0 22264 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_238
timestamp 1
transform 1 0 23000 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1636968456
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1636968456
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 1636968456
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 1636968456
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 1
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1636968456
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 1636968456
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_333
timestamp 1
transform 1 0 31740 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_341
timestamp 1
transform 1 0 32476 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_6
timestamp 1
transform 1 0 1656 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_14
timestamp 1
transform 1 0 2392 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_21
timestamp 1
transform 1 0 3036 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_25
timestamp 1
transform 1 0 3404 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_35
timestamp 1
transform 1 0 4324 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_48
timestamp 1
transform 1 0 5520 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_57
timestamp 1
transform 1 0 6348 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_63
timestamp 1
transform 1 0 6900 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_76
timestamp 1
transform 1 0 8096 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_91
timestamp 1
transform 1 0 9476 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_116
timestamp 1
transform 1 0 11776 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_130
timestamp 1636968456
transform 1 0 13064 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_142
timestamp 1636968456
transform 1 0 14168 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_154
timestamp 1
transform 1 0 15272 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_160
timestamp 1
transform 1 0 15824 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_166
timestamp 1
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_176
timestamp 1
transform 1 0 17296 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_189
timestamp 1636968456
transform 1 0 18492 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_201
timestamp 1
transform 1 0 19596 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_210
timestamp 1636968456
transform 1 0 20424 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_222
timestamp 1
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_225
timestamp 1
transform 1 0 21804 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_233
timestamp 1
transform 1 0 22540 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_241
timestamp 1
transform 1 0 23276 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_246
timestamp 1
transform 1 0 23736 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_263
timestamp 1636968456
transform 1 0 25300 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_275
timestamp 1
transform 1 0 26404 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1636968456
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1636968456
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 1636968456
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 1636968456
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 1
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_337
timestamp 1
transform 1 0 32108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_341
timestamp 1
transform 1 0 32476 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1636968456
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_15
timestamp 1
transform 1 0 2484 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_19
timestamp 1
transform 1 0 2852 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_26
timestamp 1
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1636968456
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1636968456
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1636968456
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1636968456
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_85
timestamp 1
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_90
timestamp 1
transform 1 0 9384 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_94
timestamp 1
transform 1 0 9752 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_106
timestamp 1636968456
transform 1 0 10856 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_118
timestamp 1636968456
transform 1 0 11960 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_130
timestamp 1
transform 1 0 13064 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_138
timestamp 1
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1636968456
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_153
timestamp 1
transform 1 0 15180 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_192
timestamp 1
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1636968456
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_209
timestamp 1
transform 1 0 20332 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_220
timestamp 1
transform 1 0 21344 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_269
timestamp 1636968456
transform 1 0 25852 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_281
timestamp 1636968456
transform 1 0 26956 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_293
timestamp 1636968456
transform 1 0 28060 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_305
timestamp 1
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1636968456
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 1636968456
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_333
timestamp 1
transform 1 0 31740 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_341
timestamp 1
transform 1 0 32476 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1636968456
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1636968456
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1636968456
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1636968456
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1636968456
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1636968456
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1636968456
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1636968456
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1636968456
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1636968456
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1636968456
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1636968456
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_169
timestamp 1
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_201
timestamp 1
transform 1 0 19596 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_207
timestamp 1
transform 1 0 20148 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_236
timestamp 1636968456
transform 1 0 22816 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_248
timestamp 1636968456
transform 1 0 23920 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_260
timestamp 1636968456
transform 1 0 25024 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_272
timestamp 1
transform 1 0 26128 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1636968456
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1636968456
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 1636968456
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 1636968456
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 1
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_337
timestamp 1
transform 1 0 32108 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_341
timestamp 1
transform 1 0 32476 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1636968456
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1636968456
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1636968456
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1636968456
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1636968456
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1636968456
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1636968456
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1636968456
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 1636968456
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1636968456
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1636968456
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 1636968456
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 1636968456
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 1636968456
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 1
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1636968456
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1636968456
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 1636968456
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 1636968456
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 1
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1636968456
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1636968456
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 1636968456
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 1636968456
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 1
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1636968456
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1636968456
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_333
timestamp 1
transform 1 0 31740 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_341
timestamp 1
transform 1 0 32476 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1636968456
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1636968456
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_27
timestamp 1
transform 1 0 3588 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_29
timestamp 1636968456
transform 1 0 3772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_41
timestamp 1636968456
transform 1 0 4876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_53
timestamp 1
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1636968456
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1636968456
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_81
timestamp 1
transform 1 0 8556 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_85
timestamp 1636968456
transform 1 0 8924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_97
timestamp 1636968456
transform 1 0 10028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_109
timestamp 1
transform 1 0 11132 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1636968456
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1636968456
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_137
timestamp 1
transform 1 0 13708 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_141
timestamp 1636968456
transform 1 0 14076 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_153
timestamp 1636968456
transform 1 0 15180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_165
timestamp 1
transform 1 0 16284 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_169
timestamp 1
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_177
timestamp 1636968456
transform 1 0 17388 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_189
timestamp 1
transform 1 0 18492 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_195
timestamp 1
transform 1 0 19044 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_203
timestamp 1636968456
transform 1 0 19780 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_215
timestamp 1
transform 1 0 20884 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_231
timestamp 1
transform 1 0 22356 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_239
timestamp 1
transform 1 0 23092 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_247
timestamp 1
transform 1 0 23828 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_251
timestamp 1
transform 1 0 24196 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_253
timestamp 1
transform 1 0 24380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_261
timestamp 1
transform 1 0 25116 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_268
timestamp 1636968456
transform 1 0 25760 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1636968456
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 1636968456
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_305
timestamp 1
transform 1 0 29164 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_309
timestamp 1636968456
transform 1 0 29532 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_321
timestamp 1636968456
transform 1 0 30636 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_333
timestamp 1
transform 1 0 31740 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_337
timestamp 1
transform 1 0 32108 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_341
timestamp 1
transform 1 0 32476 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 19964 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform -1 0 32016 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 32016 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 32016 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform -1 0 32384 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform -1 0 32476 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform -1 0 32016 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 32016 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform -1 0 32292 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform -1 0 32568 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform -1 0 32568 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform -1 0 32292 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform -1 0 32016 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform -1 0 32568 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform -1 0 32384 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 32384 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 31556 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform -1 0 23736 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform -1 0 17572 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform -1 0 30820 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform -1 0 25852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform 1 0 20884 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform -1 0 26036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform -1 0 31648 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform -1 0 32016 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 22540 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform -1 0 25300 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform -1 0 31096 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform -1 0 24196 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform -1 0 18124 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform -1 0 19596 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform -1 0 1656 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform -1 0 1656 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform -1 0 1656 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform -1 0 1656 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform -1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform -1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1
transform -1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1
transform 1 0 32292 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1
transform -1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1
transform 1 0 32200 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1
transform 1 0 32200 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1
transform -1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1
transform 1 0 32200 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1
transform -1 0 32568 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1
transform -1 0 17388 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1
transform 1 0 32200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1
transform 1 0 32200 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1
transform 1 0 32200 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1
transform 1 0 32200 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1
transform -1 0 32568 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1
transform 1 0 32108 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1
transform 1 0 32200 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1
transform 1 0 32200 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1
transform 1 0 32200 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1
transform 1 0 32200 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1
transform 1 0 32200 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1
transform 1 0 32200 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1
transform 1 0 32200 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1
transform 1 0 19228 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1
transform -1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1
transform 1 0 32200 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1
transform -1 0 31096 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1
transform 1 0 21804 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1
transform -1 0 24932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1
transform -1 0 23828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1
transform 1 0 25208 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1
transform 1 0 32200 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_54
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 32844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_55
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 32844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_56
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_57
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 32844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_58
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 32844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_59
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 32844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_60
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 32844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_61
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 32844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_62
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 32844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_63
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 32844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_64
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 32844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_65
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 32844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_66
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 32844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_67
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 32844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_68
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 32844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_69
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 32844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_70
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 32844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_71
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 32844 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_72
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 32844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_73
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 32844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_74
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 32844 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_75
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 32844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_76
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 32844 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_77
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 32844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_78
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 32844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_79
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 32844 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_80
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 32844 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_81
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 32844 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_82
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 32844 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_83
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 32844 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_84
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 32844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_85
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 32844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_86
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 32844 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_87
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 32844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_88
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 32844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_89
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 32844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_90
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 32844 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_91
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 32844 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_92
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 32844 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_93
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1
transform -1 0 32844 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_94
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1
transform -1 0 32844 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_95
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1
transform -1 0 32844 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_96
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1
transform -1 0 32844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_97
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1
transform -1 0 32844 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_98
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1
transform -1 0 32844 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_99
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1
transform -1 0 32844 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_100
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1
transform -1 0 32844 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_101
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1
transform -1 0 32844 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_102
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1
transform -1 0 32844 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_103
timestamp 1
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1
transform -1 0 32844 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_104
timestamp 1
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1
transform -1 0 32844 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_105
timestamp 1
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1
transform -1 0 32844 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_106
timestamp 1
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1
transform -1 0 32844 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_107
timestamp 1
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1
transform -1 0 32844 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_108
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_109
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_110
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_111
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_112
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_113
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_114
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_115
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_116
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_117
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_118
timestamp 1
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_119
timestamp 1
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_120
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_121
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_122
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_123
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_124
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_125
timestamp 1
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_126
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_127
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_128
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_129
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_130
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_131
timestamp 1
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_132
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_133
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_134
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_135
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_136
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_137
timestamp 1
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_138
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_139
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_140
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_141
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_142
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_143
timestamp 1
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_144
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_145
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_146
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_147
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_148
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_149
timestamp 1
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_150
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_151
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_152
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_153
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_154
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_155
timestamp 1
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_156
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_157
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_158
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_159
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_160
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_161
timestamp 1
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_162
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_163
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_164
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_165
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_166
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_167
timestamp 1
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_168
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_169
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_170
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_171
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_172
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_173
timestamp 1
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_174
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_175
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_176
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_177
timestamp 1
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_178
timestamp 1
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_179
timestamp 1
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_180
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_181
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_182
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_183
timestamp 1
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_184
timestamp 1
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_185
timestamp 1
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_186
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_187
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_188
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_189
timestamp 1
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_190
timestamp 1
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_191
timestamp 1
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_192
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_193
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_194
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_195
timestamp 1
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_196
timestamp 1
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_197
timestamp 1
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_198
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_199
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_200
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_201
timestamp 1
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_202
timestamp 1
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_203
timestamp 1
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_204
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_205
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_206
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_207
timestamp 1
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_208
timestamp 1
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_209
timestamp 1
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_210
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_211
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_212
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_213
timestamp 1
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_214
timestamp 1
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_215
timestamp 1
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_216
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_217
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_218
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_219
timestamp 1
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_220
timestamp 1
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_221
timestamp 1
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_222
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_223
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_224
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_225
timestamp 1
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_226
timestamp 1
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_227
timestamp 1
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_228
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_229
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_230
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_231
timestamp 1
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_232
timestamp 1
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_233
timestamp 1
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_234
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_235
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_236
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_237
timestamp 1
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_238
timestamp 1
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_239
timestamp 1
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_240
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_241
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_242
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_243
timestamp 1
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_244
timestamp 1
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_245
timestamp 1
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_246
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_247
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_248
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_249
timestamp 1
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_250
timestamp 1
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_251
timestamp 1
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_252
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_253
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_254
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_255
timestamp 1
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_256
timestamp 1
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_257
timestamp 1
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_258
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_259
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_260
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_261
timestamp 1
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_262
timestamp 1
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_263
timestamp 1
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_264
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_265
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_266
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_267
timestamp 1
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_268
timestamp 1
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_269
timestamp 1
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_270
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_271
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_272
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_273
timestamp 1
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_274
timestamp 1
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_275
timestamp 1
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_276
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_277
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_278
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_279
timestamp 1
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_280
timestamp 1
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_281
timestamp 1
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_282
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_283
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_284
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_285
timestamp 1
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_286
timestamp 1
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_287
timestamp 1
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_288
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_289
timestamp 1
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_290
timestamp 1
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_291
timestamp 1
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_292
timestamp 1
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_293
timestamp 1
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_294
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_295
timestamp 1
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_296
timestamp 1
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_297
timestamp 1
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_298
timestamp 1
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_299
timestamp 1
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_300
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_301
timestamp 1
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_302
timestamp 1
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_303
timestamp 1
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_304
timestamp 1
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_305
timestamp 1
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_306
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_307
timestamp 1
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_308
timestamp 1
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_309
timestamp 1
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_310
timestamp 1
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_311
timestamp 1
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_312
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_313
timestamp 1
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_314
timestamp 1
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_315
timestamp 1
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_316
timestamp 1
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_317
timestamp 1
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_318
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_319
timestamp 1
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_320
timestamp 1
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_321
timestamp 1
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_322
timestamp 1
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_323
timestamp 1
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_324
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_325
timestamp 1
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_326
timestamp 1
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_327
timestamp 1
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_328
timestamp 1
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_329
timestamp 1
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_330
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_331
timestamp 1
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_332
timestamp 1
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_333
timestamp 1
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_334
timestamp 1
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_335
timestamp 1
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_336
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_337
timestamp 1
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_338
timestamp 1
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_339
timestamp 1
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_340
timestamp 1
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_341
timestamp 1
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_342
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_343
timestamp 1
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_344
timestamp 1
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_345
timestamp 1
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_346
timestamp 1
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_347
timestamp 1
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_348
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_349
timestamp 1
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_350
timestamp 1
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_351
timestamp 1
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_352
timestamp 1
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_353
timestamp 1
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_354
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_355
timestamp 1
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_356
timestamp 1
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_357
timestamp 1
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_358
timestamp 1
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_359
timestamp 1
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_360
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_361
timestamp 1
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_362
timestamp 1
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_363
timestamp 1
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_364
timestamp 1
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_365
timestamp 1
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_366
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_367
timestamp 1
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_368
timestamp 1
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_369
timestamp 1
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_370
timestamp 1
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_371
timestamp 1
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_372
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_373
timestamp 1
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_374
timestamp 1
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_375
timestamp 1
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_376
timestamp 1
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_377
timestamp 1
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_378
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_379
timestamp 1
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_380
timestamp 1
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_381
timestamp 1
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_382
timestamp 1
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_383
timestamp 1
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_384
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_385
timestamp 1
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_386
timestamp 1
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_387
timestamp 1
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_388
timestamp 1
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_389
timestamp 1
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_390
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_391
timestamp 1
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_392
timestamp 1
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_393
timestamp 1
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_394
timestamp 1
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_395
timestamp 1
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_396
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_397
timestamp 1
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_398
timestamp 1
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_399
timestamp 1
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_400
timestamp 1
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_401
timestamp 1
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_402
timestamp 1
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_403
timestamp 1
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_404
timestamp 1
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_405
timestamp 1
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_406
timestamp 1
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_407
timestamp 1
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_408
timestamp 1
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_409
timestamp 1
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_410
timestamp 1
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_411
timestamp 1
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_412
timestamp 1
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_413
timestamp 1
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_414
timestamp 1
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_415
timestamp 1
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_416
timestamp 1
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_417
timestamp 1
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_418
timestamp 1
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_419
timestamp 1
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_420
timestamp 1
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_421
timestamp 1
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_422
timestamp 1
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_423
timestamp 1
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_424
timestamp 1
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_425
timestamp 1
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_426
timestamp 1
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_427
timestamp 1
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_428
timestamp 1
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_429
timestamp 1
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_430
timestamp 1
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_431
timestamp 1
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_432
timestamp 1
transform 1 0 3680 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_433
timestamp 1
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_434
timestamp 1
transform 1 0 8832 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_435
timestamp 1
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_436
timestamp 1
transform 1 0 13984 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_437
timestamp 1
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_438
timestamp 1
transform 1 0 19136 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_439
timestamp 1
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_440
timestamp 1
transform 1 0 24288 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_441
timestamp 1
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_442
timestamp 1
transform 1 0 29440 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_443
timestamp 1
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire57
timestamp 1
transform -1 0 25760 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  wire274
timestamp 1
transform 1 0 13432 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire465
timestamp 1
transform -1 0 3772 0 -1 29376
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 addr0[0]
port 0 nsew signal input
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 addr0[1]
port 1 nsew signal input
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 addr0[2]
port 2 nsew signal input
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 addr0[3]
port 3 nsew signal input
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 addr0[4]
port 4 nsew signal input
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 addr0[5]
port 5 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 addr0[6]
port 6 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 addr0[7]
port 7 nsew signal input
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 clk0
port 8 nsew signal input
flabel metal3 s 33200 12928 34000 13048 0 FreeSans 480 0 0 0 cs0
port 9 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 dout0[0]
port 10 nsew signal output
flabel metal3 s 33200 23128 34000 23248 0 FreeSans 480 0 0 0 dout0[10]
port 11 nsew signal output
flabel metal3 s 33200 20408 34000 20528 0 FreeSans 480 0 0 0 dout0[11]
port 12 nsew signal output
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 dout0[12]
port 13 nsew signal output
flabel metal3 s 33200 8168 34000 8288 0 FreeSans 480 0 0 0 dout0[13]
port 14 nsew signal output
flabel metal3 s 33200 25848 34000 25968 0 FreeSans 480 0 0 0 dout0[14]
port 15 nsew signal output
flabel metal2 s 16762 33200 16818 34000 0 FreeSans 224 90 0 0 dout0[15]
port 16 nsew signal output
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 dout0[16]
port 17 nsew signal output
flabel metal3 s 33200 10208 34000 10328 0 FreeSans 480 0 0 0 dout0[17]
port 18 nsew signal output
flabel metal3 s 33200 14968 34000 15088 0 FreeSans 480 0 0 0 dout0[18]
port 19 nsew signal output
flabel metal3 s 33200 13608 34000 13728 0 FreeSans 480 0 0 0 dout0[19]
port 20 nsew signal output
flabel metal3 s 33200 23808 34000 23928 0 FreeSans 480 0 0 0 dout0[1]
port 21 nsew signal output
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 dout0[20]
port 22 nsew signal output
flabel metal3 s 33200 9528 34000 9648 0 FreeSans 480 0 0 0 dout0[21]
port 23 nsew signal output
flabel metal3 s 33200 6808 34000 6928 0 FreeSans 480 0 0 0 dout0[22]
port 24 nsew signal output
flabel metal3 s 33200 17688 34000 17808 0 FreeSans 480 0 0 0 dout0[23]
port 25 nsew signal output
flabel metal3 s 33200 7488 34000 7608 0 FreeSans 480 0 0 0 dout0[24]
port 26 nsew signal output
flabel metal3 s 33200 15648 34000 15768 0 FreeSans 480 0 0 0 dout0[25]
port 27 nsew signal output
flabel metal3 s 33200 22448 34000 22568 0 FreeSans 480 0 0 0 dout0[26]
port 28 nsew signal output
flabel metal3 s 33200 19048 34000 19168 0 FreeSans 480 0 0 0 dout0[27]
port 29 nsew signal output
flabel metal3 s 33200 17008 34000 17128 0 FreeSans 480 0 0 0 dout0[28]
port 30 nsew signal output
flabel metal3 s 33200 11568 34000 11688 0 FreeSans 480 0 0 0 dout0[29]
port 31 nsew signal output
flabel metal2 s 18694 33200 18750 34000 0 FreeSans 224 90 0 0 dout0[2]
port 32 nsew signal output
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 dout0[30]
port 33 nsew signal output
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 dout0[31]
port 34 nsew signal output
flabel metal3 s 33200 19728 34000 19848 0 FreeSans 480 0 0 0 dout0[3]
port 35 nsew signal output
flabel metal3 s 33200 24488 34000 24608 0 FreeSans 480 0 0 0 dout0[4]
port 36 nsew signal output
flabel metal2 s 21270 33200 21326 34000 0 FreeSans 224 90 0 0 dout0[5]
port 37 nsew signal output
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 dout0[6]
port 38 nsew signal output
flabel metal2 s 23202 33200 23258 34000 0 FreeSans 224 90 0 0 dout0[7]
port 39 nsew signal output
flabel metal2 s 25134 33200 25190 34000 0 FreeSans 224 90 0 0 dout0[8]
port 40 nsew signal output
flabel metal3 s 33200 21088 34000 21208 0 FreeSans 480 0 0 0 dout0[9]
port 41 nsew signal output
flabel metal4 s 4208 2128 4528 31600 0 FreeSans 1920 90 0 0 vccd1
port 42 nsew power bidirectional
flabel metal4 s 4868 2128 5188 31600 0 FreeSans 1920 90 0 0 vssd1
port 43 nsew ground bidirectional
rlabel metal1 16974 31008 16974 31008 0 vccd1
rlabel metal1 16974 31552 16974 31552 0 vssd1
rlabel metal2 18814 3876 18814 3876 0 _0000_
rlabel metal2 30498 23970 30498 23970 0 _0001_
rlabel metal2 18722 30022 18722 30022 0 _0002_
rlabel metal1 30482 22678 30482 22678 0 _0003_
rlabel metal1 30114 23766 30114 23766 0 _0004_
rlabel metal1 20654 29818 20654 29818 0 _0005_
rlabel metal1 25060 4590 25060 4590 0 _0006_
rlabel metal2 22494 29410 22494 29410 0 _0007_
rlabel metal2 24518 29410 24518 29410 0 _0008_
rlabel metal2 31326 21318 31326 21318 0 _0009_
rlabel metal1 30390 25942 30390 25942 0 _0010_
rlabel metal1 31316 19822 31316 19822 0 _0011_
rlabel via1 22489 4114 22489 4114 0 _0012_
rlabel metal1 31316 7854 31316 7854 0 _0013_
rlabel via1 31413 25262 31413 25262 0 _0014_
rlabel metal2 17250 29274 17250 29274 0 _0015_
rlabel via1 24145 4114 24145 4114 0 _0016_
rlabel metal1 30304 9554 30304 9554 0 _0017_
rlabel metal2 31786 13702 31786 13702 0 _0018_
rlabel metal1 31040 11118 31040 11118 0 _0019_
rlabel metal1 21532 3502 21532 3502 0 _0020_
rlabel metal1 31080 8874 31080 8874 0 _0021_
rlabel metal1 31218 6698 31218 6698 0 _0022_
rlabel metal1 31316 18734 31316 18734 0 _0023_
rlabel metal1 29608 7786 29608 7786 0 _0024_
rlabel metal1 31316 15470 31316 15470 0 _0025_
rlabel metal2 31510 22610 31510 22610 0 _0026_
rlabel metal1 31464 17850 31464 17850 0 _0027_
rlabel metal2 31602 16966 31602 16966 0 _0028_
rlabel metal1 31183 11798 31183 11798 0 _0029_
rlabel metal2 16790 3876 16790 3876 0 _0030_
rlabel metal1 7084 28730 7084 28730 0 _0031_
rlabel metal1 19274 19210 19274 19210 0 _0032_
rlabel via2 12190 18411 12190 18411 0 _0033_
rlabel metal2 23782 25143 23782 25143 0 _0034_
rlabel metal1 23460 17850 23460 17850 0 _0035_
rlabel metal2 21850 18564 21850 18564 0 _0036_
rlabel metal2 21850 8092 21850 8092 0 _0037_
rlabel metal1 26450 16966 26450 16966 0 _0038_
rlabel metal2 2162 25075 2162 25075 0 _0039_
rlabel metal2 5382 25279 5382 25279 0 _0040_
rlabel metal2 11086 24786 11086 24786 0 _0041_
rlabel metal2 13202 23970 13202 23970 0 _0042_
rlabel metal2 21022 25823 21022 25823 0 _0043_
rlabel metal2 14674 23018 14674 23018 0 _0044_
rlabel metal2 10258 24684 10258 24684 0 _0045_
rlabel metal1 13340 23494 13340 23494 0 _0046_
rlabel metal1 23966 25296 23966 25296 0 _0047_
rlabel metal1 23000 26554 23000 26554 0 _0048_
rlabel metal1 25852 17646 25852 17646 0 _0049_
rlabel metal1 3450 28390 3450 28390 0 _0050_
rlabel metal1 18262 27982 18262 27982 0 _0051_
rlabel metal2 12006 22236 12006 22236 0 _0052_
rlabel metal2 14306 28322 14306 28322 0 _0053_
rlabel metal1 18768 28390 18768 28390 0 _0054_
rlabel via2 19366 7429 19366 7429 0 _0055_
rlabel metal2 18630 27761 18630 27761 0 _0056_
rlabel metal1 13892 25874 13892 25874 0 _0057_
rlabel metal1 13202 25908 13202 25908 0 _0058_
rlabel metal3 14628 17952 14628 17952 0 _0059_
rlabel metal2 13754 26180 13754 26180 0 _0060_
rlabel metal2 10442 24497 10442 24497 0 _0061_
rlabel metal1 23046 7378 23046 7378 0 _0062_
rlabel metal1 7406 24072 7406 24072 0 _0063_
rlabel metal1 14168 19822 14168 19822 0 _0064_
rlabel metal1 14306 19482 14306 19482 0 _0065_
rlabel metal3 18492 24072 18492 24072 0 _0066_
rlabel metal2 14306 23902 14306 23902 0 _0067_
rlabel metal1 21574 22406 21574 22406 0 _0068_
rlabel metal1 27692 24038 27692 24038 0 _0069_
rlabel metal2 13478 28543 13478 28543 0 _0070_
rlabel metal2 14122 30464 14122 30464 0 _0071_
rlabel metal2 14030 28067 14030 28067 0 _0072_
rlabel metal3 29233 20468 29233 20468 0 _0073_
rlabel metal2 8234 19907 8234 19907 0 _0074_
rlabel metal1 28152 19686 28152 19686 0 _0075_
rlabel metal1 9200 18394 9200 18394 0 _0076_
rlabel metal1 28612 17646 28612 17646 0 _0077_
rlabel metal2 3358 19482 3358 19482 0 _0078_
rlabel metal2 3450 19754 3450 19754 0 _0079_
rlabel metal1 6026 9350 6026 9350 0 _0080_
rlabel metal3 17388 18768 17388 18768 0 _0081_
rlabel via2 7682 18581 7682 18581 0 _0082_
rlabel metal1 4830 23528 4830 23528 0 _0083_
rlabel metal2 6900 17170 6900 17170 0 _0084_
rlabel metal2 23230 26588 23230 26588 0 _0085_
rlabel metal1 27324 21318 27324 21318 0 _0086_
rlabel metal2 2346 15028 2346 15028 0 _0087_
rlabel metal1 16928 8806 16928 8806 0 _0088_
rlabel metal2 14398 4862 14398 4862 0 _0089_
rlabel metal1 17250 9146 17250 9146 0 _0090_
rlabel metal2 32706 11356 32706 11356 0 _0091_
rlabel metal1 20286 8840 20286 8840 0 _0092_
rlabel metal1 26588 17170 26588 17170 0 _0093_
rlabel metal1 2990 15130 2990 15130 0 _0094_
rlabel via2 24150 13685 24150 13685 0 _0095_
rlabel metal2 19458 22423 19458 22423 0 _0096_
rlabel via2 17618 23035 17618 23035 0 _0097_
rlabel metal1 23690 14348 23690 14348 0 _0098_
rlabel metal3 17089 11900 17089 11900 0 _0099_
rlabel metal2 25254 14178 25254 14178 0 _0100_
rlabel metal1 6716 9078 6716 9078 0 _0101_
rlabel metal2 15134 11407 15134 11407 0 _0102_
rlabel metal2 2530 11764 2530 11764 0 _0103_
rlabel metal1 9062 5712 9062 5712 0 _0104_
rlabel metal2 23046 6052 23046 6052 0 _0105_
rlabel metal1 23138 16014 23138 16014 0 _0106_
rlabel metal1 17480 11050 17480 11050 0 _0107_
rlabel metal1 27140 21114 27140 21114 0 _0108_
rlabel metal1 12834 24718 12834 24718 0 _0109_
rlabel via2 21942 25245 21942 25245 0 _0110_
rlabel metal1 16192 26962 16192 26962 0 _0111_
rlabel metal1 21758 25160 21758 25160 0 _0112_
rlabel metal1 25806 15334 25806 15334 0 _0113_
rlabel metal2 20930 23341 20930 23341 0 _0114_
rlabel metal1 14950 28526 14950 28526 0 _0115_
rlabel metal2 22034 15589 22034 15589 0 _0116_
rlabel metal1 25576 22066 25576 22066 0 _0117_
rlabel metal1 4784 23290 4784 23290 0 _0118_
rlabel metal1 5796 22634 5796 22634 0 _0119_
rlabel metal2 8234 21182 8234 21182 0 _0120_
rlabel metal1 3726 20026 3726 20026 0 _0121_
rlabel metal1 12558 18088 12558 18088 0 _0122_
rlabel metal1 17020 10574 17020 10574 0 _0123_
rlabel via3 5405 21420 5405 21420 0 _0124_
rlabel metal1 9522 21012 9522 21012 0 _0125_
rlabel via3 21643 21012 21643 21012 0 _0126_
rlabel metal1 18170 18122 18170 18122 0 _0127_
rlabel metal1 7820 17646 7820 17646 0 _0128_
rlabel metal3 14329 18564 14329 18564 0 _0129_
rlabel metal1 15778 16626 15778 16626 0 _0130_
rlabel metal2 15594 20740 15594 20740 0 _0131_
rlabel metal1 5198 15028 5198 15028 0 _0132_
rlabel metal1 20286 16456 20286 16456 0 _0133_
rlabel metal4 2300 15028 2300 15028 0 _0134_
rlabel metal1 10902 15504 10902 15504 0 _0135_
rlabel metal1 6026 13294 6026 13294 0 _0136_
rlabel metal1 9522 16524 9522 16524 0 _0137_
rlabel metal1 22126 7208 22126 7208 0 _0138_
rlabel metal1 9476 16966 9476 16966 0 _0139_
rlabel via2 24242 17187 24242 17187 0 _0140_
rlabel metal1 4508 22474 4508 22474 0 _0141_
rlabel metal1 4554 22134 4554 22134 0 _0142_
rlabel metal2 13294 17221 13294 17221 0 _0143_
rlabel metal1 4876 14994 4876 14994 0 _0144_
rlabel metal1 14536 17646 14536 17646 0 _0145_
rlabel metal1 7452 11254 7452 11254 0 _0146_
rlabel metal1 9844 10642 9844 10642 0 _0147_
rlabel metal1 18906 21590 18906 21590 0 _0148_
rlabel metal1 17342 8568 17342 8568 0 _0149_
rlabel metal1 19642 9452 19642 9452 0 _0150_
rlabel metal1 12098 22100 12098 22100 0 _0151_
rlabel metal2 21298 18887 21298 18887 0 _0152_
rlabel metal2 19642 22644 19642 22644 0 _0153_
rlabel metal2 13018 7684 13018 7684 0 _0154_
rlabel metal1 12926 10472 12926 10472 0 _0155_
rlabel metal1 8464 16762 8464 16762 0 _0156_
rlabel metal1 26864 10438 26864 10438 0 _0157_
rlabel metal1 28336 13498 28336 13498 0 _0158_
rlabel metal1 3772 21658 3772 21658 0 _0159_
rlabel metal1 4002 20468 4002 20468 0 _0160_
rlabel metal1 13248 13906 13248 13906 0 _0161_
rlabel metal1 7912 8330 7912 8330 0 _0162_
rlabel metal1 20378 7854 20378 7854 0 _0163_
rlabel metal2 14582 8704 14582 8704 0 _0164_
rlabel metal2 1150 9843 1150 9843 0 _0165_
rlabel metal1 15686 13906 15686 13906 0 _0166_
rlabel metal1 15916 14246 15916 14246 0 _0167_
rlabel metal1 21666 21012 21666 21012 0 _0168_
rlabel metal2 9890 14705 9890 14705 0 _0169_
rlabel metal2 14950 13872 14950 13872 0 _0170_
rlabel metal2 21482 13855 21482 13855 0 _0171_
rlabel metal2 21482 9163 21482 9163 0 _0172_
rlabel metal1 21965 14246 21965 14246 0 _0173_
rlabel metal1 25208 14382 25208 14382 0 _0174_
rlabel metal1 15870 6740 15870 6740 0 _0175_
rlabel metal2 8970 8772 8970 8772 0 _0176_
rlabel metal1 9890 7412 9890 7412 0 _0177_
rlabel via2 9154 22491 9154 22491 0 _0178_
rlabel metal2 25254 5916 25254 5916 0 _0179_
rlabel metal2 15778 7446 15778 7446 0 _0180_
rlabel metal1 26818 6426 26818 6426 0 _0181_
rlabel metal2 2714 20808 2714 20808 0 _0182_
rlabel metal3 16629 12716 16629 12716 0 _0183_
rlabel metal1 17618 6222 17618 6222 0 _0184_
rlabel via2 19458 12155 19458 12155 0 _0185_
rlabel metal1 24012 12818 24012 12818 0 _0186_
rlabel metal2 21758 13311 21758 13311 0 _0187_
rlabel via2 24794 12835 24794 12835 0 _0188_
rlabel metal2 19458 18836 19458 18836 0 _0189_
rlabel metal1 25990 12886 25990 12886 0 _0190_
rlabel metal1 28428 12818 28428 12818 0 _0191_
rlabel metal1 3956 12818 3956 12818 0 _0192_
rlabel metal3 17388 6528 17388 6528 0 _0193_
rlabel via2 22034 10659 22034 10659 0 _0194_
rlabel metal2 6946 10880 6946 10880 0 _0195_
rlabel metal1 8050 13192 8050 13192 0 _0196_
rlabel metal2 18446 16558 18446 16558 0 _0197_
rlabel via1 21114 13906 21114 13906 0 _0198_
rlabel metal3 18745 12716 18745 12716 0 _0199_
rlabel metal2 5290 14144 5290 14144 0 _0200_
rlabel metal2 10442 8806 10442 8806 0 _0201_
rlabel metal1 11178 6086 11178 6086 0 _0202_
rlabel metal1 4462 7208 4462 7208 0 _0203_
rlabel metal3 4439 6732 4439 6732 0 _0204_
rlabel metal2 20746 5100 20746 5100 0 _0205_
rlabel metal2 20746 15640 20746 15640 0 _0206_
rlabel metal1 27922 13362 27922 13362 0 _0207_
rlabel metal1 12374 20400 12374 20400 0 _0208_
rlabel metal1 9660 20434 9660 20434 0 _0209_
rlabel metal2 8372 22950 8372 22950 0 _0210_
rlabel metal1 5290 15538 5290 15538 0 _0211_
rlabel metal2 11914 14688 11914 14688 0 _0212_
rlabel metal1 15548 6698 15548 6698 0 _0213_
rlabel metal1 16514 23290 16514 23290 0 _0214_
rlabel metal1 12926 12648 12926 12648 0 _0215_
rlabel metal1 4830 23834 4830 23834 0 _0216_
rlabel via3 12949 21420 12949 21420 0 _0217_
rlabel metal2 20194 29019 20194 29019 0 _0218_
rlabel metal1 7544 19414 7544 19414 0 _0219_
rlabel metal1 17986 29104 17986 29104 0 _0220_
rlabel metal1 10212 16762 10212 16762 0 _0221_
rlabel metal2 20286 21369 20286 21369 0 _0222_
rlabel metal2 13018 27710 13018 27710 0 _0223_
rlabel metal1 19366 28050 19366 28050 0 _0224_
rlabel metal1 20424 23018 20424 23018 0 _0225_
rlabel metal3 7475 20740 7475 20740 0 _0226_
rlabel metal3 4531 16524 4531 16524 0 _0227_
rlabel metal2 16238 25398 16238 25398 0 _0228_
rlabel metal1 25944 26962 25944 26962 0 _0229_
rlabel metal1 14812 18938 14812 18938 0 _0230_
rlabel metal2 25622 27778 25622 27778 0 _0231_
rlabel metal1 15042 27540 15042 27540 0 _0232_
rlabel metal4 12972 15368 12972 15368 0 _0233_
rlabel metal2 11086 28441 11086 28441 0 _0234_
rlabel metal2 10258 27829 10258 27829 0 _0235_
rlabel metal1 27370 21012 27370 21012 0 _0236_
rlabel metal1 16238 26520 16238 26520 0 _0237_
rlabel viali 12834 8466 12834 8466 0 _0238_
rlabel metal2 21574 25976 21574 25976 0 _0239_
rlabel metal1 8694 25704 8694 25704 0 _0240_
rlabel metal2 15042 29291 15042 29291 0 _0241_
rlabel metal2 18538 7378 18538 7378 0 _0242_
rlabel metal1 25622 27472 25622 27472 0 _0243_
rlabel metal1 27784 15402 27784 15402 0 _0244_
rlabel metal1 11684 7854 11684 7854 0 _0245_
rlabel metal2 11362 8772 11362 8772 0 _0246_
rlabel metal1 15502 12750 15502 12750 0 _0247_
rlabel metal1 5658 11016 5658 11016 0 _0248_
rlabel metal1 4738 14348 4738 14348 0 _0249_
rlabel metal1 18814 21420 18814 21420 0 _0250_
rlabel metal2 7176 12988 7176 12988 0 _0251_
rlabel metal1 16698 11696 16698 11696 0 _0252_
rlabel metal2 17158 12002 17158 12002 0 _0253_
rlabel metal2 15134 9333 15134 9333 0 _0254_
rlabel metal1 8740 14382 8740 14382 0 _0255_
rlabel metal1 11178 6732 11178 6732 0 _0256_
rlabel metal1 6578 19686 6578 19686 0 _0257_
rlabel metal1 18630 13940 18630 13940 0 _0258_
rlabel metal2 20378 5950 20378 5950 0 _0259_
rlabel metal2 3910 15521 3910 15521 0 _0260_
rlabel metal1 7912 21658 7912 21658 0 _0261_
rlabel metal1 20516 15878 20516 15878 0 _0262_
rlabel metal1 15042 12206 15042 12206 0 _0263_
rlabel via2 6946 10149 6946 10149 0 _0264_
rlabel metal2 3266 13634 3266 13634 0 _0265_
rlabel metal1 14536 13498 14536 13498 0 _0266_
rlabel metal2 18354 16796 18354 16796 0 _0267_
rlabel metal1 25208 16490 25208 16490 0 _0268_
rlabel metal2 28106 16864 28106 16864 0 _0269_
rlabel metal1 28612 17510 28612 17510 0 _0270_
rlabel metal1 11730 21114 11730 21114 0 _0271_
rlabel metal2 14674 18105 14674 18105 0 _0272_
rlabel metal1 28566 16558 28566 16558 0 _0273_
rlabel metal1 28704 13498 28704 13498 0 _0274_
rlabel metal2 27462 13260 27462 13260 0 _0275_
rlabel metal1 28658 13430 28658 13430 0 _0276_
rlabel metal1 26910 12614 26910 12614 0 _0277_
rlabel metal2 17250 12189 17250 12189 0 _0278_
rlabel metal1 27140 12410 27140 12410 0 _0279_
rlabel metal1 28290 12954 28290 12954 0 _0280_
rlabel metal1 29854 13498 29854 13498 0 _0281_
rlabel metal1 10672 14518 10672 14518 0 _0282_
rlabel metal1 14582 8908 14582 8908 0 _0283_
rlabel metal2 17618 25534 17618 25534 0 _0284_
rlabel metal1 17848 23766 17848 23766 0 _0285_
rlabel metal3 18377 22644 18377 22644 0 _0286_
rlabel metal2 13386 10540 13386 10540 0 _0287_
rlabel metal1 13248 8262 13248 8262 0 _0288_
rlabel metal1 14306 27846 14306 27846 0 _0289_
rlabel metal2 24794 7650 24794 7650 0 _0290_
rlabel metal2 13754 6885 13754 6885 0 _0291_
rlabel metal1 14030 11322 14030 11322 0 _0292_
rlabel metal2 13202 14450 13202 14450 0 _0293_
rlabel metal1 13570 9520 13570 9520 0 _0294_
rlabel metal2 18538 10047 18538 10047 0 _0295_
rlabel metal1 13478 25364 13478 25364 0 _0296_
rlabel metal1 13294 22746 13294 22746 0 _0297_
rlabel metal3 15732 13668 15732 13668 0 _0298_
rlabel metal1 14214 8602 14214 8602 0 _0299_
rlabel metal2 14122 9146 14122 9146 0 _0300_
rlabel metal1 18446 8976 18446 8976 0 _0301_
rlabel metal2 18262 6154 18262 6154 0 _0302_
rlabel via2 16790 15691 16790 15691 0 _0303_
rlabel metal2 25898 19040 25898 19040 0 _0304_
rlabel metal1 17848 5746 17848 5746 0 _0305_
rlabel metal2 31786 9129 31786 9129 0 _0306_
rlabel via2 18814 14875 18814 14875 0 _0307_
rlabel metal2 26818 17986 26818 17986 0 _0308_
rlabel metal2 16790 14671 16790 14671 0 _0309_
rlabel metal2 14674 21029 14674 21029 0 _0310_
rlabel metal2 24748 14382 24748 14382 0 _0311_
rlabel metal4 22172 18836 22172 18836 0 _0312_
rlabel metal1 19458 26962 19458 26962 0 _0313_
rlabel metal1 17296 24582 17296 24582 0 _0314_
rlabel metal1 29026 16728 29026 16728 0 _0315_
rlabel metal1 29072 19346 29072 19346 0 _0316_
rlabel metal2 18998 18870 18998 18870 0 _0317_
rlabel metal1 30360 13906 30360 13906 0 _0318_
rlabel metal2 29394 19652 29394 19652 0 _0319_
rlabel metal1 30314 19924 30314 19924 0 _0320_
rlabel metal1 24932 14586 24932 14586 0 _0321_
rlabel metal1 19550 18700 19550 18700 0 _0322_
rlabel metal1 23368 19346 23368 19346 0 _0323_
rlabel metal2 23138 21726 23138 21726 0 _0324_
rlabel metal2 24426 20230 24426 20230 0 _0325_
rlabel metal1 24610 19414 24610 19414 0 _0326_
rlabel metal2 18906 16014 18906 16014 0 _0327_
rlabel metal1 25714 19482 25714 19482 0 _0328_
rlabel metal1 26312 19346 26312 19346 0 _0329_
rlabel metal2 26082 17238 26082 17238 0 _0330_
rlabel metal1 27416 19482 27416 19482 0 _0331_
rlabel metal1 29992 23698 29992 23698 0 _0332_
rlabel metal2 20746 12784 20746 12784 0 _0333_
rlabel metal2 16790 25483 16790 25483 0 _0334_
rlabel metal2 14490 22236 14490 22236 0 _0335_
rlabel metal1 22494 14994 22494 14994 0 _0336_
rlabel metal1 15962 20536 15962 20536 0 _0337_
rlabel metal1 20010 25908 20010 25908 0 _0338_
rlabel metal2 13662 6851 13662 6851 0 _0339_
rlabel metal1 7636 18394 7636 18394 0 _0340_
rlabel metal1 10350 21522 10350 21522 0 _0341_
rlabel metal2 10258 21046 10258 21046 0 _0342_
rlabel metal1 10166 21420 10166 21420 0 _0343_
rlabel metal1 9062 21556 9062 21556 0 _0344_
rlabel metal2 16698 25092 16698 25092 0 _0345_
rlabel metal1 9016 9146 9016 9146 0 _0346_
rlabel metal1 16928 25466 16928 25466 0 _0347_
rlabel metal2 9522 20060 9522 20060 0 _0348_
rlabel metal2 1334 12036 1334 12036 0 _0349_
rlabel metal1 9338 18836 9338 18836 0 _0350_
rlabel metal1 9200 10234 9200 10234 0 _0351_
rlabel metal2 16422 25024 16422 25024 0 _0352_
rlabel metal1 17848 29614 17848 29614 0 _0353_
rlabel metal1 18078 11594 18078 11594 0 _0354_
rlabel metal1 18492 11730 18492 11730 0 _0355_
rlabel metal1 20976 19822 20976 19822 0 _0356_
rlabel metal1 27876 7378 27876 7378 0 _0357_
rlabel metal1 18906 18326 18906 18326 0 _0358_
rlabel metal2 27922 18207 27922 18207 0 _0359_
rlabel metal1 28658 18394 28658 18394 0 _0360_
rlabel metal1 27784 23290 27784 23290 0 _0361_
rlabel metal2 16514 9826 16514 9826 0 _0362_
rlabel metal2 32706 22627 32706 22627 0 _0363_
rlabel metal1 28658 23154 28658 23154 0 _0364_
rlabel metal1 29762 22984 29762 22984 0 _0365_
rlabel metal2 18538 23324 18538 23324 0 _0366_
rlabel metal1 18446 23154 18446 23154 0 _0367_
rlabel metal2 18906 22797 18906 22797 0 _0368_
rlabel metal1 29808 22610 29808 22610 0 _0369_
rlabel metal1 20700 25466 20700 25466 0 _0370_
rlabel metal3 26657 18020 26657 18020 0 _0371_
rlabel metal1 13248 16762 13248 16762 0 _0372_
rlabel metal2 25806 23392 25806 23392 0 _0373_
rlabel metal1 17894 17510 17894 17510 0 _0374_
rlabel metal1 26634 20026 26634 20026 0 _0375_
rlabel metal1 19964 20366 19964 20366 0 _0376_
rlabel metal4 20884 11956 20884 11956 0 _0377_
rlabel metal1 20884 21522 20884 21522 0 _0378_
rlabel metal1 27094 19720 27094 19720 0 _0379_
rlabel metal1 19780 21658 19780 21658 0 _0380_
rlabel metal2 20746 21760 20746 21760 0 _0381_
rlabel via2 19366 21675 19366 21675 0 _0382_
rlabel metal2 23506 21216 23506 21216 0 _0383_
rlabel metal2 13846 21913 13846 21913 0 _0384_
rlabel metal1 26128 23290 26128 23290 0 _0385_
rlabel metal1 15134 17816 15134 17816 0 _0386_
rlabel metal1 14904 17646 14904 17646 0 _0387_
rlabel metal1 15456 17510 15456 17510 0 _0388_
rlabel metal1 21896 18938 21896 18938 0 _0389_
rlabel metal2 22494 15776 22494 15776 0 _0390_
rlabel metal2 22218 15759 22218 15759 0 _0391_
rlabel metal1 22448 15402 22448 15402 0 _0392_
rlabel metal1 21896 15674 21896 15674 0 _0393_
rlabel metal1 21758 17646 21758 17646 0 _0394_
rlabel metal1 19274 25364 19274 25364 0 _0395_
rlabel metal1 20102 25670 20102 25670 0 _0396_
rlabel metal2 20746 24990 20746 24990 0 _0397_
rlabel metal2 7314 14178 7314 14178 0 _0398_
rlabel metal1 8096 14586 8096 14586 0 _0399_
rlabel metal1 8648 14790 8648 14790 0 _0400_
rlabel metal1 6670 15504 6670 15504 0 _0401_
rlabel metal2 8418 15164 8418 15164 0 _0402_
rlabel metal1 9338 14008 9338 14008 0 _0403_
rlabel metal4 1012 23188 1012 23188 0 _0404_
rlabel metal1 21206 24650 21206 24650 0 _0405_
rlabel metal2 23966 27370 23966 27370 0 _0406_
rlabel metal1 27324 15470 27324 15470 0 _0407_
rlabel metal1 6578 12954 6578 12954 0 _0408_
rlabel metal2 9430 9877 9430 9877 0 _0409_
rlabel metal2 11270 9945 11270 9945 0 _0410_
rlabel metal1 20010 8602 20010 8602 0 _0411_
rlabel metal1 20332 8398 20332 8398 0 _0412_
rlabel metal2 20930 9044 20930 9044 0 _0413_
rlabel via2 16330 10421 16330 10421 0 _0414_
rlabel metal1 22264 8942 22264 8942 0 _0415_
rlabel via2 19918 25891 19918 25891 0 _0416_
rlabel metal1 26174 11118 26174 11118 0 _0417_
rlabel metal1 23368 11118 23368 11118 0 _0418_
rlabel metal1 25806 9350 25806 9350 0 _0419_
rlabel metal1 24150 8262 24150 8262 0 _0420_
rlabel metal1 24334 8364 24334 8364 0 _0421_
rlabel metal1 24242 8568 24242 8568 0 _0422_
rlabel metal2 24702 9044 24702 9044 0 _0423_
rlabel metal1 26312 9622 26312 9622 0 _0424_
rlabel metal2 24518 7310 24518 7310 0 _0425_
rlabel metal2 21758 19023 21758 19023 0 _0426_
rlabel metal1 17342 18598 17342 18598 0 _0427_
rlabel metal1 16882 18938 16882 18938 0 _0428_
rlabel metal1 11178 22406 11178 22406 0 _0429_
rlabel metal1 21068 18666 21068 18666 0 _0430_
rlabel metal2 20746 18989 20746 18989 0 _0431_
rlabel metal1 18768 7990 18768 7990 0 _0432_
rlabel metal2 2484 13906 2484 13906 0 _0433_
rlabel metal1 21942 18734 21942 18734 0 _0434_
rlabel metal2 18722 18496 18722 18496 0 _0435_
rlabel metal1 16468 22406 16468 22406 0 _0436_
rlabel metal3 19067 18020 19067 18020 0 _0437_
rlabel metal1 22126 18904 22126 18904 0 _0438_
rlabel metal1 22034 18666 22034 18666 0 _0439_
rlabel via2 22494 18955 22494 18955 0 _0440_
rlabel metal1 9890 14042 9890 14042 0 _0441_
rlabel metal1 9936 14586 9936 14586 0 _0442_
rlabel metal1 10074 14484 10074 14484 0 _0443_
rlabel metal1 9614 11866 9614 11866 0 _0444_
rlabel metal2 10442 14297 10442 14297 0 _0445_
rlabel metal1 29670 21522 29670 21522 0 _0446_
rlabel metal1 23782 14790 23782 14790 0 _0447_
rlabel metal1 22862 18666 22862 18666 0 _0448_
rlabel metal1 23000 15402 23000 15402 0 _0449_
rlabel metal1 23414 14926 23414 14926 0 _0450_
rlabel metal1 28198 14586 28198 14586 0 _0451_
rlabel via2 12650 4709 12650 4709 0 _0452_
rlabel metal1 22632 7854 22632 7854 0 _0453_
rlabel via2 23874 21301 23874 21301 0 _0454_
rlabel metal1 23828 15130 23828 15130 0 _0455_
rlabel metal1 23966 29104 23966 29104 0 _0456_
rlabel via2 3634 12835 3634 12835 0 _0457_
rlabel metal1 21344 12138 21344 12138 0 _0458_
rlabel metal1 26358 21046 26358 21046 0 _0459_
rlabel metal2 29854 15776 29854 15776 0 _0460_
rlabel metal1 29716 16082 29716 16082 0 _0461_
rlabel metal1 3128 12682 3128 12682 0 _0462_
rlabel metal1 15778 19346 15778 19346 0 _0463_
rlabel metal2 15226 15759 15226 15759 0 _0464_
rlabel via1 15781 19414 15781 19414 0 _0465_
rlabel metal2 16238 20043 16238 20043 0 _0466_
rlabel metal2 30038 20502 30038 20502 0 _0467_
rlabel metal2 30222 17510 30222 17510 0 _0468_
rlabel metal1 30590 20570 30590 20570 0 _0469_
rlabel via3 28221 23460 28221 23460 0 _0470_
rlabel metal1 29164 24650 29164 24650 0 _0471_
rlabel metal1 21390 20434 21390 20434 0 _0472_
rlabel metal2 28244 12750 28244 12750 0 _0473_
rlabel metal1 26864 21386 26864 21386 0 _0474_
rlabel metal1 29394 21658 29394 21658 0 _0475_
rlabel metal1 12650 21386 12650 21386 0 _0476_
rlabel metal3 13938 15028 13938 15028 0 _0477_
rlabel via2 19642 22083 19642 22083 0 _0478_
rlabel metal1 23690 25908 23690 25908 0 _0479_
rlabel metal2 23690 27081 23690 27081 0 _0480_
rlabel metal1 23552 25874 23552 25874 0 _0481_
rlabel metal1 29532 25262 29532 25262 0 _0482_
rlabel metal1 29808 25466 29808 25466 0 _0483_
rlabel metal2 16054 16864 16054 16864 0 _0484_
rlabel metal3 15479 16796 15479 16796 0 _0485_
rlabel metal1 16422 20230 16422 20230 0 _0486_
rlabel metal2 15686 20060 15686 20060 0 _0487_
rlabel metal1 9338 6630 9338 6630 0 _0488_
rlabel metal2 10258 19142 10258 19142 0 _0489_
rlabel metal1 12466 19142 12466 19142 0 _0490_
rlabel metal2 12098 19074 12098 19074 0 _0491_
rlabel metal1 12006 19448 12006 19448 0 _0492_
rlabel metal1 12788 19210 12788 19210 0 _0493_
rlabel metal2 16514 20230 16514 20230 0 _0494_
rlabel via2 17158 20315 17158 20315 0 _0495_
rlabel metal1 11362 20434 11362 20434 0 _0496_
rlabel metal1 21620 6222 21620 6222 0 _0497_
rlabel metal1 22770 10234 22770 10234 0 _0498_
rlabel metal1 22402 9996 22402 9996 0 _0499_
rlabel metal2 22586 10268 22586 10268 0 _0500_
rlabel metal1 12374 17068 12374 17068 0 _0501_
rlabel metal1 20562 13906 20562 13906 0 _0502_
rlabel metal2 22218 9860 22218 9860 0 _0503_
rlabel metal1 22908 6426 22908 6426 0 _0504_
rlabel metal1 22218 9384 22218 9384 0 _0505_
rlabel metal1 12236 17238 12236 17238 0 _0506_
rlabel metal3 13225 14756 13225 14756 0 _0507_
rlabel metal1 22356 7990 22356 7990 0 _0508_
rlabel metal2 21942 9350 21942 9350 0 _0509_
rlabel metal1 22264 4590 22264 4590 0 _0510_
rlabel metal1 27462 14042 27462 14042 0 _0511_
rlabel metal2 24150 7293 24150 7293 0 _0512_
rlabel metal4 21804 15232 21804 15232 0 _0513_
rlabel metal1 20470 9044 20470 9044 0 _0514_
rlabel metal1 24196 20366 24196 20366 0 _0515_
rlabel metal2 22954 10489 22954 10489 0 _0516_
rlabel metal2 25990 8636 25990 8636 0 _0517_
rlabel metal2 20562 6681 20562 6681 0 _0518_
rlabel metal1 13248 6766 13248 6766 0 _0519_
rlabel metal2 26082 7446 26082 7446 0 _0520_
rlabel metal1 24150 7310 24150 7310 0 _0521_
rlabel metal1 13892 6902 13892 6902 0 _0522_
rlabel metal1 25898 7412 25898 7412 0 _0523_
rlabel metal1 26956 7514 26956 7514 0 _0524_
rlabel metal3 22839 19380 22839 19380 0 _0525_
rlabel metal2 24518 20060 24518 20060 0 _0526_
rlabel metal1 10166 17000 10166 17000 0 _0527_
rlabel metal2 8418 16762 8418 16762 0 _0528_
rlabel metal2 8050 17034 8050 17034 0 _0529_
rlabel metal1 10810 15130 10810 15130 0 _0530_
rlabel metal1 10350 16218 10350 16218 0 _0531_
rlabel metal1 10856 17306 10856 17306 0 _0532_
rlabel metal1 21114 15878 21114 15878 0 _0533_
rlabel metal1 23506 18734 23506 18734 0 _0534_
rlabel metal2 24150 19380 24150 19380 0 _0535_
rlabel via2 24794 20043 24794 20043 0 _0536_
rlabel metal2 13018 16949 13018 16949 0 _0537_
rlabel metal2 15226 26996 15226 26996 0 _0538_
rlabel metal2 14950 27234 14950 27234 0 _0539_
rlabel metal1 16054 27540 16054 27540 0 _0540_
rlabel metal1 15594 16660 15594 16660 0 _0541_
rlabel metal1 15456 12954 15456 12954 0 _0542_
rlabel metal2 15962 16473 15962 16473 0 _0543_
rlabel metal1 24058 27404 24058 27404 0 _0544_
rlabel metal1 23966 25126 23966 25126 0 _0545_
rlabel metal1 22770 27642 22770 27642 0 _0546_
rlabel metal2 16330 28356 16330 28356 0 _0547_
rlabel via2 26542 17765 26542 17765 0 _0548_
rlabel metal1 18952 5610 18952 5610 0 _0549_
rlabel metal1 22448 6426 22448 6426 0 _0550_
rlabel metal2 14490 17884 14490 17884 0 _0551_
rlabel metal1 14306 17578 14306 17578 0 _0552_
rlabel metal2 14858 17697 14858 17697 0 _0553_
rlabel metal1 21022 10608 21022 10608 0 _0554_
rlabel metal2 20562 11356 20562 11356 0 _0555_
rlabel metal1 26220 10506 26220 10506 0 _0556_
rlabel metal2 22494 9010 22494 9010 0 _0557_
rlabel metal1 22310 7276 22310 7276 0 _0558_
rlabel via1 9157 12206 9157 12206 0 _0559_
rlabel metal2 18814 7667 18814 7667 0 _0560_
rlabel metal1 22356 6698 22356 6698 0 _0561_
rlabel metal2 23598 5916 23598 5916 0 _0562_
rlabel metal2 7498 10914 7498 10914 0 _0563_
rlabel metal2 25622 11118 25622 11118 0 _0564_
rlabel metal1 29256 15470 29256 15470 0 _0565_
rlabel metal2 28474 11798 28474 11798 0 _0566_
rlabel via3 28635 12036 28635 12036 0 _0567_
rlabel metal2 28106 11526 28106 11526 0 _0568_
rlabel metal2 29118 10234 29118 10234 0 _0569_
rlabel metal1 14766 6426 14766 6426 0 _0570_
rlabel metal1 8050 11220 8050 11220 0 _0571_
rlabel metal1 15364 8058 15364 8058 0 _0572_
rlabel metal1 14950 8568 14950 8568 0 _0573_
rlabel via2 15410 8347 15410 8347 0 _0574_
rlabel metal2 29302 9350 29302 9350 0 _0575_
rlabel metal1 29946 13872 29946 13872 0 _0576_
rlabel metal2 20930 10761 20930 10761 0 _0577_
rlabel metal1 19320 10642 19320 10642 0 _0578_
rlabel metal1 29946 13736 29946 13736 0 _0579_
rlabel metal2 29854 14076 29854 14076 0 _0580_
rlabel metal1 18814 24786 18814 24786 0 _0581_
rlabel metal2 19274 10149 19274 10149 0 _0582_
rlabel metal1 18906 5882 18906 5882 0 _0583_
rlabel metal1 17710 10710 17710 10710 0 _0584_
rlabel metal1 18998 10744 18998 10744 0 _0585_
rlabel metal1 29394 13838 29394 13838 0 _0586_
rlabel metal2 30958 13668 30958 13668 0 _0587_
rlabel metal1 22678 10472 22678 10472 0 _0588_
rlabel metal1 17526 11526 17526 11526 0 _0589_
rlabel metal2 17342 27166 17342 27166 0 _0590_
rlabel metal3 17825 15028 17825 15028 0 _0591_
rlabel metal1 18538 13498 18538 13498 0 _0592_
rlabel metal1 18262 11798 18262 11798 0 _0593_
rlabel metal1 20562 11084 20562 11084 0 _0594_
rlabel metal1 19826 7752 19826 7752 0 _0595_
rlabel metal1 22264 10642 22264 10642 0 _0596_
rlabel metal1 23598 10778 23598 10778 0 _0597_
rlabel metal1 11270 12138 11270 12138 0 _0598_
rlabel metal2 12190 11798 12190 11798 0 _0599_
rlabel metal1 11270 11322 11270 11322 0 _0600_
rlabel metal1 12236 11730 12236 11730 0 _0601_
rlabel metal1 21068 11118 21068 11118 0 _0602_
rlabel metal1 20194 11050 20194 11050 0 _0603_
rlabel metal1 20930 11220 20930 11220 0 _0604_
rlabel metal1 25392 21862 25392 21862 0 _0605_
rlabel metal2 22034 22576 22034 22576 0 _0606_
rlabel metal2 22218 21556 22218 21556 0 _0607_
rlabel metal1 22356 21998 22356 21998 0 _0608_
rlabel metal1 21666 21862 21666 21862 0 _0609_
rlabel metal1 20930 11322 20930 11322 0 _0610_
rlabel metal1 24196 5882 24196 5882 0 _0611_
rlabel metal1 22954 12818 22954 12818 0 _0612_
rlabel metal1 24150 12274 24150 12274 0 _0613_
rlabel metal1 23966 12138 23966 12138 0 _0614_
rlabel metal2 26818 11424 26818 11424 0 _0615_
rlabel metal1 24702 10744 24702 10744 0 _0616_
rlabel metal1 25530 10744 25530 10744 0 _0617_
rlabel metal1 26404 10778 26404 10778 0 _0618_
rlabel metal1 30222 10098 30222 10098 0 _0619_
rlabel metal1 17204 14450 17204 14450 0 _0620_
rlabel metal1 16790 14314 16790 14314 0 _0621_
rlabel metal2 17710 11356 17710 11356 0 _0622_
rlabel metal2 17526 7174 17526 7174 0 _0623_
rlabel metal2 16330 6290 16330 6290 0 _0624_
rlabel metal2 17158 8262 17158 8262 0 _0625_
rlabel metal1 24058 8398 24058 8398 0 _0626_
rlabel metal2 20976 16252 20976 16252 0 _0627_
rlabel metal2 29946 9078 29946 9078 0 _0628_
rlabel metal1 31050 12954 31050 12954 0 _0629_
rlabel metal1 29118 12206 29118 12206 0 _0630_
rlabel metal1 29854 11560 29854 11560 0 _0631_
rlabel metal2 32062 19720 32062 19720 0 _0632_
rlabel metal1 26220 11662 26220 11662 0 _0633_
rlabel metal1 29486 11798 29486 11798 0 _0634_
rlabel metal1 29900 8466 29900 8466 0 _0635_
rlabel metal1 30314 6766 30314 6766 0 _0636_
rlabel metal2 21114 16932 21114 16932 0 _0637_
rlabel metal2 20746 20128 20746 20128 0 _0638_
rlabel metal2 6578 24378 6578 24378 0 _0639_
rlabel metal1 20930 20332 20930 20332 0 _0640_
rlabel metal1 5428 14518 5428 14518 0 _0641_
rlabel metal1 6210 14484 6210 14484 0 _0642_
rlabel metal2 6072 14042 6072 14042 0 _0643_
rlabel metal2 17802 19958 17802 19958 0 _0644_
rlabel metal1 18262 20366 18262 20366 0 _0645_
rlabel metal1 15456 20026 15456 20026 0 _0646_
rlabel metal1 20838 20536 20838 20536 0 _0647_
rlabel metal1 26358 20536 26358 20536 0 _0648_
rlabel metal1 5520 23698 5520 23698 0 _0649_
rlabel metal2 12190 16864 12190 16864 0 _0650_
rlabel metal1 12512 14042 12512 14042 0 _0651_
rlabel metal1 12926 16218 12926 16218 0 _0652_
rlabel metal2 15732 15674 15732 15674 0 _0653_
rlabel metal1 14444 11186 14444 11186 0 _0654_
rlabel metal1 13984 24786 13984 24786 0 _0655_
rlabel metal3 14559 11764 14559 11764 0 _0656_
rlabel metal1 15134 11322 15134 11322 0 _0657_
rlabel metal1 15318 11152 15318 11152 0 _0658_
rlabel metal2 15686 9469 15686 9469 0 _0659_
rlabel metal1 6509 24786 6509 24786 0 _0660_
rlabel metal1 30314 15572 30314 15572 0 _0661_
rlabel metal1 19320 16082 19320 16082 0 _0662_
rlabel metal1 19964 15878 19964 15878 0 _0663_
rlabel metal1 3910 14382 3910 14382 0 _0664_
rlabel metal1 19780 16150 19780 16150 0 _0665_
rlabel metal2 20010 16286 20010 16286 0 _0666_
rlabel metal1 23414 16184 23414 16184 0 _0667_
rlabel metal1 27784 21454 27784 21454 0 _0668_
rlabel metal2 27094 15062 27094 15062 0 _0669_
rlabel metal1 6486 23698 6486 23698 0 _0670_
rlabel metal1 17250 12682 17250 12682 0 _0671_
rlabel metal1 30130 15470 30130 15470 0 _0672_
rlabel metal2 30590 15810 30590 15810 0 _0673_
rlabel metal1 25714 26860 25714 26860 0 _0674_
rlabel metal1 26128 26554 26128 26554 0 _0675_
rlabel metal2 26082 25228 26082 25228 0 _0676_
rlabel metal1 28106 21624 28106 21624 0 _0677_
rlabel metal1 27554 17850 27554 17850 0 _0678_
rlabel metal2 27830 22950 27830 22950 0 _0679_
rlabel metal1 19734 23052 19734 23052 0 _0680_
rlabel metal2 27646 22134 27646 22134 0 _0681_
rlabel metal1 30866 21998 30866 21998 0 _0682_
rlabel metal1 28244 15334 28244 15334 0 _0683_
rlabel metal1 25760 16762 25760 16762 0 _0684_
rlabel metal1 25622 17272 25622 17272 0 _0685_
rlabel metal1 28198 17000 28198 17000 0 _0686_
rlabel metal1 27784 16626 27784 16626 0 _0687_
rlabel metal1 28198 17272 28198 17272 0 _0688_
rlabel metal1 29808 17306 29808 17306 0 _0689_
rlabel metal1 5290 27846 5290 27846 0 _0690_
rlabel metal1 27324 16558 27324 16558 0 _0691_
rlabel metal1 28474 16762 28474 16762 0 _0692_
rlabel metal1 30682 16558 30682 16558 0 _0693_
rlabel metal1 29808 12614 29808 12614 0 _0694_
rlabel metal1 5704 21998 5704 21998 0 _0695_
rlabel metal1 17572 20570 17572 20570 0 _0696_
rlabel via1 15326 19346 15326 19346 0 _0697_
rlabel metal2 4094 25228 4094 25228 0 _0698_
rlabel metal2 3542 25840 3542 25840 0 _0699_
rlabel metal2 14490 24905 14490 24905 0 _0700_
rlabel metal1 3818 26214 3818 26214 0 _0701_
rlabel metal1 6532 28458 6532 28458 0 _0702_
rlabel metal1 7682 24582 7682 24582 0 _0703_
rlabel metal2 31786 6289 31786 6289 0 _0704_
rlabel metal1 4370 25738 4370 25738 0 _0705_
rlabel via2 2622 26877 2622 26877 0 _0706_
rlabel metal1 5934 16150 5934 16150 0 _0707_
rlabel metal2 21022 17306 21022 17306 0 _0708_
rlabel metal1 3634 27574 3634 27574 0 _0709_
rlabel metal2 2254 28322 2254 28322 0 _0710_
rlabel metal1 10166 23630 10166 23630 0 _0711_
rlabel metal1 7682 29478 7682 29478 0 _0712_
rlabel metal1 8096 29682 8096 29682 0 _0713_
rlabel metal3 12420 18224 12420 18224 0 _0714_
rlabel metal1 5934 27982 5934 27982 0 _0715_
rlabel metal3 751 25908 751 25908 0 addr0[0]
rlabel metal3 1050 28628 1050 28628 0 addr0[1]
rlabel metal3 1096 27948 1096 27948 0 addr0[2]
rlabel metal3 751 23868 751 23868 0 addr0[3]
rlabel metal3 751 14348 751 14348 0 addr0[4]
rlabel metal3 1004 19108 1004 19108 0 addr0[5]
rlabel metal3 1050 10948 1050 10948 0 addr0[6]
rlabel metal3 751 16388 751 16388 0 addr0[7]
rlabel metal1 3312 26554 3312 26554 0 addr0_reg\[0\]
rlabel metal1 3726 28662 3726 28662 0 addr0_reg\[1\]
rlabel metal1 3036 28186 3036 28186 0 addr0_reg\[2\]
rlabel metal1 3358 25466 3358 25466 0 addr0_reg\[3\]
rlabel metal2 2070 21828 2070 21828 0 addr0_reg\[4\]
rlabel metal1 4002 19856 4002 19856 0 addr0_reg\[5\]
rlabel metal2 2070 19924 2070 19924 0 addr0_reg\[6\]
rlabel metal2 2346 22916 2346 22916 0 addr0_reg\[7\]
rlabel metal1 17342 17238 17342 17238 0 clk0
rlabel metal1 18032 17306 18032 17306 0 clknet_0_clk0
rlabel via2 1426 21539 1426 21539 0 clknet_2_0__leaf_clk0
rlabel metal1 18630 3978 18630 3978 0 clknet_2_1__leaf_clk0
rlabel metal1 31970 12852 31970 12852 0 clknet_2_2__leaf_clk0
rlabel metal1 30912 18802 30912 18802 0 clknet_2_3__leaf_clk0
rlabel metal2 32522 12903 32522 12903 0 cs0
rlabel metal2 30314 13056 30314 13056 0 cs0_reg
rlabel metal2 19366 1520 19366 1520 0 dout0[0]
rlabel metal1 32476 24582 32476 24582 0 dout0[10]
rlabel metal2 32430 20893 32430 20893 0 dout0[11]
rlabel metal2 22586 1520 22586 1520 0 dout0[12]
rlabel metal2 32430 8279 32430 8279 0 dout0[13]
rlabel metal2 31694 26333 31694 26333 0 dout0[14]
rlabel metal1 16836 31382 16836 31382 0 dout0[15]
rlabel metal2 25806 1520 25806 1520 0 dout0[16]
rlabel metal2 32430 10353 32430 10353 0 dout0[17]
rlabel metal2 32430 15079 32430 15079 0 dout0[18]
rlabel metal2 32430 13855 32430 13855 0 dout0[19]
rlabel metal1 32108 25670 32108 25670 0 dout0[1]
rlabel metal2 21298 1520 21298 1520 0 dout0[20]
rlabel metal2 32338 9503 32338 9503 0 dout0[21]
rlabel metal3 32852 6868 32852 6868 0 dout0[22]
rlabel metal2 32430 17901 32430 17901 0 dout0[23]
rlabel metal2 31694 6987 31694 6987 0 dout0[24]
rlabel metal2 32430 15793 32430 15793 0 dout0[25]
rlabel metal2 32430 23001 32430 23001 0 dout0[26]
rlabel metal2 32430 19295 32430 19295 0 dout0[27]
rlabel via2 32430 17051 32430 17051 0 dout0[28]
rlabel via2 32430 11611 32430 11611 0 dout0[29]
rlabel metal1 19090 31450 19090 31450 0 dout0[2]
rlabel metal2 17434 1520 17434 1520 0 dout0[30]
rlabel metal2 32430 20009 32430 20009 0 dout0[3]
rlabel metal2 30866 24837 30866 24837 0 dout0[4]
rlabel metal2 21298 32344 21298 32344 0 dout0[5]
rlabel metal2 24518 1520 24518 1520 0 dout0[6]
rlabel metal1 23276 31382 23276 31382 0 dout0[7]
rlabel metal1 25300 31450 25300 31450 0 dout0[8]
rlabel metal1 32476 22406 32476 22406 0 dout0[9]
rlabel metal1 1656 26010 1656 26010 0 net1
rlabel metal1 19780 4590 19780 4590 0 net10
rlabel metal2 15686 14212 15686 14212 0 net100
rlabel metal2 22310 27234 22310 27234 0 net101
rlabel metal2 32292 17612 32292 17612 0 net102
rlabel via2 20286 6851 20286 6851 0 net103
rlabel metal2 14582 27914 14582 27914 0 net104
rlabel metal2 22126 6460 22126 6460 0 net105
rlabel metal2 22448 25908 22448 25908 0 net106
rlabel metal1 16882 27370 16882 27370 0 net107
rlabel metal1 22448 26486 22448 26486 0 net108
rlabel metal2 21712 16796 21712 16796 0 net109
rlabel metal2 32246 25262 32246 25262 0 net11
rlabel metal1 1242 21318 1242 21318 0 net110
rlabel metal1 23230 18938 23230 18938 0 net111
rlabel metal2 12558 6562 12558 6562 0 net112
rlabel metal1 22356 25874 22356 25874 0 net113
rlabel metal2 12650 7361 12650 7361 0 net114
rlabel metal1 15594 27302 15594 27302 0 net115
rlabel metal1 18446 29002 18446 29002 0 net116
rlabel metal1 7774 19346 7774 19346 0 net117
rlabel metal2 17342 28594 17342 28594 0 net118
rlabel metal2 23782 28288 23782 28288 0 net119
rlabel metal1 32246 20366 32246 20366 0 net12
rlabel metal1 17434 29274 17434 29274 0 net120
rlabel metal4 644 24208 644 24208 0 net121
rlabel metal1 19642 23494 19642 23494 0 net122
rlabel metal1 20792 13498 20792 13498 0 net123
rlabel metal1 20378 19346 20378 19346 0 net124
rlabel metal1 18124 28390 18124 28390 0 net125
rlabel metal2 18446 28798 18446 28798 0 net126
rlabel via2 18170 29019 18170 29019 0 net127
rlabel metal1 20056 28594 20056 28594 0 net128
rlabel metal2 17802 27676 17802 27676 0 net129
rlabel metal1 23276 2414 23276 2414 0 net13
rlabel metal2 920 23732 920 23732 0 net130
rlabel metal1 21160 9554 21160 9554 0 net131
rlabel metal1 19872 27846 19872 27846 0 net132
rlabel metal1 20194 15368 20194 15368 0 net133
rlabel metal2 12834 21403 12834 21403 0 net134
rlabel metal1 18998 20230 18998 20230 0 net135
rlabel metal2 16192 19380 16192 19380 0 net136
rlabel metal1 16284 23290 16284 23290 0 net137
rlabel metal3 13984 6868 13984 6868 0 net138
rlabel metal4 14444 17272 14444 17272 0 net139
rlabel metal2 32246 8262 32246 8262 0 net14
rlabel metal1 6486 12852 6486 12852 0 net140
rlabel metal1 10304 17102 10304 17102 0 net141
rlabel metal2 19458 9843 19458 9843 0 net142
rlabel metal2 18170 24582 18170 24582 0 net143
rlabel metal1 11086 6664 11086 6664 0 net144
rlabel metal1 5336 15130 5336 15130 0 net145
rlabel metal1 10166 4624 10166 4624 0 net146
rlabel metal1 6026 12614 6026 12614 0 net147
rlabel metal1 10672 7174 10672 7174 0 net148
rlabel metal2 12742 10421 12742 10421 0 net149
rlabel metal2 32522 26656 32522 26656 0 net15
rlabel metal1 5520 15674 5520 15674 0 net150
rlabel metal1 19918 12920 19918 12920 0 net151
rlabel metal2 16790 10285 16790 10285 0 net152
rlabel metal1 17480 10438 17480 10438 0 net153
rlabel metal4 20884 16592 20884 16592 0 net154
rlabel metal2 20102 12614 20102 12614 0 net155
rlabel metal1 21482 10676 21482 10676 0 net156
rlabel metal1 25484 12954 25484 12954 0 net157
rlabel metal1 20332 20230 20332 20230 0 net158
rlabel metal2 19734 20825 19734 20825 0 net159
rlabel metal1 17986 29750 17986 29750 0 net16
rlabel metal1 22862 12274 22862 12274 0 net160
rlabel metal1 24380 12614 24380 12614 0 net161
rlabel metal1 14996 12750 14996 12750 0 net162
rlabel metal2 17618 13311 17618 13311 0 net163
rlabel metal2 15134 12716 15134 12716 0 net164
rlabel via2 17802 6069 17802 6069 0 net165
rlabel metal1 11546 6222 11546 6222 0 net166
rlabel metal1 17986 13430 17986 13430 0 net167
rlabel metal1 25668 19686 25668 19686 0 net168
rlabel metal1 15272 6290 15272 6290 0 net169
rlabel metal2 25254 3978 25254 3978 0 net17
rlabel metal1 20516 6970 20516 6970 0 net170
rlabel metal1 26450 6936 26450 6936 0 net171
rlabel metal1 18170 13464 18170 13464 0 net172
rlabel metal3 9131 13804 9131 13804 0 net173
rlabel metal1 26450 6222 26450 6222 0 net174
rlabel metal2 20470 25959 20470 25959 0 net175
rlabel metal1 13340 14382 13340 14382 0 net176
rlabel metal2 22034 9248 22034 9248 0 net177
rlabel metal1 9154 14314 9154 14314 0 net178
rlabel metal1 21022 13770 21022 13770 0 net179
rlabel metal2 31510 10336 31510 10336 0 net18
rlabel metal2 13570 15232 13570 15232 0 net180
rlabel metal2 20470 14637 20470 14637 0 net181
rlabel metal1 15870 4624 15870 4624 0 net182
rlabel metal2 9338 21471 9338 21471 0 net183
rlabel metal1 14950 13294 14950 13294 0 net184
rlabel via2 12650 7157 12650 7157 0 net185
rlabel metal1 15824 11322 15824 11322 0 net186
rlabel metal1 15180 12614 15180 12614 0 net187
rlabel metal2 13478 13940 13478 13940 0 net188
rlabel metal2 13018 9486 13018 9486 0 net189
rlabel metal1 32108 14042 32108 14042 0 net19
rlabel metal1 13754 7378 13754 7378 0 net190
rlabel via2 15042 15453 15042 15453 0 net191
rlabel metal1 13018 10642 13018 10642 0 net192
rlabel metal2 15042 21471 15042 21471 0 net193
rlabel metal3 18722 19108 18722 19108 0 net194
rlabel metal2 14582 10370 14582 10370 0 net195
rlabel metal2 12926 8721 12926 8721 0 net196
rlabel metal1 16928 8602 16928 8602 0 net197
rlabel metal1 7682 18088 7682 18088 0 net198
rlabel metal1 15778 10234 15778 10234 0 net199
rlabel via1 1697 28526 1697 28526 0 net2
rlabel metal1 32200 11322 32200 11322 0 net20
rlabel metal1 13110 17544 13110 17544 0 net200
rlabel metal1 7590 18258 7590 18258 0 net201
rlabel metal1 16468 9350 16468 9350 0 net202
rlabel metal1 8372 17102 8372 17102 0 net203
rlabel metal1 9798 16422 9798 16422 0 net204
rlabel metal2 18262 9724 18262 9724 0 net205
rlabel metal1 14628 17170 14628 17170 0 net206
rlabel metal1 9936 10234 9936 10234 0 net207
rlabel metal1 9062 11764 9062 11764 0 net208
rlabel metal2 18538 5440 18538 5440 0 net209
rlabel metal2 32154 25058 32154 25058 0 net21
rlabel metal1 10028 19754 10028 19754 0 net210
rlabel metal1 17848 9554 17848 9554 0 net211
rlabel metal1 13616 14042 13616 14042 0 net212
rlabel metal2 13800 13906 13800 13906 0 net213
rlabel metal1 15134 17612 15134 17612 0 net214
rlabel metal2 17158 24514 17158 24514 0 net215
rlabel metal2 6394 16167 6394 16167 0 net216
rlabel metal2 15042 16439 15042 16439 0 net217
rlabel metal1 19044 6902 19044 6902 0 net218
rlabel metal1 5842 13940 5842 13940 0 net219
rlabel metal1 20976 3366 20976 3366 0 net22
rlabel metal1 16928 18326 16928 18326 0 net220
rlabel metal1 16928 18190 16928 18190 0 net221
rlabel metal1 17618 21998 17618 21998 0 net222
rlabel metal1 17572 22610 17572 22610 0 net223
rlabel metal2 11638 11186 11638 11186 0 net224
rlabel metal3 22080 17000 22080 17000 0 net225
rlabel metal1 18032 18598 18032 18598 0 net226
rlabel metal1 11086 9996 11086 9996 0 net227
rlabel metal1 11454 17782 11454 17782 0 net228
rlabel metal2 14858 12206 14858 12206 0 net229
rlabel metal2 32522 9792 32522 9792 0 net23
rlabel metal1 23644 18666 23644 18666 0 net230
rlabel metal2 31418 6035 31418 6035 0 net231
rlabel metal2 13938 27761 13938 27761 0 net232
rlabel metal1 17158 12750 17158 12750 0 net233
rlabel metal1 19136 22746 19136 22746 0 net234
rlabel metal2 16054 26503 16054 26503 0 net235
rlabel metal2 19550 21165 19550 21165 0 net236
rlabel metal1 18354 24820 18354 24820 0 net237
rlabel metal1 22448 24854 22448 24854 0 net238
rlabel metal2 16330 25568 16330 25568 0 net239
rlabel metal1 32338 7378 32338 7378 0 net24
rlabel metal1 24380 25466 24380 25466 0 net240
rlabel metal3 24679 22236 24679 22236 0 net241
rlabel metal1 27600 14314 27600 14314 0 net242
rlabel metal1 24932 6426 24932 6426 0 net243
rlabel metal4 12236 6544 12236 6544 0 net244
rlabel metal2 2116 13124 2116 13124 0 net245
rlabel metal1 26312 13702 26312 13702 0 net246
rlabel metal1 17250 16422 17250 16422 0 net247
rlabel metal2 26634 13651 26634 13651 0 net248
rlabel metal3 20447 14484 20447 14484 0 net249
rlabel metal1 32706 18938 32706 18938 0 net25
rlabel metal1 7682 10982 7682 10982 0 net250
rlabel metal1 19090 14892 19090 14892 0 net251
rlabel metal2 18906 15079 18906 15079 0 net252
rlabel metal1 18722 14382 18722 14382 0 net253
rlabel metal1 21022 11832 21022 11832 0 net254
rlabel metal1 19458 21522 19458 21522 0 net255
rlabel metal3 23069 15300 23069 15300 0 net256
rlabel metal1 24610 16966 24610 16966 0 net257
rlabel metal2 21482 16847 21482 16847 0 net258
rlabel metal2 25116 15844 25116 15844 0 net259
rlabel metal2 32246 6800 32246 6800 0 net26
rlabel metal3 15916 9452 15916 9452 0 net260
rlabel metal2 9154 9180 9154 9180 0 net261
rlabel metal1 26542 9384 26542 9384 0 net262
rlabel metal1 17986 8942 17986 8942 0 net263
rlabel metal2 18446 21148 18446 21148 0 net264
rlabel metal1 15272 12818 15272 12818 0 net265
rlabel metal1 17342 14790 17342 14790 0 net266
rlabel metal2 18170 21046 18170 21046 0 net267
rlabel metal1 17894 19346 17894 19346 0 net268
rlabel metal1 25898 21080 25898 21080 0 net269
rlabel metal2 32246 15878 32246 15878 0 net27
rlabel metal1 7176 17306 7176 17306 0 net270
rlabel metal1 9338 10098 9338 10098 0 net271
rlabel metal1 26818 21454 26818 21454 0 net272
rlabel metal2 23782 26588 23782 26588 0 net273
rlabel metal1 14352 20774 14352 20774 0 net274
rlabel metal1 26818 20774 26818 20774 0 net275
rlabel metal2 13018 19499 13018 19499 0 net276
rlabel metal2 7498 18972 7498 18972 0 net277
rlabel metal1 20240 16626 20240 16626 0 net278
rlabel metal1 25576 21114 25576 21114 0 net279
rlabel metal1 32568 22950 32568 22950 0 net28
rlabel metal1 18860 13906 18860 13906 0 net280
rlabel metal3 25645 10948 25645 10948 0 net281
rlabel via2 15042 26571 15042 26571 0 net282
rlabel metal1 9246 19856 9246 19856 0 net283
rlabel metal1 14260 26554 14260 26554 0 net284
rlabel metal1 8142 19856 8142 19856 0 net285
rlabel metal1 27646 26520 27646 26520 0 net286
rlabel via2 6670 17187 6670 17187 0 net287
rlabel metal2 28382 25347 28382 25347 0 net288
rlabel metal2 12742 22304 12742 22304 0 net289
rlabel metal1 32108 18394 32108 18394 0 net29
rlabel metal1 29624 18190 29624 18190 0 net290
rlabel metal1 14168 23494 14168 23494 0 net291
rlabel metal2 21942 24089 21942 24089 0 net292
rlabel metal1 28106 24242 28106 24242 0 net293
rlabel metal2 28658 19482 28658 19482 0 net294
rlabel metal1 28014 24650 28014 24650 0 net295
rlabel metal2 23874 20128 23874 20128 0 net296
rlabel metal1 13524 19278 13524 19278 0 net297
rlabel metal1 27692 19278 27692 19278 0 net298
rlabel via2 17710 21301 17710 21301 0 net299
rlabel metal1 1656 27642 1656 27642 0 net3
rlabel metal1 32108 17170 32108 17170 0 net30
rlabel metal1 24932 23834 24932 23834 0 net300
rlabel metal1 13984 21998 13984 21998 0 net301
rlabel via1 18262 24854 18262 24854 0 net302
rlabel metal1 25346 26962 25346 26962 0 net303
rlabel metal1 23138 23596 23138 23596 0 net304
rlabel metal2 13110 23783 13110 23783 0 net305
rlabel metal1 22356 23086 22356 23086 0 net306
rlabel metal1 13800 23698 13800 23698 0 net307
rlabel metal1 14076 28050 14076 28050 0 net308
rlabel metal1 18124 27846 18124 27846 0 net309
rlabel metal2 32246 11968 32246 11968 0 net31
rlabel metal2 414 16320 414 16320 0 net310
rlabel metal1 1150 23630 1150 23630 0 net311
rlabel metal1 22448 23018 22448 23018 0 net312
rlabel metal2 21482 26316 21482 26316 0 net313
rlabel metal2 19918 25092 19918 25092 0 net314
rlabel metal1 12604 23698 12604 23698 0 net315
rlabel metal1 20056 24718 20056 24718 0 net316
rlabel metal1 21114 25670 21114 25670 0 net317
rlabel metal1 21482 25262 21482 25262 0 net318
rlabel metal1 21160 22202 21160 22202 0 net319
rlabel metal1 19412 30226 19412 30226 0 net32
rlabel metal1 21988 24922 21988 24922 0 net320
rlabel metal1 21298 24786 21298 24786 0 net321
rlabel metal2 19366 22491 19366 22491 0 net322
rlabel metal2 16790 22032 16790 22032 0 net323
rlabel metal1 20378 16694 20378 16694 0 net324
rlabel metal1 17940 24786 17940 24786 0 net325
rlabel metal3 15249 21284 15249 21284 0 net326
rlabel metal1 22678 20366 22678 20366 0 net327
rlabel metal3 12098 30260 12098 30260 0 net328
rlabel metal1 20746 17646 20746 17646 0 net329
rlabel metal1 17756 2414 17756 2414 0 net33
rlabel metal2 23460 24786 23460 24786 0 net330
rlabel metal3 2116 19312 2116 19312 0 net331
rlabel metal2 20746 23664 20746 23664 0 net332
rlabel metal1 23092 21998 23092 21998 0 net333
rlabel metal1 12558 17646 12558 17646 0 net334
rlabel metal2 20654 16354 20654 16354 0 net335
rlabel metal1 12144 14926 12144 14926 0 net336
rlabel metal2 6578 25942 6578 25942 0 net337
rlabel metal1 5842 25874 5842 25874 0 net338
rlabel metal1 10718 28424 10718 28424 0 net339
rlabel metal2 31786 21420 31786 21420 0 net34
rlabel metal2 11546 28730 11546 28730 0 net340
rlabel metal2 8786 28322 8786 28322 0 net341
rlabel metal2 10074 28628 10074 28628 0 net342
rlabel metal1 5934 24038 5934 24038 0 net343
rlabel metal2 4738 7174 4738 7174 0 net344
rlabel metal1 4048 7446 4048 7446 0 net345
rlabel metal2 2990 10234 2990 10234 0 net346
rlabel metal1 4738 21114 4738 21114 0 net347
rlabel metal2 2208 13396 2208 13396 0 net348
rlabel metal2 9706 8704 9706 8704 0 net349
rlabel metal2 31878 24990 31878 24990 0 net35
rlabel metal2 10350 9010 10350 9010 0 net350
rlabel metal1 9062 13226 9062 13226 0 net351
rlabel metal1 8786 13872 8786 13872 0 net352
rlabel metal1 5014 18292 5014 18292 0 net353
rlabel metal1 8096 21318 8096 21318 0 net354
rlabel metal1 4002 20230 4002 20230 0 net355
rlabel metal2 9890 8636 9890 8636 0 net356
rlabel metal2 10534 8942 10534 8942 0 net357
rlabel metal2 10994 9282 10994 9282 0 net358
rlabel metal2 9890 14059 9890 14059 0 net359
rlabel metal1 21804 30362 21804 30362 0 net36
rlabel metal2 4278 21369 4278 21369 0 net360
rlabel metal2 4094 21675 4094 21675 0 net361
rlabel metal2 8142 7820 8142 7820 0 net362
rlabel metal1 8050 8500 8050 8500 0 net363
rlabel metal1 7268 8806 7268 8806 0 net364
rlabel metal1 7107 8942 7107 8942 0 net365
rlabel metal1 8510 11628 8510 11628 0 net366
rlabel metal1 7544 20502 7544 20502 0 net367
rlabel metal2 6578 22729 6578 22729 0 net368
rlabel metal1 8832 7854 8832 7854 0 net369
rlabel metal1 25300 2414 25300 2414 0 net37
rlabel metal1 8280 8466 8280 8466 0 net370
rlabel metal2 7774 7786 7774 7786 0 net371
rlabel metal1 4738 10744 4738 10744 0 net372
rlabel metal1 5014 10982 5014 10982 0 net373
rlabel metal1 6762 22644 6762 22644 0 net374
rlabel metal2 8326 18751 8326 18751 0 net375
rlabel metal1 5980 23834 5980 23834 0 net376
rlabel metal2 6762 7616 6762 7616 0 net377
rlabel via2 4278 7395 4278 7395 0 net378
rlabel metal1 4048 12410 4048 12410 0 net379
rlabel metal1 23552 29818 23552 29818 0 net38
rlabel metal1 6302 21318 6302 21318 0 net380
rlabel metal1 6072 21046 6072 21046 0 net381
rlabel via2 5474 20893 5474 20893 0 net382
rlabel metal1 4186 17680 4186 17680 0 net383
rlabel metal1 4278 18768 4278 18768 0 net384
rlabel metal1 6992 22746 6992 22746 0 net385
rlabel metal1 5152 22474 5152 22474 0 net386
rlabel metal1 5934 18768 5934 18768 0 net387
rlabel metal1 5704 17170 5704 17170 0 net388
rlabel metal2 7360 19822 7360 19822 0 net389
rlabel metal1 25300 29138 25300 29138 0 net39
rlabel metal1 7544 22746 7544 22746 0 net390
rlabel metal1 7498 22406 7498 22406 0 net391
rlabel metal1 5980 23086 5980 23086 0 net392
rlabel metal2 5382 23358 5382 23358 0 net393
rlabel via1 6486 9146 6486 9146 0 net394
rlabel metal1 5566 9656 5566 9656 0 net395
rlabel metal2 4002 10438 4002 10438 0 net396
rlabel metal2 3542 9214 3542 9214 0 net397
rlabel metal1 2760 16490 2760 16490 0 net398
rlabel metal1 3312 17238 3312 17238 0 net399
rlabel metal1 1656 24378 1656 24378 0 net4
rlabel metal1 32108 21658 32108 21658 0 net40
rlabel metal1 2622 18224 2622 18224 0 net400
rlabel metal2 6670 9146 6670 9146 0 net401
rlabel metal1 5796 9554 5796 9554 0 net402
rlabel metal1 4554 10642 4554 10642 0 net403
rlabel metal1 3726 9520 3726 9520 0 net404
rlabel metal2 3542 11900 3542 11900 0 net405
rlabel metal2 2254 15708 2254 15708 0 net406
rlabel metal1 3358 17170 3358 17170 0 net407
rlabel metal1 5796 19822 5796 19822 0 net408
rlabel metal1 3450 14926 3450 14926 0 net409
rlabel metal1 18446 3400 18446 3400 0 net41
rlabel metal2 9614 22049 9614 22049 0 net410
rlabel metal1 7222 26248 7222 26248 0 net411
rlabel metal1 8878 26010 8878 26010 0 net412
rlabel metal1 7682 25262 7682 25262 0 net413
rlabel metal1 9338 27336 9338 27336 0 net414
rlabel metal1 11684 29002 11684 29002 0 net415
rlabel metal1 9890 25976 9890 25976 0 net416
rlabel metal1 8326 28186 8326 28186 0 net417
rlabel metal2 9706 25670 9706 25670 0 net418
rlabel metal1 7268 26350 7268 26350 0 net419
rlabel metal1 23874 4590 23874 4590 0 net42
rlabel metal1 7728 26010 7728 26010 0 net420
rlabel metal1 9568 27438 9568 27438 0 net421
rlabel metal1 12880 28186 12880 28186 0 net422
rlabel metal1 11362 26282 11362 26282 0 net423
rlabel metal1 9844 28050 9844 28050 0 net424
rlabel metal1 9522 29206 9522 29206 0 net425
rlabel metal1 6578 10166 6578 10166 0 net426
rlabel metal1 9062 8364 9062 8364 0 net427
rlabel metal1 7774 7854 7774 7854 0 net428
rlabel metal1 10442 24208 10442 24208 0 net429
rlabel metal2 29026 7242 29026 7242 0 net43
rlabel metal2 6670 28492 6670 28492 0 net430
rlabel metal1 6900 29002 6900 29002 0 net431
rlabel metal3 943 20740 943 20740 0 net432
rlabel metal2 5658 8432 5658 8432 0 net433
rlabel via2 9246 8228 9246 8228 0 net434
rlabel metal2 6026 11441 6026 11441 0 net435
rlabel metal1 10672 29478 10672 29478 0 net436
rlabel metal1 10626 29580 10626 29580 0 net437
rlabel metal1 7038 28526 7038 28526 0 net438
rlabel metal2 7498 29359 7498 29359 0 net439
rlabel metal1 30636 10438 30636 10438 0 net44
rlabel metal2 5566 8772 5566 8772 0 net440
rlabel metal2 8234 7463 8234 7463 0 net441
rlabel metal2 10166 13532 10166 13532 0 net442
rlabel metal2 9982 27676 9982 27676 0 net443
rlabel metal2 9798 28356 9798 28356 0 net444
rlabel metal1 8326 28084 8326 28084 0 net445
rlabel metal4 2668 23732 2668 23732 0 net446
rlabel metal2 9890 29087 9890 29087 0 net447
rlabel metal2 6394 7310 6394 7310 0 net448
rlabel metal1 7912 7378 7912 7378 0 net449
rlabel metal2 30452 10642 30452 10642 0 net45
rlabel metal2 8510 11900 8510 11900 0 net450
rlabel metal2 10166 26350 10166 26350 0 net451
rlabel metal1 10166 26248 10166 26248 0 net452
rlabel metal1 10534 26350 10534 26350 0 net453
rlabel metal1 7820 17510 7820 17510 0 net454
rlabel metal2 11086 26911 11086 26911 0 net455
rlabel metal1 2898 11152 2898 11152 0 net456
rlabel metal1 3818 13362 3818 13362 0 net457
rlabel metal1 4784 13906 4784 13906 0 net458
rlabel metal1 2438 17238 2438 17238 0 net459
rlabel metal1 30498 14586 30498 14586 0 net46
rlabel metal1 9154 24072 9154 24072 0 net460
rlabel metal1 9154 28424 9154 28424 0 net461
rlabel metal2 9246 27642 9246 27642 0 net462
rlabel metal2 9430 29019 9430 29019 0 net463
rlabel metal4 2484 23528 2484 23528 0 net464
rlabel metal1 8970 29206 8970 29206 0 net465
rlabel metal1 2714 11118 2714 11118 0 net466
rlabel metal1 3680 12206 3680 12206 0 net467
rlabel metal1 5106 13294 5106 13294 0 net468
rlabel metal1 3082 17510 3082 17510 0 net469
rlabel metal1 31096 14586 31096 14586 0 net47
rlabel metal2 9338 24276 9338 24276 0 net470
rlabel metal1 8924 28662 8924 28662 0 net471
rlabel metal1 8280 28390 8280 28390 0 net472
rlabel metal1 8142 28526 8142 28526 0 net473
rlabel metal2 8878 29478 8878 29478 0 net474
rlabel metal2 2714 18054 2714 18054 0 net475
rlabel metal1 5244 18326 5244 18326 0 net476
rlabel metal2 4370 20978 4370 20978 0 net477
rlabel metal1 5014 25942 5014 25942 0 net478
rlabel metal2 5566 26146 5566 26146 0 net479
rlabel metal1 31096 14858 31096 14858 0 net48
rlabel metal1 5014 26384 5014 26384 0 net480
rlabel metal2 6302 24956 6302 24956 0 net481
rlabel metal1 6118 27472 6118 27472 0 net482
rlabel metal2 2714 16796 2714 16796 0 net483
rlabel metal1 3634 18360 3634 18360 0 net484
rlabel metal1 3772 18258 3772 18258 0 net485
rlabel metal1 5934 24786 5934 24786 0 net486
rlabel metal2 6394 26180 6394 26180 0 net487
rlabel metal1 5750 25296 5750 25296 0 net488
rlabel metal2 5290 25092 5290 25092 0 net489
rlabel via2 30866 14773 30866 14773 0 net49
rlabel metal1 5520 26554 5520 26554 0 net490
rlabel metal1 4600 9622 4600 9622 0 net491
rlabel metal1 7590 9588 7590 9588 0 net492
rlabel metal2 4094 10880 4094 10880 0 net493
rlabel metal2 5658 16099 5658 16099 0 net494
rlabel metal1 8326 26894 8326 26894 0 net495
rlabel metal1 7268 26962 7268 26962 0 net496
rlabel metal1 6900 27438 6900 27438 0 net497
rlabel metal1 7912 27846 7912 27846 0 net498
rlabel via3 6509 17884 6509 17884 0 net499
rlabel metal1 1564 14586 1564 14586 0 net5
rlabel metal1 30958 20944 30958 20944 0 net50
rlabel metal2 5014 12308 5014 12308 0 net500
rlabel metal1 5750 9622 5750 9622 0 net501
rlabel metal2 5382 15232 5382 15232 0 net502
rlabel metal2 7866 25670 7866 25670 0 net503
rlabel metal1 7452 27030 7452 27030 0 net504
rlabel metal1 7268 27438 7268 27438 0 net505
rlabel metal1 7452 21590 7452 21590 0 net506
rlabel metal3 6785 19108 6785 19108 0 net507
rlabel metal1 6670 25840 6670 25840 0 net508
rlabel metal1 6624 27098 6624 27098 0 net509
rlabel metal2 30866 20774 30866 20774 0 net51
rlabel metal1 12374 28560 12374 28560 0 net510
rlabel metal1 10258 27370 10258 27370 0 net511
rlabel metal2 10810 28628 10810 28628 0 net512
rlabel metal1 11132 27574 11132 27574 0 net513
rlabel metal1 6394 26928 6394 26928 0 net514
rlabel metal1 7682 21488 7682 21488 0 net515
rlabel metal1 4600 23698 4600 23698 0 net516
rlabel metal2 4370 24769 4370 24769 0 net517
rlabel metal1 5704 19754 5704 19754 0 net518
rlabel metal2 8234 20706 8234 20706 0 net519
rlabel metal2 31878 19924 31878 19924 0 net52
rlabel metal1 6394 21658 6394 21658 0 net520
rlabel metal1 8602 22644 8602 22644 0 net521
rlabel metal2 11730 26078 11730 26078 0 net522
rlabel metal1 12466 28016 12466 28016 0 net523
rlabel via2 5934 22117 5934 22117 0 net524
rlabel metal1 6210 20230 6210 20230 0 net525
rlabel metal1 6900 20434 6900 20434 0 net526
rlabel via1 5290 21862 5290 21862 0 net527
rlabel metal1 4968 21998 4968 21998 0 net528
rlabel metal2 11454 26146 11454 26146 0 net529
rlabel metal1 29854 25976 29854 25976 0 net53
rlabel metal1 11500 28050 11500 28050 0 net530
rlabel metal2 6210 21777 6210 21777 0 net531
rlabel metal1 4094 8568 4094 8568 0 net532
rlabel metal1 10442 9520 10442 9520 0 net533
rlabel via3 5451 8364 5451 8364 0 net534
rlabel metal2 12282 25058 12282 25058 0 net535
rlabel metal2 12926 28577 12926 28577 0 net536
rlabel metal1 12627 29274 12627 29274 0 net537
rlabel metal2 13294 27047 13294 27047 0 net538
rlabel metal3 2093 19652 2093 19652 0 net539
rlabel metal1 31142 18598 31142 18598 0 net54
rlabel metal1 8694 24650 8694 24650 0 net540
rlabel metal1 10810 25296 10810 25296 0 net541
rlabel metal1 12466 25330 12466 25330 0 net542
rlabel metal1 10902 24140 10902 24140 0 net543
rlabel metal1 6026 24684 6026 24684 0 net544
rlabel metal2 4830 7548 4830 7548 0 net545
rlabel metal1 10166 9588 10166 9588 0 net546
rlabel metal1 4324 11866 4324 11866 0 net547
rlabel metal1 12420 28458 12420 28458 0 net548
rlabel metal1 12650 28560 12650 28560 0 net549
rlabel metal1 17848 29546 17848 29546 0 net55
rlabel metal1 13156 28730 13156 28730 0 net550
rlabel metal1 7268 23086 7268 23086 0 net551
rlabel metal2 5474 22729 5474 22729 0 net552
rlabel metal1 9890 24208 9890 24208 0 net553
rlabel metal1 11408 24378 11408 24378 0 net554
rlabel metal1 11132 25126 11132 25126 0 net555
rlabel via2 9522 24565 9522 24565 0 net556
rlabel metal2 6946 24412 6946 24412 0 net557
rlabel metal1 18630 3536 18630 3536 0 net558
rlabel metal2 24242 5100 24242 5100 0 net559
rlabel metal1 31004 18734 31004 18734 0 net56
rlabel metal1 29118 7752 29118 7752 0 net560
rlabel metal1 31924 9554 31924 9554 0 net561
rlabel metal2 31602 7684 31602 7684 0 net562
rlabel metal2 30314 14807 30314 14807 0 net563
rlabel metal1 30728 14586 30728 14586 0 net564
rlabel metal1 31096 14246 31096 14246 0 net565
rlabel metal2 30912 14382 30912 14382 0 net566
rlabel metal1 31142 20842 31142 20842 0 net567
rlabel metal1 30912 20026 30912 20026 0 net568
rlabel metal1 30360 19482 30360 19482 0 net569
rlabel metal2 27830 13906 27830 13906 0 net57
rlabel metal2 29946 27574 29946 27574 0 net570
rlabel metal1 29900 19346 29900 19346 0 net571
rlabel metal2 18446 29376 18446 29376 0 net572
rlabel metal2 31786 15334 31786 15334 0 net573
rlabel metal1 2070 20570 2070 20570 0 net574
rlabel metal1 1518 20944 1518 20944 0 net575
rlabel metal2 3910 21284 3910 21284 0 net576
rlabel metal1 2898 24140 2898 24140 0 net577
rlabel metal1 4186 24242 4186 24242 0 net578
rlabel metal1 2691 23222 2691 23222 0 net579
rlabel metal2 13984 9316 13984 9316 0 net58
rlabel metal1 2116 23290 2116 23290 0 net580
rlabel metal2 3266 20672 3266 20672 0 net581
rlabel metal1 3174 21658 3174 21658 0 net582
rlabel metal2 2714 21845 2714 21845 0 net583
rlabel metal2 4462 20774 4462 20774 0 net584
rlabel metal1 2714 24038 2714 24038 0 net585
rlabel metal2 1886 23970 1886 23970 0 net586
rlabel metal1 3726 24718 3726 24718 0 net587
rlabel metal2 2438 24310 2438 24310 0 net588
rlabel metal1 2300 20910 2300 20910 0 net589
rlabel metal2 14766 11645 14766 11645 0 net59
rlabel metal2 2622 20706 2622 20706 0 net590
rlabel metal1 2208 21046 2208 21046 0 net591
rlabel metal1 2898 24344 2898 24344 0 net592
rlabel metal1 4324 24650 4324 24650 0 net593
rlabel metal1 4278 24854 4278 24854 0 net594
rlabel metal2 3082 24548 3082 24548 0 net595
rlabel metal1 2254 20808 2254 20808 0 net596
rlabel metal2 2346 20060 2346 20060 0 net597
rlabel metal1 3496 21454 3496 21454 0 net598
rlabel metal1 2530 22032 2530 22032 0 net599
rlabel metal1 1656 19482 1656 19482 0 net6
rlabel metal1 26312 25194 26312 25194 0 net60
rlabel metal1 4968 24106 4968 24106 0 net600
rlabel metal1 3358 25160 3358 25160 0 net601
rlabel metal1 2990 24650 2990 24650 0 net602
rlabel metal1 2438 23562 2438 23562 0 net603
rlabel metal2 2254 22610 2254 22610 0 net604
rlabel metal1 2254 26928 2254 26928 0 net605
rlabel metal1 2622 27540 2622 27540 0 net606
rlabel metal1 5980 27914 5980 27914 0 net607
rlabel metal2 5382 28424 5382 28424 0 net608
rlabel metal2 4922 26758 4922 26758 0 net609
rlabel via2 11178 15861 11178 15861 0 net61
rlabel metal1 2070 27030 2070 27030 0 net610
rlabel metal1 3128 26418 3128 26418 0 net611
rlabel metal2 3726 25772 3726 25772 0 net612
rlabel metal1 3174 29478 3174 29478 0 net613
rlabel metal1 5244 28390 5244 28390 0 net614
rlabel metal1 4876 28050 4876 28050 0 net615
rlabel metal1 4002 29172 4002 29172 0 net616
rlabel metal1 3542 25942 3542 25942 0 net617
rlabel metal1 2944 27370 2944 27370 0 net618
rlabel metal1 4968 28594 4968 28594 0 net619
rlabel metal2 20930 7140 20930 7140 0 net62
rlabel metal1 4324 29002 4324 29002 0 net620
rlabel metal1 4416 29138 4416 29138 0 net621
rlabel metal2 2806 29121 2806 29121 0 net622
rlabel metal1 3174 25840 3174 25840 0 net623
rlabel metal1 2438 27370 2438 27370 0 net624
rlabel metal1 2944 28730 2944 28730 0 net625
rlabel metal1 4784 27914 4784 27914 0 net626
rlabel metal2 4370 28322 4370 28322 0 net627
rlabel metal1 4692 27098 4692 27098 0 net628
rlabel metal1 2530 29206 2530 29206 0 net629
rlabel metal2 25070 12172 25070 12172 0 net63
rlabel metal2 29670 1588 29670 1588 0 net630
rlabel metal2 18538 3978 18538 3978 0 net631
rlabel metal2 30866 6970 30866 6970 0 net632
rlabel metal1 31188 16082 31188 16082 0 net633
rlabel metal1 31188 8466 31188 8466 0 net634
rlabel metal1 31510 12206 31510 12206 0 net635
rlabel metal1 31602 16558 31602 16558 0 net636
rlabel metal1 31188 19346 31188 19346 0 net637
rlabel metal2 29210 24378 29210 24378 0 net638
rlabel metal2 30314 23868 30314 23868 0 net639
rlabel metal1 18998 21352 18998 21352 0 net64
rlabel metal1 31602 21998 31602 21998 0 net640
rlabel metal2 31326 26758 31326 26758 0 net641
rlabel metal1 31372 20910 31372 20910 0 net642
rlabel metal1 31188 20434 31188 20434 0 net643
rlabel metal1 30590 10064 30590 10064 0 net644
rlabel metal1 31510 17646 31510 17646 0 net645
rlabel metal1 31510 13294 31510 13294 0 net646
rlabel metal1 29946 9588 29946 9588 0 net647
rlabel metal1 22862 4590 22862 4590 0 net648
rlabel metal1 16744 3502 16744 3502 0 net649
rlabel metal1 18768 16762 18768 16762 0 net65
rlabel metal2 29210 7684 29210 7684 0 net650
rlabel metal1 25024 5202 25024 5202 0 net651
rlabel metal2 21206 4420 21206 4420 0 net652
rlabel metal2 23966 4726 23966 4726 0 net653
rlabel metal1 30498 25874 30498 25874 0 net654
rlabel metal2 30590 10948 30590 10948 0 net655
rlabel metal2 20930 29818 20930 29818 0 net656
rlabel metal1 24472 29138 24472 29138 0 net657
rlabel metal2 30130 22780 30130 22780 0 net658
rlabel metal1 22356 29138 22356 29138 0 net659
rlabel metal2 19458 16014 19458 16014 0 net66
rlabel metal1 17250 29138 17250 29138 0 net660
rlabel metal1 18722 29614 18722 29614 0 net661
rlabel metal1 20792 8466 20792 8466 0 net67
rlabel metal1 22862 18292 22862 18292 0 net68
rlabel metal2 16054 9299 16054 9299 0 net69
rlabel via1 1697 18666 1697 18666 0 net7
rlabel metal1 16146 11254 16146 11254 0 net70
rlabel metal2 16514 11169 16514 11169 0 net71
rlabel metal2 2530 13498 2530 13498 0 net72
rlabel metal1 16284 12750 16284 12750 0 net73
rlabel metal1 16606 14586 16606 14586 0 net74
rlabel metal1 29716 13430 29716 13430 0 net75
rlabel metal1 16376 12818 16376 12818 0 net76
rlabel metal1 10948 11866 10948 11866 0 net77
rlabel metal2 4094 13503 4094 13503 0 net78
rlabel metal1 3956 15674 3956 15674 0 net79
rlabel metal2 1610 19251 1610 19251 0 net8
rlabel metal2 9338 5899 9338 5899 0 net80
rlabel metal1 19826 6358 19826 6358 0 net81
rlabel metal1 19780 6222 19780 6222 0 net82
rlabel metal1 11086 14280 11086 14280 0 net83
rlabel metal2 20102 6426 20102 6426 0 net84
rlabel metal1 19458 9588 19458 9588 0 net85
rlabel metal2 17434 5899 17434 5899 0 net86
rlabel metal1 14812 26282 14812 26282 0 net87
rlabel metal2 20010 6562 20010 6562 0 net88
rlabel metal1 20838 6358 20838 6358 0 net89
rlabel metal1 31878 12784 31878 12784 0 net9
rlabel metal1 13110 9486 13110 9486 0 net90
rlabel metal1 16652 9690 16652 9690 0 net91
rlabel metal3 16813 11492 16813 11492 0 net92
rlabel metal2 17250 8313 17250 8313 0 net93
rlabel metal1 15272 15334 15272 15334 0 net94
rlabel metal2 10534 16983 10534 16983 0 net95
rlabel metal1 16284 15470 16284 15470 0 net96
rlabel metal1 7360 14926 7360 14926 0 net97
rlabel metal1 11408 8058 11408 8058 0 net98
rlabel metal1 15456 12818 15456 12818 0 net99
<< properties >>
string FIXED_BBOX 0 0 34000 34000
<< end >>
