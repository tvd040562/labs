assign table2[0] = 32'h00000000;
assign table2[1] = 32'hff36f078;
assign table2[2] = 32'hfe6de2e0;
assign table2[3] = 32'hfda4d929;
assign table2[4] = 32'hfcdbd541;
assign table2[5] = 32'hfc12d91a;
assign table2[6] = 32'hfb49e6a3;
assign table2[7] = 32'hfa80ffcb;
assign table2[8] = 32'hf9b82684;
assign table2[9] = 32'hf8ef5cbb;
assign table2[10] = 32'hf826a462;
assign table2[11] = 32'hf75dff66;
assign table2[12] = 32'hf6956fb7;
assign table2[13] = 32'hf5ccf744;
assign table2[14] = 32'hf50497fb;
assign table2[15] = 32'hf43c53cb;
assign table2[16] = 32'hf3742ca2;
assign table2[17] = 32'hf2ac246e;
assign table2[18] = 32'hf1e43d1c;
assign table2[19] = 32'hf11c789a;
assign table2[20] = 32'hf054d8d5;
assign table2[21] = 32'hef8d5fb8;
assign table2[22] = 32'heec60f31;
assign table2[23] = 32'hedfee92b;
assign table2[24] = 32'hed37ef92;
assign table2[25] = 32'hec71244f;
assign table2[26] = 32'hebaa894f;
assign table2[27] = 32'heae4207b;
assign table2[28] = 32'hea1debbc;
assign table2[29] = 32'he957ecfb;
assign table2[30] = 32'he8922622;
assign table2[31] = 32'he7cc9918;
assign table2[32] = 32'he70747c4;
assign table2[33] = 32'he642340d;
assign table2[34] = 32'he57d5fdb;
assign table2[35] = 32'he4b8cd11;
assign table2[36] = 32'he3f47d96;
assign table2[37] = 32'he330734d;
assign table2[38] = 32'he26cb01b;
assign table2[39] = 32'he1a935e2;
assign table2[40] = 32'he0e60685;
assign table2[41] = 32'he02323e5;
assign table2[42] = 32'hdf608fe4;
assign table2[43] = 32'hde9e4c61;
assign table2[44] = 32'hdddc5b3b;
assign table2[45] = 32'hdd1abe51;
assign table2[46] = 32'hdc597782;
assign table2[47] = 32'hdb9888a9;
assign table2[48] = 32'hdad7f3a3;
assign table2[49] = 32'hda17ba4a;
assign table2[50] = 32'hd957de7b;
assign table2[51] = 32'hd898620c;
assign table2[52] = 32'hd7d946d8;
assign table2[53] = 32'hd71a8eb6;
assign table2[54] = 32'hd65c3b7b;
assign table2[55] = 32'hd59e4eff;
assign table2[56] = 32'hd4e0cb15;
assign table2[57] = 32'hd423b191;
assign table2[58] = 32'hd3670446;
assign table2[59] = 32'hd2aac505;
assign table2[60] = 32'hd1eef59e;
assign table2[61] = 32'hd13397e2;
assign table2[62] = 32'hd078ad9e;
assign table2[63] = 32'hcfbe38a0;
assign table2[64] = 32'hcf043ab3;
assign table2[65] = 32'hce4ab5a3;
assign table2[66] = 32'hcd91ab39;
assign table2[67] = 32'hccd91d3e;
assign table2[68] = 32'hcc210d79;
assign table2[69] = 32'hcb697db1;
assign table2[70] = 32'hcab26faa;
assign table2[71] = 32'hc9fbe527;
assign table2[72] = 32'hc945dfed;
assign table2[73] = 32'hc89061ba;
assign table2[74] = 32'hc7db6c50;
assign table2[75] = 32'hc727016d;
assign table2[76] = 32'hc67322ce;
assign table2[77] = 32'hc5bfd22f;
assign table2[78] = 32'hc50d1149;
assign table2[79] = 32'hc45ae1d7;
assign table2[80] = 32'hc3a94590;
assign table2[81] = 32'hc2f83e2b;
assign table2[82] = 32'hc247cd5b;
assign table2[83] = 32'hc197f4d4;
assign table2[84] = 32'hc0e8b649;
assign table2[85] = 32'hc03a1369;
assign table2[86] = 32'hbf8c0de3;
assign table2[87] = 32'hbedea766;
assign table2[88] = 32'hbe31e19c;
assign table2[89] = 32'hbd85be30;
assign table2[90] = 32'hbcda3ecb;
assign table2[91] = 32'hbc2f6514;
assign table2[92] = 32'hbb8532b0;
assign table2[93] = 32'hbadba944;
assign table2[94] = 32'hba32ca71;
assign table2[95] = 32'hb98a97d9;
assign table2[96] = 32'hb8e3131a;
assign table2[97] = 32'hb83c3dd2;
assign table2[98] = 32'hb796199c;
assign table2[99] = 32'hb6f0a812;
assign table2[100] = 32'hb64beacd;
assign table2[101] = 32'hb5a7e363;
assign table2[102] = 32'hb5049369;
assign table2[103] = 32'hb461fc71;
assign table2[104] = 32'hb3c0200d;
assign table2[105] = 32'hb31effcc;
assign table2[106] = 32'hb27e9d3d;
assign table2[107] = 32'hb1def9e9;
assign table2[108] = 32'hb140175c;
assign table2[109] = 32'hb0a1f71e;
assign table2[110] = 32'hb0049ab4;
assign table2[111] = 32'haf6803a2;
assign table2[112] = 32'haecc336c;
assign table2[113] = 32'hae312b92;
assign table2[114] = 32'had96ed92;
assign table2[115] = 32'hacfd7ae9;
assign table2[116] = 32'hac64d511;
assign table2[117] = 32'habccfd83;
assign table2[118] = 32'hab35f5b6;
assign table2[119] = 32'haa9fbf1e;
assign table2[120] = 32'haa0a5b2e;
assign table2[121] = 32'ha975cb57;
assign table2[122] = 32'ha8e21107;
assign table2[123] = 32'ha84f2dab;
assign table2[124] = 32'ha7bd22ac;
assign table2[125] = 32'ha72bf174;
assign table2[126] = 32'ha69b9b69;
assign table2[127] = 32'ha60c21ee;
assign table2[128] = 32'ha57d8667;
assign table2[129] = 32'ha4efca32;
assign table2[130] = 32'ha462eead;
assign table2[131] = 32'ha3d6f534;
assign table2[132] = 32'ha34bdf21;
assign table2[133] = 32'ha2c1adca;
assign table2[134] = 32'ha2386285;
assign table2[135] = 32'ha1affea3;
assign table2[136] = 32'ha1288377;
assign table2[137] = 32'ha0a1f24e;
assign table2[138] = 32'ha01c4c73;
assign table2[139] = 32'h9f979332;
assign table2[140] = 32'h9f13c7d1;
assign table2[141] = 32'h9e90eb95;
assign table2[142] = 32'h9e0effc2;
assign table2[143] = 32'h9d8e0598;
assign table2[144] = 32'h9d0dfe54;
assign table2[145] = 32'h9c8eeb34;
assign table2[146] = 32'h9c10cd71;
assign table2[147] = 32'h9b93a641;
assign table2[148] = 32'h9b1776db;
assign table2[149] = 32'h9a9c406f;
assign table2[150] = 32'h9a22042e;
assign table2[151] = 32'h99a8c345;
assign table2[152] = 32'h99307ee1;
assign table2[153] = 32'h98b93829;
assign table2[154] = 32'h9842f044;
assign table2[155] = 32'h97cda856;
assign table2[156] = 32'h97596180;
assign table2[157] = 32'h96e61ce1;
assign table2[158] = 32'h9673db95;
assign table2[159] = 32'h96029eb6;
assign table2[160] = 32'h9592675d;
assign table2[161] = 32'h9523369c;
assign table2[162] = 32'h94b50d88;
assign table2[163] = 32'h9447ed30;
assign table2[164] = 32'h93dbd6a1;
assign table2[165] = 32'h9370cae5;
assign table2[166] = 32'h9306cb05;
assign table2[167] = 32'h929dd807;
assign table2[168] = 32'h9235f2ec;
assign table2[169] = 32'h91cf1cb7;
assign table2[170] = 32'h91695664;
assign table2[171] = 32'h9104a0ef;
assign table2[172] = 32'h90a0fd4f;
assign table2[173] = 32'h903e6c7c;
assign table2[174] = 32'h8fdcef67;
assign table2[175] = 32'h8f7c8702;
assign table2[176] = 32'h8f1d343b;
assign table2[177] = 32'h8ebef7fc;
assign table2[178] = 32'h8e61d32f;
assign table2[179] = 32'h8e05c6b8;
assign table2[180] = 32'h8daad37c;
assign table2[181] = 32'h8d50fa5a;
assign table2[182] = 32'h8cf83c31;
assign table2[183] = 32'h8ca099db;
assign table2[184] = 32'h8c4a1430;
assign table2[185] = 32'h8bf4ac06;
assign table2[186] = 32'h8ba06230;
assign table2[187] = 32'h8b4d377d;
assign table2[188] = 32'h8afb2cbc;
assign table2[189] = 32'h8aaa42b5;
assign table2[190] = 32'h8a5a7a32;
assign table2[191] = 32'h8a0bd3f6;
assign table2[192] = 32'h89be50c4;
assign table2[193] = 32'h8971f15b;
assign table2[194] = 32'h8926b678;
assign table2[195] = 32'h88dca0d4;
assign table2[196] = 32'h8893b126;
assign table2[197] = 32'h884be821;
assign table2[198] = 32'h88054678;
assign table2[199] = 32'h87bfccd8;
assign table2[200] = 32'h877b7bed;
assign table2[201] = 32'h8738545f;
assign table2[202] = 32'h86f656d4;
assign table2[203] = 32'h86b583ef;
assign table2[204] = 32'h8675dc50;
assign table2[205] = 32'h86376093;
assign table2[206] = 32'h85fa1154;
assign table2[207] = 32'h85bdef28;
assign table2[208] = 32'h8582faa6;
assign table2[209] = 32'h8549345d;
assign table2[210] = 32'h85109cdd;
assign table2[211] = 32'h84d934b2;
assign table2[212] = 32'h84a2fc63;
assign table2[213] = 32'h846df478;
assign table2[214] = 32'h843a1d71;
assign table2[215] = 32'h840777d1;
assign table2[216] = 32'h83d60413;
assign table2[217] = 32'h83a5c2b1;
assign table2[218] = 32'h8376b423;
assign table2[219] = 32'h8348d8dd;
assign table2[220] = 32'h831c314f;
assign table2[221] = 32'h82f0bde9;
assign table2[222] = 32'h82c67f15;
assign table2[223] = 32'h829d753b;
assign table2[224] = 32'h8275a0c1;
assign table2[225] = 32'h824f0209;
assign table2[226] = 32'h82299972;
assign table2[227] = 32'h82056759;
assign table2[228] = 32'h81e26c17;
assign table2[229] = 32'h81c0a802;
assign table2[230] = 32'h81a01b6e;
assign table2[231] = 32'h8180c6aa;
assign table2[232] = 32'h8162aa05;
assign table2[233] = 32'h8145c5c8;
assign table2[234] = 32'h812a1a3b;
assign table2[235] = 32'h810fa7a1;
assign table2[236] = 32'h80f66e3d;
assign table2[237] = 32'h80de6e4d;
assign table2[238] = 32'h80c7a80b;
assign table2[239] = 32'h80b21bb0;
assign table2[240] = 32'h809dc972;
assign table2[241] = 32'h808ab181;
assign table2[242] = 32'h8078d40e;
assign table2[243] = 32'h80683144;
assign table2[244] = 32'h8058c94d;
assign table2[245] = 32'h804a9c4e;
assign table2[246] = 32'h803daa6b;
assign table2[247] = 32'h8031f3c3;
assign table2[248] = 32'h80277873;
assign table2[249] = 32'h801e3896;
assign table2[250] = 32'h80163441;
assign table2[251] = 32'h800f6b89;
assign table2[252] = 32'h8009de7f;
assign table2[253] = 32'h80058d30;
assign table2[254] = 32'h800277a7;
assign table2[255] = 32'h80009deb;
