module cust_rom (clk0,
    cs0,
    addr0,
    dout0);
 input clk0;
 input cs0;
 input [7:0] addr0;
 output [31:0] dout0;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire \addr0_reg[0] ;
 wire \addr0_reg[1] ;
 wire \addr0_reg[2] ;
 wire \addr0_reg[3] ;
 wire \addr0_reg[4] ;
 wire \addr0_reg[5] ;
 wire \addr0_reg[6] ;
 wire \addr0_reg[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire clknet_0_clk0;
 wire clknet_2_0__leaf_clk0;
 wire clknet_2_1__leaf_clk0;
 wire clknet_2_2__leaf_clk0;
 wire clknet_2_3__leaf_clk0;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;

 sky130_fd_sc_hd__clkinv_4 _0809_ (.A(net94),
    .Y(_0652_));
 sky130_fd_sc_hd__inv_2 _0810_ (.A(net102),
    .Y(_0662_));
 sky130_fd_sc_hd__inv_2 _0811_ (.A(net103),
    .Y(_0673_));
 sky130_fd_sc_hd__inv_2 _0812_ (.A(net118),
    .Y(_0683_));
 sky130_fd_sc_hd__inv_2 _0813_ (.A(net133),
    .Y(_0694_));
 sky130_fd_sc_hd__inv_2 _0814_ (.A(net144),
    .Y(_0704_));
 sky130_fd_sc_hd__inv_2 _0815_ (.A(net169),
    .Y(_0715_));
 sky130_fd_sc_hd__inv_2 _0816_ (.A(net175),
    .Y(_0725_));
 sky130_fd_sc_hd__and2_2 _0817_ (.A(net156),
    .B(net164),
    .X(_0736_));
 sky130_fd_sc_hd__nand2_1 _0818_ (.A(net156),
    .B(net164),
    .Y(_0746_));
 sky130_fd_sc_hd__nor2_4 _0819_ (.A(net153),
    .B(net162),
    .Y(_0757_));
 sky130_fd_sc_hd__xor2_2 _0820_ (.A(net160),
    .B(net167),
    .X(_0767_));
 sky130_fd_sc_hd__xnor2_2 _0821_ (.A(net153),
    .B(net162),
    .Y(_0777_));
 sky130_fd_sc_hd__and2b_1 _0822_ (.A_N(net158),
    .B(net165),
    .X(_0787_));
 sky130_fd_sc_hd__nand2b_4 _0823_ (.A_N(net158),
    .B(net165),
    .Y(_0796_));
 sky130_fd_sc_hd__and2b_2 _0824_ (.A_N(net153),
    .B(net144),
    .X(_0798_));
 sky130_fd_sc_hd__nand2b_1 _0825_ (.A_N(net160),
    .B(net150),
    .Y(_0799_));
 sky130_fd_sc_hd__nand2_4 _0826_ (.A(net148),
    .B(net165),
    .Y(_0800_));
 sky130_fd_sc_hd__and2b_4 _0827_ (.A_N(net162),
    .B(net153),
    .X(_0801_));
 sky130_fd_sc_hd__nand2b_2 _0828_ (.A_N(net163),
    .B(net155),
    .Y(_0802_));
 sky130_fd_sc_hd__nand2_1 _0829_ (.A(net65),
    .B(_0800_),
    .Y(_0803_));
 sky130_fd_sc_hd__nand2_4 _0830_ (.A(net133),
    .B(_0796_),
    .Y(_0804_));
 sky130_fd_sc_hd__and3_2 _0831_ (.A(net137),
    .B(net146),
    .C(net67),
    .X(_0805_));
 sky130_fd_sc_hd__or3_2 _0832_ (.A(net73),
    .B(_0704_),
    .C(net69),
    .X(_0806_));
 sky130_fd_sc_hd__o21a_2 _0833_ (.A1(net156),
    .A2(net164),
    .B1(net137),
    .X(_0807_));
 sky130_fd_sc_hd__o21ai_4 _0834_ (.A1(net161),
    .A2(net168),
    .B1(net140),
    .Y(_0808_));
 sky130_fd_sc_hd__and2b_1 _0835_ (.A_N(net147),
    .B(net164),
    .X(_0032_));
 sky130_fd_sc_hd__nand2b_2 _0836_ (.A_N(net146),
    .B(net164),
    .Y(_0033_));
 sky130_fd_sc_hd__and2b_1 _0837_ (.A_N(net144),
    .B(net153),
    .X(_0034_));
 sky130_fd_sc_hd__nand2b_1 _0838_ (.A_N(net144),
    .B(net154),
    .Y(_0035_));
 sky130_fd_sc_hd__nand2b_1 _0839_ (.A_N(net148),
    .B(net133),
    .Y(_0036_));
 sky130_fd_sc_hd__nor2_2 _0840_ (.A(net147),
    .B(_0808_),
    .Y(_0037_));
 sky130_fd_sc_hd__nand2_1 _0841_ (.A(_0704_),
    .B(_0807_),
    .Y(_0038_));
 sky130_fd_sc_hd__nand2_1 _0842_ (.A(net72),
    .B(net65),
    .Y(_0039_));
 sky130_fd_sc_hd__and2b_4 _0843_ (.A_N(net139),
    .B(net167),
    .X(_0040_));
 sky130_fd_sc_hd__nand2b_2 _0844_ (.A_N(net141),
    .B(net168),
    .Y(_0041_));
 sky130_fd_sc_hd__nand2_1 _0845_ (.A(net65),
    .B(_0040_),
    .Y(_0042_));
 sky130_fd_sc_hd__nor2_2 _0846_ (.A(net140),
    .B(net160),
    .Y(_0043_));
 sky130_fd_sc_hd__or2_4 _0847_ (.A(net139),
    .B(net160),
    .X(_0044_));
 sky130_fd_sc_hd__nor2_4 _0848_ (.A(net133),
    .B(net148),
    .Y(_0045_));
 sky130_fd_sc_hd__or2_4 _0849_ (.A(net138),
    .B(net146),
    .X(_0046_));
 sky130_fd_sc_hd__nor2_1 _0850_ (.A(net147),
    .B(_0044_),
    .Y(_0047_));
 sky130_fd_sc_hd__or3_2 _0851_ (.A(net137),
    .B(net146),
    .C(net156),
    .X(_0048_));
 sky130_fd_sc_hd__nand2_2 _0852_ (.A(net123),
    .B(_0042_),
    .Y(_0049_));
 sky130_fd_sc_hd__nor2_2 _0853_ (.A(net131),
    .B(_0801_),
    .Y(_0050_));
 sky130_fd_sc_hd__or3_1 _0854_ (.A(net130),
    .B(_0798_),
    .C(_0801_),
    .X(_0051_));
 sky130_fd_sc_hd__or4b_1 _0855_ (.A(net74),
    .B(_0805_),
    .C(_0037_),
    .D_N(_0051_),
    .X(_0052_));
 sky130_fd_sc_hd__nor2_1 _0856_ (.A(net86),
    .B(net82),
    .Y(_0053_));
 sky130_fd_sc_hd__nand2_1 _0857_ (.A(net107),
    .B(net118),
    .Y(_0054_));
 sky130_fd_sc_hd__a21bo_4 _0858_ (.A1(net148),
    .A2(net165),
    .B1_N(net133),
    .X(_0055_));
 sky130_fd_sc_hd__nand2_1 _0859_ (.A(net71),
    .B(_0035_),
    .Y(_0056_));
 sky130_fd_sc_hd__nor2_2 _0860_ (.A(net138),
    .B(net61),
    .Y(_0057_));
 sky130_fd_sc_hd__nor2_1 _0861_ (.A(net150),
    .B(net167),
    .Y(_0058_));
 sky130_fd_sc_hd__or2_2 _0862_ (.A(net144),
    .B(net162),
    .X(_0059_));
 sky130_fd_sc_hd__xor2_2 _0863_ (.A(net144),
    .B(net162),
    .X(_0060_));
 sky130_fd_sc_hd__xnor2_1 _0864_ (.A(net144),
    .B(net162),
    .Y(_0061_));
 sky130_fd_sc_hd__and3_1 _0865_ (.A(net71),
    .B(_0035_),
    .C(_0059_),
    .X(_0062_));
 sky130_fd_sc_hd__or3_2 _0866_ (.A(net130),
    .B(net60),
    .C(net51),
    .X(_0063_));
 sky130_fd_sc_hd__nand2_1 _0867_ (.A(net132),
    .B(net60),
    .Y(_0064_));
 sky130_fd_sc_hd__nand2_4 _0868_ (.A(net132),
    .B(_0801_),
    .Y(_0065_));
 sky130_fd_sc_hd__a31o_1 _0869_ (.A1(_0063_),
    .A2(_0064_),
    .A3(_0065_),
    .B1(net116),
    .X(_0066_));
 sky130_fd_sc_hd__and2_2 _0870_ (.A(net145),
    .B(net155),
    .X(_0067_));
 sky130_fd_sc_hd__nand2_4 _0871_ (.A(net148),
    .B(net158),
    .Y(_0068_));
 sky130_fd_sc_hd__xor2_4 _0872_ (.A(net144),
    .B(net153),
    .X(_0069_));
 sky130_fd_sc_hd__xnor2_1 _0873_ (.A(net144),
    .B(net153),
    .Y(_0070_));
 sky130_fd_sc_hd__nand2_2 _0874_ (.A(net162),
    .B(net48),
    .Y(_0071_));
 sky130_fd_sc_hd__and2b_4 _0875_ (.A_N(net163),
    .B(net145),
    .X(_0072_));
 sky130_fd_sc_hd__nand2b_1 _0876_ (.A_N(net167),
    .B(net150),
    .Y(_0073_));
 sky130_fd_sc_hd__nor2_1 _0877_ (.A(net135),
    .B(_0072_),
    .Y(_0074_));
 sky130_fd_sc_hd__nand2_4 _0878_ (.A(net139),
    .B(net65),
    .Y(_0075_));
 sky130_fd_sc_hd__or3_1 _0879_ (.A(net71),
    .B(net66),
    .C(_0798_),
    .X(_0076_));
 sky130_fd_sc_hd__a21boi_1 _0880_ (.A1(_0071_),
    .A2(_0074_),
    .B1_N(_0076_),
    .Y(_0077_));
 sky130_fd_sc_hd__nand2_2 _0881_ (.A(net154),
    .B(net51),
    .Y(_0078_));
 sky130_fd_sc_hd__a21oi_1 _0882_ (.A1(net155),
    .A2(net51),
    .B1(net131),
    .Y(_0079_));
 sky130_fd_sc_hd__nand2_1 _0883_ (.A(net120),
    .B(_0055_),
    .Y(_0080_));
 sky130_fd_sc_hd__o221a_1 _0884_ (.A1(net121),
    .A2(_0077_),
    .B1(_0079_),
    .B2(_0080_),
    .C1(net84),
    .X(_0081_));
 sky130_fd_sc_hd__a311o_1 _0885_ (.A1(net103),
    .A2(_0052_),
    .A3(_0066_),
    .B1(_0081_),
    .C1(net97),
    .X(_0082_));
 sky130_fd_sc_hd__and2b_1 _0886_ (.A_N(net158),
    .B(net133),
    .X(_0083_));
 sky130_fd_sc_hd__or2_1 _0887_ (.A(net72),
    .B(net158),
    .X(_0084_));
 sky130_fd_sc_hd__and2_2 _0888_ (.A(net133),
    .B(net165),
    .X(_0085_));
 sky130_fd_sc_hd__nand2_4 _0889_ (.A(net139),
    .B(net167),
    .Y(_0086_));
 sky130_fd_sc_hd__or2_1 _0890_ (.A(_0055_),
    .B(net56),
    .X(_0087_));
 sky130_fd_sc_hd__nand2_1 _0891_ (.A(net53),
    .B(net46),
    .Y(_0088_));
 sky130_fd_sc_hd__a221o_1 _0892_ (.A1(net64),
    .A2(net46),
    .B1(_0088_),
    .B2(_0071_),
    .C1(net115),
    .X(_0089_));
 sky130_fd_sc_hd__nand2_1 _0893_ (.A(net66),
    .B(_0045_),
    .Y(_0090_));
 sky130_fd_sc_hd__a221o_1 _0894_ (.A1(net66),
    .A2(_0045_),
    .B1(_0048_),
    .B2(net51),
    .C1(net78),
    .X(_0091_));
 sky130_fd_sc_hd__nor2_1 _0895_ (.A(net88),
    .B(net83),
    .Y(_0092_));
 sky130_fd_sc_hd__nand2_4 _0896_ (.A(net102),
    .B(net113),
    .Y(_0093_));
 sky130_fd_sc_hd__a21o_1 _0897_ (.A1(_0089_),
    .A2(_0091_),
    .B1(_0093_),
    .X(_0094_));
 sky130_fd_sc_hd__o21a_2 _0898_ (.A1(net145),
    .A2(net154),
    .B1(net70),
    .X(_0095_));
 sky130_fd_sc_hd__o21bai_2 _0899_ (.A1(net150),
    .A2(net160),
    .B1_N(net139),
    .Y(_0096_));
 sky130_fd_sc_hd__nand2_1 _0900_ (.A(net124),
    .B(_0073_),
    .Y(_0097_));
 sky130_fd_sc_hd__nor2_1 _0901_ (.A(net137),
    .B(net48),
    .Y(_0098_));
 sky130_fd_sc_hd__a21oi_2 _0902_ (.A1(net54),
    .A2(_0098_),
    .B1(net77),
    .Y(_0099_));
 sky130_fd_sc_hd__o21a_1 _0903_ (.A1(net53),
    .A2(_0095_),
    .B1(_0099_),
    .X(_0100_));
 sky130_fd_sc_hd__a21oi_4 _0904_ (.A1(net156),
    .A2(net164),
    .B1(net146),
    .Y(_0101_));
 sky130_fd_sc_hd__nor2_2 _0905_ (.A(_0736_),
    .B(net59),
    .Y(_0102_));
 sky130_fd_sc_hd__nor3b_2 _0906_ (.A(net157),
    .B(net164),
    .C_N(net146),
    .Y(_0103_));
 sky130_fd_sc_hd__or3b_1 _0907_ (.A(net156),
    .B(net164),
    .C_N(net146),
    .X(_0104_));
 sky130_fd_sc_hd__o21ai_2 _0908_ (.A1(_0101_),
    .A2(_0103_),
    .B1(net132),
    .Y(_0105_));
 sky130_fd_sc_hd__o21a_1 _0909_ (.A1(_0101_),
    .A2(_0103_),
    .B1(net138),
    .X(_0106_));
 sky130_fd_sc_hd__a21oi_2 _0910_ (.A1(net146),
    .A2(net164),
    .B1(net137),
    .Y(_0107_));
 sky130_fd_sc_hd__a21o_1 _0911_ (.A1(net144),
    .A2(net162),
    .B1(net130),
    .X(_0108_));
 sky130_fd_sc_hd__o211a_1 _0912_ (.A1(net50),
    .A2(_0108_),
    .B1(_0105_),
    .C1(net74),
    .X(_0109_));
 sky130_fd_sc_hd__nand2_2 _0913_ (.A(net98),
    .B(net85),
    .Y(_0110_));
 sky130_fd_sc_hd__o311a_1 _0914_ (.A1(_0100_),
    .A2(_0109_),
    .A3(_0110_),
    .B1(_0094_),
    .C1(net173),
    .X(_0111_));
 sky130_fd_sc_hd__nand2_2 _0915_ (.A(net73),
    .B(net62),
    .Y(_0112_));
 sky130_fd_sc_hd__nor2_1 _0916_ (.A(net134),
    .B(net53),
    .Y(_0113_));
 sky130_fd_sc_hd__o2bb2a_1 _0917_ (.A1_N(_0082_),
    .A2_N(_0111_),
    .B1(net202),
    .B2(net173),
    .X(_0000_));
 sky130_fd_sc_hd__a21bo_4 _0918_ (.A1(net153),
    .A2(net162),
    .B1_N(net130),
    .X(_0114_));
 sky130_fd_sc_hd__or2_1 _0919_ (.A(net60),
    .B(_0114_),
    .X(_0115_));
 sky130_fd_sc_hd__or3_2 _0920_ (.A(net60),
    .B(_0103_),
    .C(_0114_),
    .X(_0116_));
 sky130_fd_sc_hd__nor2_2 _0921_ (.A(_0715_),
    .B(net48),
    .Y(_0117_));
 sky130_fd_sc_hd__nor3_2 _0922_ (.A(net148),
    .B(net158),
    .C(net165),
    .Y(_0118_));
 sky130_fd_sc_hd__a211o_2 _0923_ (.A1(net165),
    .A2(net50),
    .B1(_0118_),
    .C1(net133),
    .X(_0119_));
 sky130_fd_sc_hd__or3b_2 _0924_ (.A(net151),
    .B(net168),
    .C_N(net157),
    .X(_0120_));
 sky130_fd_sc_hd__and4_1 _0925_ (.A(net121),
    .B(_0796_),
    .C(_0075_),
    .D(_0120_),
    .X(_0121_));
 sky130_fd_sc_hd__or3_1 _0926_ (.A(net134),
    .B(_0798_),
    .C(net56),
    .X(_0122_));
 sky130_fd_sc_hd__xnor2_1 _0927_ (.A(net159),
    .B(net53),
    .Y(_0123_));
 sky130_fd_sc_hd__xnor2_4 _0928_ (.A(net153),
    .B(net51),
    .Y(_0124_));
 sky130_fd_sc_hd__o21a_1 _0929_ (.A1(net70),
    .A2(_0123_),
    .B1(_0122_),
    .X(_0125_));
 sky130_fd_sc_hd__nor2_4 _0930_ (.A(net83),
    .B(net123),
    .Y(_0126_));
 sky130_fd_sc_hd__nand2_4 _0931_ (.A(net112),
    .B(net81),
    .Y(_0127_));
 sky130_fd_sc_hd__o21a_2 _0932_ (.A1(net146),
    .A2(net157),
    .B1(net138),
    .X(_0128_));
 sky130_fd_sc_hd__o21ai_4 _0933_ (.A1(net147),
    .A2(net157),
    .B1(net138),
    .Y(_0129_));
 sky130_fd_sc_hd__nor2_1 _0934_ (.A(_0715_),
    .B(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__or2_1 _0935_ (.A(net79),
    .B(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__and3_1 _0936_ (.A(net70),
    .B(net149),
    .C(_0802_),
    .X(_0132_));
 sky130_fd_sc_hd__o221a_1 _0937_ (.A1(net121),
    .A2(_0125_),
    .B1(_0131_),
    .B2(_0132_),
    .C1(net109),
    .X(_0133_));
 sky130_fd_sc_hd__a31o_1 _0938_ (.A1(net79),
    .A2(_0116_),
    .A3(_0119_),
    .B1(_0121_),
    .X(_0134_));
 sky130_fd_sc_hd__a211o_1 _0939_ (.A1(net87),
    .A2(_0134_),
    .B1(_0133_),
    .C1(net101),
    .X(_0135_));
 sky130_fd_sc_hd__and3b_1 _0940_ (.A_N(net167),
    .B(net160),
    .C(net151),
    .X(_0136_));
 sky130_fd_sc_hd__or3_2 _0941_ (.A(net140),
    .B(_0118_),
    .C(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__nor2_1 _0942_ (.A(net63),
    .B(_0137_),
    .Y(_0138_));
 sky130_fd_sc_hd__nor2_2 _0943_ (.A(net148),
    .B(net68),
    .Y(_0139_));
 sky130_fd_sc_hd__a21o_1 _0944_ (.A1(_0704_),
    .A2(net69),
    .B1(_0072_),
    .X(_0140_));
 sky130_fd_sc_hd__o211a_1 _0945_ (.A1(net150),
    .A2(net67),
    .B1(_0073_),
    .C1(net135),
    .X(_0141_));
 sky130_fd_sc_hd__nor2_1 _0946_ (.A(net67),
    .B(net59),
    .Y(_0142_));
 sky130_fd_sc_hd__or3b_2 _0947_ (.A(net136),
    .B(net63),
    .C_N(net156),
    .X(_0143_));
 sky130_fd_sc_hd__or2_1 _0948_ (.A(net135),
    .B(_0078_),
    .X(_0144_));
 sky130_fd_sc_hd__nor2_1 _0949_ (.A(net131),
    .B(net66),
    .Y(_0145_));
 sky130_fd_sc_hd__or3_1 _0950_ (.A(net132),
    .B(net66),
    .C(net48),
    .X(_0146_));
 sky130_fd_sc_hd__o211a_1 _0951_ (.A1(net56),
    .A2(_0075_),
    .B1(_0146_),
    .C1(net121),
    .X(_0147_));
 sky130_fd_sc_hd__a311o_1 _0952_ (.A1(net79),
    .A2(_0076_),
    .A3(_0144_),
    .B1(_0147_),
    .C1(net84),
    .X(_0148_));
 sky130_fd_sc_hd__o211a_1 _0953_ (.A1(net68),
    .A2(net59),
    .B1(_0042_),
    .C1(net80),
    .X(_0149_));
 sky130_fd_sc_hd__o21a_1 _0954_ (.A1(_0138_),
    .A2(_0141_),
    .B1(net124),
    .X(_0150_));
 sky130_fd_sc_hd__o311a_1 _0955_ (.A1(net109),
    .A2(_0149_),
    .A3(_0150_),
    .B1(_0148_),
    .C1(net101),
    .X(_0151_));
 sky130_fd_sc_hd__or3b_1 _0956_ (.A(net93),
    .B(_0151_),
    .C_N(_0135_),
    .X(_0152_));
 sky130_fd_sc_hd__o21a_1 _0957_ (.A1(_0075_),
    .A2(_0139_),
    .B1(_0143_),
    .X(_0153_));
 sky130_fd_sc_hd__a21o_1 _0958_ (.A1(net139),
    .A2(net61),
    .B1(net127),
    .X(_0154_));
 sky130_fd_sc_hd__nor2_1 _0959_ (.A(net61),
    .B(_0041_),
    .Y(_0155_));
 sky130_fd_sc_hd__a31o_1 _0960_ (.A1(net139),
    .A2(_0799_),
    .A3(_0800_),
    .B1(_0155_),
    .X(_0156_));
 sky130_fd_sc_hd__o32a_1 _0961_ (.A1(net167),
    .A2(_0057_),
    .A3(_0154_),
    .B1(_0156_),
    .B2(net82),
    .X(_0157_));
 sky130_fd_sc_hd__o21bai_4 _0962_ (.A1(net159),
    .A2(net165),
    .B1_N(net133),
    .Y(_0158_));
 sky130_fd_sc_hd__a211o_1 _0963_ (.A1(net54),
    .A2(_0158_),
    .B1(_0127_),
    .C1(_0736_),
    .X(_0159_));
 sky130_fd_sc_hd__nor2_1 _0964_ (.A(net132),
    .B(net68),
    .Y(_0160_));
 sky130_fd_sc_hd__nand2_1 _0965_ (.A(net72),
    .B(net69),
    .Y(_0161_));
 sky130_fd_sc_hd__o211a_1 _0966_ (.A1(net57),
    .A2(_0153_),
    .B1(_0159_),
    .C1(net88),
    .X(_0162_));
 sky130_fd_sc_hd__o21a_1 _0967_ (.A1(net113),
    .A2(_0157_),
    .B1(_0162_),
    .X(_0163_));
 sky130_fd_sc_hd__nand2_2 _0968_ (.A(net94),
    .B(net88),
    .Y(_0164_));
 sky130_fd_sc_hd__nand2_2 _0969_ (.A(net71),
    .B(_0757_),
    .Y(_0165_));
 sky130_fd_sc_hd__or2_1 _0970_ (.A(net142),
    .B(_0139_),
    .X(_0166_));
 sky130_fd_sc_hd__o221a_1 _0971_ (.A1(net166),
    .A2(_0084_),
    .B1(_0139_),
    .B2(_0039_),
    .C1(net80),
    .X(_0167_));
 sky130_fd_sc_hd__o21a_1 _0972_ (.A1(net61),
    .A2(_0113_),
    .B1(net123),
    .X(_0168_));
 sky130_fd_sc_hd__o21a_1 _0973_ (.A1(_0167_),
    .A2(_0168_),
    .B1(net83),
    .X(_0169_));
 sky130_fd_sc_hd__o211a_1 _0974_ (.A1(net165),
    .A2(_0039_),
    .B1(net42),
    .C1(_0806_),
    .X(_0170_));
 sky130_fd_sc_hd__or2_1 _0975_ (.A(net66),
    .B(_0055_),
    .X(_0171_));
 sky130_fd_sc_hd__o211a_1 _0976_ (.A1(net68),
    .A2(_0046_),
    .B1(_0126_),
    .C1(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__o31a_1 _0977_ (.A1(_0169_),
    .A2(_0170_),
    .A3(_0172_),
    .B1(net101),
    .X(_0173_));
 sky130_fd_sc_hd__o31a_1 _0978_ (.A1(_0652_),
    .A2(_0163_),
    .A3(_0173_),
    .B1(net176),
    .X(_0174_));
 sky130_fd_sc_hd__a22o_1 _0979_ (.A1(net171),
    .A2(net200),
    .B1(_0152_),
    .B2(_0174_),
    .X(_0001_));
 sky130_fd_sc_hd__nor2_1 _0980_ (.A(net94),
    .B(net102),
    .Y(_0175_));
 sky130_fd_sc_hd__or2_2 _0981_ (.A(net90),
    .B(net98),
    .X(_0176_));
 sky130_fd_sc_hd__or3b_2 _0982_ (.A(net151),
    .B(net160),
    .C_N(net139),
    .X(_0177_));
 sky130_fd_sc_hd__or4_1 _0983_ (.A(net127),
    .B(_0040_),
    .C(_0043_),
    .D(_0045_),
    .X(_0178_));
 sky130_fd_sc_hd__and3b_1 _0984_ (.A_N(_0178_),
    .B(_0177_),
    .C(_0086_),
    .X(_0179_));
 sky130_fd_sc_hd__o311a_1 _0985_ (.A1(net135),
    .A2(_0803_),
    .A3(_0101_),
    .B1(_0806_),
    .C1(net124),
    .X(_0180_));
 sky130_fd_sc_hd__nand2_1 _0986_ (.A(net131),
    .B(_0802_),
    .Y(_0181_));
 sky130_fd_sc_hd__or3_1 _0987_ (.A(net46),
    .B(_0085_),
    .C(_0178_),
    .X(_0182_));
 sky130_fd_sc_hd__and3_4 _0988_ (.A(net149),
    .B(net158),
    .C(net166),
    .X(_0183_));
 sky130_fd_sc_hd__nand3_4 _0989_ (.A(net150),
    .B(net160),
    .C(net167),
    .Y(_0184_));
 sky130_fd_sc_hd__nor2_1 _0990_ (.A(net73),
    .B(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__o31a_2 _0991_ (.A1(net139),
    .A2(net161),
    .A3(net168),
    .B1(net128),
    .X(_0186_));
 sky130_fd_sc_hd__o21ai_1 _0992_ (.A1(net73),
    .A2(_0184_),
    .B1(_0186_),
    .Y(_0187_));
 sky130_fd_sc_hd__nor2_2 _0993_ (.A(net70),
    .B(_0183_),
    .Y(_0188_));
 sky130_fd_sc_hd__o311a_1 _0994_ (.A1(net72),
    .A2(_0118_),
    .A3(_0183_),
    .B1(_0158_),
    .C1(net123),
    .X(_0189_));
 sky130_fd_sc_hd__nand3_4 _0995_ (.A(net135),
    .B(net148),
    .C(net158),
    .Y(_0190_));
 sky130_fd_sc_hd__and3_1 _0996_ (.A(net80),
    .B(_0065_),
    .C(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__a221o_1 _0997_ (.A1(net65),
    .A2(_0807_),
    .B1(_0059_),
    .B2(_0160_),
    .C1(net115),
    .X(_0192_));
 sky130_fd_sc_hd__nand2_1 _0998_ (.A(_0131_),
    .B(_0192_),
    .Y(_0193_));
 sky130_fd_sc_hd__o31a_1 _0999_ (.A1(net83),
    .A2(_0189_),
    .A3(_0191_),
    .B1(net93),
    .X(_0194_));
 sky130_fd_sc_hd__o21ai_1 _1000_ (.A1(net110),
    .A2(_0193_),
    .B1(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__nor2_1 _1001_ (.A(_0114_),
    .B(_0118_),
    .Y(_0196_));
 sky130_fd_sc_hd__o31a_1 _1002_ (.A1(_0040_),
    .A2(_0057_),
    .A3(_0196_),
    .B1(_0126_),
    .X(_0197_));
 sky130_fd_sc_hd__or3_1 _1003_ (.A(net141),
    .B(net168),
    .C(_0067_),
    .X(_0198_));
 sky130_fd_sc_hd__nand2_1 _1004_ (.A(net55),
    .B(net47),
    .Y(_0199_));
 sky130_fd_sc_hd__nand2_1 _1005_ (.A(_0198_),
    .B(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__a21o_1 _1006_ (.A1(_0767_),
    .A2(net54),
    .B1(net140),
    .X(_0201_));
 sky130_fd_sc_hd__nand2_2 _1007_ (.A(net137),
    .B(net55),
    .Y(_0202_));
 sky130_fd_sc_hd__nand2_1 _1008_ (.A(net128),
    .B(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__nor2_1 _1009_ (.A(net128),
    .B(net55),
    .Y(_0204_));
 sky130_fd_sc_hd__nor2_1 _1010_ (.A(net55),
    .B(_0158_),
    .Y(_0205_));
 sky130_fd_sc_hd__a21o_1 _1011_ (.A1(_0799_),
    .A2(_0807_),
    .B1(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__a31o_1 _1012_ (.A1(net127),
    .A2(_0201_),
    .A3(_0202_),
    .B1(net111),
    .X(_0207_));
 sky130_fd_sc_hd__a21oi_1 _1013_ (.A1(net81),
    .A2(_0206_),
    .B1(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__a2111o_1 _1014_ (.A1(net42),
    .A2(_0200_),
    .B1(_0208_),
    .C1(_0197_),
    .D1(net95),
    .X(_0209_));
 sky130_fd_sc_hd__nand2_1 _1015_ (.A(_0050_),
    .B(_0071_),
    .Y(_0210_));
 sky130_fd_sc_hd__or3b_1 _1016_ (.A(net121),
    .B(_0188_),
    .C_N(_0112_),
    .X(_0211_));
 sky130_fd_sc_hd__or2_1 _1017_ (.A(_0055_),
    .B(net44),
    .X(_0212_));
 sky130_fd_sc_hd__nor2_1 _1018_ (.A(_0055_),
    .B(net44),
    .Y(_0213_));
 sky130_fd_sc_hd__a21o_1 _1019_ (.A1(net149),
    .A2(_0145_),
    .B1(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__o21ai_2 _1020_ (.A1(net149),
    .A2(_0796_),
    .B1(_0050_),
    .Y(_0215_));
 sky130_fd_sc_hd__and3_1 _1021_ (.A(net126),
    .B(_0086_),
    .C(_0177_),
    .X(_0216_));
 sky130_fd_sc_hd__a21oi_1 _1022_ (.A1(_0182_),
    .A2(_0187_),
    .B1(net110),
    .Y(_0217_));
 sky130_fd_sc_hd__o21a_1 _1023_ (.A1(_0084_),
    .A2(_0097_),
    .B1(net110),
    .X(_0218_));
 sky130_fd_sc_hd__o211a_1 _1024_ (.A1(net80),
    .A2(_0210_),
    .B1(_0211_),
    .C1(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__a221o_1 _1025_ (.A1(net80),
    .A2(_0214_),
    .B1(_0215_),
    .B2(_0216_),
    .C1(net86),
    .X(_0220_));
 sky130_fd_sc_hd__o311a_1 _1026_ (.A1(net113),
    .A2(_0179_),
    .A3(_0180_),
    .B1(_0220_),
    .C1(_0175_),
    .X(_0221_));
 sky130_fd_sc_hd__o31ai_1 _1027_ (.A1(_0164_),
    .A2(_0217_),
    .A3(_0219_),
    .B1(net176),
    .Y(_0222_));
 sky130_fd_sc_hd__a31o_1 _1028_ (.A1(net101),
    .A2(_0195_),
    .A3(_0209_),
    .B1(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__o22a_1 _1029_ (.A1(net176),
    .A2(net178),
    .B1(_0221_),
    .B2(_0223_),
    .X(_0002_));
 sky130_fd_sc_hd__nand2_1 _1030_ (.A(net142),
    .B(net62),
    .Y(_0224_));
 sky130_fd_sc_hd__a21oi_1 _1031_ (.A1(net62),
    .A2(_0051_),
    .B1(net116),
    .Y(_0225_));
 sky130_fd_sc_hd__nand2_4 _1032_ (.A(net137),
    .B(net50),
    .Y(_0226_));
 sky130_fd_sc_hd__or2_1 _1033_ (.A(net164),
    .B(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__a21o_1 _1034_ (.A1(_0068_),
    .A2(_0140_),
    .B1(net132),
    .X(_0228_));
 sky130_fd_sc_hd__a311o_1 _1035_ (.A1(net116),
    .A2(_0227_),
    .A3(_0228_),
    .B1(_0225_),
    .C1(net103),
    .X(_0229_));
 sky130_fd_sc_hd__nor2_1 _1036_ (.A(net159),
    .B(net53),
    .Y(_0230_));
 sky130_fd_sc_hd__o2bb2a_1 _1037_ (.A1_N(_0078_),
    .A2_N(_0128_),
    .B1(_0230_),
    .B2(net135),
    .X(_0231_));
 sky130_fd_sc_hd__nor2_1 _1038_ (.A(net66),
    .B(net59),
    .Y(_0232_));
 sky130_fd_sc_hd__or2_1 _1039_ (.A(_0787_),
    .B(net59),
    .X(_0233_));
 sky130_fd_sc_hd__o22a_2 _1040_ (.A1(net66),
    .A2(_0036_),
    .B1(_0129_),
    .B2(net67),
    .X(_0234_));
 sky130_fd_sc_hd__o21a_1 _1041_ (.A1(_0800_),
    .A2(_0044_),
    .B1(net122),
    .X(_0235_));
 sky130_fd_sc_hd__a221o_1 _1042_ (.A1(net79),
    .A2(_0231_),
    .B1(_0234_),
    .B2(_0235_),
    .C1(net83),
    .X(_0236_));
 sky130_fd_sc_hd__a21oi_1 _1043_ (.A1(_0229_),
    .A2(_0236_),
    .B1(_0176_),
    .Y(_0237_));
 sky130_fd_sc_hd__a21o_1 _1044_ (.A1(_0746_),
    .A2(_0107_),
    .B1(net77),
    .X(_0238_));
 sky130_fd_sc_hd__and3b_2 _1045_ (.A_N(net148),
    .B(net158),
    .C(net166),
    .X(_0239_));
 sky130_fd_sc_hd__nand2_1 _1046_ (.A(net136),
    .B(net67),
    .Y(_0240_));
 sky130_fd_sc_hd__nand2_1 _1047_ (.A(net151),
    .B(net69),
    .Y(_0241_));
 sky130_fd_sc_hd__a21o_2 _1048_ (.A1(net151),
    .A2(net69),
    .B1(net73),
    .X(_0242_));
 sky130_fd_sc_hd__nor2_1 _1049_ (.A(_0805_),
    .B(_0102_),
    .Y(_0243_));
 sky130_fd_sc_hd__or3_1 _1050_ (.A(_0805_),
    .B(_0102_),
    .C(_0238_),
    .X(_0244_));
 sky130_fd_sc_hd__nand2_1 _1051_ (.A(_0046_),
    .B(_0158_),
    .Y(_0245_));
 sky130_fd_sc_hd__or3_4 _1052_ (.A(net137),
    .B(net45),
    .C(_0183_),
    .X(_0246_));
 sky130_fd_sc_hd__a31o_1 _1053_ (.A1(_0202_),
    .A2(_0226_),
    .A3(_0246_),
    .B1(net118),
    .X(_0247_));
 sky130_fd_sc_hd__a21oi_1 _1054_ (.A1(net150),
    .A2(net67),
    .B1(net55),
    .Y(_0248_));
 sky130_fd_sc_hd__a211o_2 _1055_ (.A1(net150),
    .A2(net69),
    .B1(net63),
    .C1(_0096_),
    .X(_0249_));
 sky130_fd_sc_hd__inv_2 _1056_ (.A(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__and3_1 _1057_ (.A(net138),
    .B(net65),
    .C(_0120_),
    .X(_0251_));
 sky130_fd_sc_hd__o32a_1 _1058_ (.A1(net118),
    .A2(_0250_),
    .A3(_0251_),
    .B1(_0106_),
    .B2(_0238_),
    .X(_0252_));
 sky130_fd_sc_hd__a31o_1 _1059_ (.A1(net90),
    .A2(_0244_),
    .A3(_0247_),
    .B1(_0093_),
    .X(_0253_));
 sky130_fd_sc_hd__o21ba_1 _1060_ (.A1(net90),
    .A2(_0252_),
    .B1_N(_0253_),
    .X(_0254_));
 sky130_fd_sc_hd__a211o_1 _1061_ (.A1(_0796_),
    .A2(_0078_),
    .B1(_0040_),
    .C1(net115),
    .X(_0255_));
 sky130_fd_sc_hd__nor2_1 _1062_ (.A(net168),
    .B(_0075_),
    .Y(_0256_));
 sky130_fd_sc_hd__or3b_1 _1063_ (.A(_0256_),
    .B(net81),
    .C_N(_0800_),
    .X(_0257_));
 sky130_fd_sc_hd__nor2_1 _1064_ (.A(_0108_),
    .B(net44),
    .Y(_0258_));
 sky130_fd_sc_hd__a21o_1 _1065_ (.A1(net131),
    .A2(_0120_),
    .B1(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__a211oi_1 _1066_ (.A1(net119),
    .A2(_0259_),
    .B1(_0225_),
    .C1(net105),
    .Y(_0260_));
 sky130_fd_sc_hd__a311o_1 _1067_ (.A1(net105),
    .A2(_0255_),
    .A3(_0257_),
    .B1(_0260_),
    .C1(_0164_),
    .X(_0261_));
 sky130_fd_sc_hd__nor2_1 _1068_ (.A(_0039_),
    .B(_0072_),
    .Y(_0262_));
 sky130_fd_sc_hd__or3b_1 _1069_ (.A(_0262_),
    .B(_0203_),
    .C_N(_0226_),
    .X(_0263_));
 sky130_fd_sc_hd__a221o_1 _1070_ (.A1(net63),
    .A2(net46),
    .B1(_0107_),
    .B2(_0120_),
    .C1(net119),
    .X(_0264_));
 sky130_fd_sc_hd__a21o_1 _1071_ (.A1(_0043_),
    .A2(_0059_),
    .B1(net75),
    .X(_0265_));
 sky130_fd_sc_hd__nor2_1 _1072_ (.A(net64),
    .B(_0145_),
    .Y(_0266_));
 sky130_fd_sc_hd__o32a_1 _1073_ (.A1(net115),
    .A2(net60),
    .A3(_0266_),
    .B1(_0265_),
    .B2(_0805_),
    .X(_0267_));
 sky130_fd_sc_hd__nor2_1 _1074_ (.A(_0652_),
    .B(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__a21oi_1 _1075_ (.A1(_0263_),
    .A2(_0264_),
    .B1(net91),
    .Y(_0269_));
 sky130_fd_sc_hd__o311ai_2 _1076_ (.A1(_0110_),
    .A2(_0268_),
    .A3(_0269_),
    .B1(_0261_),
    .C1(net173),
    .Y(_0270_));
 sky130_fd_sc_hd__o32a_1 _1077_ (.A1(_0237_),
    .A2(_0254_),
    .A3(_0270_),
    .B1(net185),
    .B2(net173),
    .X(_0003_));
 sky130_fd_sc_hd__o21ai_1 _1078_ (.A1(net153),
    .A2(net53),
    .B1(_0068_),
    .Y(_0271_));
 sky130_fd_sc_hd__o211a_1 _1079_ (.A1(net156),
    .A2(net54),
    .B1(_0068_),
    .C1(net136),
    .X(_0272_));
 sky130_fd_sc_hd__a21o_1 _1080_ (.A1(net62),
    .A2(_0095_),
    .B1(net85),
    .X(_0273_));
 sky130_fd_sc_hd__o21a_1 _1081_ (.A1(_0272_),
    .A2(_0273_),
    .B1(net57),
    .X(_0274_));
 sky130_fd_sc_hd__o31a_1 _1082_ (.A1(_0801_),
    .A2(_0804_),
    .A3(_0067_),
    .B1(_0099_),
    .X(_0275_));
 sky130_fd_sc_hd__nand2_2 _1083_ (.A(_0802_),
    .B(_0107_),
    .Y(_0276_));
 sky130_fd_sc_hd__nand2_2 _1084_ (.A(net141),
    .B(net69),
    .Y(_0277_));
 sky130_fd_sc_hd__a21o_1 _1085_ (.A1(net147),
    .A2(net67),
    .B1(_0129_),
    .X(_0278_));
 sky130_fd_sc_hd__or3_1 _1086_ (.A(net70),
    .B(net60),
    .C(_0072_),
    .X(_0279_));
 sky130_fd_sc_hd__a41o_1 _1087_ (.A1(net117),
    .A2(_0190_),
    .A3(_0246_),
    .A4(_0279_),
    .B1(net108),
    .X(_0280_));
 sky130_fd_sc_hd__a31o_1 _1088_ (.A1(net78),
    .A2(_0276_),
    .A3(_0278_),
    .B1(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__o21ai_1 _1089_ (.A1(_0274_),
    .A2(_0275_),
    .B1(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__a21oi_1 _1090_ (.A1(_0046_),
    .A2(_0158_),
    .B1(_0239_),
    .Y(_0283_));
 sky130_fd_sc_hd__or3_1 _1091_ (.A(net143),
    .B(net45),
    .C(_0239_),
    .X(_0284_));
 sky130_fd_sc_hd__a21oi_1 _1092_ (.A1(_0277_),
    .A2(_0284_),
    .B1(net77),
    .Y(_0285_));
 sky130_fd_sc_hd__a2bb2o_1 _1093_ (.A1_N(_0034_),
    .A2_N(_0242_),
    .B1(_0095_),
    .B2(net69),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _1094_ (.A0(_0214_),
    .A1(_0286_),
    .S(net74),
    .X(_0287_));
 sky130_fd_sc_hd__o221a_1 _1095_ (.A1(_0274_),
    .A2(_0285_),
    .B1(_0287_),
    .B2(net108),
    .C1(net91),
    .X(_0288_));
 sky130_fd_sc_hd__a211o_1 _1096_ (.A1(_0652_),
    .A2(_0282_),
    .B1(_0288_),
    .C1(net89),
    .X(_0289_));
 sky130_fd_sc_hd__or4_4 _1097_ (.A(net136),
    .B(_0736_),
    .C(net60),
    .D(_0103_),
    .X(_0290_));
 sky130_fd_sc_hd__o21ai_4 _1098_ (.A1(_0055_),
    .A2(net56),
    .B1(net75),
    .Y(_0291_));
 sky130_fd_sc_hd__nor2_1 _1099_ (.A(net47),
    .B(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__a32o_1 _1100_ (.A1(net117),
    .A2(_0276_),
    .A3(_0278_),
    .B1(_0290_),
    .B2(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__o21a_1 _1101_ (.A1(_0801_),
    .A2(_0056_),
    .B1(_0115_),
    .X(_0294_));
 sky130_fd_sc_hd__a21o_1 _1102_ (.A1(net48),
    .A2(_0107_),
    .B1(net77),
    .X(_0295_));
 sky130_fd_sc_hd__nor2_1 _1103_ (.A(net55),
    .B(_0129_),
    .Y(_0296_));
 sky130_fd_sc_hd__nor2_1 _1104_ (.A(_0808_),
    .B(_0101_),
    .Y(_0297_));
 sky130_fd_sc_hd__o221a_1 _1105_ (.A1(net119),
    .A2(_0294_),
    .B1(_0295_),
    .B2(_0297_),
    .C1(net86),
    .X(_0298_));
 sky130_fd_sc_hd__o21ai_1 _1106_ (.A1(net86),
    .A2(_0293_),
    .B1(_0175_),
    .Y(_0299_));
 sky130_fd_sc_hd__o221a_1 _1107_ (.A1(net160),
    .A2(_0055_),
    .B1(_0096_),
    .B2(_0777_),
    .C1(net128),
    .X(_0300_));
 sky130_fd_sc_hd__a31o_1 _1108_ (.A1(_0184_),
    .A2(_0201_),
    .A3(_0204_),
    .B1(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__a21oi_1 _1109_ (.A1(net113),
    .A2(_0301_),
    .B1(_0298_),
    .Y(_0302_));
 sky130_fd_sc_hd__o221a_1 _1110_ (.A1(_0298_),
    .A2(_0299_),
    .B1(_0302_),
    .B2(_0164_),
    .C1(net175),
    .X(_0303_));
 sky130_fd_sc_hd__a22o_1 _1111_ (.A1(net171),
    .A2(net201),
    .B1(_0289_),
    .B2(_0303_),
    .X(_0004_));
 sky130_fd_sc_hd__or3_2 _1112_ (.A(net134),
    .B(_0072_),
    .C(_0239_),
    .X(_0304_));
 sky130_fd_sc_hd__o31a_1 _1113_ (.A1(net70),
    .A2(_0798_),
    .A3(_0801_),
    .B1(net104),
    .X(_0305_));
 sky130_fd_sc_hd__a21oi_1 _1114_ (.A1(_0304_),
    .A2(_0305_),
    .B1(net42),
    .Y(_0306_));
 sky130_fd_sc_hd__a31o_1 _1115_ (.A1(net122),
    .A2(_0065_),
    .A3(_0144_),
    .B1(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__and2_1 _1116_ (.A(net123),
    .B(net59),
    .X(_0308_));
 sky130_fd_sc_hd__nand2_1 _1117_ (.A(net127),
    .B(net59),
    .Y(_0309_));
 sky130_fd_sc_hd__a31oi_1 _1118_ (.A1(net65),
    .A2(_0078_),
    .A3(_0308_),
    .B1(net109),
    .Y(_0310_));
 sky130_fd_sc_hd__a221o_1 _1119_ (.A1(\addr0_reg[3] ),
    .A2(net52),
    .B1(net46),
    .B2(_0715_),
    .C1(net122),
    .X(_0311_));
 sky130_fd_sc_hd__o21ai_1 _1120_ (.A1(_0262_),
    .A2(_0311_),
    .B1(_0310_),
    .Y(_0312_));
 sky130_fd_sc_hd__a21oi_1 _1121_ (.A1(_0307_),
    .A2(_0312_),
    .B1(net93),
    .Y(_0313_));
 sky130_fd_sc_hd__a41o_1 _1122_ (.A1(net121),
    .A2(_0065_),
    .A3(_0144_),
    .A4(_0190_),
    .B1(_0306_),
    .X(_0314_));
 sky130_fd_sc_hd__o21ai_1 _1123_ (.A1(_0045_),
    .A2(_0311_),
    .B1(_0310_),
    .Y(_0315_));
 sky130_fd_sc_hd__a311o_1 _1124_ (.A1(net93),
    .A2(_0314_),
    .A3(_0315_),
    .B1(net88),
    .C1(_0313_),
    .X(_0316_));
 sky130_fd_sc_hd__o211a_1 _1125_ (.A1(net149),
    .A2(net68),
    .B1(_0073_),
    .C1(net71),
    .X(_0317_));
 sky130_fd_sc_hd__or2_1 _1126_ (.A(net58),
    .B(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__or2_1 _1127_ (.A(_0102_),
    .B(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__a211o_1 _1128_ (.A1(net71),
    .A2(net148),
    .B1(_0040_),
    .C1(_0124_),
    .X(_0320_));
 sky130_fd_sc_hd__nand2_1 _1129_ (.A(_0126_),
    .B(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__or2_1 _1130_ (.A(_0158_),
    .B(_0183_),
    .X(_0322_));
 sky130_fd_sc_hd__nor2_1 _1131_ (.A(net56),
    .B(_0114_),
    .Y(_0323_));
 sky130_fd_sc_hd__o221a_1 _1132_ (.A1(net56),
    .A2(_0114_),
    .B1(_0158_),
    .B2(_0101_),
    .C1(net124),
    .X(_0324_));
 sky130_fd_sc_hd__a41o_1 _1133_ (.A1(net80),
    .A2(_0808_),
    .A3(net59),
    .A4(_0322_),
    .B1(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__nand2_1 _1134_ (.A(net83),
    .B(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__a31o_1 _1135_ (.A1(_0319_),
    .A2(_0321_),
    .A3(_0326_),
    .B1(_0164_),
    .X(_0327_));
 sky130_fd_sc_hd__a21boi_1 _1136_ (.A1(_0078_),
    .A2(_0128_),
    .B1_N(_0119_),
    .Y(_0328_));
 sky130_fd_sc_hd__o2111a_1 _1137_ (.A1(net58),
    .A2(_0328_),
    .B1(_0326_),
    .C1(_0321_),
    .D1(_0175_),
    .X(_0329_));
 sky130_fd_sc_hd__nor2_1 _1138_ (.A(net171),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__a32o_1 _1139_ (.A1(_0316_),
    .A2(_0327_),
    .A3(_0330_),
    .B1(net177),
    .B2(net171),
    .X(_0005_));
 sky130_fd_sc_hd__and2_1 _1140_ (.A(net171),
    .B(net205),
    .X(_0331_));
 sky130_fd_sc_hd__and3_1 _1141_ (.A(net143),
    .B(_0068_),
    .C(_0140_),
    .X(_0332_));
 sky130_fd_sc_hd__o21ba_1 _1142_ (.A1(net146),
    .A2(_0757_),
    .B1_N(_0246_),
    .X(_0333_));
 sky130_fd_sc_hd__or3_1 _1143_ (.A(net78),
    .B(_0332_),
    .C(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__and4b_1 _1144_ (.A_N(net139),
    .B(net151),
    .C(net160),
    .D(net167),
    .X(_0335_));
 sky130_fd_sc_hd__o31a_1 _1145_ (.A1(net127),
    .A2(_0130_),
    .A3(_0335_),
    .B1(net102),
    .X(_0336_));
 sky130_fd_sc_hd__nand2_1 _1146_ (.A(net67),
    .B(_0057_),
    .Y(_0337_));
 sky130_fd_sc_hd__a32o_1 _1147_ (.A1(_0086_),
    .A2(_0226_),
    .A3(_0337_),
    .B1(_0241_),
    .B2(_0204_),
    .X(_0338_));
 sky130_fd_sc_hd__a221o_1 _1148_ (.A1(_0334_),
    .A2(_0336_),
    .B1(_0338_),
    .B2(net88),
    .C1(net111),
    .X(_0339_));
 sky130_fd_sc_hd__o211a_1 _1149_ (.A1(_0044_),
    .A2(net52),
    .B1(_0190_),
    .C1(net127),
    .X(_0340_));
 sky130_fd_sc_hd__a311o_1 _1150_ (.A1(net82),
    .A2(_0065_),
    .A3(_0137_),
    .B1(_0340_),
    .C1(_0093_),
    .X(_0341_));
 sky130_fd_sc_hd__nor2_2 _1151_ (.A(net98),
    .B(net85),
    .Y(_0342_));
 sky130_fd_sc_hd__nand2_4 _1152_ (.A(net89),
    .B(net112),
    .Y(_0343_));
 sky130_fd_sc_hd__nor2_1 _1153_ (.A(net49),
    .B(_0112_),
    .Y(_0344_));
 sky130_fd_sc_hd__nor2_1 _1154_ (.A(net72),
    .B(net50),
    .Y(_0345_));
 sky130_fd_sc_hd__or3_1 _1155_ (.A(net126),
    .B(_0344_),
    .C(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__a21o_1 _1156_ (.A1(_0049_),
    .A2(_0346_),
    .B1(_0343_),
    .X(_0347_));
 sky130_fd_sc_hd__a31o_1 _1157_ (.A1(_0339_),
    .A2(_0341_),
    .A3(_0347_),
    .B1(net95),
    .X(_0348_));
 sky130_fd_sc_hd__a21oi_4 _1158_ (.A1(net72),
    .A2(net63),
    .B1(net81),
    .Y(_0349_));
 sky130_fd_sc_hd__a21boi_1 _1159_ (.A1(_0184_),
    .A2(_0349_),
    .B1_N(_0346_),
    .Y(_0350_));
 sky130_fd_sc_hd__o211a_1 _1160_ (.A1(net150),
    .A2(net161),
    .B1(_0073_),
    .C1(net127),
    .X(_0351_));
 sky130_fd_sc_hd__a211o_1 _1161_ (.A1(_0065_),
    .A2(_0137_),
    .B1(_0351_),
    .C1(_0093_),
    .X(_0352_));
 sky130_fd_sc_hd__o2111ai_1 _1162_ (.A1(_0343_),
    .A2(_0350_),
    .B1(_0352_),
    .C1(_0339_),
    .D1(net95),
    .Y(_0353_));
 sky130_fd_sc_hd__a31o_1 _1163_ (.A1(net175),
    .A2(_0348_),
    .A3(_0353_),
    .B1(_0331_),
    .X(_0006_));
 sky130_fd_sc_hd__a31o_1 _1164_ (.A1(net72),
    .A2(net62),
    .A3(_0104_),
    .B1(net117),
    .X(_0354_));
 sky130_fd_sc_hd__o211a_1 _1165_ (.A1(net45),
    .A2(_0112_),
    .B1(_0234_),
    .C1(net77),
    .X(_0355_));
 sky130_fd_sc_hd__a41o_1 _1166_ (.A1(net119),
    .A2(_0041_),
    .A3(_0048_),
    .A4(_0226_),
    .B1(net107),
    .X(_0356_));
 sky130_fd_sc_hd__o21a_1 _1167_ (.A1(_0355_),
    .A2(_0356_),
    .B1(net88),
    .X(_0357_));
 sky130_fd_sc_hd__a41o_1 _1168_ (.A1(net76),
    .A2(_0048_),
    .A3(_0143_),
    .A4(_0227_),
    .B1(net85),
    .X(_0358_));
 sky130_fd_sc_hd__and4_1 _1169_ (.A(net136),
    .B(_0796_),
    .C(_0059_),
    .D(_0068_),
    .X(_0359_));
 sky130_fd_sc_hd__nor2_1 _1170_ (.A(_0295_),
    .B(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__o21ai_1 _1171_ (.A1(_0358_),
    .A2(_0360_),
    .B1(_0357_),
    .Y(_0361_));
 sky130_fd_sc_hd__o31a_1 _1172_ (.A1(_0805_),
    .A2(_0037_),
    .A3(_0057_),
    .B1(net76),
    .X(_0362_));
 sky130_fd_sc_hd__o211a_1 _1173_ (.A1(net63),
    .A2(_0115_),
    .B1(_0249_),
    .C1(net118),
    .X(_0363_));
 sky130_fd_sc_hd__o31a_1 _1174_ (.A1(net107),
    .A2(_0362_),
    .A3(_0363_),
    .B1(net98),
    .X(_0364_));
 sky130_fd_sc_hd__or3b_1 _1175_ (.A(net85),
    .B(_0805_),
    .C_N(_0202_),
    .X(_0365_));
 sky130_fd_sc_hd__o21ai_1 _1176_ (.A1(_0333_),
    .A2(_0365_),
    .B1(net57),
    .Y(_0366_));
 sky130_fd_sc_hd__nor2_1 _1177_ (.A(net61),
    .B(_0055_),
    .Y(_0367_));
 sky130_fd_sc_hd__nor2_1 _1178_ (.A(net163),
    .B(_0056_),
    .Y(_0368_));
 sky130_fd_sc_hd__or3_1 _1179_ (.A(_0049_),
    .B(_0367_),
    .C(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__a21bo_1 _1180_ (.A1(_0366_),
    .A2(_0369_),
    .B1_N(_0364_),
    .X(_0370_));
 sky130_fd_sc_hd__a21oi_1 _1181_ (.A1(_0361_),
    .A2(_0370_),
    .B1(net90),
    .Y(_0371_));
 sky130_fd_sc_hd__or3_2 _1182_ (.A(net136),
    .B(_0736_),
    .C(net53),
    .X(_0372_));
 sky130_fd_sc_hd__or3_1 _1183_ (.A(net132),
    .B(net68),
    .C(net53),
    .X(_0373_));
 sky130_fd_sc_hd__a211o_1 _1184_ (.A1(_0226_),
    .A2(_0372_),
    .B1(net76),
    .C1(_0757_),
    .X(_0374_));
 sky130_fd_sc_hd__a21bo_1 _1185_ (.A1(_0366_),
    .A2(_0374_),
    .B1_N(_0364_),
    .X(_0375_));
 sky130_fd_sc_hd__a21oi_1 _1186_ (.A1(net67),
    .A2(_0128_),
    .B1(_0295_),
    .Y(_0376_));
 sky130_fd_sc_hd__o21ai_1 _1187_ (.A1(_0358_),
    .A2(_0376_),
    .B1(_0357_),
    .Y(_0377_));
 sky130_fd_sc_hd__a31o_1 _1188_ (.A1(net90),
    .A2(_0375_),
    .A3(_0377_),
    .B1(net170),
    .X(_0378_));
 sky130_fd_sc_hd__a2bb2o_1 _1189_ (.A1_N(_0378_),
    .A2_N(_0371_),
    .B1(net197),
    .B2(net170),
    .X(_0007_));
 sky130_fd_sc_hd__o21ai_1 _1190_ (.A1(net158),
    .A2(net51),
    .B1(net133),
    .Y(_0379_));
 sky130_fd_sc_hd__and3_1 _1191_ (.A(net123),
    .B(_0119_),
    .C(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__or2_1 _1192_ (.A(_0158_),
    .B(_0239_),
    .X(_0381_));
 sky130_fd_sc_hd__and4_1 _1193_ (.A(net82),
    .B(_0086_),
    .C(_0226_),
    .D(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__o31a_1 _1194_ (.A1(net102),
    .A2(_0380_),
    .A3(_0382_),
    .B1(_0343_),
    .X(_0383_));
 sky130_fd_sc_hd__a21oi_1 _1195_ (.A1(_0800_),
    .A2(net47),
    .B1(_0178_),
    .Y(_0384_));
 sky130_fd_sc_hd__o21a_1 _1196_ (.A1(net67),
    .A2(_0075_),
    .B1(_0349_),
    .X(_0385_));
 sky130_fd_sc_hd__o21a_1 _1197_ (.A1(_0384_),
    .A2(_0385_),
    .B1(net113),
    .X(_0386_));
 sky130_fd_sc_hd__nand2_1 _1198_ (.A(_0068_),
    .B(_0085_),
    .Y(_0387_));
 sky130_fd_sc_hd__a221o_1 _1199_ (.A1(net62),
    .A2(_0043_),
    .B1(net50),
    .B2(_0085_),
    .C1(net127),
    .X(_0388_));
 sky130_fd_sc_hd__a21o_1 _1200_ (.A1(_0199_),
    .A2(_0276_),
    .B1(net82),
    .X(_0389_));
 sky130_fd_sc_hd__a21oi_1 _1201_ (.A1(_0388_),
    .A2(_0389_),
    .B1(net113),
    .Y(_0390_));
 sky130_fd_sc_hd__a211o_1 _1202_ (.A1(_0087_),
    .A2(_0372_),
    .B1(_0127_),
    .C1(_0757_),
    .X(_0391_));
 sky130_fd_sc_hd__nand2_1 _1203_ (.A(net102),
    .B(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__and3_1 _1204_ (.A(net42),
    .B(_0084_),
    .C(_0137_),
    .X(_0393_));
 sky130_fd_sc_hd__o32a_1 _1205_ (.A1(_0390_),
    .A2(_0392_),
    .A3(_0393_),
    .B1(_0386_),
    .B2(_0383_),
    .X(_0394_));
 sky130_fd_sc_hd__o21ai_1 _1206_ (.A1(net167),
    .A2(net50),
    .B1(net59),
    .Y(_0395_));
 sky130_fd_sc_hd__and3_1 _1207_ (.A(net42),
    .B(_0084_),
    .C(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__nor3_1 _1208_ (.A(_0390_),
    .B(_0392_),
    .C(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__o211a_1 _1209_ (.A1(_0069_),
    .A2(_0086_),
    .B1(_0349_),
    .C1(_0065_),
    .X(_0398_));
 sky130_fd_sc_hd__o21a_1 _1210_ (.A1(_0384_),
    .A2(_0398_),
    .B1(net113),
    .X(_0399_));
 sky130_fd_sc_hd__o21ai_1 _1211_ (.A1(_0383_),
    .A2(_0399_),
    .B1(net95),
    .Y(_0400_));
 sky130_fd_sc_hd__o221a_1 _1212_ (.A1(net95),
    .A2(_0394_),
    .B1(_0397_),
    .B2(_0400_),
    .C1(net175),
    .X(_0401_));
 sky130_fd_sc_hd__o21ba_1 _1213_ (.A1(net9),
    .A2(net184),
    .B1_N(_0401_),
    .X(_0008_));
 sky130_fd_sc_hd__and2_1 _1214_ (.A(net171),
    .B(net203),
    .X(_0402_));
 sky130_fd_sc_hd__o221a_1 _1215_ (.A1(net142),
    .A2(net50),
    .B1(_0242_),
    .B2(net61),
    .C1(_0041_),
    .X(_0403_));
 sky130_fd_sc_hd__nand2b_1 _1216_ (.A_N(net131),
    .B(net115),
    .Y(_0404_));
 sky130_fd_sc_hd__a21o_1 _1217_ (.A1(net135),
    .A2(_0798_),
    .B1(net79),
    .X(_0405_));
 sky130_fd_sc_hd__o21ai_1 _1218_ (.A1(net45),
    .A2(_0112_),
    .B1(_0087_),
    .Y(_0406_));
 sky130_fd_sc_hd__o22a_1 _1219_ (.A1(net126),
    .A2(_0403_),
    .B1(_0405_),
    .B2(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__or2_1 _1220_ (.A(_0093_),
    .B(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__o21a_1 _1221_ (.A1(_0256_),
    .A2(_0344_),
    .B1(net42),
    .X(_0409_));
 sky130_fd_sc_hd__a211o_1 _1222_ (.A1(net151),
    .A2(_0767_),
    .B1(net63),
    .C1(_0129_),
    .X(_0410_));
 sky130_fd_sc_hd__nand3_1 _1223_ (.A(net125),
    .B(_0276_),
    .C(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__or3_1 _1224_ (.A(net125),
    .B(_0074_),
    .C(_0367_),
    .X(_0412_));
 sky130_fd_sc_hd__a21oi_1 _1225_ (.A1(_0201_),
    .A2(_0234_),
    .B1(_0127_),
    .Y(_0413_));
 sky130_fd_sc_hd__a311o_1 _1226_ (.A1(net86),
    .A2(_0411_),
    .A3(_0412_),
    .B1(_0413_),
    .C1(net102),
    .X(_0414_));
 sky130_fd_sc_hd__or2_1 _1227_ (.A(_0409_),
    .B(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__a31o_1 _1228_ (.A1(net117),
    .A2(net65),
    .A3(_0059_),
    .B1(_0110_),
    .X(_0416_));
 sky130_fd_sc_hd__or3_1 _1229_ (.A(_0332_),
    .B(_0368_),
    .C(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__a31o_1 _1230_ (.A1(_0408_),
    .A2(_0415_),
    .A3(_0417_),
    .B1(net94),
    .X(_0418_));
 sky130_fd_sc_hd__o21a_1 _1231_ (.A1(net55),
    .A2(_0276_),
    .B1(_0202_),
    .X(_0419_));
 sky130_fd_sc_hd__o22a_1 _1232_ (.A1(_0127_),
    .A2(_0403_),
    .B1(_0419_),
    .B2(net58),
    .X(_0420_));
 sky130_fd_sc_hd__nor2_1 _1233_ (.A(net63),
    .B(_0075_),
    .Y(_0421_));
 sky130_fd_sc_hd__o21a_1 _1234_ (.A1(_0344_),
    .A2(_0421_),
    .B1(net43),
    .X(_0422_));
 sky130_fd_sc_hd__o211a_1 _1235_ (.A1(net89),
    .A2(_0420_),
    .B1(_0417_),
    .C1(net94),
    .X(_0423_));
 sky130_fd_sc_hd__o21ai_1 _1236_ (.A1(_0414_),
    .A2(_0422_),
    .B1(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__a31o_1 _1237_ (.A1(net175),
    .A2(_0418_),
    .A3(_0424_),
    .B1(_0402_),
    .X(_0009_));
 sky130_fd_sc_hd__o31a_1 _1238_ (.A1(net75),
    .A2(net155),
    .A3(net53),
    .B1(_0404_),
    .X(_0425_));
 sky130_fd_sc_hd__or2_1 _1239_ (.A(_0095_),
    .B(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__a21o_1 _1240_ (.A1(_0050_),
    .A2(net48),
    .B1(_0291_),
    .X(_0427_));
 sky130_fd_sc_hd__a31o_1 _1241_ (.A1(net84),
    .A2(_0426_),
    .A3(_0427_),
    .B1(net100),
    .X(_0428_));
 sky130_fd_sc_hd__a21oi_1 _1242_ (.A1(_0119_),
    .A2(_0181_),
    .B1(net114),
    .Y(_0429_));
 sky130_fd_sc_hd__a21o_1 _1243_ (.A1(_0119_),
    .A2(_0181_),
    .B1(net114),
    .X(_0430_));
 sky130_fd_sc_hd__o21ai_2 _1244_ (.A1(net130),
    .A2(_0271_),
    .B1(net114),
    .Y(_0431_));
 sky130_fd_sc_hd__a221oi_1 _1245_ (.A1(net114),
    .A2(_0188_),
    .B1(_0430_),
    .B2(_0431_),
    .C1(net84),
    .Y(_0432_));
 sky130_fd_sc_hd__o21a_1 _1246_ (.A1(_0808_),
    .A2(net51),
    .B1(_0186_),
    .X(_0433_));
 sky130_fd_sc_hd__a31o_1 _1247_ (.A1(net75),
    .A2(net48),
    .A3(_0108_),
    .B1(net88),
    .X(_0434_));
 sky130_fd_sc_hd__o21a_1 _1248_ (.A1(_0433_),
    .A2(_0434_),
    .B1(_0093_),
    .X(_0435_));
 sky130_fd_sc_hd__or3_1 _1249_ (.A(net142),
    .B(net68),
    .C(net52),
    .X(_0436_));
 sky130_fd_sc_hd__o211ai_4 _1250_ (.A1(net154),
    .A2(net162),
    .B1(net130),
    .C1(net145),
    .Y(_0437_));
 sky130_fd_sc_hd__o311a_1 _1251_ (.A1(net131),
    .A2(net68),
    .A3(net51),
    .B1(_0437_),
    .C1(net75),
    .X(_0438_));
 sky130_fd_sc_hd__o211a_1 _1252_ (.A1(_0055_),
    .A2(_0067_),
    .B1(_0063_),
    .C1(net114),
    .X(_0439_));
 sky130_fd_sc_hd__o21a_1 _1253_ (.A1(_0438_),
    .A2(_0439_),
    .B1(net104),
    .X(_0440_));
 sky130_fd_sc_hd__o22a_1 _1254_ (.A1(_0428_),
    .A2(_0432_),
    .B1(_0435_),
    .B2(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__and3_1 _1255_ (.A(net114),
    .B(net70),
    .C(_0271_),
    .X(_0442_));
 sky130_fd_sc_hd__o21a_1 _1256_ (.A1(_0429_),
    .A2(_0442_),
    .B1(net104),
    .X(_0443_));
 sky130_fd_sc_hd__a31o_1 _1257_ (.A1(net115),
    .A2(_0063_),
    .A3(_0242_),
    .B1(_0438_),
    .X(_0444_));
 sky130_fd_sc_hd__a21o_1 _1258_ (.A1(net104),
    .A2(_0444_),
    .B1(_0435_),
    .X(_0445_));
 sky130_fd_sc_hd__o211ai_1 _1259_ (.A1(_0428_),
    .A2(_0443_),
    .B1(_0445_),
    .C1(net92),
    .Y(_0446_));
 sky130_fd_sc_hd__o211a_1 _1260_ (.A1(net92),
    .A2(_0441_),
    .B1(_0446_),
    .C1(net173),
    .X(_0447_));
 sky130_fd_sc_hd__o21ba_1 _1261_ (.A1(net173),
    .A2(net192),
    .B1_N(_0447_),
    .X(_0010_));
 sky130_fd_sc_hd__a211o_1 _1262_ (.A1(net64),
    .A2(net46),
    .B1(_0095_),
    .C1(net120),
    .X(_0448_));
 sky130_fd_sc_hd__or3_1 _1263_ (.A(net44),
    .B(_0183_),
    .C(_0405_),
    .X(_0449_));
 sky130_fd_sc_hd__a31o_1 _1264_ (.A1(net84),
    .A2(_0448_),
    .A3(_0449_),
    .B1(net88),
    .X(_0450_));
 sky130_fd_sc_hd__and3_1 _1265_ (.A(net131),
    .B(_0802_),
    .C(_0068_),
    .X(_0451_));
 sky130_fd_sc_hd__or2_1 _1266_ (.A(_0067_),
    .B(_0181_),
    .X(_0452_));
 sky130_fd_sc_hd__o21ai_2 _1267_ (.A1(_0757_),
    .A2(_0304_),
    .B1(net120),
    .Y(_0453_));
 sky130_fd_sc_hd__o221a_1 _1268_ (.A1(_0291_),
    .A2(_0333_),
    .B1(_0451_),
    .B2(_0453_),
    .C1(net104),
    .X(_0454_));
 sky130_fd_sc_hd__a211o_1 _1269_ (.A1(_0071_),
    .A2(_0074_),
    .B1(_0345_),
    .C1(net79),
    .X(_0455_));
 sky130_fd_sc_hd__a21o_1 _1270_ (.A1(_0076_),
    .A2(_0165_),
    .B1(net121),
    .X(_0456_));
 sky130_fd_sc_hd__a21oi_1 _1271_ (.A1(net166),
    .A2(_0069_),
    .B1(_0158_),
    .Y(_0457_));
 sky130_fd_sc_hd__nor2_1 _1272_ (.A(net165),
    .B(_0190_),
    .Y(_0458_));
 sky130_fd_sc_hd__o21a_1 _1273_ (.A1(_0457_),
    .A2(_0458_),
    .B1(_0126_),
    .X(_0459_));
 sky130_fd_sc_hd__a311o_1 _1274_ (.A1(net87),
    .A2(_0455_),
    .A3(_0456_),
    .B1(_0459_),
    .C1(net101),
    .X(_0460_));
 sky130_fd_sc_hd__and3_1 _1275_ (.A(net42),
    .B(_0108_),
    .C(_0437_),
    .X(_0461_));
 sky130_fd_sc_hd__o221a_1 _1276_ (.A1(_0450_),
    .A2(_0454_),
    .B1(_0460_),
    .B2(_0461_),
    .C1(net93),
    .X(_0462_));
 sky130_fd_sc_hd__or2_1 _1277_ (.A(net134),
    .B(_0800_),
    .X(_0463_));
 sky130_fd_sc_hd__a21oi_1 _1278_ (.A1(_0242_),
    .A2(_0463_),
    .B1(net58),
    .Y(_0464_));
 sky130_fd_sc_hd__o21ai_1 _1279_ (.A1(_0757_),
    .A2(_0304_),
    .B1(_0181_),
    .Y(_0465_));
 sky130_fd_sc_hd__o221a_1 _1280_ (.A1(_0291_),
    .A2(_0333_),
    .B1(_0465_),
    .B2(net75),
    .C1(net104),
    .X(_0466_));
 sky130_fd_sc_hd__o22a_1 _1281_ (.A1(_0460_),
    .A2(_0464_),
    .B1(_0466_),
    .B2(_0450_),
    .X(_0467_));
 sky130_fd_sc_hd__o21ai_1 _1282_ (.A1(net93),
    .A2(_0467_),
    .B1(net176),
    .Y(_0468_));
 sky130_fd_sc_hd__o22a_1 _1283_ (.A1(net176),
    .A2(net193),
    .B1(_0462_),
    .B2(_0468_),
    .X(_0011_));
 sky130_fd_sc_hd__nor2_1 _1284_ (.A(net122),
    .B(_0062_),
    .Y(_0469_));
 sky130_fd_sc_hd__a22o_1 _1285_ (.A1(_0215_),
    .A2(_0308_),
    .B1(_0469_),
    .B2(_0234_),
    .X(_0470_));
 sky130_fd_sc_hd__a21o_1 _1286_ (.A1(net83),
    .A2(_0470_),
    .B1(net88),
    .X(_0471_));
 sky130_fd_sc_hd__and2_1 _1287_ (.A(net134),
    .B(_0071_),
    .X(_0472_));
 sky130_fd_sc_hd__a2111o_1 _1288_ (.A1(net163),
    .A2(net48),
    .B1(_0757_),
    .C1(net70),
    .D1(net56),
    .X(_0473_));
 sky130_fd_sc_hd__nand2_1 _1289_ (.A(net71),
    .B(_0124_),
    .Y(_0474_));
 sky130_fd_sc_hd__a21oi_1 _1290_ (.A1(_0473_),
    .A2(_0474_),
    .B1(net120),
    .Y(_0475_));
 sky130_fd_sc_hd__or3_1 _1291_ (.A(net134),
    .B(_0803_),
    .C(_0139_),
    .X(_0476_));
 sky130_fd_sc_hd__and3_1 _1292_ (.A(net120),
    .B(_0181_),
    .C(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__o21a_1 _1293_ (.A1(_0475_),
    .A2(_0477_),
    .B1(net104),
    .X(_0478_));
 sky130_fd_sc_hd__o211a_2 _1294_ (.A1(net163),
    .A2(net50),
    .B1(net62),
    .C1(net131),
    .X(_0479_));
 sky130_fd_sc_hd__o21a_1 _1295_ (.A1(_0075_),
    .A2(_0139_),
    .B1(_0322_),
    .X(_0480_));
 sky130_fd_sc_hd__o32a_1 _1296_ (.A1(_0047_),
    .A2(_0049_),
    .A3(_0479_),
    .B1(_0480_),
    .B2(net121),
    .X(_0481_));
 sky130_fd_sc_hd__a221o_1 _1297_ (.A1(_0800_),
    .A2(_0807_),
    .B1(_0059_),
    .B2(_0095_),
    .C1(net119),
    .X(_0482_));
 sky130_fd_sc_hd__nand2_1 _1298_ (.A(net105),
    .B(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__nand2_2 _1299_ (.A(net54),
    .B(_0128_),
    .Y(_0484_));
 sky130_fd_sc_hd__a21oi_1 _1300_ (.A1(_0373_),
    .A2(_0484_),
    .B1(net74),
    .Y(_0485_));
 sky130_fd_sc_hd__o22a_1 _1301_ (.A1(net105),
    .A2(_0481_),
    .B1(_0483_),
    .B2(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__o221a_1 _1302_ (.A1(_0471_),
    .A2(_0478_),
    .B1(_0486_),
    .B2(net100),
    .C1(net92),
    .X(_0487_));
 sky130_fd_sc_hd__nor2_1 _1303_ (.A(_0072_),
    .B(_0114_),
    .Y(_0488_));
 sky130_fd_sc_hd__or2_1 _1304_ (.A(_0072_),
    .B(_0114_),
    .X(_0489_));
 sky130_fd_sc_hd__o311a_1 _1305_ (.A1(_0049_),
    .A2(_0368_),
    .A3(_0488_),
    .B1(_0482_),
    .C1(net105),
    .X(_0490_));
 sky130_fd_sc_hd__o21ba_1 _1306_ (.A1(net105),
    .A2(_0481_),
    .B1_N(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__a31o_1 _1307_ (.A1(net120),
    .A2(_0452_),
    .A3(_0476_),
    .B1(_0475_),
    .X(_0492_));
 sky130_fd_sc_hd__a211oi_1 _1308_ (.A1(net104),
    .A2(_0492_),
    .B1(_0471_),
    .C1(net92),
    .Y(_0493_));
 sky130_fd_sc_hd__o21ai_1 _1309_ (.A1(_0176_),
    .A2(_0491_),
    .B1(net173),
    .Y(_0494_));
 sky130_fd_sc_hd__o32a_1 _1310_ (.A1(_0487_),
    .A2(_0493_),
    .A3(_0494_),
    .B1(net182),
    .B2(net174),
    .X(_0012_));
 sky130_fd_sc_hd__a221o_1 _1311_ (.A1(net71),
    .A2(net64),
    .B1(net48),
    .B2(_0085_),
    .C1(net122),
    .X(_0495_));
 sky130_fd_sc_hd__nand2_1 _1312_ (.A(net62),
    .B(net46),
    .Y(_0496_));
 sky130_fd_sc_hd__nand2_1 _1313_ (.A(_0040_),
    .B(_0068_),
    .Y(_0497_));
 sky130_fd_sc_hd__a21o_1 _1314_ (.A1(_0496_),
    .A2(_0497_),
    .B1(net79),
    .X(_0498_));
 sky130_fd_sc_hd__a31o_1 _1315_ (.A1(net83),
    .A2(_0495_),
    .A3(_0498_),
    .B1(net101),
    .X(_0499_));
 sky130_fd_sc_hd__a21oi_1 _1316_ (.A1(_0090_),
    .A2(_0473_),
    .B1(net120),
    .Y(_0500_));
 sky130_fd_sc_hd__o21bai_1 _1317_ (.A1(_0431_),
    .A2(_0472_),
    .B1_N(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__a21o_1 _1318_ (.A1(net109),
    .A2(_0501_),
    .B1(_0499_),
    .X(_0502_));
 sky130_fd_sc_hd__a221o_1 _1319_ (.A1(net134),
    .A2(_0069_),
    .B1(_0463_),
    .B2(_0055_),
    .C1(net120),
    .X(_0503_));
 sky130_fd_sc_hd__a21o_1 _1320_ (.A1(net62),
    .A2(_0095_),
    .B1(_0080_),
    .X(_0504_));
 sky130_fd_sc_hd__a31oi_1 _1321_ (.A1(net101),
    .A2(_0503_),
    .A3(_0504_),
    .B1(_0092_),
    .Y(_0505_));
 sky130_fd_sc_hd__nand2b_1 _1322_ (.A_N(_0130_),
    .B(_0235_),
    .Y(_0506_));
 sky130_fd_sc_hd__o211ai_2 _1323_ (.A1(net66),
    .A2(_0224_),
    .B1(_0215_),
    .C1(net79),
    .Y(_0507_));
 sky130_fd_sc_hd__a31o_1 _1324_ (.A1(net109),
    .A2(_0506_),
    .A3(_0507_),
    .B1(_0505_),
    .X(_0508_));
 sky130_fd_sc_hd__a21oi_1 _1325_ (.A1(_0502_),
    .A2(_0508_),
    .B1(net93),
    .Y(_0509_));
 sky130_fd_sc_hd__a311o_1 _1326_ (.A1(net120),
    .A2(net64),
    .A3(net46),
    .B1(_0442_),
    .C1(_0500_),
    .X(_0510_));
 sky130_fd_sc_hd__a21o_1 _1327_ (.A1(net109),
    .A2(_0510_),
    .B1(_0499_),
    .X(_0511_));
 sky130_fd_sc_hd__o21ai_1 _1328_ (.A1(net48),
    .A2(_0086_),
    .B1(_0235_),
    .Y(_0512_));
 sky130_fd_sc_hd__a31o_1 _1329_ (.A1(net109),
    .A2(_0507_),
    .A3(_0512_),
    .B1(_0505_),
    .X(_0513_));
 sky130_fd_sc_hd__a31o_1 _1330_ (.A1(net93),
    .A2(_0511_),
    .A3(_0513_),
    .B1(net171),
    .X(_0514_));
 sky130_fd_sc_hd__o22a_1 _1331_ (.A1(net176),
    .A2(net188),
    .B1(_0509_),
    .B2(_0514_),
    .X(_0013_));
 sky130_fd_sc_hd__o41a_1 _1332_ (.A1(net136),
    .A2(_0736_),
    .A3(net63),
    .A4(net60),
    .B1(net76),
    .X(_0515_));
 sky130_fd_sc_hd__nand2_1 _1333_ (.A(_0473_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__a31o_1 _1334_ (.A1(net132),
    .A2(net68),
    .A3(_0035_),
    .B1(_0265_),
    .X(_0517_));
 sky130_fd_sc_hd__a21oi_1 _1335_ (.A1(_0516_),
    .A2(_0517_),
    .B1(net106),
    .Y(_0518_));
 sky130_fd_sc_hd__and3b_1 _1336_ (.A_N(_0102_),
    .B(net116),
    .C(_0051_),
    .X(_0519_));
 sky130_fd_sc_hd__a31o_1 _1337_ (.A1(net74),
    .A2(_0063_),
    .A3(_0279_),
    .B1(net103),
    .X(_0520_));
 sky130_fd_sc_hd__o21a_1 _1338_ (.A1(_0519_),
    .A2(_0520_),
    .B1(net97),
    .X(_0521_));
 sky130_fd_sc_hd__and3_1 _1339_ (.A(net130),
    .B(_0796_),
    .C(_0120_),
    .X(_0522_));
 sky130_fd_sc_hd__o21a_1 _1340_ (.A1(_0050_),
    .A2(_0522_),
    .B1(net75),
    .X(_0523_));
 sky130_fd_sc_hd__nand2_1 _1341_ (.A(_0802_),
    .B(_0045_),
    .Y(_0524_));
 sky130_fd_sc_hd__or2_1 _1342_ (.A(_0075_),
    .B(_0239_),
    .X(_0525_));
 sky130_fd_sc_hd__a31o_1 _1343_ (.A1(net114),
    .A2(_0524_),
    .A3(_0525_),
    .B1(_0523_),
    .X(_0526_));
 sky130_fd_sc_hd__a21bo_1 _1344_ (.A1(net103),
    .A2(_0526_),
    .B1_N(_0521_),
    .X(_0527_));
 sky130_fd_sc_hd__a21o_1 _1345_ (.A1(_0046_),
    .A2(_0105_),
    .B1(net116),
    .X(_0528_));
 sky130_fd_sc_hd__a221o_1 _1346_ (.A1(net130),
    .A2(net51),
    .B1(_0160_),
    .B2(_0059_),
    .C1(net74),
    .X(_0529_));
 sky130_fd_sc_hd__a31o_1 _1347_ (.A1(net103),
    .A2(_0528_),
    .A3(_0529_),
    .B1(net97),
    .X(_0530_));
 sky130_fd_sc_hd__a32o_1 _1348_ (.A1(net130),
    .A2(net51),
    .A3(_0068_),
    .B1(_0160_),
    .B2(_0059_),
    .X(_0531_));
 sky130_fd_sc_hd__o211a_1 _1349_ (.A1(net74),
    .A2(_0531_),
    .B1(_0528_),
    .C1(net103),
    .X(_0532_));
 sky130_fd_sc_hd__or3_1 _1350_ (.A(net97),
    .B(_0518_),
    .C(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__o211a_1 _1351_ (.A1(net145),
    .A2(net154),
    .B1(_0065_),
    .C1(_0349_),
    .X(_0534_));
 sky130_fd_sc_hd__o21ai_1 _1352_ (.A1(_0523_),
    .A2(_0534_),
    .B1(net104),
    .Y(_0535_));
 sky130_fd_sc_hd__o2bb2a_1 _1353_ (.A1_N(_0521_),
    .A2_N(_0535_),
    .B1(_0530_),
    .B2(_0518_),
    .X(_0536_));
 sky130_fd_sc_hd__nor2_1 _1354_ (.A(net92),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__a31o_1 _1355_ (.A1(net92),
    .A2(_0527_),
    .A3(_0533_),
    .B1(net170),
    .X(_0538_));
 sky130_fd_sc_hd__o22a_1 _1356_ (.A1(net173),
    .A2(net190),
    .B1(_0537_),
    .B2(_0538_),
    .X(_0014_));
 sky130_fd_sc_hd__and2_1 _1357_ (.A(net170),
    .B(net206),
    .X(_0539_));
 sky130_fd_sc_hd__nand2_1 _1358_ (.A(_0078_),
    .B(_0095_),
    .Y(_0540_));
 sky130_fd_sc_hd__a21o_1 _1359_ (.A1(_0105_),
    .A2(_0540_),
    .B1(net57),
    .X(_0541_));
 sky130_fd_sc_hd__and3_1 _1360_ (.A(net136),
    .B(net62),
    .C(net49),
    .X(_0542_));
 sky130_fd_sc_hd__o32a_1 _1361_ (.A1(net76),
    .A2(_0245_),
    .A3(_0542_),
    .B1(_0359_),
    .B2(_0354_),
    .X(_0543_));
 sky130_fd_sc_hd__or2_1 _1362_ (.A(net107),
    .B(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__o21ai_1 _1363_ (.A1(_0155_),
    .A2(_0479_),
    .B1(_0126_),
    .Y(_0545_));
 sky130_fd_sc_hd__a31o_1 _1364_ (.A1(_0541_),
    .A2(_0544_),
    .A3(_0545_),
    .B1(net98),
    .X(_0546_));
 sky130_fd_sc_hd__o211a_1 _1365_ (.A1(net130),
    .A2(_0124_),
    .B1(_0804_),
    .C1(net116),
    .X(_0547_));
 sky130_fd_sc_hd__o211a_1 _1366_ (.A1(_0704_),
    .A2(_0114_),
    .B1(_0051_),
    .C1(net74),
    .X(_0548_));
 sky130_fd_sc_hd__o31ai_2 _1367_ (.A1(net103),
    .A2(_0547_),
    .A3(_0548_),
    .B1(net97),
    .Y(_0549_));
 sky130_fd_sc_hd__nor2_1 _1368_ (.A(net50),
    .B(_0112_),
    .Y(_0550_));
 sky130_fd_sc_hd__o31a_1 _1369_ (.A1(net46),
    .A2(_0291_),
    .A3(_0550_),
    .B1(net107),
    .X(_0551_));
 sky130_fd_sc_hd__a22o_1 _1370_ (.A1(_0746_),
    .A2(_0057_),
    .B1(net50),
    .B2(_0807_),
    .X(_0552_));
 sky130_fd_sc_hd__nand2_1 _1371_ (.A(net118),
    .B(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__a21o_1 _1372_ (.A1(_0551_),
    .A2(_0553_),
    .B1(_0549_),
    .X(_0554_));
 sky130_fd_sc_hd__nand3_1 _1373_ (.A(net90),
    .B(_0546_),
    .C(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__or3b_1 _1374_ (.A(net136),
    .B(_0072_),
    .C_N(net156),
    .X(_0556_));
 sky130_fd_sc_hd__or3b_1 _1375_ (.A(net76),
    .B(_0367_),
    .C_N(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__a211o_1 _1376_ (.A1(_0551_),
    .A2(_0557_),
    .B1(net90),
    .C1(_0549_),
    .X(_0558_));
 sky130_fd_sc_hd__nand2_1 _1377_ (.A(net174),
    .B(_0176_),
    .Y(_0559_));
 sky130_fd_sc_hd__a21o_1 _1378_ (.A1(_0243_),
    .A2(_0540_),
    .B1(net57),
    .X(_0560_));
 sky130_fd_sc_hd__a31o_1 _1379_ (.A1(_0544_),
    .A2(_0545_),
    .A3(_0560_),
    .B1(_0176_),
    .X(_0561_));
 sky130_fd_sc_hd__a41o_1 _1380_ (.A1(net174),
    .A2(_0555_),
    .A3(_0558_),
    .A4(_0561_),
    .B1(_0539_),
    .X(_0015_));
 sky130_fd_sc_hd__o221a_1 _1381_ (.A1(_0258_),
    .A2(_0311_),
    .B1(_0425_),
    .B2(_0079_),
    .C1(net84),
    .X(_0562_));
 sky130_fd_sc_hd__or2_1 _1382_ (.A(net99),
    .B(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__nor2_1 _1383_ (.A(net55),
    .B(_0246_),
    .Y(_0564_));
 sky130_fd_sc_hd__o211ai_1 _1384_ (.A1(_0804_),
    .A2(net55),
    .B1(_0143_),
    .C1(net126),
    .Y(_0565_));
 sky130_fd_sc_hd__o311a_1 _1385_ (.A1(net126),
    .A2(_0037_),
    .A3(_0564_),
    .B1(_0565_),
    .C1(net111),
    .X(_0566_));
 sky130_fd_sc_hd__o21a_1 _1386_ (.A1(net169),
    .A2(_0129_),
    .B1(_0048_),
    .X(_0567_));
 sky130_fd_sc_hd__o311a_1 _1387_ (.A1(_0040_),
    .A2(_0045_),
    .A3(net47),
    .B1(_0796_),
    .C1(net77),
    .X(_0568_));
 sky130_fd_sc_hd__a31oi_1 _1388_ (.A1(net117),
    .A2(_0143_),
    .A3(_0567_),
    .B1(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__a221o_1 _1389_ (.A1(net65),
    .A2(_0062_),
    .B1(_0072_),
    .B2(net46),
    .C1(_0127_),
    .X(_0570_));
 sky130_fd_sc_hd__o211a_1 _1390_ (.A1(net108),
    .A2(_0569_),
    .B1(_0570_),
    .C1(net99),
    .X(_0571_));
 sky130_fd_sc_hd__a31o_1 _1391_ (.A1(net142),
    .A2(net69),
    .A3(net54),
    .B1(_0318_),
    .X(_0572_));
 sky130_fd_sc_hd__a2bb2o_1 _1392_ (.A1_N(_0563_),
    .A2_N(_0566_),
    .B1(_0571_),
    .B2(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__nand2_1 _1393_ (.A(_0652_),
    .B(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__nand3_1 _1394_ (.A(net126),
    .B(_0143_),
    .C(_0484_),
    .Y(_0575_));
 sky130_fd_sc_hd__o311a_1 _1395_ (.A1(net126),
    .A2(_0037_),
    .A3(_0564_),
    .B1(_0575_),
    .C1(net111),
    .X(_0576_));
 sky130_fd_sc_hd__nor2_1 _1396_ (.A(_0563_),
    .B(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__o221a_1 _1397_ (.A1(net58),
    .A2(_0202_),
    .B1(_0318_),
    .B2(_0345_),
    .C1(_0571_),
    .X(_0578_));
 sky130_fd_sc_hd__o31a_1 _1398_ (.A1(_0652_),
    .A2(_0577_),
    .A3(_0578_),
    .B1(net175),
    .X(_0579_));
 sky130_fd_sc_hd__o2bb2a_1 _1399_ (.A1_N(_0574_),
    .A2_N(_0579_),
    .B1(net175),
    .B2(net199),
    .X(_0016_));
 sky130_fd_sc_hd__o311a_1 _1400_ (.A1(_0736_),
    .A2(net45),
    .A3(_0112_),
    .B1(_0278_),
    .C1(net77),
    .X(_0580_));
 sky130_fd_sc_hd__o211a_1 _1401_ (.A1(net136),
    .A2(_0117_),
    .B1(_0115_),
    .C1(net117),
    .X(_0581_));
 sky130_fd_sc_hd__o31ai_2 _1402_ (.A1(net108),
    .A2(_0580_),
    .A3(_0581_),
    .B1(net99),
    .Y(_0582_));
 sky130_fd_sc_hd__a221o_1 _1403_ (.A1(net151),
    .A2(_0807_),
    .B1(_0045_),
    .B2(net69),
    .C1(net80),
    .X(_0583_));
 sky130_fd_sc_hd__o311a_1 _1404_ (.A1(net126),
    .A2(_0062_),
    .A3(_0213_),
    .B1(_0583_),
    .C1(net111),
    .X(_0584_));
 sky130_fd_sc_hd__o211a_1 _1405_ (.A1(_0804_),
    .A2(_0058_),
    .B1(_0436_),
    .C1(net128),
    .X(_0585_));
 sky130_fd_sc_hd__a31o_1 _1406_ (.A1(net82),
    .A2(_0075_),
    .A3(_0096_),
    .B1(net102),
    .X(_0586_));
 sky130_fd_sc_hd__o21a_1 _1407_ (.A1(_0585_),
    .A2(_0586_),
    .B1(_0343_),
    .X(_0587_));
 sky130_fd_sc_hd__o21a_1 _1408_ (.A1(net64),
    .A2(_0114_),
    .B1(_0284_),
    .X(_0588_));
 sky130_fd_sc_hd__nor2_1 _1409_ (.A(_0127_),
    .B(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__o221a_1 _1410_ (.A1(_0808_),
    .A2(net49),
    .B1(_0112_),
    .B2(_0757_),
    .C1(net43),
    .X(_0590_));
 sky130_fd_sc_hd__o32a_1 _1411_ (.A1(_0587_),
    .A2(_0589_),
    .A3(_0590_),
    .B1(_0584_),
    .B2(_0582_),
    .X(_0591_));
 sky130_fd_sc_hd__or2_1 _1412_ (.A(net94),
    .B(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__o21a_1 _1413_ (.A1(_0062_),
    .A2(_0213_),
    .B1(net81),
    .X(_0593_));
 sky130_fd_sc_hd__a31o_1 _1414_ (.A1(net126),
    .A2(_0166_),
    .A3(_0242_),
    .B1(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__a21oi_1 _1415_ (.A1(net111),
    .A2(_0594_),
    .B1(_0582_),
    .Y(_0595_));
 sky130_fd_sc_hd__nand2_1 _1416_ (.A(net81),
    .B(_0588_),
    .Y(_0596_));
 sky130_fd_sc_hd__or3b_1 _1417_ (.A(_0367_),
    .B(net81),
    .C_N(_0276_),
    .X(_0597_));
 sky130_fd_sc_hd__a31oi_1 _1418_ (.A1(net112),
    .A2(_0596_),
    .A3(_0597_),
    .B1(_0587_),
    .Y(_0598_));
 sky130_fd_sc_hd__o31a_1 _1419_ (.A1(_0652_),
    .A2(_0595_),
    .A3(_0598_),
    .B1(net175),
    .X(_0599_));
 sky130_fd_sc_hd__o2bb2a_1 _1420_ (.A1_N(_0592_),
    .A2_N(_0599_),
    .B1(net175),
    .B2(net198),
    .X(_0017_));
 sky130_fd_sc_hd__and2_1 _1421_ (.A(net171),
    .B(net204),
    .X(_0600_));
 sky130_fd_sc_hd__a31o_1 _1422_ (.A1(net142),
    .A2(_0068_),
    .A3(_0140_),
    .B1(_0283_),
    .X(_0601_));
 sky130_fd_sc_hd__o211ai_1 _1423_ (.A1(_0096_),
    .A2(_0136_),
    .B1(_0177_),
    .C1(_0086_),
    .Y(_0602_));
 sky130_fd_sc_hd__a21o_1 _1424_ (.A1(net82),
    .A2(_0602_),
    .B1(net113),
    .X(_0603_));
 sky130_fd_sc_hd__a21o_1 _1425_ (.A1(net128),
    .A2(_0601_),
    .B1(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__or3_1 _1426_ (.A(net86),
    .B(_0138_),
    .C(_0142_),
    .X(_0605_));
 sky130_fd_sc_hd__o21a_1 _1427_ (.A1(_0585_),
    .A2(_0605_),
    .B1(_0604_),
    .X(_0606_));
 sky130_fd_sc_hd__or2_1 _1428_ (.A(_0164_),
    .B(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__or4_1 _1429_ (.A(net111),
    .B(_0132_),
    .C(_0332_),
    .D(_0593_),
    .X(_0608_));
 sky130_fd_sc_hd__and3_1 _1430_ (.A(net65),
    .B(_0107_),
    .C(_0120_),
    .X(_0609_));
 sky130_fd_sc_hd__o21ai_1 _1431_ (.A1(_0154_),
    .A2(_0609_),
    .B1(net111),
    .Y(_0610_));
 sky130_fd_sc_hd__a211o_1 _1432_ (.A1(net59),
    .A2(_0277_),
    .B1(net63),
    .C1(net61),
    .X(_0611_));
 sky130_fd_sc_hd__a31o_1 _1433_ (.A1(net125),
    .A2(_0198_),
    .A3(_0611_),
    .B1(_0610_),
    .X(_0612_));
 sky130_fd_sc_hd__a21oi_1 _1434_ (.A1(_0608_),
    .A2(_0612_),
    .B1(net94),
    .Y(_0613_));
 sky130_fd_sc_hd__o21a_1 _1435_ (.A1(_0205_),
    .A2(_0272_),
    .B1(net125),
    .X(_0614_));
 sky130_fd_sc_hd__o211a_1 _1436_ (.A1(_0610_),
    .A2(_0614_),
    .B1(net94),
    .C1(_0608_),
    .X(_0615_));
 sky130_fd_sc_hd__or3_1 _1437_ (.A(net89),
    .B(_0613_),
    .C(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__a32o_1 _1438_ (.A1(net128),
    .A2(_0436_),
    .A3(_0484_),
    .B1(_0605_),
    .B2(net58),
    .X(_0617_));
 sky130_fd_sc_hd__nand3_1 _1439_ (.A(_0175_),
    .B(_0604_),
    .C(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__a41o_1 _1440_ (.A1(net176),
    .A2(_0607_),
    .A3(_0616_),
    .A4(_0618_),
    .B1(_0600_),
    .X(_0018_));
 sky130_fd_sc_hd__o211a_1 _1441_ (.A1(_0807_),
    .A2(_0183_),
    .B1(_0035_),
    .C1(net74),
    .X(_0619_));
 sky130_fd_sc_hd__a31o_1 _1442_ (.A1(net115),
    .A2(_0190_),
    .A3(_0373_),
    .B1(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__a21o_1 _1443_ (.A1(net84),
    .A2(_0620_),
    .B1(net97),
    .X(_0621_));
 sky130_fd_sc_hd__o21ai_1 _1444_ (.A1(_0251_),
    .A2(_0273_),
    .B1(net57),
    .Y(_0622_));
 sky130_fd_sc_hd__o21ai_1 _1445_ (.A1(_0804_),
    .A2(net49),
    .B1(_0284_),
    .Y(_0623_));
 sky130_fd_sc_hd__nand2_1 _1446_ (.A(net116),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__a21o_1 _1447_ (.A1(_0622_),
    .A2(_0624_),
    .B1(_0621_),
    .X(_0625_));
 sky130_fd_sc_hd__a21oi_1 _1448_ (.A1(_0064_),
    .A2(_0290_),
    .B1(net116),
    .Y(_0626_));
 sky130_fd_sc_hd__a311oi_2 _1449_ (.A1(net116),
    .A2(_0228_),
    .A3(_0243_),
    .B1(_0626_),
    .C1(net106),
    .Y(_0627_));
 sky130_fd_sc_hd__a21oi_1 _1450_ (.A1(_0043_),
    .A2(net56),
    .B1(net115),
    .Y(_0628_));
 sky130_fd_sc_hd__a21oi_1 _1451_ (.A1(_0088_),
    .A2(_0628_),
    .B1(net84),
    .Y(_0629_));
 sky130_fd_sc_hd__o31a_1 _1452_ (.A1(net60),
    .A2(_0097_),
    .A3(_0188_),
    .B1(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__o21ai_1 _1453_ (.A1(_0627_),
    .A2(_0630_),
    .B1(net97),
    .Y(_0631_));
 sky130_fd_sc_hd__a21oi_1 _1454_ (.A1(_0625_),
    .A2(_0631_),
    .B1(net92),
    .Y(_0632_));
 sky130_fd_sc_hd__o21a_1 _1455_ (.A1(_0056_),
    .A2(_0097_),
    .B1(_0629_),
    .X(_0633_));
 sky130_fd_sc_hd__o21ai_1 _1456_ (.A1(_0627_),
    .A2(_0633_),
    .B1(net97),
    .Y(_0634_));
 sky130_fd_sc_hd__nand2_1 _1457_ (.A(_0099_),
    .B(_0116_),
    .Y(_0635_));
 sky130_fd_sc_hd__a21o_1 _1458_ (.A1(_0622_),
    .A2(_0635_),
    .B1(_0621_),
    .X(_0636_));
 sky130_fd_sc_hd__a31o_1 _1459_ (.A1(net92),
    .A2(_0634_),
    .A3(_0636_),
    .B1(net170),
    .X(_0637_));
 sky130_fd_sc_hd__o22a_1 _1460_ (.A1(net173),
    .A2(net183),
    .B1(_0632_),
    .B2(_0637_),
    .X(_0019_));
 sky130_fd_sc_hd__a21oi_1 _1461_ (.A1(_0116_),
    .A2(_0497_),
    .B1(net122),
    .Y(_0638_));
 sky130_fd_sc_hd__a21oi_1 _1462_ (.A1(_0804_),
    .A2(_0201_),
    .B1(_0309_),
    .Y(_0639_));
 sky130_fd_sc_hd__o31a_1 _1463_ (.A1(net109),
    .A2(_0638_),
    .A3(_0639_),
    .B1(net88),
    .X(_0640_));
 sky130_fd_sc_hd__o21a_1 _1464_ (.A1(net159),
    .A2(net52),
    .B1(_0451_),
    .X(_0641_));
 sky130_fd_sc_hd__o31ai_1 _1465_ (.A1(net120),
    .A2(_0145_),
    .A3(_0641_),
    .B1(net109),
    .Y(_0642_));
 sky130_fd_sc_hd__a21oi_1 _1466_ (.A1(_0474_),
    .A2(_0489_),
    .B1(net79),
    .Y(_0643_));
 sky130_fd_sc_hd__o21ai_1 _1467_ (.A1(_0642_),
    .A2(_0643_),
    .B1(_0640_),
    .Y(_0644_));
 sky130_fd_sc_hd__o211a_1 _1468_ (.A1(_0039_),
    .A2(net53),
    .B1(_0212_),
    .C1(net80),
    .X(_0645_));
 sky130_fd_sc_hd__a31o_1 _1469_ (.A1(net123),
    .A2(_0290_),
    .A3(_0387_),
    .B1(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__or3_1 _1470_ (.A(net121),
    .B(_0062_),
    .C(_0479_),
    .X(_0647_));
 sky130_fd_sc_hd__a21o_1 _1471_ (.A1(_0122_),
    .A2(_0171_),
    .B1(net79),
    .X(_0648_));
 sky130_fd_sc_hd__a31oi_1 _1472_ (.A1(net101),
    .A2(_0647_),
    .A3(_0648_),
    .B1(_0092_),
    .Y(_0649_));
 sky130_fd_sc_hd__a21o_1 _1473_ (.A1(net110),
    .A2(_0646_),
    .B1(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__a21oi_1 _1474_ (.A1(_0644_),
    .A2(_0650_),
    .B1(net93),
    .Y(_0651_));
 sky130_fd_sc_hd__o211a_1 _1475_ (.A1(net134),
    .A2(_0124_),
    .B1(_0484_),
    .C1(net123),
    .X(_0653_));
 sky130_fd_sc_hd__o21ai_1 _1476_ (.A1(_0642_),
    .A2(_0653_),
    .B1(_0640_),
    .Y(_0654_));
 sky130_fd_sc_hd__a31o_1 _1477_ (.A1(net123),
    .A2(_0086_),
    .A3(_0290_),
    .B1(_0645_),
    .X(_0655_));
 sky130_fd_sc_hd__a21o_1 _1478_ (.A1(net110),
    .A2(_0655_),
    .B1(_0649_),
    .X(_0656_));
 sky130_fd_sc_hd__a31o_1 _1479_ (.A1(net93),
    .A2(_0654_),
    .A3(_0656_),
    .B1(net171),
    .X(_0657_));
 sky130_fd_sc_hd__o22a_1 _1480_ (.A1(net176),
    .A2(net187),
    .B1(_0651_),
    .B2(_0657_),
    .X(_0020_));
 sky130_fd_sc_hd__a21oi_2 _1481_ (.A1(net70),
    .A2(_0124_),
    .B1(net75),
    .Y(_0658_));
 sky130_fd_sc_hd__o211ai_2 _1482_ (.A1(net135),
    .A2(_0123_),
    .B1(_0242_),
    .C1(net121),
    .Y(_0659_));
 sky130_fd_sc_hd__a21o_1 _1483_ (.A1(_0161_),
    .A2(_0184_),
    .B1(net125),
    .X(_0660_));
 sky130_fd_sc_hd__a31o_1 _1484_ (.A1(net89),
    .A2(_0659_),
    .A3(_0660_),
    .B1(_0342_),
    .X(_0661_));
 sky130_fd_sc_hd__a31o_1 _1485_ (.A1(_0806_),
    .A2(_0038_),
    .A3(_0137_),
    .B1(net127),
    .X(_0663_));
 sky130_fd_sc_hd__o21a_1 _1486_ (.A1(_0106_),
    .A2(_0453_),
    .B1(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__o21ai_1 _1487_ (.A1(net85),
    .A2(_0664_),
    .B1(_0661_),
    .Y(_0665_));
 sky130_fd_sc_hd__o32a_1 _1488_ (.A1(net72),
    .A2(net66),
    .A3(_0798_),
    .B1(_0801_),
    .B2(_0046_),
    .X(_0666_));
 sky130_fd_sc_hd__o22a_1 _1489_ (.A1(_0295_),
    .A2(_0542_),
    .B1(_0666_),
    .B2(net117),
    .X(_0667_));
 sky130_fd_sc_hd__nor2_1 _1490_ (.A(_0047_),
    .B(_0251_),
    .Y(_0668_));
 sky130_fd_sc_hd__o221a_1 _1491_ (.A1(net107),
    .A2(_0667_),
    .B1(_0668_),
    .B2(_0127_),
    .C1(net99),
    .X(_0669_));
 sky130_fd_sc_hd__or4_1 _1492_ (.A(_0801_),
    .B(net61),
    .C(_0043_),
    .D(net57),
    .X(_0670_));
 sky130_fd_sc_hd__nand2_1 _1493_ (.A(_0669_),
    .B(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__a21oi_1 _1494_ (.A1(_0665_),
    .A2(_0671_),
    .B1(net91),
    .Y(_0672_));
 sky130_fd_sc_hd__o31a_1 _1495_ (.A1(_0805_),
    .A2(_0102_),
    .A3(_0453_),
    .B1(_0663_),
    .X(_0674_));
 sky130_fd_sc_hd__o21ai_1 _1496_ (.A1(net85),
    .A2(_0674_),
    .B1(_0661_),
    .Y(_0675_));
 sky130_fd_sc_hd__nor2_1 _1497_ (.A(net47),
    .B(_0335_),
    .Y(_0676_));
 sky130_fd_sc_hd__o21ai_1 _1498_ (.A1(net57),
    .A2(_0676_),
    .B1(_0669_),
    .Y(_0677_));
 sky130_fd_sc_hd__a31o_1 _1499_ (.A1(net91),
    .A2(_0675_),
    .A3(_0677_),
    .B1(net170),
    .X(_0678_));
 sky130_fd_sc_hd__o22a_1 _1500_ (.A1(net174),
    .A2(net180),
    .B1(_0672_),
    .B2(_0678_),
    .X(_0021_));
 sky130_fd_sc_hd__a21o_1 _1501_ (.A1(_0304_),
    .A2(_0496_),
    .B1(net122),
    .X(_0679_));
 sky130_fd_sc_hd__a31o_1 _1502_ (.A1(net71),
    .A2(_0796_),
    .A3(_0033_),
    .B1(net80),
    .X(_0680_));
 sky130_fd_sc_hd__a31o_1 _1503_ (.A1(net101),
    .A2(_0679_),
    .A3(_0680_),
    .B1(_0092_),
    .X(_0681_));
 sky130_fd_sc_hd__o31a_1 _1504_ (.A1(net83),
    .A2(_0232_),
    .A3(_0317_),
    .B1(net58),
    .X(_0682_));
 sky130_fd_sc_hd__nor2_1 _1505_ (.A(_0309_),
    .B(_0335_),
    .Y(_0684_));
 sky130_fd_sc_hd__o21ai_1 _1506_ (.A1(_0682_),
    .A2(_0684_),
    .B1(_0681_),
    .Y(_0685_));
 sky130_fd_sc_hd__o32a_1 _1507_ (.A1(net142),
    .A2(_0787_),
    .A3(net55),
    .B1(net52),
    .B2(_0808_),
    .X(_0686_));
 sky130_fd_sc_hd__o221a_1 _1508_ (.A1(net150),
    .A2(_0736_),
    .B1(_0183_),
    .B2(net72),
    .C1(net81),
    .X(_0687_));
 sky130_fd_sc_hd__a21o_1 _1509_ (.A1(net127),
    .A2(_0686_),
    .B1(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__o21ai_1 _1510_ (.A1(net135),
    .A2(_0183_),
    .B1(_0387_),
    .Y(_0689_));
 sky130_fd_sc_hd__a221o_1 _1511_ (.A1(net83),
    .A2(_0688_),
    .B1(_0689_),
    .B2(_0126_),
    .C1(net101),
    .X(_0690_));
 sky130_fd_sc_hd__o21a_1 _1512_ (.A1(_0323_),
    .A2(_0457_),
    .B1(net42),
    .X(_0691_));
 sky130_fd_sc_hd__o211a_1 _1513_ (.A1(_0690_),
    .A2(_0691_),
    .B1(net96),
    .C1(_0685_),
    .X(_0692_));
 sky130_fd_sc_hd__a21o_1 _1514_ (.A1(_0184_),
    .A2(_0308_),
    .B1(_0682_),
    .X(_0693_));
 sky130_fd_sc_hd__and3_1 _1515_ (.A(net42),
    .B(_0210_),
    .C(_0233_),
    .X(_0695_));
 sky130_fd_sc_hd__a2bb2o_1 _1516_ (.A1_N(_0690_),
    .A2_N(_0695_),
    .B1(_0693_),
    .B2(_0681_),
    .X(_0696_));
 sky130_fd_sc_hd__a21o_1 _1517_ (.A1(_0652_),
    .A2(_0696_),
    .B1(net171),
    .X(_0697_));
 sky130_fd_sc_hd__o22a_1 _1518_ (.A1(net176),
    .A2(net181),
    .B1(_0692_),
    .B2(_0697_),
    .X(_0022_));
 sky130_fd_sc_hd__a21o_1 _1519_ (.A1(net151),
    .A2(_0767_),
    .B1(net141),
    .X(_0698_));
 sky130_fd_sc_hd__a21oi_1 _1520_ (.A1(_0715_),
    .A2(_0128_),
    .B1(net125),
    .Y(_0699_));
 sky130_fd_sc_hd__a22o_1 _1521_ (.A1(net129),
    .A2(_0044_),
    .B1(_0698_),
    .B2(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__o21ai_1 _1522_ (.A1(net111),
    .A2(_0700_),
    .B1(net102),
    .Y(_0701_));
 sky130_fd_sc_hd__a211o_1 _1523_ (.A1(_0033_),
    .A2(_0043_),
    .B1(_0141_),
    .C1(net123),
    .X(_0702_));
 sky130_fd_sc_hd__nand2b_1 _1524_ (.A_N(_0680_),
    .B(_0387_),
    .Y(_0703_));
 sky130_fd_sc_hd__a21oi_1 _1525_ (.A1(_0702_),
    .A2(_0703_),
    .B1(net87),
    .Y(_0705_));
 sky130_fd_sc_hd__o221a_1 _1526_ (.A1(_0808_),
    .A2(_0117_),
    .B1(_0158_),
    .B2(net52),
    .C1(net126),
    .X(_0706_));
 sky130_fd_sc_hd__o211a_1 _1527_ (.A1(_0787_),
    .A2(_0224_),
    .B1(_0041_),
    .C1(net81),
    .X(_0707_));
 sky130_fd_sc_hd__o31a_1 _1528_ (.A1(net102),
    .A2(_0706_),
    .A3(_0707_),
    .B1(_0343_),
    .X(_0708_));
 sky130_fd_sc_hd__nor2_1 _1529_ (.A(_0127_),
    .B(_0277_),
    .Y(_0709_));
 sky130_fd_sc_hd__o211a_1 _1530_ (.A1(_0058_),
    .A2(_0246_),
    .B1(_0177_),
    .C1(net43),
    .X(_0710_));
 sky130_fd_sc_hd__o32a_1 _1531_ (.A1(_0708_),
    .A2(_0709_),
    .A3(_0710_),
    .B1(_0705_),
    .B2(_0701_),
    .X(_0711_));
 sky130_fd_sc_hd__nor2_1 _1532_ (.A(net94),
    .B(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__nand2_1 _1533_ (.A(_0128_),
    .B(_0184_),
    .Y(_0713_));
 sky130_fd_sc_hd__o21ai_1 _1534_ (.A1(net141),
    .A2(_0248_),
    .B1(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__a211o_1 _1535_ (.A1(net43),
    .A2(_0714_),
    .B1(_0709_),
    .C1(_0708_),
    .X(_0716_));
 sky130_fd_sc_hd__o21ai_1 _1536_ (.A1(_0085_),
    .A2(_0680_),
    .B1(_0702_),
    .Y(_0717_));
 sky130_fd_sc_hd__a21o_1 _1537_ (.A1(net111),
    .A2(_0717_),
    .B1(_0701_),
    .X(_0718_));
 sky130_fd_sc_hd__a31o_1 _1538_ (.A1(net94),
    .A2(_0716_),
    .A3(_0718_),
    .B1(net172),
    .X(_0719_));
 sky130_fd_sc_hd__o22a_1 _1539_ (.A1(net175),
    .A2(net179),
    .B1(_0712_),
    .B2(_0719_),
    .X(_0023_));
 sky130_fd_sc_hd__nor2_1 _1540_ (.A(net125),
    .B(_0676_),
    .Y(_0720_));
 sky130_fd_sc_hd__a211o_1 _1541_ (.A1(_0086_),
    .A2(_0658_),
    .B1(_0720_),
    .C1(net112),
    .X(_0721_));
 sky130_fd_sc_hd__a21oi_1 _1542_ (.A1(net77),
    .A2(_0129_),
    .B1(net85),
    .Y(_0722_));
 sky130_fd_sc_hd__a21bo_1 _1543_ (.A1(_0044_),
    .A2(_0277_),
    .B1_N(_0722_),
    .X(_0723_));
 sky130_fd_sc_hd__o2111ai_2 _1544_ (.A1(_0127_),
    .A2(_0249_),
    .B1(_0721_),
    .C1(_0723_),
    .D1(net99),
    .Y(_0724_));
 sky130_fd_sc_hd__o211a_1 _1545_ (.A1(net61),
    .A2(_0698_),
    .B1(_0410_),
    .C1(net125),
    .X(_0726_));
 sky130_fd_sc_hd__a311oi_1 _1546_ (.A1(net81),
    .A2(_0044_),
    .A3(_0277_),
    .B1(_0726_),
    .C1(net112),
    .Y(_0727_));
 sky130_fd_sc_hd__a21o_1 _1547_ (.A1(_0161_),
    .A2(_0184_),
    .B1(net77),
    .X(_0728_));
 sky130_fd_sc_hd__o311a_1 _1548_ (.A1(net125),
    .A2(_0040_),
    .A3(_0479_),
    .B1(_0728_),
    .C1(net107),
    .X(_0729_));
 sky130_fd_sc_hd__or3_1 _1549_ (.A(net99),
    .B(_0727_),
    .C(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__and3_1 _1550_ (.A(net118),
    .B(net137),
    .C(_0183_),
    .X(_0731_));
 sky130_fd_sc_hd__nand2_1 _1551_ (.A(net117),
    .B(_0185_),
    .Y(_0732_));
 sky130_fd_sc_hd__nor2_1 _1552_ (.A(net91),
    .B(_0731_),
    .Y(_0733_));
 sky130_fd_sc_hd__a21oi_1 _1553_ (.A1(_0724_),
    .A2(_0730_),
    .B1(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__a31o_1 _1554_ (.A1(_0652_),
    .A2(_0724_),
    .A3(_0730_),
    .B1(net170),
    .X(_0735_));
 sky130_fd_sc_hd__a2bb2o_1 _1555_ (.A1_N(_0735_),
    .A2_N(_0734_),
    .B1(net196),
    .B2(net170),
    .X(_0024_));
 sky130_fd_sc_hd__and2_1 _1556_ (.A(net170),
    .B(net208),
    .X(_0737_));
 sky130_fd_sc_hd__a32o_1 _1557_ (.A1(_0240_),
    .A2(_0349_),
    .A3(_0556_),
    .B1(_0226_),
    .B2(net74),
    .X(_0738_));
 sky130_fd_sc_hd__o21ai_1 _1558_ (.A1(net103),
    .A2(_0738_),
    .B1(net97),
    .Y(_0739_));
 sky130_fd_sc_hd__nand2_1 _1559_ (.A(_0803_),
    .B(_0804_),
    .Y(_0740_));
 sky130_fd_sc_hd__a41o_1 _1560_ (.A1(net109),
    .A2(_0090_),
    .A3(_0233_),
    .A4(_0740_),
    .B1(net42),
    .X(_0741_));
 sky130_fd_sc_hd__o31ai_1 _1561_ (.A1(net70),
    .A2(net56),
    .A3(_0117_),
    .B1(_0658_),
    .Y(_0742_));
 sky130_fd_sc_hd__a21oi_1 _1562_ (.A1(_0741_),
    .A2(_0742_),
    .B1(_0739_),
    .Y(_0743_));
 sky130_fd_sc_hd__a21o_1 _1563_ (.A1(_0044_),
    .A2(_0525_),
    .B1(net114),
    .X(_0744_));
 sky130_fd_sc_hd__a21oi_1 _1564_ (.A1(net114),
    .A2(_0188_),
    .B1(_0442_),
    .Y(_0745_));
 sky130_fd_sc_hd__nand2_1 _1565_ (.A(_0744_),
    .B(_0745_),
    .Y(_0747_));
 sky130_fd_sc_hd__nand2_1 _1566_ (.A(net115),
    .B(_0372_),
    .Y(_0748_));
 sky130_fd_sc_hd__o32a_1 _1567_ (.A1(net114),
    .A2(_0113_),
    .A3(_0479_),
    .B1(_0522_),
    .B2(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__nor2_1 _1568_ (.A(net98),
    .B(net107),
    .Y(_0750_));
 sky130_fd_sc_hd__o31ai_1 _1569_ (.A1(net97),
    .A2(net103),
    .A3(_0749_),
    .B1(net92),
    .Y(_0751_));
 sky130_fd_sc_hd__a211o_1 _1570_ (.A1(_0342_),
    .A2(_0747_),
    .B1(_0751_),
    .C1(_0743_),
    .X(_0752_));
 sky130_fd_sc_hd__o21ai_1 _1571_ (.A1(net60),
    .A2(_0087_),
    .B1(_0658_),
    .Y(_0753_));
 sky130_fd_sc_hd__a211o_1 _1572_ (.A1(_0741_),
    .A2(_0753_),
    .B1(net92),
    .C1(_0739_),
    .X(_0754_));
 sky130_fd_sc_hd__a21o_1 _1573_ (.A1(net84),
    .A2(_0749_),
    .B1(_0176_),
    .X(_0755_));
 sky130_fd_sc_hd__a31o_1 _1574_ (.A1(net104),
    .A2(_0431_),
    .A3(_0744_),
    .B1(_0755_),
    .X(_0756_));
 sky130_fd_sc_hd__a41o_1 _1575_ (.A1(net173),
    .A2(_0752_),
    .A3(_0754_),
    .A4(_0756_),
    .B1(_0737_),
    .X(_0025_));
 sky130_fd_sc_hd__and2_1 _1576_ (.A(net170),
    .B(net207),
    .X(_0758_));
 sky130_fd_sc_hd__and4_1 _1577_ (.A(net76),
    .B(net137),
    .C(net147),
    .D(net156),
    .X(_0759_));
 sky130_fd_sc_hd__o21a_1 _1578_ (.A1(_0045_),
    .A2(_0272_),
    .B1(net119),
    .X(_0760_));
 sky130_fd_sc_hd__or3_1 _1579_ (.A(net107),
    .B(_0759_),
    .C(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__nor2_1 _1580_ (.A(net76),
    .B(_0623_),
    .Y(_0762_));
 sky130_fd_sc_hd__o21a_1 _1581_ (.A1(_0804_),
    .A2(net49),
    .B1(_0515_),
    .X(_0763_));
 sky130_fd_sc_hd__o311a_1 _1582_ (.A1(net85),
    .A2(_0762_),
    .A3(_0763_),
    .B1(_0761_),
    .C1(net98),
    .X(_0764_));
 sky130_fd_sc_hd__or4_1 _1583_ (.A(_0040_),
    .B(net57),
    .C(_0095_),
    .D(_0188_),
    .X(_0765_));
 sky130_fd_sc_hd__o21ai_1 _1584_ (.A1(_0098_),
    .A2(_0296_),
    .B1(_0126_),
    .Y(_0766_));
 sky130_fd_sc_hd__a21oi_1 _1585_ (.A1(_0765_),
    .A2(_0766_),
    .B1(net98),
    .Y(_0768_));
 sky130_fd_sc_hd__and3_1 _1586_ (.A(net119),
    .B(_0146_),
    .C(_0525_),
    .X(_0769_));
 sky130_fd_sc_hd__and4_1 _1587_ (.A(net76),
    .B(_0104_),
    .C(_0115_),
    .D(_0556_),
    .X(_0770_));
 sky130_fd_sc_hd__o21a_1 _1588_ (.A1(_0769_),
    .A2(_0770_),
    .B1(_0750_),
    .X(_0771_));
 sky130_fd_sc_hd__or4_1 _1589_ (.A(net90),
    .B(_0764_),
    .C(_0768_),
    .D(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__o32ai_1 _1590_ (.A1(_0764_),
    .A2(_0768_),
    .A3(_0771_),
    .B1(_0731_),
    .B2(net90),
    .Y(_0773_));
 sky130_fd_sc_hd__a31o_1 _1591_ (.A1(net174),
    .A2(_0772_),
    .A3(_0773_),
    .B1(_0758_),
    .X(_0026_));
 sky130_fd_sc_hd__nand2_1 _1592_ (.A(_0046_),
    .B(_0186_),
    .Y(_0774_));
 sky130_fd_sc_hd__a31o_1 _1593_ (.A1(_0046_),
    .A2(_0165_),
    .A3(_0713_),
    .B1(net125),
    .X(_0775_));
 sky130_fd_sc_hd__o211a_1 _1594_ (.A1(_0296_),
    .A2(_0774_),
    .B1(_0775_),
    .C1(_0750_),
    .X(_0776_));
 sky130_fd_sc_hd__a21oi_1 _1595_ (.A1(net117),
    .A2(_0437_),
    .B1(net107),
    .Y(_0778_));
 sky130_fd_sc_hd__a31o_1 _1596_ (.A1(_0046_),
    .A2(_0129_),
    .A3(_0165_),
    .B1(net57),
    .X(_0779_));
 sky130_fd_sc_hd__o311a_1 _1597_ (.A1(_0045_),
    .A2(_0722_),
    .A3(_0778_),
    .B1(_0779_),
    .C1(net99),
    .X(_0780_));
 sky130_fd_sc_hd__o311a_1 _1598_ (.A1(net117),
    .A2(_0047_),
    .A3(_0296_),
    .B1(_0342_),
    .C1(_0732_),
    .X(_0781_));
 sky130_fd_sc_hd__o31a_1 _1599_ (.A1(_0776_),
    .A2(_0780_),
    .A3(_0781_),
    .B1(_0652_),
    .X(_0782_));
 sky130_fd_sc_hd__nor2_1 _1600_ (.A(net91),
    .B(_0185_),
    .Y(_0783_));
 sky130_fd_sc_hd__or4_1 _1601_ (.A(_0776_),
    .B(_0780_),
    .C(_0781_),
    .D(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__nand2_1 _1602_ (.A(net174),
    .B(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__a2bb2o_1 _1603_ (.A1_N(_0785_),
    .A2_N(_0782_),
    .B1(net195),
    .B2(net172),
    .X(_0027_));
 sky130_fd_sc_hd__o211a_1 _1604_ (.A1(net118),
    .A2(_0048_),
    .B1(_0342_),
    .C1(_0732_),
    .X(_0786_));
 sky130_fd_sc_hd__o211a_1 _1605_ (.A1(net76),
    .A2(_0437_),
    .B1(net98),
    .C1(net85),
    .X(_0788_));
 sky130_fd_sc_hd__o2111a_1 _1606_ (.A1(net118),
    .A2(_0128_),
    .B1(_0343_),
    .C1(_0774_),
    .D1(_0110_),
    .X(_0789_));
 sky130_fd_sc_hd__or3_1 _1607_ (.A(_0786_),
    .B(_0788_),
    .C(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__a21oi_1 _1608_ (.A1(net43),
    .A2(_0185_),
    .B1(net91),
    .Y(_0791_));
 sky130_fd_sc_hd__mux2_1 _1609_ (.A0(_0791_),
    .A1(net90),
    .S(_0790_),
    .X(_0792_));
 sky130_fd_sc_hd__mux2_1 _1610_ (.A0(net186),
    .A1(_0792_),
    .S(net174),
    .X(_0028_));
 sky130_fd_sc_hd__nor2_1 _1611_ (.A(_0343_),
    .B(_0732_),
    .Y(_0793_));
 sky130_fd_sc_hd__a221o_1 _1612_ (.A1(net98),
    .A2(_0722_),
    .B1(_0750_),
    .B2(_0774_),
    .C1(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _1613_ (.A0(net91),
    .A1(_0733_),
    .S(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__mux2_1 _1614_ (.A0(net194),
    .A1(_0795_),
    .S(net174),
    .X(_0029_));
 sky130_fd_sc_hd__or2_1 _1615_ (.A(net172),
    .B(_0791_),
    .X(_0797_));
 sky130_fd_sc_hd__o22a_1 _1616_ (.A1(net174),
    .A2(net189),
    .B1(_0793_),
    .B2(_0797_),
    .X(_0030_));
 sky130_fd_sc_hd__o22a_1 _1617_ (.A1(net9),
    .A2(net191),
    .B1(_0559_),
    .B2(_0791_),
    .X(_0031_));
 sky130_fd_sc_hd__dfxtp_1 _1618_ (.CLK(clknet_2_0__leaf_clk0),
    .D(_0000_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_1 _1619_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0001_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_1 _1620_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0002_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _1621_ (.CLK(clknet_2_0__leaf_clk0),
    .D(_0003_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _1622_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0004_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _1623_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0005_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _1624_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0006_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _1625_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0007_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _1626_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0008_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _1627_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0009_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _1628_ (.CLK(clknet_2_0__leaf_clk0),
    .D(_0010_),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_1 _1629_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0011_),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_1 _1630_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0012_),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_1 _1631_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0013_),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_1 _1632_ (.CLK(clknet_2_0__leaf_clk0),
    .D(_0014_),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_1 _1633_ (.CLK(clknet_2_0__leaf_clk0),
    .D(_0015_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_1 _1634_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0016_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_1 _1635_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0017_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_1 _1636_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0018_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_1 _1637_ (.CLK(clknet_2_0__leaf_clk0),
    .D(_0019_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_1 _1638_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0020_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_1 _1639_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0021_),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_1 _1640_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0022_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_1 _1641_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0023_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_1 _1642_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0024_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_1 _1643_ (.CLK(clknet_2_0__leaf_clk0),
    .D(_0025_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_1 _1644_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0026_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _1645_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0027_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_1 _1646_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0028_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _1647_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0029_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _1648_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0030_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _1649_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0031_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _1650_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net1),
    .Q(\addr0_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1651_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net2),
    .Q(\addr0_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1652_ (.CLK(clknet_2_1__leaf_clk0),
    .D(net3),
    .Q(\addr0_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1653_ (.CLK(clknet_2_1__leaf_clk0),
    .D(net4),
    .Q(\addr0_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1654_ (.CLK(clknet_2_1__leaf_clk0),
    .D(net5),
    .Q(\addr0_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _1655_ (.CLK(clknet_2_1__leaf_clk0),
    .D(net6),
    .Q(\addr0_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1656_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net7),
    .Q(\addr0_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1657_ (.CLK(clknet_2_1__leaf_clk0),
    .D(net8),
    .Q(\addr0_reg[7] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_373 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(addr0[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(addr0[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(addr0[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(addr0[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(addr0[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(addr0[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(addr0[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(addr0[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(cs0),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(dout0[0]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(dout0[10]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(dout0[11]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(dout0[12]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(dout0[13]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(dout0[14]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(dout0[15]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(dout0[16]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(dout0[17]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(dout0[18]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(dout0[19]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(dout0[1]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(dout0[20]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(dout0[21]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(dout0[22]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(dout0[23]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(dout0[24]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(dout0[25]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(dout0[26]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(dout0[27]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(dout0[28]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(dout0[29]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(dout0[2]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(dout0[30]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(dout0[31]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(dout0[3]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(dout0[4]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(dout0[5]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(dout0[6]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(dout0[7]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(dout0[8]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(dout0[9]));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(_0053_),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 fanout43 (.A(_0053_),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 max_cap44 (.A(_0118_),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 max_cap45 (.A(_0103_),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(_0083_),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 fanout47 (.A(_0083_),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 fanout48 (.A(_0070_),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 fanout49 (.A(_0070_),
    .X(net49));
 sky130_fd_sc_hd__buf_4 fanout50 (.A(_0069_),
    .X(net50));
 sky130_fd_sc_hd__buf_4 fanout51 (.A(_0061_),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 fanout52 (.A(_0061_),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 fanout53 (.A(_0060_),
    .X(net53));
 sky130_fd_sc_hd__buf_2 fanout54 (.A(_0060_),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 fanout56 (.A(_0058_),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 fanout57 (.A(_0054_),
    .X(net57));
 sky130_fd_sc_hd__buf_2 fanout58 (.A(_0054_),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 fanout59 (.A(_0036_),
    .X(net59));
 sky130_fd_sc_hd__buf_2 fanout60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__buf_4 fanout61 (.A(_0034_),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(_0033_),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net64),
    .X(net63));
 sky130_fd_sc_hd__buf_2 fanout64 (.A(_0032_),
    .X(net64));
 sky130_fd_sc_hd__buf_4 fanout65 (.A(_0799_),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 fanout66 (.A(_0787_),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 fanout68 (.A(_0777_),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_4 fanout69 (.A(_0767_),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 fanout71 (.A(net72),
    .X(net71));
 sky130_fd_sc_hd__buf_4 fanout72 (.A(_0694_),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 fanout73 (.A(_0694_),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 fanout74 (.A(net78),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_4 fanout75 (.A(net78),
    .X(net75));
 sky130_fd_sc_hd__buf_2 fanout76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_4 fanout77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 fanout78 (.A(_0683_),
    .X(net78));
 sky130_fd_sc_hd__buf_2 fanout79 (.A(net80),
    .X(net79));
 sky130_fd_sc_hd__buf_2 fanout80 (.A(_0683_),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 fanout81 (.A(_0683_),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 fanout82 (.A(_0683_),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 fanout83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 fanout84 (.A(net87),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 fanout85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 fanout87 (.A(_0673_),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 fanout88 (.A(_0662_),
    .X(net88));
 sky130_fd_sc_hd__buf_2 fanout89 (.A(_0662_),
    .X(net89));
 sky130_fd_sc_hd__buf_2 fanout90 (.A(net96),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 fanout91 (.A(net96),
    .X(net91));
 sky130_fd_sc_hd__buf_2 fanout92 (.A(net96),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 fanout93 (.A(net96),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_4 fanout94 (.A(net96),
    .X(net94));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_4 fanout96 (.A(\addr0_reg[7] ),
    .X(net96));
 sky130_fd_sc_hd__buf_2 fanout97 (.A(net100),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 fanout98 (.A(net100),
    .X(net98));
 sky130_fd_sc_hd__buf_2 fanout99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 fanout100 (.A(\addr0_reg[6] ),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_4 fanout101 (.A(\addr0_reg[6] ),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_4 fanout102 (.A(\addr0_reg[6] ),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 fanout103 (.A(net106),
    .X(net103));
 sky130_fd_sc_hd__buf_2 fanout104 (.A(net106),
    .X(net104));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 fanout106 (.A(net108),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 fanout107 (.A(net108),
    .X(net107));
 sky130_fd_sc_hd__buf_2 fanout108 (.A(\addr0_reg[5] ),
    .X(net108));
 sky130_fd_sc_hd__buf_2 fanout109 (.A(\addr0_reg[5] ),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 fanout110 (.A(\addr0_reg[5] ),
    .X(net110));
 sky130_fd_sc_hd__buf_2 fanout111 (.A(net113),
    .X(net111));
 sky130_fd_sc_hd__buf_2 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 fanout113 (.A(\addr0_reg[5] ),
    .X(net113));
 sky130_fd_sc_hd__buf_2 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__buf_2 fanout115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__buf_2 fanout116 (.A(net119),
    .X(net116));
 sky130_fd_sc_hd__buf_2 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__buf_2 fanout118 (.A(net119),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 fanout119 (.A(\addr0_reg[4] ),
    .X(net119));
 sky130_fd_sc_hd__buf_2 fanout120 (.A(net122),
    .X(net120));
 sky130_fd_sc_hd__buf_2 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__buf_2 fanout122 (.A(net124),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_4 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 fanout124 (.A(\addr0_reg[4] ),
    .X(net124));
 sky130_fd_sc_hd__buf_2 fanout125 (.A(net129),
    .X(net125));
 sky130_fd_sc_hd__buf_2 fanout126 (.A(net129),
    .X(net126));
 sky130_fd_sc_hd__buf_2 fanout127 (.A(net129),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 fanout129 (.A(\addr0_reg[4] ),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(net132),
    .X(net130));
 sky130_fd_sc_hd__buf_2 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(\addr0_reg[3] ),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_4 fanout135 (.A(\addr0_reg[3] ),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 fanout136 (.A(net143),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(net138),
    .X(net137));
 sky130_fd_sc_hd__buf_2 fanout138 (.A(net143),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__buf_2 fanout140 (.A(net141),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_2 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__buf_2 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 fanout143 (.A(\addr0_reg[3] ),
    .X(net143));
 sky130_fd_sc_hd__buf_4 fanout144 (.A(net152),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 fanout145 (.A(net152),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_4 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__buf_2 fanout147 (.A(net152),
    .X(net147));
 sky130_fd_sc_hd__buf_4 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 fanout149 (.A(net152),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__buf_2 fanout151 (.A(net152),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 fanout152 (.A(\addr0_reg[2] ),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_8 fanout153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__buf_2 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 fanout155 (.A(\addr0_reg[1] ),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__buf_2 fanout157 (.A(\addr0_reg[1] ),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__buf_2 fanout159 (.A(net161),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_4 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__buf_2 fanout161 (.A(\addr0_reg[1] ),
    .X(net161));
 sky130_fd_sc_hd__buf_4 fanout162 (.A(net169),
    .X(net162));
 sky130_fd_sc_hd__buf_1 fanout163 (.A(net169),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_4 fanout164 (.A(net169),
    .X(net164));
 sky130_fd_sc_hd__buf_4 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout166 (.A(net169),
    .X(net166));
 sky130_fd_sc_hd__buf_4 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_4 fanout169 (.A(\addr0_reg[0] ),
    .X(net169));
 sky130_fd_sc_hd__buf_2 fanout170 (.A(net172),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_4 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 fanout172 (.A(_0725_),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_4 fanout174 (.A(net9),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_4 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_4 fanout176 (.A(net9),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk0 (.A(clk0),
    .X(clknet_0_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_0__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_1__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_2__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_3__leaf_clk0));
 sky130_fd_sc_hd__bufinv_16 clkload0 (.A(clknet_2_0__leaf_clk0));
 sky130_fd_sc_hd__clkinv_4 clkload1 (.A(clknet_2_2__leaf_clk0));
 sky130_fd_sc_hd__clkinv_4 clkload2 (.A(clknet_2_3__leaf_clk0));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net37),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net32),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net25),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net23),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net24),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net13),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net20),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net40),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net35),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net30),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net22),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net14),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net33),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net15),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net34),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net11),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net12),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net31),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net29),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net26),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net39),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net18),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net17),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net21),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net36),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net10),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net41),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net19),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net38),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net16),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net28),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net27),
    .X(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0044_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0065_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0658_));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
endmodule
