VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rom5
  CLASS BLOCK ;
  FOREIGN rom5 ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 236.880 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 236.880 ;
    END
  END VPWR
  PIN addr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 34.040 250.000 34.640 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 246.000 37.440 250.000 38.040 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 40.840 250.000 41.440 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 44.240 250.000 44.840 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 47.640 250.000 48.240 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END addr0[8]
  PIN clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END clk0
  PIN dout0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 119.040 250.000 119.640 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 142.840 250.000 143.440 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 109.570 246.000 109.850 250.000 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 128.890 246.000 129.170 250.000 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 151.430 246.000 151.710 250.000 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 170.750 246.000 171.030 250.000 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 67.710 246.000 67.990 250.000 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 199.730 246.000 200.010 250.000 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 144.990 246.000 145.270 250.000 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 96.690 246.000 96.970 250.000 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 77.370 246.000 77.650 250.000 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.950 246.000 42.230 250.000 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 64.490 246.000 64.770 250.000 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 51.610 246.000 51.890 250.000 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 81.640 250.000 82.240 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END dout0[31]
  PIN dout0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END dout0[3]
  PIN dout0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 246.000 98.640 250.000 99.240 ;
    END
  END dout0[4]
  PIN dout0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END dout0[5]
  PIN dout0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END dout0[9]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 244.450 236.830 ;
      LAYER li1 ;
        RECT 5.520 10.795 244.260 236.725 ;
      LAYER met1 ;
        RECT 1.450 6.160 248.330 242.380 ;
      LAYER met2 ;
        RECT 1.470 245.720 41.670 246.685 ;
        RECT 42.510 245.720 51.330 246.685 ;
        RECT 52.170 245.720 64.210 246.685 ;
        RECT 65.050 245.720 67.430 246.685 ;
        RECT 68.270 245.720 77.090 246.685 ;
        RECT 77.930 245.720 96.410 246.685 ;
        RECT 97.250 245.720 109.290 246.685 ;
        RECT 110.130 245.720 128.610 246.685 ;
        RECT 129.450 245.720 144.710 246.685 ;
        RECT 145.550 245.720 151.150 246.685 ;
        RECT 151.990 245.720 170.470 246.685 ;
        RECT 171.310 245.720 199.450 246.685 ;
        RECT 200.290 245.720 248.310 246.685 ;
        RECT 1.470 4.280 248.310 245.720 ;
        RECT 1.470 4.000 35.230 4.280 ;
        RECT 36.070 4.000 83.530 4.280 ;
        RECT 84.370 4.000 118.950 4.280 ;
        RECT 119.790 4.000 122.170 4.280 ;
        RECT 123.010 4.000 144.710 4.280 ;
        RECT 145.550 4.000 157.590 4.280 ;
        RECT 158.430 4.000 173.690 4.280 ;
        RECT 174.530 4.000 248.310 4.280 ;
      LAYER met3 ;
        RECT 1.445 222.040 248.335 246.665 ;
        RECT 4.400 220.640 248.335 222.040 ;
        RECT 1.445 215.240 248.335 220.640 ;
        RECT 4.400 213.840 248.335 215.240 ;
        RECT 1.445 211.840 248.335 213.840 ;
        RECT 4.400 210.440 248.335 211.840 ;
        RECT 1.445 208.440 248.335 210.440 ;
        RECT 4.400 207.040 248.335 208.440 ;
        RECT 1.445 205.040 248.335 207.040 ;
        RECT 4.400 203.640 248.335 205.040 ;
        RECT 1.445 201.640 248.335 203.640 ;
        RECT 4.400 200.240 248.335 201.640 ;
        RECT 1.445 198.240 248.335 200.240 ;
        RECT 4.400 196.840 248.335 198.240 ;
        RECT 1.445 191.440 248.335 196.840 ;
        RECT 4.400 190.040 248.335 191.440 ;
        RECT 1.445 164.240 248.335 190.040 ;
        RECT 4.400 162.840 248.335 164.240 ;
        RECT 1.445 143.840 248.335 162.840 ;
        RECT 1.445 142.440 245.600 143.840 ;
        RECT 1.445 137.040 248.335 142.440 ;
        RECT 4.400 135.640 248.335 137.040 ;
        RECT 1.445 126.840 248.335 135.640 ;
        RECT 4.400 125.440 248.335 126.840 ;
        RECT 1.445 120.040 248.335 125.440 ;
        RECT 1.445 118.640 245.600 120.040 ;
        RECT 1.445 113.240 248.335 118.640 ;
        RECT 4.400 111.840 248.335 113.240 ;
        RECT 1.445 99.640 248.335 111.840 ;
        RECT 1.445 98.240 245.600 99.640 ;
        RECT 1.445 96.240 248.335 98.240 ;
        RECT 4.400 94.840 248.335 96.240 ;
        RECT 1.445 89.440 248.335 94.840 ;
        RECT 4.400 88.040 248.335 89.440 ;
        RECT 1.445 82.640 248.335 88.040 ;
        RECT 1.445 81.240 245.600 82.640 ;
        RECT 1.445 48.640 248.335 81.240 ;
        RECT 1.445 47.240 245.600 48.640 ;
        RECT 1.445 45.240 248.335 47.240 ;
        RECT 1.445 43.840 245.600 45.240 ;
        RECT 1.445 41.840 248.335 43.840 ;
        RECT 1.445 40.440 245.600 41.840 ;
        RECT 1.445 38.440 248.335 40.440 ;
        RECT 1.445 37.040 245.600 38.440 ;
        RECT 1.445 35.040 248.335 37.040 ;
        RECT 1.445 33.640 245.600 35.040 ;
        RECT 1.445 4.255 248.335 33.640 ;
      LAYER met4 ;
        RECT 2.135 237.280 245.345 246.665 ;
        RECT 2.135 10.240 20.640 237.280 ;
        RECT 23.040 10.240 23.940 237.280 ;
        RECT 26.340 10.240 174.240 237.280 ;
        RECT 176.640 10.240 177.540 237.280 ;
        RECT 179.940 10.240 245.345 237.280 ;
        RECT 2.135 4.255 245.345 10.240 ;
  END
END rom5
END LIBRARY

