logic [0:ROM_DEPTH-1] [DATA_WIDTH-1:0] table_ = {
32'h00000000,
32'h006487c4,
32'h00c90e90,
32'h012d936c,
32'h0192155f,
32'h01f69373,
32'h025b0caf,
32'h02bf801a,
32'h0323ecbe,
32'h038851a2,
32'h03ecadcf,
32'h0451004d,
32'h04b54825,
32'h0519845e,
32'h057db403,
32'h05e1d61b,
32'h0645e9af,
32'h06a9edc9,
32'h070de172,
32'h0771c3b3,
32'h07d59396,
32'h08395024,
32'h089cf867,
32'h09008b6a,
32'h09640837,
32'h09c76dd8,
32'h0a2abb59,
32'h0a8defc3,
32'h0af10a22,
32'h0b540982,
32'h0bb6ecef,
32'h0c19b374,
32'h0c7c5c1e,
32'h0cdee5f9,
32'h0d415013,
32'h0da39978,
32'h0e05c135,
32'h0e67c65a,
32'h0ec9a7f3,
32'h0f2b650f,
32'h0f8cfcbe,
32'h0fee6e0d,
32'h104fb80e,
32'h10b0d9d0,
32'h1111d263,
32'h1172a0d7,
32'h11d3443f,
32'h1233bbac,
32'h1294062f,
32'h12f422db,
32'h135410c3,
32'h13b3cefa,
32'h14135c94,
32'h1472b8a5,
32'h14d1e242,
32'h1530d881,
32'h158f9a76,
32'h15ee2738,
32'h164c7ddd,
32'h16aa9d7e,
32'h17088531,
32'h1766340f,
32'h17c3a931,
32'h1820e3b0,
32'h187de2a7,
32'h18daa52f,
32'h19372a64,
32'h19937161,
32'h19ef7944,
32'h1a4b4128,
32'h1aa6c82b,
32'h1b020d6c,
32'h1b5d100a,
32'h1bb7cf23,
32'h1c1249d8,
32'h1c6c7f4a,
32'h1cc66e99,
32'h1d2016e9,
32'h1d79775c,
32'h1dd28f15,
32'h1e2b5d38,
32'h1e83e0eb,
32'h1edc1953,
32'h1f340596,
32'h1f8ba4dc,
32'h1fe2f64c,
32'h2039f90f,
32'h2090ac4d,
32'h20e70f32,
32'h213d20e8,
32'h2192e09b,
32'h21e84d76,
32'h223d66a8,
32'h22922b5e,
32'h22e69ac8,
32'h233ab414,
32'h238e7673,
32'h23e1e117,
32'h2434f332,
32'h2487abf7,
32'h24da0a9a,
32'h252c0e4f,
32'h257db64c,
32'h25cf01c8,
32'h261feffa,
32'h2670801a,
32'h26c0b162,
32'h2710830c,
32'h275ff452,
32'h27af0472,
32'h27fdb2a7,
32'h284bfe2f,
32'h2899e64a,
32'h28e76a37,
32'h29348937,
32'h2981428c,
32'h29cd9578,
32'h2a19813f,
32'h2a650525,
32'h2ab02071,
32'h2afad269,
32'h2b451a55,
32'h2b8ef77d,
32'h2bd8692b,
32'h2c216eaa,
32'h2c6a0746,
32'h2cb2324c,
32'h2cf9ef09,
32'h2d413ccd,
32'h2d881ae8,
32'h2dce88aa,
32'h2e148566,
32'h2e5a1070,
32'h2e9f291b,
32'h2ee3cebe,
32'h2f2800af,
32'h2f6bbe45,
32'h2faf06da,
32'h2ff1d9c7,
32'h30343667,
32'h30761c18,
32'h30b78a36,
32'h30f8801f,
32'h3138fd35,
32'h317900d6,
32'h31b88a66,
32'h31f79948,
32'h32362ce0,
32'h32744493,
32'h32b1dfc9,
32'h32eefdea,
32'h332b9e5e,
32'h3367c090,
32'h33a363ec,
32'h33de87de,
32'h34192bd5,
32'h34534f41,
32'h348cf190,
32'h34c61236,
32'h34feb0a5,
32'h3536cc52,
32'h356e64b2,
32'h35a5793c,
32'h35dc0968,
32'h361214b0,
32'h36479a8e,
32'h367c9a7e,
32'h36b113fd,
32'h36e5068a,
32'h371871a5,
32'h374b54ce,
32'h377daf89,
32'h37af8159,
32'h37e0c9c3,
32'h3811884d,
32'h3841bc7f,
32'h387165e3,
32'h38a08402,
32'h38cf1669,
32'h38fd1ca4,
32'h392a9642,
32'h395782d3,
32'h3983e1e8,
32'h39afb313,
32'h39daf5e8,
32'h3a05a9fd,
32'h3a2fcee8,
32'h3a596442,
32'h3a8269a3,
32'h3aaadea6,
32'h3ad2c2e8,
32'h3afa1605,
32'h3b20d79e,
32'h3b470753,
32'h3b6ca4c4,
32'h3b91af97,
32'h3bb6276e,
32'h3bda0bf0,
32'h3bfd5cc4,
32'h3c201994,
32'h3c42420a,
32'h3c63d5d1,
32'h3c84d496,
32'h3ca53e09,
32'h3cc511d9,
32'h3ce44fb7,
32'h3d02f757,
32'h3d21086c,
32'h3d3e82ae,
32'h3d5b65d2,
32'h3d77b192,
32'h3d9365a8,
32'h3dae81cf,
32'h3dc905c5,
32'h3de2f148,
32'h3dfc4418,
32'h3e14fdf7,
32'h3e2d1ea8,
32'h3e44a5ef,
32'h3e5b9392,
32'h3e71e759,
32'h3e87a10c,
32'h3e9cc076,
32'h3eb14563,
32'h3ec52fa0,
32'h3ed87efc,
32'h3eeb3347,
32'h3efd4c54,
32'h3f0ec9f5,
32'h3f1fabff,
32'h3f2ff24a,
32'h3f3f9cab,
32'h3f4eaafe,
32'h3f5d1d1d,
32'h3f6af2e3,
32'h3f782c30,
32'h3f84c8e2,
32'h3f90c8da,
32'h3f9c2bfb,
32'h3fa6f228,
32'h3fb11b48,
32'h3fbaa740,
32'h3fc395f9,
32'h3fcbe75e,
32'h3fd39b5a,
32'h3fdab1d9,
32'h3fe12acb,
32'h3fe7061f,
32'h3fec43c7,
32'h3ff0e3b6,
32'h3ff4e5e0,
32'h3ff84a3c,
32'h3ffb10c1,
32'h3ffd3969,
32'h3ffec42d,
32'h3fffb10b,
32'h40000000,
32'h3fffb10b,
32'h3ffec42d,
32'h3ffd3969,
32'h3ffb10c1,
32'h3ff84a3c,
32'h3ff4e5e0,
32'h3ff0e3b6,
32'h3fec43c7,
32'h3fe7061f,
32'h3fe12acb,
32'h3fdab1d9,
32'h3fd39b5a,
32'h3fcbe75e,
32'h3fc395f9,
32'h3fbaa740,
32'h3fb11b48,
32'h3fa6f228,
32'h3f9c2bfb,
32'h3f90c8da,
32'h3f84c8e2,
32'h3f782c30,
32'h3f6af2e3,
32'h3f5d1d1d,
32'h3f4eaafe,
32'h3f3f9cab,
32'h3f2ff24a,
32'h3f1fabff,
32'h3f0ec9f5,
32'h3efd4c54,
32'h3eeb3347,
32'h3ed87efc,
32'h3ec52fa0,
32'h3eb14563,
32'h3e9cc076,
32'h3e87a10c,
32'h3e71e759,
32'h3e5b9392,
32'h3e44a5ef,
32'h3e2d1ea8,
32'h3e14fdf7,
32'h3dfc4418,
32'h3de2f148,
32'h3dc905c5,
32'h3dae81cf,
32'h3d9365a8,
32'h3d77b192,
32'h3d5b65d2,
32'h3d3e82ae,
32'h3d21086c,
32'h3d02f757,
32'h3ce44fb7,
32'h3cc511d9,
32'h3ca53e09,
32'h3c84d496,
32'h3c63d5d1,
32'h3c42420a,
32'h3c201994,
32'h3bfd5cc4,
32'h3bda0bf0,
32'h3bb6276e,
32'h3b91af97,
32'h3b6ca4c4,
32'h3b470753,
32'h3b20d79e,
32'h3afa1605,
32'h3ad2c2e8,
32'h3aaadea6,
32'h3a8269a3,
32'h3a596442,
32'h3a2fcee8,
32'h3a05a9fd,
32'h39daf5e8,
32'h39afb313,
32'h3983e1e8,
32'h395782d3,
32'h392a9642,
32'h38fd1ca4,
32'h38cf1669,
32'h38a08402,
32'h387165e3,
32'h3841bc7f,
32'h3811884d,
32'h37e0c9c3,
32'h37af8159,
32'h377daf89,
32'h374b54ce,
32'h371871a5,
32'h36e5068a,
32'h36b113fd,
32'h367c9a7e,
32'h36479a8e,
32'h361214b0,
32'h35dc0968,
32'h35a5793c,
32'h356e64b2,
32'h3536cc52,
32'h34feb0a5,
32'h34c61236,
32'h348cf190,
32'h34534f41,
32'h34192bd5,
32'h33de87de,
32'h33a363ec,
32'h3367c090,
32'h332b9e5e,
32'h32eefdea,
32'h32b1dfc9,
32'h32744493,
32'h32362ce0,
32'h31f79948,
32'h31b88a66,
32'h317900d6,
32'h3138fd35,
32'h30f8801f,
32'h30b78a36,
32'h30761c18,
32'h30343667,
32'h2ff1d9c7,
32'h2faf06da,
32'h2f6bbe45,
32'h2f2800af,
32'h2ee3cebe,
32'h2e9f291b,
32'h2e5a1070,
32'h2e148566,
32'h2dce88aa,
32'h2d881ae8,
32'h2d413ccd,
32'h2cf9ef09,
32'h2cb2324c,
32'h2c6a0746,
32'h2c216eaa,
32'h2bd8692b,
32'h2b8ef77d,
32'h2b451a55,
32'h2afad269,
32'h2ab02071,
32'h2a650525,
32'h2a19813f,
32'h29cd9578,
32'h2981428c,
32'h29348937,
32'h28e76a37,
32'h2899e64a,
32'h284bfe2f,
32'h27fdb2a7,
32'h27af0472,
32'h275ff452,
32'h2710830c,
32'h26c0b162,
32'h2670801a,
32'h261feffa,
32'h25cf01c8,
32'h257db64c,
32'h252c0e4f,
32'h24da0a9a,
32'h2487abf7,
32'h2434f332,
32'h23e1e117,
32'h238e7673,
32'h233ab414,
32'h22e69ac8,
32'h22922b5e,
32'h223d66a8,
32'h21e84d76,
32'h2192e09b,
32'h213d20e8,
32'h20e70f32,
32'h2090ac4d,
32'h2039f90f,
32'h1fe2f64c,
32'h1f8ba4dc,
32'h1f340596,
32'h1edc1953,
32'h1e83e0eb,
32'h1e2b5d38,
32'h1dd28f15,
32'h1d79775c,
32'h1d2016e9,
32'h1cc66e99,
32'h1c6c7f4a,
32'h1c1249d8,
32'h1bb7cf23,
32'h1b5d100a,
32'h1b020d6c,
32'h1aa6c82b,
32'h1a4b4128,
32'h19ef7944,
32'h19937161,
32'h19372a64,
32'h18daa52f,
32'h187de2a7,
32'h1820e3b0,
32'h17c3a931,
32'h1766340f,
32'h17088531,
32'h16aa9d7e,
32'h164c7ddd,
32'h15ee2738,
32'h158f9a76,
32'h1530d881,
32'h14d1e242,
32'h1472b8a5,
32'h14135c94,
32'h13b3cefa,
32'h135410c3,
32'h12f422db,
32'h1294062f,
32'h1233bbac,
32'h11d3443f,
32'h1172a0d7,
32'h1111d263,
32'h10b0d9d0,
32'h104fb80e,
32'h0fee6e0d,
32'h0f8cfcbe,
32'h0f2b650f,
32'h0ec9a7f3,
32'h0e67c65a,
32'h0e05c135,
32'h0da39978,
32'h0d415013,
32'h0cdee5f9,
32'h0c7c5c1e,
32'h0c19b374,
32'h0bb6ecef,
32'h0b540982,
32'h0af10a22,
32'h0a8defc3,
32'h0a2abb59,
32'h09c76dd8,
32'h09640837,
32'h09008b6a,
32'h089cf867,
32'h08395024,
32'h07d59396,
32'h0771c3b3,
32'h070de172,
32'h06a9edc9,
32'h0645e9af,
32'h05e1d61b,
32'h057db403,
32'h0519845e,
32'h04b54825,
32'h0451004d,
32'h03ecadcf,
32'h038851a2,
32'h0323ecbe,
32'h02bf801a,
32'h025b0caf,
32'h01f69373,
32'h0192155f,
32'h012d936c,
32'h00c90e90,
32'h006487c4,
32'h00000000,
32'hff9b783c,
32'hff36f170,
32'hfed26c94,
32'hfe6deaa1,
32'hfe096c8d,
32'hfda4f351,
32'hfd407fe6,
32'hfcdc1342,
32'hfc77ae5e,
32'hfc135231,
32'hfbaeffb3,
32'hfb4ab7db,
32'hfae67ba2,
32'hfa824bfd,
32'hfa1e29e5,
32'hf9ba1651,
32'hf9561237,
32'hf8f21e8e,
32'hf88e3c4d,
32'hf82a6c6a,
32'hf7c6afdc,
32'hf7630799,
32'hf6ff7496,
32'hf69bf7c9,
32'hf6389228,
32'hf5d544a7,
32'hf572103d,
32'hf50ef5de,
32'hf4abf67e,
32'hf4491311,
32'hf3e64c8c,
32'hf383a3e2,
32'hf3211a07,
32'hf2beafed,
32'hf25c6688,
32'hf1fa3ecb,
32'hf19839a6,
32'hf136580d,
32'hf0d49af1,
32'hf0730342,
32'hf01191f3,
32'hefb047f2,
32'hef4f2630,
32'heeee2d9d,
32'hee8d5f29,
32'hee2cbbc1,
32'hedcc4454,
32'hed6bf9d1,
32'hed0bdd25,
32'hecabef3d,
32'hec4c3106,
32'hebeca36c,
32'heb8d475b,
32'heb2e1dbe,
32'heacf277f,
32'hea70658a,
32'hea11d8c8,
32'he9b38223,
32'he9556282,
32'he8f77acf,
32'he899cbf1,
32'he83c56cf,
32'he7df1c50,
32'he7821d59,
32'he7255ad1,
32'he6c8d59c,
32'he66c8e9f,
32'he61086bc,
32'he5b4bed8,
32'he55937d5,
32'he4fdf294,
32'he4a2eff6,
32'he44830dd,
32'he3edb628,
32'he39380b6,
32'he3399167,
32'he2dfe917,
32'he28688a4,
32'he22d70eb,
32'he1d4a2c8,
32'he17c1f15,
32'he123e6ad,
32'he0cbfa6a,
32'he0745b24,
32'he01d09b4,
32'hdfc606f1,
32'hdf6f53b3,
32'hdf18f0ce,
32'hdec2df18,
32'hde6d1f65,
32'hde17b28a,
32'hddc29958,
32'hdd6dd4a2,
32'hdd196538,
32'hdcc54bec,
32'hdc71898d,
32'hdc1e1ee9,
32'hdbcb0cce,
32'hdb785409,
32'hdb25f566,
32'hdad3f1b1,
32'hda8249b4,
32'hda30fe38,
32'hd9e01006,
32'hd98f7fe6,
32'hd93f4e9e,
32'hd8ef7cf4,
32'hd8a00bae,
32'hd850fb8e,
32'hd8024d59,
32'hd7b401d1,
32'hd76619b6,
32'hd71895c9,
32'hd6cb76c9,
32'hd67ebd74,
32'hd6326a88,
32'hd5e67ec1,
32'hd59afadb,
32'hd54fdf8f,
32'hd5052d97,
32'hd4bae5ab,
32'hd4710883,
32'hd42796d5,
32'hd3de9156,
32'hd395f8ba,
32'hd34dcdb4,
32'hd30610f7,
32'hd2bec333,
32'hd277e518,
32'hd2317756,
32'hd1eb7a9a,
32'hd1a5ef90,
32'hd160d6e5,
32'hd11c3142,
32'hd0d7ff51,
32'hd09441bb,
32'hd050f926,
32'hd00e2639,
32'hcfcbc999,
32'hcf89e3e8,
32'hcf4875ca,
32'hcf077fe1,
32'hcec702cb,
32'hce86ff2a,
32'hce47759a,
32'hce0866b8,
32'hcdc9d320,
32'hcd8bbb6d,
32'hcd4e2037,
32'hcd110216,
32'hccd461a2,
32'hcc983f70,
32'hcc5c9c14,
32'hcc217822,
32'hcbe6d42b,
32'hcbacb0bf,
32'hcb730e70,
32'hcb39edca,
32'hcb014f5b,
32'hcac933ae,
32'hca919b4e,
32'hca5a86c4,
32'hca23f698,
32'hc9edeb50,
32'hc9b86572,
32'hc9836582,
32'hc94eec03,
32'hc91af976,
32'hc8e78e5b,
32'hc8b4ab32,
32'hc8825077,
32'hc8507ea7,
32'hc81f363d,
32'hc7ee77b3,
32'hc7be4381,
32'hc78e9a1d,
32'hc75f7bfe,
32'hc730e997,
32'hc702e35c,
32'hc6d569be,
32'hc6a87d2d,
32'hc67c1e18,
32'hc6504ced,
32'hc6250a18,
32'hc5fa5603,
32'hc5d03118,
32'hc5a69bbe,
32'hc57d965d,
32'hc555215a,
32'hc52d3d18,
32'hc505e9fb,
32'hc4df2862,
32'hc4b8f8ad,
32'hc4935b3c,
32'hc46e5069,
32'hc449d892,
32'hc425f410,
32'hc402a33c,
32'hc3dfe66c,
32'hc3bdbdf6,
32'hc39c2a2f,
32'hc37b2b6a,
32'hc35ac1f7,
32'hc33aee27,
32'hc31bb049,
32'hc2fd08a9,
32'hc2def794,
32'hc2c17d52,
32'hc2a49a2e,
32'hc2884e6e,
32'hc26c9a58,
32'hc2517e31,
32'hc236fa3b,
32'hc21d0eb8,
32'hc203bbe8,
32'hc1eb0209,
32'hc1d2e158,
32'hc1bb5a11,
32'hc1a46c6e,
32'hc18e18a7,
32'hc1785ef4,
32'hc1633f8a,
32'hc14eba9d,
32'hc13ad060,
32'hc1278104,
32'hc114ccb9,
32'hc102b3ac,
32'hc0f1360b,
32'hc0e05401,
32'hc0d00db6,
32'hc0c06355,
32'hc0b15502,
32'hc0a2e2e3,
32'hc0950d1d,
32'hc087d3d0,
32'hc07b371e,
32'hc06f3726,
32'hc063d405,
32'hc0590dd8,
32'hc04ee4b8,
32'hc04558c0,
32'hc03c6a07,
32'hc03418a2,
32'hc02c64a6,
32'hc0254e27,
32'hc01ed535,
32'hc018f9e1,
32'hc013bc39,
32'hc00f1c4a,
32'hc00b1a20,
32'hc007b5c4,
32'hc004ef3f,
32'hc002c697,
32'hc0013bd3,
32'hc0004ef5,
32'hc0000000,
32'hc0004ef5,
32'hc0013bd3,
32'hc002c697,
32'hc004ef3f,
32'hc007b5c4,
32'hc00b1a20,
32'hc00f1c4a,
32'hc013bc39,
32'hc018f9e1,
32'hc01ed535,
32'hc0254e27,
32'hc02c64a6,
32'hc03418a2,
32'hc03c6a07,
32'hc04558c0,
32'hc04ee4b8,
32'hc0590dd8,
32'hc063d405,
32'hc06f3726,
32'hc07b371e,
32'hc087d3d0,
32'hc0950d1d,
32'hc0a2e2e3,
32'hc0b15502,
32'hc0c06355,
32'hc0d00db6,
32'hc0e05401,
32'hc0f1360b,
32'hc102b3ac,
32'hc114ccb9,
32'hc1278104,
32'hc13ad060,
32'hc14eba9d,
32'hc1633f8a,
32'hc1785ef4,
32'hc18e18a7,
32'hc1a46c6e,
32'hc1bb5a11,
32'hc1d2e158,
32'hc1eb0209,
32'hc203bbe8,
32'hc21d0eb8,
32'hc236fa3b,
32'hc2517e31,
32'hc26c9a58,
32'hc2884e6e,
32'hc2a49a2e,
32'hc2c17d52,
32'hc2def794,
32'hc2fd08a9,
32'hc31bb049,
32'hc33aee27,
32'hc35ac1f7,
32'hc37b2b6a,
32'hc39c2a2f,
32'hc3bdbdf6,
32'hc3dfe66c,
32'hc402a33c,
32'hc425f410,
32'hc449d892,
32'hc46e5069,
32'hc4935b3c,
32'hc4b8f8ad,
32'hc4df2862,
32'hc505e9fb,
32'hc52d3d18,
32'hc555215a,
32'hc57d965d,
32'hc5a69bbe,
32'hc5d03118,
32'hc5fa5603,
32'hc6250a18,
32'hc6504ced,
32'hc67c1e18,
32'hc6a87d2d,
32'hc6d569be,
32'hc702e35c,
32'hc730e997,
32'hc75f7bfe,
32'hc78e9a1d,
32'hc7be4381,
32'hc7ee77b3,
32'hc81f363d,
32'hc8507ea7,
32'hc8825077,
32'hc8b4ab32,
32'hc8e78e5b,
32'hc91af976,
32'hc94eec03,
32'hc9836582,
32'hc9b86572,
32'hc9edeb50,
32'hca23f698,
32'hca5a86c4,
32'hca919b4e,
32'hcac933ae,
32'hcb014f5b,
32'hcb39edca,
32'hcb730e70,
32'hcbacb0bf,
32'hcbe6d42b,
32'hcc217822,
32'hcc5c9c14,
32'hcc983f70,
32'hccd461a2,
32'hcd110216,
32'hcd4e2037,
32'hcd8bbb6d,
32'hcdc9d320,
32'hce0866b8,
32'hce47759a,
32'hce86ff2a,
32'hcec702cb,
32'hcf077fe1,
32'hcf4875ca,
32'hcf89e3e8,
32'hcfcbc999,
32'hd00e2639,
32'hd050f926,
32'hd09441bb,
32'hd0d7ff51,
32'hd11c3142,
32'hd160d6e5,
32'hd1a5ef90,
32'hd1eb7a9a,
32'hd2317756,
32'hd277e518,
32'hd2bec333,
32'hd30610f7,
32'hd34dcdb4,
32'hd395f8ba,
32'hd3de9156,
32'hd42796d5,
32'hd4710883,
32'hd4bae5ab,
32'hd5052d97,
32'hd54fdf8f,
32'hd59afadb,
32'hd5e67ec1,
32'hd6326a88,
32'hd67ebd74,
32'hd6cb76c9,
32'hd71895c9,
32'hd76619b6,
32'hd7b401d1,
32'hd8024d59,
32'hd850fb8e,
32'hd8a00bae,
32'hd8ef7cf4,
32'hd93f4e9e,
32'hd98f7fe6,
32'hd9e01006,
32'hda30fe38,
32'hda8249b4,
32'hdad3f1b1,
32'hdb25f566,
32'hdb785409,
32'hdbcb0cce,
32'hdc1e1ee9,
32'hdc71898d,
32'hdcc54bec,
32'hdd196538,
32'hdd6dd4a2,
32'hddc29958,
32'hde17b28a,
32'hde6d1f65,
32'hdec2df18,
32'hdf18f0ce,
32'hdf6f53b3,
32'hdfc606f1,
32'he01d09b4,
32'he0745b24,
32'he0cbfa6a,
32'he123e6ad,
32'he17c1f15,
32'he1d4a2c8,
32'he22d70eb,
32'he28688a4,
32'he2dfe917,
32'he3399167,
32'he39380b6,
32'he3edb628,
32'he44830dd,
32'he4a2eff6,
32'he4fdf294,
32'he55937d5,
32'he5b4bed8,
32'he61086bc,
32'he66c8e9f,
32'he6c8d59c,
32'he7255ad1,
32'he7821d59,
32'he7df1c50,
32'he83c56cf,
32'he899cbf1,
32'he8f77acf,
32'he9556282,
32'he9b38223,
32'hea11d8c8,
32'hea70658a,
32'heacf277f,
32'heb2e1dbe,
32'heb8d475b,
32'hebeca36c,
32'hec4c3106,
32'hecabef3d,
32'hed0bdd25,
32'hed6bf9d1,
32'hedcc4454,
32'hee2cbbc1,
32'hee8d5f29,
32'heeee2d9d,
32'hef4f2630,
32'hefb047f2,
32'hf01191f3,
32'hf0730342,
32'hf0d49af1,
32'hf136580d,
32'hf19839a6,
32'hf1fa3ecb,
32'hf25c6688,
32'hf2beafed,
32'hf3211a07,
32'hf383a3e2,
32'hf3e64c8c,
32'hf4491311,
32'hf4abf67e,
32'hf50ef5de,
32'hf572103d,
32'hf5d544a7,
32'hf6389228,
32'hf69bf7c9,
32'hf6ff7496,
32'hf7630799,
32'hf7c6afdc,
32'hf82a6c6a,
32'hf88e3c4d,
32'hf8f21e8e,
32'hf9561237,
32'hf9ba1651,
32'hfa1e29e5,
32'hfa824bfd,
32'hfae67ba2,
32'hfb4ab7db,
32'hfbaeffb3,
32'hfc135231,
32'hfc77ae5e,
32'hfcdc1342,
32'hfd407fe6,
32'hfda4f351,
32'hfe096c8d,
32'hfe6deaa1,
32'hfed26c94,
32'hff36f170,
32'hff9b783c
};
