logic [0:ROM_DEPTH-1] [DATA_WIDTH-1:0] table_ = {
32'hc0000000,
32'hc00004ef,
32'hc00013bd,
32'hc0002c6a,
32'hc0004ef5,
32'hc0007b5f,
32'hc000b1a7,
32'hc000f1ce,
32'hc0013bd3,
32'hc0018fb6,
32'hc001ed78,
32'hc0025519,
32'hc002c697,
32'hc00341f4,
32'hc003c72f,
32'hc0045648,
32'hc004ef3f,
32'hc0059214,
32'hc0063ec6,
32'hc006f556,
32'hc007b5c4,
32'hc008800f,
32'hc0095438,
32'hc00a323d,
32'hc00b1a20,
32'hc00c0be0,
32'hc00d077c,
32'hc00e0cf5,
32'hc00f1c4a,
32'hc010357c,
32'hc011588a,
32'hc0128574,
32'hc013bc39,
32'hc014fcda,
32'hc0164757,
32'hc0179bae,
32'hc018f9e1,
32'hc01a61ee,
32'hc01bd3d6,
32'hc01d4f99,
32'hc01ed535,
32'hc02064ab,
32'hc021fdfb,
32'hc023a124,
32'hc0254e27,
32'hc0270502,
32'hc028c5b6,
32'hc02a9042,
32'hc02c64a6,
32'hc02e42e2,
32'hc0302af5,
32'hc0321ce0,
32'hc03418a2,
32'hc0361e3a,
32'hc0382da8,
32'hc03a46ed,
32'hc03c6a07,
32'hc03e96f6,
32'hc040cdba,
32'hc0430e53,
32'hc04558c0,
32'hc047ad01,
32'hc04a0b16,
32'hc04c72fe,
32'hc04ee4b8,
32'hc0516045,
32'hc053e5a5,
32'hc05674d6,
32'hc0590dd8,
32'hc05bb0ab,
32'hc05e5d4e,
32'hc06113c2,
32'hc063d405,
32'hc0669e18,
32'hc06971f9,
32'hc06c4fa8,
32'hc06f3726,
32'hc0722871,
32'hc0752389,
32'hc078286e,
32'hc07b371e,
32'hc07e4f9b,
32'hc08171e2,
32'hc0849df4,
32'hc087d3d0,
32'hc08b1376,
32'hc08e5ce5,
32'hc091b01d,
32'hc0950d1d,
32'hc09873e4,
32'hc09be473,
32'hc09f5ec8,
32'hc0a2e2e3,
32'hc0a670c4,
32'hc0aa086a,
32'hc0ada9d4,
32'hc0b15502,
32'hc0b509f3,
32'hc0b8c8a7,
32'hc0bc911d,
32'hc0c06355,
32'hc0c43f4d,
32'hc0c82506,
32'hc0cc147f,
32'hc0d00db6,
32'hc0d410ad,
32'hc0d81d61,
32'hc0dc33d2,
32'hc0e05401,
32'hc0e47deb,
32'hc0e8b190,
32'hc0eceef1,
32'hc0f1360b,
32'hc0f586df,
32'hc0f9e16b,
32'hc0fe45b0,
32'hc102b3ac,
32'hc1072b5f,
32'hc10bacc8,
32'hc11037e6,
32'hc114ccb9,
32'hc1196b3f,
32'hc11e1379,
32'hc122c566,
32'hc1278104,
32'hc12c4653,
32'hc1311553,
32'hc135ee02,
32'hc13ad060,
32'hc13fbc6c,
32'hc144b225,
32'hc149b18b,
32'hc14eba9d,
32'hc153cd5a,
32'hc158e9c1,
32'hc15e0fd1,
32'hc1633f8a,
32'hc16878eb,
32'hc16dbbf3,
32'hc17308a1,
32'hc1785ef4,
32'hc17dbeec,
32'hc1832888,
32'hc1889bc6,
32'hc18e18a7,
32'hc1939f29,
32'hc1992f4c,
32'hc19ec90d,
32'hc1a46c6e,
32'hc1aa196c,
32'hc1afd007,
32'hc1b5903f,
32'hc1bb5a11,
32'hc1c12d7e,
32'hc1c70a84,
32'hc1ccf122,
32'hc1d2e158,
32'hc1d8db25,
32'hc1dede87,
32'hc1e4eb7e,
32'hc1eb0209,
32'hc1f12227,
32'hc1f74bd6,
32'hc1fd7f17,
32'hc203bbe8,
32'hc20a0248,
32'hc2105236,
32'hc216abb1,
32'hc21d0eb8,
32'hc2237b4b,
32'hc229f167,
32'hc230710d,
32'hc236fa3b,
32'hc23d8cf1,
32'hc244292c,
32'hc24aceed,
32'hc2517e31,
32'hc25836f9,
32'hc25ef943,
32'hc265c50e,
32'hc26c9a58,
32'hc2737922,
32'hc27a616a,
32'hc281532e,
32'hc2884e6e,
32'hc28f5329,
32'hc296615d,
32'hc29d790a,
32'hc2a49a2e,
32'hc2abc4c9,
32'hc2b2f8d8,
32'hc2ba365c,
32'hc2c17d52,
32'hc2c8cdbb,
32'hc2d02794,
32'hc2d78add,
32'hc2def794,
32'hc2e66db8,
32'hc2eded49,
32'hc2f57644,
32'hc2fd08a9,
32'hc304a477,
32'hc30c49ad,
32'hc313f848,
32'hc31bb049,
32'hc32371ae,
32'hc32b3c75,
32'hc333109e,
32'hc33aee27,
32'hc342d510,
32'hc34ac556,
32'hc352bef9,
32'hc35ac1f7,
32'hc362ce50,
32'hc36ae401,
32'hc373030a,
32'hc37b2b6a,
32'hc3835d1e,
32'hc38b9827,
32'hc393dc82,
32'hc39c2a2f,
32'hc3a4812c,
32'hc3ace178,
32'hc3b54b11,
32'hc3bdbdf6,
32'hc3c63a26,
32'hc3cebfa0,
32'hc3d74e62,
32'hc3dfe66c,
32'hc3e887bb,
32'hc3f1324e,
32'hc3f9e624,
32'hc402a33c,
32'hc40b6994,
32'hc414392b,
32'hc41d11ff,
32'hc425f410,
32'hc42edf5c,
32'hc437d3e1,
32'hc440d19e,
32'hc449d892,
32'hc452e8bc,
32'hc45c0219,
32'hc46524a9,
32'hc46e5069,
32'hc477855a,
32'hc480c379,
32'hc48a0ac4,
32'hc4935b3c,
32'hc49cb4dd,
32'hc4a617a6,
32'hc4af8397,
32'hc4b8f8ad,
32'hc4c276e8,
32'hc4cbfe45,
32'hc4d58ec3,
32'hc4df2862,
32'hc4e8cb1e,
32'hc4f276f7,
32'hc4fc2bec,
32'hc505e9fb,
32'hc50fb121,
32'hc519815f,
32'hc5235ab2,
32'hc52d3d18,
32'hc5372891,
32'hc5411d1b,
32'hc54b1ab4,
32'hc555215a,
32'hc55f310d,
32'hc56949ca,
32'hc5736b90,
32'hc57d965d,
32'hc587ca31,
32'hc5920708,
32'hc59c4ce3,
32'hc5a69bbe,
32'hc5b0f399,
32'hc5bb5472,
32'hc5c5be47,
32'hc5d03118,
32'hc5daace1,
32'hc5e531a1,
32'hc5efbf58,
32'hc5fa5603,
32'hc604f5a0,
32'hc60f9e2e,
32'hc61a4fac,
32'hc6250a18,
32'hc62fcd6f,
32'hc63a99b1,
32'hc6456edb,
32'hc6504ced,
32'hc65b33e4,
32'hc66623be,
32'hc6711c7b,
32'hc67c1e18,
32'hc6872894,
32'hc6923bec,
32'hc69d5820,
32'hc6a87d2d,
32'hc6b3ab12,
32'hc6bee1cd,
32'hc6ca215c,
32'hc6d569be,
32'hc6e0baf0,
32'hc6ec14f2,
32'hc6f777c1,
32'hc702e35c,
32'hc70e57c0,
32'hc719d4ed,
32'hc7255ae0,
32'hc730e997,
32'hc73c8111,
32'hc748214c,
32'hc753ca46,
32'hc75f7bfe,
32'hc76b3671,
32'hc776f99d,
32'hc782c582,
32'hc78e9a1d,
32'hc79a776c,
32'hc7a65d6e,
32'hc7b24c20,
32'hc7be4381,
32'hc7ca438f,
32'hc7d64c47,
32'hc7e25daa,
32'hc7ee77b3,
32'hc7fa9a62,
32'hc806c5b5,
32'hc812f9a9,
32'hc81f363d,
32'hc82b7b70,
32'hc837c93e,
32'hc8441fa6,
32'hc8507ea7,
32'hc85ce63e,
32'hc869566a,
32'hc875cf28,
32'hc8825077,
32'hc88eda54,
32'hc89b6cbf,
32'hc8a807b4,
32'hc8b4ab32,
32'hc8c15736,
32'hc8ce0bc0,
32'hc8dac8cd,
32'hc8e78e5b,
32'hc8f45c68,
32'hc90132f2,
32'hc90e11f7,
32'hc91af976,
32'hc927e96b,
32'hc934e1d6,
32'hc941e2b4,
32'hc94eec03,
32'hc95bfdc1,
32'hc96917ec,
32'hc9763a83,
32'hc9836582,
32'hc99098e9,
32'hc99dd4b4,
32'hc9ab18e3,
32'hc9b86572,
32'hc9c5ba60,
32'hc9d317ab,
32'hc9e07d51,
32'hc9edeb50,
32'hc9fb61a5,
32'hca08e04f,
32'hca16674b,
32'hca23f698,
32'hca318e32,
32'hca3f2e19,
32'hca4cd64b,
32'hca5a86c4,
32'hca683f83,
32'hca760086,
32'hca83c9ca,
32'hca919b4e,
32'hca9f750f,
32'hcaad570c,
32'hcabb4141,
32'hcac933ae,
32'hcad72e4f,
32'hcae53123,
32'hcaf33c28,
32'hcb014f5b,
32'hcb0f6aba,
32'hcb1d8e43,
32'hcb2bb9f4,
32'hcb39edca,
32'hcb4829c4,
32'hcb566ddf,
32'hcb64ba19,
32'hcb730e70,
32'hcb816ae1,
32'hcb8fcf6b,
32'hcb9e3c0b,
32'hcbacb0bf,
32'hcbbb2d85,
32'hcbc9b25a,
32'hcbd83f3d,
32'hcbe6d42b,
32'hcbf57121,
32'hcc04161e,
32'hcc12c31f,
32'hcc217822,
32'hcc303524,
32'hcc3efa25,
32'hcc4dc720,
32'hcc5c9c14,
32'hcc6b78ff,
32'hcc7a5dde,
32'hcc894aaf,
32'hcc983f70,
32'hcca73c1e,
32'hccb640b8,
32'hccc54d3a,
32'hccd461a2,
32'hcce37def,
32'hccf2a21d,
32'hcd01ce2b,
32'hcd110216,
32'hcd203ddc,
32'hcd2f817b,
32'hcd3eccef,
32'hcd4e2037,
32'hcd5d7b50,
32'hcd6cde39,
32'hcd7c48ee,
32'hcd8bbb6d,
32'hcd9b35b4,
32'hcdaab7c0,
32'hcdba4190,
32'hcdc9d320,
32'hcdd96c6f,
32'hcde90d79,
32'hcdf8b63d,
32'hce0866b8,
32'hce181ee8,
32'hce27dec9,
32'hce37a65b,
32'hce47759a,
32'hce574c84,
32'hce672b16,
32'hce77114e,
32'hce86ff2a,
32'hce96f4a7,
32'hcea6f1c2,
32'hceb6f67a,
32'hcec702cb,
32'hced716b4,
32'hcee73231,
32'hcef75541,
32'hcf077fe1,
32'hcf17b20d,
32'hcf27ebc5,
32'hcf382d05,
32'hcf4875ca,
32'hcf58c613,
32'hcf691ddd,
32'hcf797d24,
32'hcf89e3e8,
32'hcf9a5225,
32'hcfaac7d8,
32'hcfbb4500,
32'hcfcbc999,
32'hcfdc55a1,
32'hcfece915,
32'hcffd83f4,
32'hd00e2639,
32'hd01ecfe4,
32'hd02f80f1,
32'hd040395d,
32'hd050f926,
32'hd061c04a,
32'hd0728ec6,
32'hd0836497,
32'hd09441bb,
32'hd0a5262f,
32'hd0b611f1,
32'hd0c704fd,
32'hd0d7ff51,
32'hd0e900ec,
32'hd0fa09c9,
32'hd10b19e7,
32'hd11c3142,
32'hd12d4fd9,
32'hd13e75a8,
32'hd14fa2ad,
32'hd160d6e5,
32'hd172124d,
32'hd18354e4,
32'hd1949ea6,
32'hd1a5ef90,
32'hd1b747a0,
32'hd1c8a6d4,
32'hd1da0d28,
32'hd1eb7a9a,
32'hd1fcef27,
32'hd20e6acc,
32'hd21fed88,
32'hd2317756,
32'hd2430835,
32'hd254a021,
32'hd2663f19,
32'hd277e518,
32'hd289921e,
32'hd29b4626,
32'hd2ad012e
};
