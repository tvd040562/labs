logic [0:ROM_DEPTH-1] [DATA_WIDTH-1:0] table_ = {
32'h00000000,
32'h0192155f,
32'h0323ecbe,
32'h04b54825,
32'h0645e9af,
32'h07d59396,
32'h09640837,
32'h0af10a22,
32'h0c7c5c1e,
32'h0e05c135,
32'h0f8cfcbe,
32'h1111d263,
32'h1294062f,
32'h14135c94,
32'h158f9a76,
32'h17088531,
32'h187de2a7,
32'h19ef7944,
32'h1b5d100a,
32'h1cc66e99,
32'h1e2b5d38,
32'h1f8ba4dc,
32'h20e70f32,
32'h223d66a8,
32'h238e7673,
32'h24da0a9a,
32'h261feffa,
32'h275ff452,
32'h2899e64a,
32'h29cd9578,
32'h2afad269,
32'h2c216eaa,
32'h2d413ccd,
32'h2e5a1070,
32'h2f6bbe45,
32'h30761c18,
32'h317900d6,
32'h32744493,
32'h3367c090,
32'h34534f41,
32'h3536cc52,
32'h361214b0,
32'h36e5068a,
32'h37af8159,
32'h387165e3,
32'h392a9642,
32'h39daf5e8,
32'h3a8269a3,
32'h3b20d79e,
32'h3bb6276e,
32'h3c42420a,
32'h3cc511d9,
32'h3d3e82ae,
32'h3dae81cf,
32'h3e14fdf7,
32'h3e71e759,
32'h3ec52fa0,
32'h3f0ec9f5,
32'h3f4eaafe,
32'h3f84c8e2,
32'h3fb11b48,
32'h3fd39b5a,
32'h3fec43c7,
32'h3ffb10c1,
32'h40000000,
32'h3ffb10c1,
32'h3fec43c7,
32'h3fd39b5a,
32'h3fb11b48,
32'h3f84c8e2,
32'h3f4eaafe,
32'h3f0ec9f5,
32'h3ec52fa0,
32'h3e71e759,
32'h3e14fdf7,
32'h3dae81cf,
32'h3d3e82ae,
32'h3cc511d9,
32'h3c42420a,
32'h3bb6276e,
32'h3b20d79e,
32'h3a8269a3,
32'h39daf5e8,
32'h392a9642,
32'h387165e3,
32'h37af8159,
32'h36e5068a,
32'h361214b0,
32'h3536cc52,
32'h34534f41,
32'h3367c090,
32'h32744493,
32'h317900d6,
32'h30761c18,
32'h2f6bbe45,
32'h2e5a1070,
32'h2d413ccd,
32'h2c216eaa,
32'h2afad269,
32'h29cd9578,
32'h2899e64a,
32'h275ff452,
32'h261feffa,
32'h24da0a9a,
32'h238e7673,
32'h223d66a8,
32'h20e70f32,
32'h1f8ba4dc,
32'h1e2b5d38,
32'h1cc66e99,
32'h1b5d100a,
32'h19ef7944,
32'h187de2a7,
32'h17088531,
32'h158f9a76,
32'h14135c94,
32'h1294062f,
32'h1111d263,
32'h0f8cfcbe,
32'h0e05c135,
32'h0c7c5c1e,
32'h0af10a22,
32'h09640837,
32'h07d59396,
32'h0645e9af,
32'h04b54825,
32'h0323ecbe,
32'h0192155f,
32'h00000000,
32'hfe6deaa1,
32'hfcdc1342,
32'hfb4ab7db,
32'hf9ba1651,
32'hf82a6c6a,
32'hf69bf7c9,
32'hf50ef5de,
32'hf383a3e2,
32'hf1fa3ecb,
32'hf0730342,
32'heeee2d9d,
32'hed6bf9d1,
32'hebeca36c,
32'hea70658a,
32'he8f77acf,
32'he7821d59,
32'he61086bc,
32'he4a2eff6,
32'he3399167,
32'he1d4a2c8,
32'he0745b24,
32'hdf18f0ce,
32'hddc29958,
32'hdc71898d,
32'hdb25f566,
32'hd9e01006,
32'hd8a00bae,
32'hd76619b6,
32'hd6326a88,
32'hd5052d97,
32'hd3de9156,
32'hd2bec333,
32'hd1a5ef90,
32'hd09441bb,
32'hcf89e3e8,
32'hce86ff2a,
32'hcd8bbb6d,
32'hcc983f70,
32'hcbacb0bf,
32'hcac933ae,
32'hc9edeb50,
32'hc91af976,
32'hc8507ea7,
32'hc78e9a1d,
32'hc6d569be,
32'hc6250a18,
32'hc57d965d,
32'hc4df2862,
32'hc449d892,
32'hc3bdbdf6,
32'hc33aee27,
32'hc2c17d52,
32'hc2517e31,
32'hc1eb0209,
32'hc18e18a7,
32'hc13ad060,
32'hc0f1360b,
32'hc0b15502,
32'hc07b371e,
32'hc04ee4b8,
32'hc02c64a6,
32'hc013bc39,
32'hc004ef3f,
32'hc0000000,
32'hc004ef3f,
32'hc013bc39,
32'hc02c64a6,
32'hc04ee4b8,
32'hc07b371e,
32'hc0b15502,
32'hc0f1360b,
32'hc13ad060,
32'hc18e18a7,
32'hc1eb0209,
32'hc2517e31,
32'hc2c17d52,
32'hc33aee27,
32'hc3bdbdf6,
32'hc449d892,
32'hc4df2862,
32'hc57d965d,
32'hc6250a18,
32'hc6d569be,
32'hc78e9a1d,
32'hc8507ea7,
32'hc91af976,
32'hc9edeb50,
32'hcac933ae,
32'hcbacb0bf,
32'hcc983f70,
32'hcd8bbb6d,
32'hce86ff2a,
32'hcf89e3e8,
32'hd09441bb,
32'hd1a5ef90,
32'hd2bec333,
32'hd3de9156,
32'hd5052d97,
32'hd6326a88,
32'hd76619b6,
32'hd8a00bae,
32'hd9e01006,
32'hdb25f566,
32'hdc71898d,
32'hddc29958,
32'hdf18f0ce,
32'he0745b24,
32'he1d4a2c8,
32'he3399167,
32'he4a2eff6,
32'he61086bc,
32'he7821d59,
32'he8f77acf,
32'hea70658a,
32'hebeca36c,
32'hed6bf9d1,
32'heeee2d9d,
32'hf0730342,
32'hf1fa3ecb,
32'hf383a3e2,
32'hf50ef5de,
32'hf69bf7c9,
32'hf82a6c6a,
32'hf9ba1651,
32'hfb4ab7db,
32'hfcdc1342,
32'hfe6deaa1
};
