VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MACRO sky130_sram_512byte_1rw1r_32x128_8
   CLASS BLOCK ;
   SIZE 480.72 BY 273.27 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  107.46 0.0 107.84 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  113.3 0.0 113.68 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  119.14 0.0 119.52 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  124.98 0.0 125.36 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  130.82 0.0 131.2 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  136.66 0.0 137.04 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  142.5 0.0 142.88 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  148.34 0.0 148.72 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  154.18 0.0 154.56 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  160.02 0.0 160.4 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  165.86 0.0 166.24 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  171.7 0.0 172.08 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  177.54 0.0 177.92 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  183.38 0.0 183.76 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  189.22 0.0 189.6 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  195.06 0.0 195.44 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  200.9 0.0 201.28 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  206.74 0.0 207.12 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  212.58 0.0 212.96 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  218.42 0.0 218.8 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  224.26 0.0 224.64 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  230.1 0.0 230.48 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  235.94 0.0 236.32 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  241.78 0.0 242.16 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  247.62 0.0 248.0 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  253.46 0.0 253.84 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  259.3 0.0 259.68 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  265.14 0.0 265.52 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  270.98 0.0 271.36 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  276.82 0.0 277.2 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  282.66 0.0 283.04 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  288.5 0.0 288.88 0.38 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  78.26 0.0 78.64 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 121.87 0.38 122.25 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 130.37 0.38 130.75 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 136.275 0.38 136.655 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 144.675 0.38 145.055 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 150.15 0.38 150.53 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 158.65 0.38 159.03 ;
      END
   END addr0[6]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  397.62 272.89 398.0 273.27 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  480.34 84.385 480.72 84.765 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  480.34 75.985 480.72 76.365 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  480.34 70.49 480.72 70.87 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  413.705 0.0 414.085 0.38 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  414.395 0.0 414.775 0.38 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  415.14 0.0 415.52 0.38 ;
      END
   END addr1[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 28.89 0.38 29.27 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  480.34 258.02 480.72 258.4 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 37.39 0.38 37.77 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  31.1 0.0 31.48 0.38 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  450.08 272.89 450.46 273.27 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  84.1 0.0 84.48 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  89.94 0.0 90.32 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  95.78 0.0 96.16 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  101.62 0.0 102.0 0.38 ;
      END
   END wmask0[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  140.12 0.0 140.5 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  146.535 0.0 146.915 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.245 0.0 155.625 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  160.71 0.0 161.09 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.55 0.0 166.93 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.585 0.0 172.965 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.825 0.0 179.205 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  185.065 0.0 185.445 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.685 0.0 193.065 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.545 0.0 197.925 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.785 0.0 204.165 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  210.025 0.0 210.405 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.265 0.0 216.645 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  222.455 0.0 222.835 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  228.06 0.0 228.44 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  234.135 0.0 234.515 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  242.605 0.0 242.985 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  248.845 0.0 249.225 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  254.15 0.0 254.53 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  260.005 0.0 260.385 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  266.185 0.0 266.565 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  272.425 0.0 272.805 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.665 0.0 279.045 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.905 0.0 285.285 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  292.525 0.0 292.905 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  297.385 0.0 297.765 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  303.625 0.0 304.005 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  309.865 0.0 310.245 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  316.105 0.0 316.485 0.38 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  322.345 0.0 322.725 0.38 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  328.585 0.0 328.965 0.38 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  334.825 0.0 335.205 0.38 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  141.445 272.89 141.825 273.27 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  147.685 272.89 148.065 273.27 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  153.925 272.89 154.305 273.27 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  160.165 272.89 160.545 273.27 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.405 272.89 166.785 273.27 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.645 272.89 173.025 273.27 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.885 272.89 179.265 273.27 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  185.125 272.89 185.505 273.27 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.365 272.89 191.745 273.27 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.605 272.89 197.985 273.27 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.845 272.89 204.225 273.27 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  210.085 272.89 210.465 273.27 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.325 272.89 216.705 273.27 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  222.565 272.89 222.945 273.27 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  228.805 272.89 229.185 273.27 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  235.045 272.89 235.425 273.27 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  241.285 272.89 241.665 273.27 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  247.525 272.89 247.905 273.27 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  253.765 272.89 254.145 273.27 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  260.005 272.89 260.385 273.27 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  266.245 272.89 266.625 273.27 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  272.485 272.89 272.865 273.27 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.725 272.89 279.105 273.27 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.965 272.89 285.345 273.27 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  291.205 272.89 291.585 273.27 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  297.445 272.89 297.825 273.27 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  303.685 272.89 304.065 273.27 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  309.925 272.89 310.305 273.27 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  316.165 272.89 316.545 273.27 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  322.405 272.89 322.785 273.27 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  328.645 272.89 329.025 273.27 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  334.885 272.89 335.265 273.27 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  0.0 0.0 480.72 1.74 ;
         LAYER met3 ;
         RECT  0.0 271.53 480.72 273.27 ;
         LAYER met4 ;
         RECT  478.98 0.0 480.72 273.27 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 273.27 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  475.5 3.48 477.24 269.79 ;
         LAYER met4 ;
         RECT  3.48 3.48 5.22 269.79 ;
         LAYER met3 ;
         RECT  3.48 268.05 477.24 269.79 ;
         LAYER met3 ;
         RECT  3.48 3.48 477.24 5.22 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 480.1 272.65 ;
   LAYER  met2 ;
      RECT  0.62 0.62 480.1 272.65 ;
   LAYER  met3 ;
      RECT  0.98 121.27 480.1 122.85 ;
      RECT  0.62 122.85 0.98 129.77 ;
      RECT  0.62 131.35 0.98 135.675 ;
      RECT  0.62 137.255 0.98 144.075 ;
      RECT  0.62 145.655 0.98 149.55 ;
      RECT  0.62 151.13 0.98 158.05 ;
      RECT  0.98 83.785 479.74 85.365 ;
      RECT  0.98 85.365 479.74 121.27 ;
      RECT  479.74 85.365 480.1 121.27 ;
      RECT  479.74 76.965 480.1 83.785 ;
      RECT  479.74 71.47 480.1 75.385 ;
      RECT  0.98 122.85 479.74 257.42 ;
      RECT  0.98 257.42 479.74 259.0 ;
      RECT  479.74 122.85 480.1 257.42 ;
      RECT  0.62 29.87 0.98 36.79 ;
      RECT  0.62 38.37 0.98 121.27 ;
      RECT  479.74 2.34 480.1 69.89 ;
      RECT  0.62 2.34 0.98 28.29 ;
      RECT  0.62 159.63 0.98 270.93 ;
      RECT  479.74 259.0 480.1 270.93 ;
      RECT  0.98 259.0 2.88 267.45 ;
      RECT  0.98 267.45 2.88 270.39 ;
      RECT  0.98 270.39 2.88 270.93 ;
      RECT  2.88 259.0 477.84 267.45 ;
      RECT  2.88 270.39 477.84 270.93 ;
      RECT  477.84 259.0 479.74 267.45 ;
      RECT  477.84 267.45 479.74 270.39 ;
      RECT  477.84 270.39 479.74 270.93 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 83.785 ;
      RECT  2.88 2.34 477.84 2.88 ;
      RECT  2.88 5.82 477.84 83.785 ;
      RECT  477.84 2.34 479.74 2.88 ;
      RECT  477.84 2.88 479.74 5.82 ;
      RECT  477.84 5.82 479.74 83.785 ;
   LAYER  met4 ;
      RECT  106.86 0.98 108.44 272.65 ;
      RECT  108.44 0.62 112.7 0.98 ;
      RECT  114.28 0.62 118.54 0.98 ;
      RECT  120.12 0.62 124.38 0.98 ;
      RECT  125.96 0.62 130.22 0.98 ;
      RECT  131.8 0.62 136.06 0.98 ;
      RECT  149.32 0.62 153.58 0.98 ;
      RECT  236.92 0.62 241.18 0.98 ;
      RECT  108.44 0.98 397.02 272.29 ;
      RECT  397.02 0.98 398.6 272.29 ;
      RECT  32.08 0.62 77.66 0.98 ;
      RECT  398.6 272.29 449.48 272.65 ;
      RECT  79.24 0.62 83.5 0.98 ;
      RECT  85.08 0.62 89.34 0.98 ;
      RECT  90.92 0.62 95.18 0.98 ;
      RECT  96.76 0.62 101.02 0.98 ;
      RECT  102.6 0.62 106.86 0.98 ;
      RECT  137.64 0.62 139.52 0.98 ;
      RECT  141.1 0.62 141.9 0.98 ;
      RECT  143.48 0.62 145.935 0.98 ;
      RECT  147.515 0.62 147.74 0.98 ;
      RECT  156.225 0.62 159.42 0.98 ;
      RECT  161.69 0.62 165.26 0.98 ;
      RECT  167.53 0.62 171.1 0.98 ;
      RECT  173.565 0.62 176.94 0.98 ;
      RECT  179.805 0.62 182.78 0.98 ;
      RECT  184.36 0.62 184.465 0.98 ;
      RECT  186.045 0.62 188.62 0.98 ;
      RECT  190.2 0.62 192.085 0.98 ;
      RECT  193.665 0.62 194.46 0.98 ;
      RECT  196.04 0.62 196.945 0.98 ;
      RECT  198.525 0.62 200.3 0.98 ;
      RECT  201.88 0.62 203.185 0.98 ;
      RECT  204.765 0.62 206.14 0.98 ;
      RECT  207.72 0.62 209.425 0.98 ;
      RECT  211.005 0.62 211.98 0.98 ;
      RECT  213.56 0.62 215.665 0.98 ;
      RECT  217.245 0.62 217.82 0.98 ;
      RECT  219.4 0.62 221.855 0.98 ;
      RECT  223.435 0.62 223.66 0.98 ;
      RECT  225.24 0.62 227.46 0.98 ;
      RECT  229.04 0.62 229.5 0.98 ;
      RECT  231.08 0.62 233.535 0.98 ;
      RECT  235.115 0.62 235.34 0.98 ;
      RECT  243.585 0.62 247.02 0.98 ;
      RECT  249.825 0.62 252.86 0.98 ;
      RECT  255.13 0.62 258.7 0.98 ;
      RECT  260.985 0.62 264.54 0.98 ;
      RECT  267.165 0.62 270.38 0.98 ;
      RECT  273.405 0.62 276.22 0.98 ;
      RECT  277.8 0.62 278.065 0.98 ;
      RECT  279.645 0.62 282.06 0.98 ;
      RECT  283.64 0.62 284.305 0.98 ;
      RECT  285.885 0.62 287.9 0.98 ;
      RECT  289.48 0.62 291.925 0.98 ;
      RECT  293.505 0.62 296.785 0.98 ;
      RECT  298.365 0.62 303.025 0.98 ;
      RECT  304.605 0.62 309.265 0.98 ;
      RECT  310.845 0.62 315.505 0.98 ;
      RECT  317.085 0.62 321.745 0.98 ;
      RECT  323.325 0.62 327.985 0.98 ;
      RECT  329.565 0.62 334.225 0.98 ;
      RECT  335.805 0.62 413.105 0.98 ;
      RECT  108.44 272.29 140.845 272.65 ;
      RECT  142.425 272.29 147.085 272.65 ;
      RECT  148.665 272.29 153.325 272.65 ;
      RECT  154.905 272.29 159.565 272.65 ;
      RECT  161.145 272.29 165.805 272.65 ;
      RECT  167.385 272.29 172.045 272.65 ;
      RECT  173.625 272.29 178.285 272.65 ;
      RECT  179.865 272.29 184.525 272.65 ;
      RECT  186.105 272.29 190.765 272.65 ;
      RECT  192.345 272.29 197.005 272.65 ;
      RECT  198.585 272.29 203.245 272.65 ;
      RECT  204.825 272.29 209.485 272.65 ;
      RECT  211.065 272.29 215.725 272.65 ;
      RECT  217.305 272.29 221.965 272.65 ;
      RECT  223.545 272.29 228.205 272.65 ;
      RECT  229.785 272.29 234.445 272.65 ;
      RECT  236.025 272.29 240.685 272.65 ;
      RECT  242.265 272.29 246.925 272.65 ;
      RECT  248.505 272.29 253.165 272.65 ;
      RECT  254.745 272.29 259.405 272.65 ;
      RECT  260.985 272.29 265.645 272.65 ;
      RECT  267.225 272.29 271.885 272.65 ;
      RECT  273.465 272.29 278.125 272.65 ;
      RECT  279.705 272.29 284.365 272.65 ;
      RECT  285.945 272.29 290.605 272.65 ;
      RECT  292.185 272.29 296.845 272.65 ;
      RECT  298.425 272.29 303.085 272.65 ;
      RECT  304.665 272.29 309.325 272.65 ;
      RECT  310.905 272.29 315.565 272.65 ;
      RECT  317.145 272.29 321.805 272.65 ;
      RECT  323.385 272.29 328.045 272.65 ;
      RECT  329.625 272.29 334.285 272.65 ;
      RECT  335.865 272.29 397.02 272.65 ;
      RECT  416.12 0.62 478.38 0.98 ;
      RECT  451.06 272.29 478.38 272.65 ;
      RECT  2.34 0.62 30.5 0.98 ;
      RECT  398.6 0.98 474.9 2.88 ;
      RECT  398.6 2.88 474.9 270.39 ;
      RECT  398.6 270.39 474.9 272.29 ;
      RECT  474.9 0.98 477.84 2.88 ;
      RECT  474.9 270.39 477.84 272.29 ;
      RECT  477.84 0.98 478.38 2.88 ;
      RECT  477.84 2.88 478.38 270.39 ;
      RECT  477.84 270.39 478.38 272.29 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 270.39 ;
      RECT  2.34 270.39 2.88 272.65 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 270.39 5.82 272.65 ;
      RECT  5.82 0.98 106.86 2.88 ;
      RECT  5.82 2.88 106.86 270.39 ;
      RECT  5.82 270.39 106.86 272.65 ;
   END
END    sky130_sram_512byte_1rw1r_32x128_8
END    LIBRARY
