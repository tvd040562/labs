* NGSPICE file created from cust_rom.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

.subckt cust_rom VGND VPWR addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6]
+ addr0[7] clk0 cs0 dout0[0] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15]
+ dout0[16] dout0[17] dout0[18] dout0[19] dout0[1] dout0[20] dout0[21] dout0[22] dout0[23]
+ dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[2] dout0[30] dout0[31]
+ dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9]
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1270_ _0076_ _0165_ net121 VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__a21o_1
X_1606_ net118 _0128_ _0343_ _0774_ _0110_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_14_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0985_ net135 _0803_ _0101_ _0806_ net124 VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__o311a_1
X_1399_ _0574_ _0579_ net175 net199 VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__o2bb2a_1
X_1537_ net111 _0717_ _0701_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__a21o_1
Xfanout138 net143 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_2
Xfanout127 net129 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__buf_2
X_1468_ _0039_ net53 _0212_ net80 VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__o211a_1
Xfanout149 net152 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
Xfanout116 net119 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__buf_2
Xfanout105 net106 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_37_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1253_ _0438_ _0439_ net104 VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__o21a_1
X_1322_ _0130_ _0235_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__nand2b_1
X_1184_ _0226_ _0372_ net76 _0757_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_20_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0968_ net94 net88 VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0899_ net150 net160 net139 VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__o21bai_2
XTAP_TAPCELL_ROW_2_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0822_ net158 net165 VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__and2b_1
XFILLER_0_51_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1236_ _0414_ _0422_ _0423_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_39_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1305_ _0049_ _0368_ _0488_ _0482_ net105 VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__o311a_1
X_1167_ _0355_ _0356_ net88 VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__o21a_1
X_1098_ _0055_ net56 net75 VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1021_ net126 _0086_ _0177_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1219_ net126 _0403_ _0405_ _0406_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold30 net16 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1570_ _0342_ _0747_ _0751_ _0743_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1004_ net55 net47 VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput31 net31 VGND VGND VPWR VPWR dout0[29] sky130_fd_sc_hd__buf_2
Xoutput20 net20 VGND VGND VPWR VPWR dout0[19] sky130_fd_sc_hd__buf_2
X_1622_ clknet_2_3__leaf_clk0 _0004_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1553_ _0724_ _0730_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__a21oi_1
X_1484_ net89 _0659_ _0660_ _0342_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0984_ _0178_ _0177_ _0086_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__and3b_1
X_1605_ net76 _0437_ net98 net85 VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1536_ _0085_ _0680_ _0702_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__o21ai_1
Xfanout139 net140 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_4
Xfanout117 net118 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_2
Xfanout128 net129 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1398_ _0652_ _0577_ _0578_ net175 VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__o31a_1
X_1467_ _0642_ _0643_ _0640_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__o21ai_1
Xfanout106 net108 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_37_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1252_ _0055_ _0067_ _0063_ net114 VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__o211a_1
X_1321_ net101 _0503_ _0504_ _0092_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__a31oi_1
X_1183_ net132 net68 net53 VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0967_ net113 _0157_ _0162_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_34_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1519_ net151 _0767_ net141 VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__a21o_1
X_0898_ net145 net154 net70 VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__o21a_2
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0821_ net153 net162 VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1235_ net89 _0420_ _0417_ net94 VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__o211a_1
X_1166_ net119 _0041_ _0048_ _0226_ net107 VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_39_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1304_ _0072_ _0114_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1097_ net136 _0736_ net60 _0103_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__or4_4
XFILLER_0_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1020_ net149 _0796_ _0050_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_44_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1149_ _0044_ net52 _0190_ net127 VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1218_ net45 _0112_ _0087_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold20 net26 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 net28 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1003_ net141 net168 _0067_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput21 net21 VGND VGND VPWR VPWR dout0[1] sky130_fd_sc_hd__buf_2
Xoutput10 net10 VGND VGND VPWR VPWR dout0[0] sky130_fd_sc_hd__buf_2
Xoutput32 net32 VGND VGND VPWR VPWR dout0[2] sky130_fd_sc_hd__buf_2
X_1552_ net91 _0731_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1621_ clknet_2_0__leaf_clk0 _0003_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dfxtp_1
X_1483_ _0161_ _0184_ net125 VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0983_ net127 _0040_ _0043_ _0045_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1535_ net43 _0714_ _0709_ _0708_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__a211o_1
Xfanout107 net108 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_4
Xfanout118 net119 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__buf_2
Xfanout129 addr0_reg\[4\] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
X_1604_ net118 _0048_ _0342_ _0732_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__o211a_1
X_1397_ net58 _0202_ _0318_ _0345_ _0571_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__o221a_1
X_1466_ _0474_ _0489_ net79 VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1320_ net62 _0095_ _0080_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__a21o_1
X_1182_ net136 _0736_ net53 VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__or3_2
X_1251_ net131 net68 net51 _0437_ net75 VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__o311a_1
XFILLER_0_24_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0966_ net57 _0153_ _0159_ net88 VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__o211a_1
X_0897_ _0089_ _0091_ _0093_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__a21o_1
X_1518_ net176 net181 _0692_ _0697_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__o22a_1
X_1449_ net116 _0228_ _0243_ _0626_ net106 VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__a311oi_2
XTAP_TAPCELL_ROW_2_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0820_ net160 net167 VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__xor2_2
XFILLER_0_36_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1303_ _0072_ _0114_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__nor2_1
X_1234_ _0344_ _0421_ net43 VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_39_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1165_ net45 _0112_ _0234_ net77 VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__o211a_1
X_1096_ _0652_ _0282_ _0288_ net89 VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0949_ net131 net66 VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1148_ _0334_ _0336_ _0338_ net88 net111 VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__a221o_1
X_1079_ net156 net54 _0068_ net136 VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__o211a_1
X_1217_ net135 _0798_ net79 VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold10 net30 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 net39 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 net27 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1002_ _0040_ _0057_ _0196_ _0126_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__o31a_1
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput33 net33 VGND VGND VPWR VPWR dout0[30] sky130_fd_sc_hd__buf_2
Xoutput11 net11 VGND VGND VPWR VPWR dout0[10] sky130_fd_sc_hd__buf_2
Xoutput22 net22 VGND VGND VPWR VPWR dout0[20] sky130_fd_sc_hd__buf_2
X_1551_ net117 _0185_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1482_ net135 _0123_ _0242_ net121 VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__o211ai_2
X_1620_ clknet_2_2__leaf_clk0 _0002_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_37_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_48_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0982_ net151 net160 net139 VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__or3b_2
XFILLER_0_14_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1603_ _0785_ _0782_ net195 net172 VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__a2bb2o_1
Xfanout108 addr0_reg\[5\] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_2
Xfanout119 addr0_reg\[4\] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_4
X_1534_ net141 _0248_ _0713_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1465_ net120 _0145_ _0641_ net109 VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__o31ai_1
X_1396_ _0563_ _0576_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1181_ _0361_ _0370_ net90 VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__a21oi_1
X_1250_ net154 net162 net130 net145 VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0896_ net102 net113 VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__nand2_4
X_0965_ net72 net69 VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1517_ _0652_ _0696_ net171 VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__a21o_1
X_1448_ _0064_ _0290_ net116 VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__a21oi_1
X_1379_ _0544_ _0545_ _0560_ _0176_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_25_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout90 net96 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_2
XFILLER_0_36_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_24_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1233_ net63 _0075_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1302_ _0471_ _0478_ _0486_ net100 net92 VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__o221a_1
X_1095_ _0274_ _0285_ _0287_ net108 net91 VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__o221a_1
X_1164_ net72 net62 _0104_ net117 VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_30_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0948_ net135 _0078_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0879_ net71 net66 _0798_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1216_ net131 net115 VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1147_ _0086_ _0226_ _0337_ _0241_ _0204_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__a32o_1
X_1078_ net153 net53 _0068_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold22 net18 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 net22 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1001_ _0114_ _0118_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput23 net23 VGND VGND VPWR VPWR dout0[21] sky130_fd_sc_hd__buf_2
Xoutput34 net34 VGND VGND VPWR VPWR dout0[31] sky130_fd_sc_hd__buf_2
XFILLER_0_43_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput12 net12 VGND VGND VPWR VPWR dout0[11] sky130_fd_sc_hd__buf_2
XFILLER_0_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1550_ net118 net137 _0183_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__and3_1
X_1481_ net70 _0124_ net75 VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_27_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0981_ net90 net98 VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__or2_2
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1602_ net174 _0784_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1533_ _0128_ _0184_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1395_ net126 _0037_ _0564_ _0575_ net111 VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__o311a_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1464_ net159 net52 _0451_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__o21a_1
Xfanout109 addr0_reg\[5\] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_2
XFILLER_0_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1180_ _0366_ _0369_ _0364_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_6_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0964_ net132 net68 VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0895_ net88 net83 VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__nor2_1
X_1516_ _0690_ _0695_ _0693_ _0681_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1447_ _0622_ _0624_ _0621_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__a21o_1
X_1378_ _0243_ _0540_ net57 VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_25_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout91 net96 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_2
Xfanout80 _0683_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_2
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1232_ _0127_ _0403_ _0419_ net58 VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_39_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1301_ net105 _0481_ _0483_ _0485_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__o22a_1
X_1163_ net175 _0348_ _0353_ _0331_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1094_ _0214_ _0286_ net74 VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0947_ net136 net63 net156 VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_30_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0878_ net139 net65 VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__nand2_4
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_41_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload0 clknet_2_0__leaf_clk0 VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_44_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1146_ net67 _0057_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__nand2_1
X_1215_ net142 net50 _0242_ net61 _0041_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1077_ _0237_ _0254_ _0270_ net185 net173 VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__o32a_1
Xhold23 net17 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 net14 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1000_ net110 _0193_ _0194_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1129_ _0126_ _0320_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput13 net13 VGND VGND VPWR VPWR dout0[12] sky130_fd_sc_hd__buf_2
Xoutput24 net24 VGND VGND VPWR VPWR dout0[22] sky130_fd_sc_hd__buf_2
Xoutput35 net35 VGND VGND VPWR VPWR dout0[3] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1480_ net176 net187 _0651_ _0657_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0980_ net94 net102 VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1532_ net94 _0711_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__nor2_1
X_1601_ _0776_ _0780_ _0781_ _0783_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1394_ net126 _0143_ _0484_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__nand3_1
X_1463_ net109 _0638_ _0639_ net88 VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__o31a_1
XFILLER_0_13_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0963_ net54 _0158_ _0127_ _0736_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0894_ net66 _0045_ _0048_ net51 net78 VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1515_ net42 _0210_ _0233_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__and3_1
X_1377_ net174 _0176_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1446_ net116 _0623_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout81 _0683_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout70 net71 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_4
Xfanout92 net96 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_2
X_1231_ net55 _0276_ _0202_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__o21a_1
X_1162_ _0343_ _0350_ _0352_ _0339_ net95 VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1300_ _0373_ _0484_ net74 VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1093_ _0034_ _0242_ _0095_ net69 VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__a2bb2o_1
X_0946_ net67 net59 VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__nor2_1
X_0877_ net135 _0072_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1429_ net111 _0132_ _0332_ _0593_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload1 clknet_2_2__leaf_clk0 VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_33_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1214_ net171 net203 VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1145_ net127 _0130_ _0335_ net102 VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__o31a_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1076_ _0110_ _0268_ _0269_ _0261_ net173 VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0929_ net70 _0123_ _0122_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__o21a_1
Xhold13 net33 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 net21 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_41_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1059_ net90 _0244_ _0247_ _0093_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__a31o_1
X_1128_ net71 net148 _0040_ _0124_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__a211o_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput36 net36 VGND VGND VPWR VPWR dout0[4] sky130_fd_sc_hd__buf_2
Xoutput25 net25 VGND VGND VPWR VPWR dout0[23] sky130_fd_sc_hd__buf_2
Xoutput14 net14 VGND VGND VPWR VPWR dout0[13] sky130_fd_sc_hd__buf_2
XFILLER_0_9_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1531_ _0708_ _0709_ _0710_ _0705_ _0701_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__o32a_1
X_1600_ net91 _0185_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__nor2_1
X_1462_ _0804_ _0201_ _0309_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1393_ _0652_ _0573_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0893_ net66 _0045_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__nand2_1
X_0962_ net159 net165 net133 VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_49_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1445_ _0804_ net49 _0284_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1514_ _0184_ _0308_ _0682_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__a21o_1
X_1376_ _0551_ _0557_ net90 _0549_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout82 _0683_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout71 net72 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_4
Xfanout93 net96 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_4
Xfanout60 net61 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
XFILLER_0_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1230_ _0408_ _0415_ _0417_ net94 VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__a31o_1
X_1092_ _0277_ _0284_ net77 VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__a21oi_1
X_1161_ _0065_ _0137_ _0351_ _0093_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0876_ net167 net150 VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0945_ net150 net67 _0073_ net135 VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__o211a_1
X_1428_ _0164_ _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__or2_1
X_1359_ _0105_ _0540_ net57 VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__a21o_1
Xclkload2 clknet_2_3__leaf_clk0 VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1213_ net9 net184 _0401_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__o21ba_1
X_1144_ net139 net151 net160 net167 VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__and4b_1
XFILLER_0_46_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1075_ _0263_ _0264_ net91 VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0928_ net153 net51 VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__xnor2_4
X_0859_ net71 _0035_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__nand2_1
Xhold25 net36 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 net15 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_41_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1058_ net118 _0250_ _0251_ _0106_ _0238_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__o32a_1
X_1127_ _0102_ _0318_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput26 net26 VGND VGND VPWR VPWR dout0[24] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR dout0[14] sky130_fd_sc_hd__buf_2
Xoutput37 net37 VGND VGND VPWR VPWR dout0[5] sky130_fd_sc_hd__buf_2
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_15_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1530_ _0058_ _0246_ _0177_ net43 VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__o211a_1
X_1392_ _0563_ _0566_ _0571_ _0572_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1461_ _0116_ _0497_ net122 VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0961_ net167 _0057_ _0154_ _0156_ net82 VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__o32a_1
XFILLER_0_40_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0892_ net64 net46 _0088_ _0071_ net115 VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1375_ net76 _0367_ _0556_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__or3b_1
XFILLER_0_10_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1513_ _0690_ _0691_ net96 _0685_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__o211a_1
X_1444_ _0251_ _0273_ net57 VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_33_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_18_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout94 net96 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_4
Xfanout83 net84 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_4
Xfanout72 _0694_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_4
Xfanout61 _0034_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_4
Xfanout50 _0069_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_4
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1091_ net143 net45 _0239_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__or3_1
X_1160_ net150 net161 _0073_ net127 VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__o211a_1
X_0944_ _0704_ net69 _0072_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0875_ net163 net145 VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__and2b_4
X_1427_ _0585_ _0605_ _0604_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_38_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1358_ _0078_ _0095_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__nand2_1
X_1289_ net71 _0124_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1212_ net95 _0394_ _0397_ _0400_ net175 VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__o221a_1
X_1143_ net78 _0332_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1074_ _0652_ _0267_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0927_ net159 net53 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_45_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0858_ net148 net165 net133 VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__a21bo_4
Xhold15 net34 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 net10 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_41_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1126_ net58 _0317_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__or2_1
X_1057_ net138 net65 _0120_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput38 net38 VGND VGND VPWR VPWR dout0[6] sky130_fd_sc_hd__buf_2
Xoutput27 net27 VGND VGND VPWR VPWR dout0[25] sky130_fd_sc_hd__buf_2
Xoutput16 net16 VGND VGND VPWR VPWR dout0[15] sky130_fd_sc_hd__buf_2
Xclkbuf_2_3__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_3__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ net113 _0301_ _0298_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1391_ net142 net69 net54 _0318_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1460_ net173 net183 _0632_ _0637_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1589_ net90 _0764_ _0768_ _0771_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_5_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0960_ net139 _0799_ _0800_ _0155_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1512_ _0323_ _0457_ net42 VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__o21a_1
X_0891_ net53 net46 VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__nand2_1
X_1443_ net84 _0620_ net97 VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__a21o_1
X_1374_ net136 _0072_ net156 VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__or3b_1
XFILLER_0_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout51 _0061_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_24_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout73 _0694_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_2
Xfanout62 _0033_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout95 net96 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout84 net87 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1090_ _0046_ _0158_ _0239_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0874_ net162 net48 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__nand2_2
X_0943_ net148 net68 VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__nor2_2
XFILLER_0_27_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1426_ net86 _0138_ _0142_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__or3_1
X_1357_ net170 net206 VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__and2_1
X_1288_ net163 net48 _0757_ net70 net56 VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1142_ net146 _0757_ _0246_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__o21ba_1
X_1211_ _0383_ _0399_ net95 VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1073_ net115 net60 _0266_ _0265_ _0805_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__o32a_1
X_0857_ net107 net118 VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__nand2_1
X_0926_ net134 _0798_ net56 VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold27 net41 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ _0127_ _0588_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__nor2_1
Xhold16 net11 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_41_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1125_ net149 net68 _0073_ net71 VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1056_ _0249_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput17 net17 VGND VGND VPWR VPWR dout0[16] sky130_fd_sc_hd__buf_2
X_0909_ _0101_ _0103_ net138 VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput28 net28 VGND VGND VPWR VPWR dout0[26] sky130_fd_sc_hd__buf_2
Xoutput39 net39 VGND VGND VPWR VPWR dout0[7] sky130_fd_sc_hd__buf_2
XFILLER_0_11_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1108_ _0184_ _0201_ _0204_ _0300_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__a31o_1
X_1039_ _0787_ net59 VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1390_ net108 _0569_ _0570_ net99 VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__o211a_1
X_1657_ clknet_2_1__leaf_clk0 net8 VGND VGND VPWR VPWR addr0_reg\[7\] sky130_fd_sc_hd__dfxtp_1
X_1588_ _0769_ _0770_ _0750_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0890_ _0055_ net56 VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1511_ net83 _0688_ _0689_ _0126_ net101 VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__a221o_1
X_1442_ net115 _0190_ _0373_ _0619_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__a31o_1
X_1373_ net90 _0546_ _0554_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_2_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout96 addr0_reg\[7\] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout63 net64 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_4
Xfanout52 _0061_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_24_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout85 net86 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_4
Xfanout74 net78 VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0942_ net63 _0137_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__nor2_1
X_0873_ net144 net153 VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1425_ net128 _0601_ _0603_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1287_ net134 _0071_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__and2_1
X_1356_ net173 net190 _0537_ _0538_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__o22a_1
XFILLER_0_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1141_ net143 _0068_ _0140_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__and3_1
X_1210_ _0384_ _0398_ net113 VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1072_ net64 _0145_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__nor2_1
X_0856_ net86 net82 VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0925_ net121 _0796_ _0075_ _0120_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__and4_1
Xhold28 net19 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ net64 _0114_ _0284_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__o21a_1
Xhold17 net12 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__dlygate4sd3_1
X_1339_ net130 _0796_ _0120_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1055_ net150 net69 net63 _0096_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__a211o_2
X_1124_ net93 _0314_ _0315_ net88 _0313_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__a311o_1
XFILLER_0_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput18 net18 VGND VGND VPWR VPWR dout0[17] sky130_fd_sc_hd__buf_2
Xoutput29 net29 VGND VGND VPWR VPWR dout0[27] sky130_fd_sc_hd__buf_2
X_0839_ net148 net133 VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__nand2b_1
X_0908_ _0101_ _0103_ net132 VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_11_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1107_ net160 _0055_ _0096_ _0777_ net128 VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1038_ net66 net59 VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1587_ net76 _0104_ _0115_ _0556_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__and4_1
X_1656_ clknet_2_0__leaf_clk0 net7 VGND VGND VPWR VPWR addr0_reg\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1510_ net135 _0183_ _0387_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__o21ai_1
X_1441_ _0807_ _0183_ _0035_ net74 VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__o211a_1
X_1372_ _0551_ _0553_ _0549_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_33_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1639_ clknet_2_1__leaf_clk0 _0021_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfxtp_1
Xfanout42 _0053_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
Xfanout64 _0032_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_2
XFILLER_0_36_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout53 _0060_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_4
Xfanout97 net100 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout75 net78 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_4
Xfanout86 net87 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0941_ net140 _0118_ _0136_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__or3_2
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0872_ net144 net153 VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__xor2_4
XPHY_EDGE_ROW_50_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1424_ net82 _0602_ net113 VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__a21o_1
X_1355_ net92 _0527_ _0533_ net170 VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_38_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1286_ net83 _0470_ net88 VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1140_ net171 net205 VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1071_ _0043_ _0059_ net75 VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__a21o_1
X_0924_ net151 net168 net157 VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__or3b_2
XFILLER_0_11_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0855_ net74 _0805_ _0037_ _0051_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__or4b_1
Xhold18 net31 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__dlygate4sd3_1
X_1407_ _0585_ _0586_ _0343_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__o21a_1
Xhold29 net38 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__dlygate4sd3_1
X_1338_ _0519_ _0520_ net97 VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__o21a_1
X_1269_ _0071_ _0074_ _0345_ net79 VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_7_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1054_ net150 net67 net55 VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__a21oi_1
X_1123_ _0045_ _0311_ _0310_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0907_ net156 net164 net146 VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__or3b_1
XFILLER_0_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput19 net19 VGND VGND VPWR VPWR dout0[18] sky130_fd_sc_hd__buf_2
XFILLER_0_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0838_ net144 net154 VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_19_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1106_ net86 _0293_ _0175_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1037_ _0078_ _0128_ _0230_ net135 VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1655_ clknet_2_1__leaf_clk0 net6 VGND VGND VPWR VPWR addr0_reg\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1586_ net119 _0146_ _0525_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_36_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1440_ net176 _0607_ _0616_ _0618_ _0600_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__a41o_1
X_1371_ net118 _0552_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1638_ clknet_2_2__leaf_clk0 _0020_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfxtp_1
X_1569_ net97 net103 _0749_ net92 VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_51_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout43 _0053_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
Xfanout76 net77 VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_2
Xfanout65 _0799_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_4
XFILLER_0_44_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout54 _0060_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_2
Xfanout98 net100 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_4
Xfanout87 _0673_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0940_ net167 net160 net151 VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__and3b_1
XFILLER_0_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0871_ net148 net158 VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__nand2_4
X_1423_ _0096_ _0136_ _0177_ _0086_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__o211ai_1
X_1354_ net92 _0536_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__nor2_1
X_1285_ _0215_ _0308_ _0469_ _0234_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_39_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1070_ net63 net46 _0107_ _0120_ net119 VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0854_ net130 _0798_ _0801_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__or3_1
X_0923_ net165 net50 _0118_ net133 VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__a211o_2
XFILLER_0_15_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_23_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold19 net29 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__dlygate4sd3_1
X_1406_ net82 _0075_ _0096_ net102 VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1268_ _0291_ _0333_ _0451_ _0453_ net104 VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__o221a_1
X_1337_ net74 _0063_ _0279_ net103 VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__a31o_1
X_1199_ net62 _0043_ net50 _0085_ net127 VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1122_ net121 _0065_ _0144_ _0190_ _0306_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__a41o_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1053_ _0202_ _0226_ _0246_ net118 VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0906_ net157 net164 net146 VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0837_ net144 net153 VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__and2b_1
XFILLER_0_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1105_ net119 _0294_ _0295_ _0297_ net86 VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_16_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1036_ net159 net53 VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1654_ clknet_2_1__leaf_clk0 net5 VGND VGND VPWR VPWR addr0_reg\[4\] sky130_fd_sc_hd__dfxtp_1
X_1585_ _0765_ _0766_ net98 VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1019_ net149 _0145_ _0213_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1370_ _0746_ _0057_ net50 _0807_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__a22o_1
X_1637_ clknet_2_0__leaf_clk0 _0019_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfxtp_1
X_1499_ net91 _0675_ _0677_ net170 VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__a31o_1
X_1568_ net98 net107 VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__nor2_1
Xfanout55 net56 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
Xfanout77 net78 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout88 _0662_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_4
Xfanout99 net100 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_2
Xfanout66 _0787_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0870_ net145 net155 VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__and2_2
XFILLER_0_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1422_ net142 _0068_ _0140_ _0283_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__a31o_1
X_1353_ _0521_ _0535_ _0530_ _0518_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__o2bb2a_1
X_1284_ net122 _0062_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0999_ net83 _0189_ _0191_ net93 VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_21_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0922_ net148 net158 net165 VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__nor3_2
X_0853_ net131 _0801_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__nor2_2
X_1405_ _0804_ _0058_ _0436_ net128 VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput1 addr0[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_1198_ _0068_ _0085_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__nand2_1
X_1267_ _0757_ _0304_ net120 VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__o21ai_2
X_1336_ _0102_ net116 _0051_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__and3b_1
XFILLER_0_14_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1052_ net137 net45 _0183_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__or3_4
X_1121_ _0307_ _0312_ net93 VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0905_ _0736_ net59 VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__nor2_2
XFILLER_0_28_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0836_ net146 net164 VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1319_ net134 _0069_ _0463_ _0055_ net120 VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1104_ _0808_ _0101_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1035_ net116 _0227_ _0228_ _0225_ net103 VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a311o_1
XFILLER_0_33_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0819_ net153 net162 VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__nor2_4
XFILLER_0_16_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1653_ clknet_2_1__leaf_clk0 net4 VGND VGND VPWR VPWR addr0_reg\[3\] sky130_fd_sc_hd__dfxtp_1
X_1584_ _0098_ _0296_ _0126_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1018_ _0055_ net44 VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1636_ clknet_2_3__leaf_clk0 _0018_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1567_ net114 _0113_ _0479_ _0522_ _0748_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__o32a_1
X_1498_ net57 _0676_ _0669_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__o21ai_1
Xfanout78 _0683_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
Xfanout89 _0662_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
Xfanout56 _0058_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_4
Xfanout67 net68 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1421_ net171 net204 VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__and2_1
X_1283_ net176 net193 _0462_ _0468_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__o22a_1
X_1352_ _0523_ _0534_ net104 VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_21_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0998_ _0131_ _0192_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1619_ clknet_2_2__leaf_clk0 _0001_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0921_ _0715_ net48 VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__nor2_2
XFILLER_0_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0852_ net123 _0042_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__nand2_2
X_1335_ _0516_ _0517_ net106 VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__a21oi_1
X_1404_ net126 _0062_ _0213_ _0583_ net111 VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__o311a_1
XFILLER_0_36_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1197_ _0384_ _0385_ net113 VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__o21a_1
X_1266_ _0067_ _0181_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__or2_1
Xinput2 addr0[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1051_ _0046_ _0158_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__nand2_1
X_1120_ _0262_ _0311_ _0310_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__o21ai_1
X_0904_ net156 net164 net146 VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0835_ net147 net164 VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1318_ net109 _0501_ _0499_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__a21o_1
X_1249_ net142 net68 net52 VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1103_ net55 _0129_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__nor2_1
X_1034_ _0068_ _0140_ net132 VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__a21o_1
X_0818_ net156 net164 VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1652_ clknet_2_1__leaf_clk0 net3 VGND VGND VPWR VPWR addr0_reg\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1583_ _0040_ net57 _0095_ _0188_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1017_ _0055_ net44 VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1635_ clknet_2_3__leaf_clk0 _0017_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfxtp_1
X_1497_ net47 _0335_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__nor2_1
X_1566_ net115 _0372_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout57 _0054_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_32_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout46 _0083_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_4
Xfanout68 _0777_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_4
Xfanout79 net80 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_2
XFILLER_0_51_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1420_ _0592_ _0599_ net175 net198 VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__o2bb2a_1
X_1351_ net145 net154 _0065_ _0349_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_46_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1282_ net93 _0467_ net176 VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1618_ clknet_2_0__leaf_clk0 _0000_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfxtp_1
X_0997_ net65 _0807_ _0059_ _0160_ net115 VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__a221o_1
X_1549_ net99 _0727_ _0729_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0920_ net60 _0103_ _0114_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__or3_2
X_0851_ net137 net146 net156 VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__or3_2
XFILLER_0_23_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1265_ net131 _0802_ _0068_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1334_ net132 net68 _0035_ _0265_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__a31o_1
X_1403_ net151 _0807_ _0045_ net69 net80 VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__a221o_1
Xinput3 addr0[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_1196_ net67 _0075_ _0349_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1050_ _0805_ _0102_ _0238_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0834_ net161 net168 net140 VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__o21ai_4
X_0903_ net53 _0095_ _0099_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1317_ _0431_ _0472_ _0500_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1248_ _0433_ _0434_ _0093_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__o21a_1
X_1179_ _0049_ _0367_ _0368_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1102_ net48 _0107_ net77 VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__a21o_1
X_1033_ net164 _0226_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0817_ net156 net164 VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__and2_2
XFILLER_0_24_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1651_ clknet_2_0__leaf_clk0 net2 VGND VGND VPWR VPWR addr0_reg\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1582_ net85 _0762_ _0763_ _0761_ net98 VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__o311a_1
XFILLER_0_44_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_14_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1016_ net121 _0188_ _0112_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__or3b_1
XFILLER_0_12_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1634_ clknet_2_3__leaf_clk0 _0016_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1496_ net85 _0674_ _0661_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1565_ _0744_ _0745_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout69 _0767_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_4
Xfanout58 _0054_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_32_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout47 _0083_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1281_ _0460_ _0464_ _0466_ _0450_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__o22a_1
X_1350_ net97 _0518_ _0532_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_46_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0996_ net80 _0065_ _0190_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__and3_1
X_1617_ net9 net191 _0559_ _0791_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__o22a_1
XFILLER_0_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1548_ net125 _0040_ _0479_ _0728_ net107 VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__o311a_1
X_1479_ net93 _0654_ _0656_ net171 VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0850_ net147 _0044_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__nor2_1
X_1402_ net108 _0580_ _0581_ net99 VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_11_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput4 addr0[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1264_ net84 _0448_ _0449_ net88 VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__a31o_1
X_1333_ _0473_ _0515_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1195_ _0800_ net47 _0178_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0979_ net171 net200 _0152_ _0174_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_2_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0902_ net54 _0098_ net77 VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__a21oi_2
X_0833_ net156 net164 net137 VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__o21a_2
XFILLER_0_51_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1316_ _0090_ _0473_ net120 VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1247_ net75 net48 _0108_ net88 VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__a31o_1
X_1178_ net163 _0056_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_44_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap44 _0118_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1032_ net137 net50 VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__nand2_4
X_1101_ _0801_ _0056_ _0115_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0816_ net175 VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1581_ _0804_ net49 _0515_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__o21a_1
X_1650_ clknet_2_0__leaf_clk0 net1 VGND VGND VPWR VPWR addr0_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1015_ _0050_ _0071_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1633_ clknet_2_0__leaf_clk0 _0015_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfxtp_1
X_1564_ net114 _0188_ _0442_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1495_ _0805_ _0102_ _0453_ _0663_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__o31a_1
XFILLER_0_39_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout48 _0070_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
Xfanout59 _0036_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_4
X_1280_ _0291_ _0333_ _0465_ net75 net104 VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_46_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0995_ net135 net148 net158 VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__nand3_4
X_1616_ net174 net189 _0793_ _0797_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__o22a_1
X_1547_ _0161_ _0184_ net77 VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__a21o_1
X_1478_ net110 _0655_ _0649_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__a21o_1
X_1401_ net136 _0117_ _0115_ net117 VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__o211a_1
Xinput5 addr0[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_1332_ net136 _0736_ net63 net60 net76 VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__o41a_1
X_1194_ net102 _0380_ _0382_ _0343_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__o31a_1
X_1263_ net44 _0183_ _0405_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0978_ _0652_ _0163_ _0173_ net176 VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__o31a_1
XFILLER_0_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0901_ net137 net48 VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0832_ net73 _0704_ net69 VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__or3_2
XFILLER_0_47_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1315_ net83 _0495_ _0498_ net101 VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__a31o_1
X_1177_ net61 _0055_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1246_ _0808_ net51 _0186_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap45 _0103_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1100_ net117 _0276_ _0278_ _0290_ _0292_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__a32o_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1031_ net62 _0051_ net116 VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0815_ net169 VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1229_ _0332_ _0368_ _0416_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_2__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_2__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
X_1580_ net76 _0623_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_13_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1014_ net42 _0200_ _0208_ _0197_ net95 VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1494_ _0665_ _0671_ net91 VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1632_ clknet_2_0__leaf_clk0 _0014_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfxtp_1
X_1563_ _0044_ _0525_ net114 VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout49 _0070_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_24_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0994_ net72 _0118_ _0183_ _0158_ net123 VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__o311a_1
X_1546_ net81 _0044_ _0277_ _0726_ net112 VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__a311oi_1
X_1615_ net172 _0791_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1477_ net123 _0086_ _0290_ _0645_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_20_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1400_ _0736_ net45 _0112_ _0278_ net77 VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__o311a_1
X_1331_ net176 net188 _0509_ _0514_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__o22a_1
Xinput6 addr0[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_1193_ net82 _0086_ _0226_ _0381_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__and4_1
X_1262_ net64 net46 _0095_ net120 VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0977_ _0169_ _0170_ _0172_ net101 VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__o31a_1
X_1529_ _0127_ _0277_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0900_ net124 _0073_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0831_ net137 net146 net67 VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1314_ _0496_ _0497_ net79 VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1176_ _0333_ _0365_ net57 VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__o21ai_1
X_1245_ net114 _0188_ _0430_ _0431_ net84 VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1030_ net142 net62 VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0814_ net144 VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__inv_2
X_1228_ net117 net65 _0059_ _0110_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__a31o_1
X_1159_ _0184_ _0349_ _0346_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1013_ net81 _0206_ _0207_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1631_ clknet_2_2__leaf_clk0 _0013_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfxtp_1
X_1493_ _0669_ _0670_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1562_ _0741_ _0742_ _0739_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_1_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_22 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0993_ net70 _0183_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__nor2_2
X_1614_ net194 _0795_ net174 VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1545_ net61 _0698_ _0410_ net125 VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1476_ _0642_ _0653_ _0640_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1330_ net93 _0511_ _0513_ net171 VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__a31o_1
X_1261_ net173 net192 _0447_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__o21ba_1
X_1192_ _0158_ _0239_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__or2_1
Xinput7 addr0[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
X_0976_ net68 _0046_ _0126_ _0171_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1528_ net102 _0706_ _0707_ _0343_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__o31a_1
X_1459_ net92 _0634_ _0636_ net170 VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0830_ net133 _0796_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__nand2_4
XFILLER_0_47_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1244_ net130 _0271_ net114 VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__o21ai_2
X_1313_ _0040_ _0068_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__nand2_1
X_1175_ net85 _0805_ _0202_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__or3b_1
X_0959_ net61 _0041_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0813_ net133 VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1227_ _0409_ _0414_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__or2_1
X_1158_ net72 net63 net81 VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__a21oi_4
X_1089_ _0274_ _0275_ _0281_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_7_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1012_ net127 _0201_ _0202_ net111 VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1630_ clknet_2_2__leaf_clk0 _0012_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfxtp_1
X_1492_ _0801_ net61 _0043_ net57 VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__or4_1
X_1561_ net70 net56 _0117_ _0658_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_1_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_35_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0992_ net73 _0184_ _0186_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1613_ net91 _0733_ _0794_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__mux2_1
X_1544_ _0127_ _0249_ _0721_ _0723_ net99 VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_41_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1475_ net134 _0124_ _0484_ net123 VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput8 addr0[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
X_1191_ net123 _0119_ _0379_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__and3_1
X_1260_ net92 _0441_ _0446_ net173 VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__o211a_1
X_0975_ net66 _0055_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__or2_1
X_1527_ _0787_ _0224_ _0041_ net81 VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__o211a_1
X_1458_ _0622_ _0635_ _0621_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__a21o_1
X_1389_ net65 _0062_ _0072_ net46 _0127_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_38_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1174_ net107 _0362_ _0363_ net98 VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__o31a_1
X_1243_ _0119_ _0181_ net114 VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__a21o_1
X_1312_ net62 net46 VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_22_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0958_ net139 net61 net127 VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__a21o_1
X_0889_ net139 net167 VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__nand2_4
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0812_ net118 VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1226_ net86 _0411_ _0412_ _0413_ net102 VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__a311o_1
X_1157_ _0339_ _0341_ _0347_ net95 VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__a31o_1
X_1088_ net78 _0276_ _0278_ _0280_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1011_ _0799_ _0807_ _0205_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1209_ _0069_ _0086_ _0349_ _0065_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_35_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1560_ net109 _0090_ _0233_ _0740_ net42 VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__a41o_1
X_1491_ net107 _0667_ _0668_ _0127_ net99 VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_49_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0991_ net139 net161 net168 net128 VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__o31a_2
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1612_ net98 _0722_ _0750_ _0774_ _0793_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__a221o_1
X_1543_ _0044_ _0277_ _0722_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_41_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1474_ _0644_ _0650_ net93 VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1190_ net158 net51 net133 VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__o21ai_1
Xinput9 cs0 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0974_ net165 _0039_ net42 _0806_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__o211a_1
X_1526_ _0808_ _0117_ _0158_ net52 net126 VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__o221a_1
X_1457_ _0099_ _0116_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__nand2_1
X_1388_ net117 _0143_ _0567_ _0568_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1311_ net71 net64 net48 _0085_ net122 VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1173_ net63 _0115_ _0249_ net118 VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__o211a_1
X_1242_ _0119_ _0181_ net114 VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0957_ _0075_ _0139_ _0143_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__o21a_1
X_0888_ net133 net165 VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__and2_2
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1509_ net127 _0686_ _0687_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0811_ net103 VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__inv_2
X_1225_ _0201_ _0234_ _0127_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__a21oi_1
X_1156_ _0049_ _0346_ _0343_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__a21o_1
X_1087_ net117 _0190_ _0246_ _0279_ net108 VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_7_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1010_ net55 _0158_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_12_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1208_ _0390_ _0392_ _0396_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__nor3_1
XFILLER_0_47_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1139_ _0316_ _0327_ _0330_ net177 net171 VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _0047_ _0251_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 net37 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1611_ _0343_ _0732_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__nor2_1
X_0990_ net73 _0184_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1542_ net77 _0129_ net85 VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__a21oi_1
X_1473_ net110 _0646_ _0649_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0973_ _0167_ _0168_ net83 VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1387_ _0040_ _0045_ net47 _0796_ net77 VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__o311a_1
X_1456_ _0627_ _0633_ net97 VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__o21ai_1
X_1525_ _0702_ _0703_ net87 VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_40_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1310_ _0487_ _0493_ _0494_ net182 net174 VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__o32a_1
X_1241_ net84 _0426_ _0427_ net100 VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__a31o_1
X_1172_ _0805_ _0037_ _0057_ net76 VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__o31a_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0956_ net93 _0151_ _0135_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__or3b_1
XFILLER_0_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0887_ net72 net158 VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__or2_1
X_1439_ _0175_ _0604_ _0617_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__nand3_1
X_1508_ net150 _0736_ _0183_ net72 net81 VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0810_ net102 VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1224_ net125 _0074_ _0367_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1155_ net126 _0344_ _0345_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__or3_1
X_1086_ net70 net60 _0072_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0939_ net87 _0134_ _0133_ net101 VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_7_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1207_ net42 _0084_ _0395_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_4_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1069_ _0262_ _0203_ _0226_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_35_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1138_ net171 _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 net32 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1610_ net186 _0792_ net174 VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1541_ _0086_ _0658_ _0720_ net112 VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1472_ net101 _0647_ _0648_ _0092_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_17_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0972_ net61 _0113_ net123 VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1524_ _0680_ _0387_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__nand2b_1
X_1386_ net169 _0129_ _0048_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__o21a_1
X_1455_ _0056_ _0097_ _0629_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1171_ _0358_ _0360_ _0357_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__o21ai_1
X_1240_ _0050_ net48 _0291_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0886_ net158 net133 VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0955_ net109 _0149_ _0150_ _0148_ net101 VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__o311a_1
X_1507_ net142 _0787_ net55 net52 _0808_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__o32a_1
X_1438_ net128 _0436_ _0484_ _0605_ net58 VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__a32o_1
X_1369_ net46 _0291_ _0550_ net107 VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__o31a_1
XFILLER_0_18_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_26_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1223_ net125 _0276_ _0410_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__nand3_1
X_1154_ net72 net50 VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__nor2_1
X_1085_ net147 net67 _0129_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0869_ _0063_ _0064_ _0065_ net116 VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__a31o_1
X_0938_ net79 _0116_ _0119_ _0121_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1206_ net167 net50 net59 VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__o21ai_1
X_1137_ net58 _0328_ _0326_ _0321_ _0175_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_35_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1068_ _0039_ _0072_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 net25 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_49_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1540_ net125 _0676_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1471_ _0122_ _0171_ net79 VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0971_ net166 _0084_ _0139_ _0039_ net80 VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__o221a_1
XFILLER_0_22_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1454_ _0625_ _0631_ net92 VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__a21oi_1
X_1523_ _0033_ _0043_ _0141_ net123 VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__a211o_1
X_1385_ net126 _0037_ _0564_ _0565_ net111 VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__o311a_1
XFILLER_0_42_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1170_ _0295_ _0359_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0885_ net103 _0052_ _0066_ _0081_ net97 VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__a311o_1
X_0954_ _0138_ _0141_ net124 VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__o21a_1
X_1437_ net89 _0613_ _0615_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__or3_1
X_1506_ _0682_ _0684_ _0681_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1368_ net50 _0112_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__nor2_1
X_1299_ net54 _0128_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__nand2_2
XFILLER_0_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1084_ net141 net69 VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__nand2_2
X_1222_ net151 _0767_ net63 _0129_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__a211o_1
X_1153_ net49 _0112_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0868_ net132 _0801_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__nand2_4
X_0937_ net121 _0125_ _0131_ _0132_ net109 VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout170 net172 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__buf_2
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1205_ _0390_ _0392_ _0393_ _0386_ _0383_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__o32a_1
X_1136_ _0078_ _0128_ _0119_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__a21boi_1
X_1067_ net105 _0255_ _0257_ _0260_ _0164_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_35_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold4 net23 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_49_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1119_ addr0_reg\[3\] net52 net46 _0715_ net122 VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1470_ net121 _0062_ _0479_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1599_ _0776_ _0780_ _0781_ _0652_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__o31a_1
XFILLER_0_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0970_ net142 _0139_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__or2_1
X_1522_ net111 _0700_ net102 VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1453_ _0627_ _0630_ net97 VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1384_ _0804_ net55 _0143_ net126 VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_45_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0884_ net121 _0077_ _0079_ _0080_ net84 VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__o221a_1
X_0953_ net68 net59 _0042_ net80 VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1436_ _0610_ _0614_ net94 _0608_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__o211a_1
X_1505_ _0309_ _0335_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__nor2_1
X_1367_ net103 _0547_ _0548_ net97 VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_37_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1298_ net105 _0482_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1221_ _0256_ _0344_ net42 VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__o21a_1
X_1152_ net89 net112 VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__nand2_4
X_1083_ _0802_ _0107_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0936_ net70 net149 _0802_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0867_ net132 net60 VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1419_ _0652_ _0595_ _0598_ net175 VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_6_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout160 net161 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_4
Xfanout171 net172 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1204_ net42 _0084_ _0137_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1066_ net119 _0259_ _0225_ net105 VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__a211oi_1
X_1135_ _0319_ _0321_ _0326_ _0164_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__a31o_1
X_0919_ net60 _0114_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__or2_1
Xhold5 net24 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1118_ net65 _0078_ _0308_ net109 VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__a31oi_1
X_1049_ _0805_ _0102_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_23_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1598_ net117 _0047_ _0296_ _0342_ _0732_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__o311a_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1521_ net129 _0044_ _0698_ _0699_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__a22o_1
X_1383_ net55 _0246_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__nor2_1
X_1452_ net60 _0097_ _0188_ _0629_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__o31a_1
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0952_ net79 _0076_ _0144_ _0147_ net84 VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__a311o_1
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0883_ net120 _0055_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__nand2_1
X_1504_ net83 _0232_ _0317_ net58 VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__o31a_1
XFILLER_0_49_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1435_ _0205_ _0272_ net125 VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__o21a_1
X_1366_ _0704_ _0114_ _0051_ net74 VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1297_ _0800_ _0807_ _0059_ _0095_ net119 VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1220_ _0093_ _0407_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__or2_1
X_1151_ net98 net85 VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__nor2_2
X_1082_ _0801_ _0804_ _0067_ _0099_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__o31a_1
X_0866_ net130 net60 net51 VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_15_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0935_ net79 _0130_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1418_ net112 _0596_ _0597_ _0587_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1349_ net74 _0531_ _0528_ net103 VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__o211a_1
Xfanout150 net151 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_4
Xfanout172 _0725_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout161 addr0_reg\[1\] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_29_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1203_ net102 _0391_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1134_ net83 _0325_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1065_ net131 _0120_ _0258_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__a21o_1
X_0849_ net138 net146 VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__or2_4
X_0918_ net153 net162 net130 VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__a21bo_4
XFILLER_0_11_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_1__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
Xhold6 net13 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dlygate4sd3_1
X_1117_ net127 net59 VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1048_ net151 net69 net73 VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__a21o_2
XFILLER_0_43_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1597_ _0045_ _0722_ _0778_ _0779_ net99 VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_51_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1520_ _0715_ _0128_ net125 VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__a21oi_1
X_1382_ net99 _0562_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__or2_1
X_1451_ _0088_ _0628_ net84 VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1649_ clknet_2_1__leaf_clk0 _0031_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0882_ net155 net51 net131 VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__a21oi_1
X_0951_ net56 _0075_ _0146_ net121 VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1503_ net101 _0679_ _0680_ _0092_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__a31o_1
X_1434_ _0608_ _0612_ net94 VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__a21oi_1
X_1365_ net130 _0124_ _0804_ net116 VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1296_ _0047_ _0049_ _0479_ _0480_ net121 VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__o32a_1
XFILLER_0_5_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1150_ net82 _0065_ _0137_ _0340_ _0093_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__a311o_1
X_1081_ _0272_ _0273_ net57 VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0934_ _0715_ _0129_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_15_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0865_ net71 _0035_ _0059_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__and3_1
X_1417_ _0367_ net81 _0276_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__or3b_1
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1279_ _0757_ _0304_ _0181_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__o21ai_1
X_1348_ net130 net51 _0068_ _0160_ _0059_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_38_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout140 net141 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__buf_2
Xfanout151 net152 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout173 net174 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_4
Xfanout162 net169 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_29_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1064_ _0108_ net44 VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__nor2_1
X_1133_ net80 _0808_ net59 _0322_ _0324_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__a41o_1
X_1202_ _0087_ _0372_ _0127_ _0757_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_47_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0848_ net133 net148 VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__nor2_4
X_0917_ _0082_ _0111_ net202 net173 VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_34_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7 net20 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1047_ net151 net69 VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1116_ net123 net59 VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_clk0 clk0 VGND VGND VPWR VPWR clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_8_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1596_ _0046_ _0129_ _0165_ net57 VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_34_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1450_ _0043_ net56 net115 VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__a21oi_1
X_1381_ _0258_ _0311_ _0425_ _0079_ net84 VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1648_ clknet_2_1__leaf_clk0 _0030_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dfxtp_1
X_1579_ net107 _0759_ _0760_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0950_ net132 net66 net48 VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__or3_1
X_0881_ net154 net51 VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__nand2_2
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1433_ net125 _0198_ _0611_ _0610_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__a31o_1
X_1502_ net71 _0796_ _0033_ net80 VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__a31o_1
X_1364_ _0541_ _0544_ _0545_ net98 VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__a31o_1
X_1295_ _0075_ _0139_ _0322_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1080_ net62 _0095_ net85 VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_15_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0933_ net147 net157 net138 VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_30_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0864_ net144 net162 VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_21_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1416_ net81 _0588_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1347_ net103 _0528_ _0529_ net97 VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__a31o_1
X_1278_ _0242_ _0463_ net58 VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout141 net142 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
Xfanout152 addr0_reg\[2\] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout174 net9 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_4
Xfanout163 net169 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__buf_1
Xfanout130 net132 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_29_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1201_ _0388_ _0389_ net113 VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1063_ _0256_ net81 _0800_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__or3b_1
XFILLER_0_34_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1132_ net56 _0114_ _0158_ _0101_ net124 VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__o221a_1
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0916_ net134 net53 VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__nor2_1
X_0847_ net139 net160 VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_3_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 net40 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1115_ net122 _0065_ _0144_ _0306_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__a31o_1
X_1046_ net136 net67 VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1595_ net117 _0437_ net107 VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1029_ net176 net178 _0221_ _0223_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1380_ net174 _0555_ _0558_ _0561_ _0539_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__a41o_1
XFILLER_0_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1647_ clknet_2_1__leaf_clk0 _0029_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dfxtp_1
X_1578_ _0045_ _0272_ net119 VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0880_ _0071_ _0074_ _0076_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1432_ net59 _0277_ net63 net61 VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__a211o_1
X_1363_ _0155_ _0479_ _0126_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__o21ai_1
X_1501_ _0304_ _0496_ net122 VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__a21o_1
X_1294_ net163 net50 net62 net131 VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__o211a_2
XFILLER_0_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0932_ net146 net157 net138 VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__o21a_2
XFILLER_0_15_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0863_ net144 net162 VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__xor2_2
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1415_ net111 _0594_ _0582_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__a21oi_1
X_1346_ net130 net51 _0160_ _0059_ net74 VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__a221o_1
X_1277_ net134 _0800_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__or2_1
Xfanout120 net122 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_2
Xfanout131 net132 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__buf_2
Xfanout142 net143 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__buf_2
Xfanout175 net176 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_29_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout153 net154 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_8
Xfanout164 net169 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1200_ _0199_ _0276_ net82 VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1062_ net168 _0075_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__nor2_1
X_1131_ net56 _0114_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0915_ net73 net62 VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__nand2_2
X_0846_ net140 net160 VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__nor2_2
XFILLER_0_11_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1329_ net109 _0507_ _0512_ _0505_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_49_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold9 net35 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_48_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1114_ _0304_ _0305_ net42 VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__a21oi_1
X_1045_ net148 net158 net166 VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__and3b_2
XFILLER_0_28_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0829_ net65 _0800_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1594_ _0296_ _0774_ _0775_ _0750_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1028_ net101 _0195_ _0209_ _0222_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1646_ clknet_2_1__leaf_clk0 _0028_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1577_ net76 net137 net147 net156 VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1500_ net174 net180 _0672_ _0678_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__o22a_1
X_1431_ _0154_ _0609_ net111 VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1293_ _0475_ _0477_ net104 VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1362_ net107 _0543_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1629_ clknet_2_2__leaf_clk0 _0011_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0931_ net112 net81 VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__nand2_4
XFILLER_0_15_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0862_ net144 net162 VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__or2_2
XFILLER_0_23_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1414_ net126 _0166_ _0242_ _0593_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1276_ _0450_ _0454_ _0460_ _0461_ net93 VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__o221a_1
X_1345_ _0046_ _0105_ net116 VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__a21o_1
Xfanout143 addr0_reg\[3\] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
Xfanout165 net166 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_4
Xfanout154 net155 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__buf_2
Xfanout110 addr0_reg\[5\] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
Xfanout132 addr0_reg\[3\] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_4
Xfanout121 net122 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_29_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout176 net9 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1130_ _0158_ _0183_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1061_ _0796_ _0078_ _0040_ net115 VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__a211o_1
X_0914_ _0100_ _0109_ _0110_ _0094_ net173 VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__o311a_1
X_0845_ net65 _0040_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1259_ _0428_ _0443_ _0445_ net92 VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_3_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1328_ net48 _0086_ _0235_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1044_ _0746_ _0107_ net77 VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_0_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1113_ net70 _0798_ _0801_ net104 VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__o31a_1
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0828_ net163 net155 VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_34_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1593_ _0046_ _0165_ _0713_ net125 VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1027_ _0164_ _0217_ _0219_ net176 VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_8_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1645_ clknet_2_1__leaf_clk0 _0027_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfxtp_1
X_1576_ net170 net207 VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1430_ net65 _0107_ _0120_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_22 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1361_ net76 _0245_ _0542_ _0359_ _0354_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__o32a_1
X_1292_ net120 _0181_ _0476_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1628_ clknet_2_0__leaf_clk0 _0010_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfxtp_1
X_1559_ _0803_ _0804_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0861_ net150 net167 VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__nor2_1
X_0930_ net83 net123 VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__nor2_4
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1413_ _0062_ _0213_ net81 VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__o21a_1
X_1275_ net42 _0108_ _0437_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__and3_1
X_1344_ net103 _0526_ _0521_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__a21bo_1
Xfanout111 net113 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_2
Xfanout166 net169 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout100 addr0_reg\[6\] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_2
Xfanout155 addr0_reg\[1\] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
Xfanout133 net134 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_4
Xfanout144 net152 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_4
Xfanout122 net124 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1060_ net90 _0252_ _0253_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_25_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0913_ net98 net85 VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__nand2_2
X_0844_ net141 net168 VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1189_ _0378_ _0371_ net197 net170 VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__a2bb2o_1
X_1327_ net109 _0510_ _0499_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__a21o_1
X_1258_ net104 _0444_ _0435_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_3_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1112_ net134 _0072_ _0239_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__or3_2
X_1043_ _0229_ _0236_ _0176_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_31_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0827_ net162 net153 VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__and2b_4
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1592_ _0046_ _0186_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__nand2_1
X_1026_ net113 _0179_ _0180_ _0220_ _0175_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__o311a_1
XPHY_EDGE_ROW_28_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1644_ clknet_2_1__leaf_clk0 _0026_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfxtp_1
X_1575_ net173 _0752_ _0754_ _0756_ _0737_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__a41o_1
XFILLER_0_21_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1009_ net128 net55 VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1360_ net136 net62 net49 VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1291_ net134 _0803_ _0139_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1627_ clknet_2_3__leaf_clk0 _0009_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1489_ _0295_ _0542_ _0666_ net117 VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__o22a_1
X_1558_ net103 _0738_ net97 VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0860_ net138 net61 VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__nor2_2
X_1412_ net94 _0591_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__or2_1
X_1343_ net114 _0524_ _0525_ _0523_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1274_ net87 _0455_ _0456_ _0459_ net101 VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__a311o_1
XFILLER_0_46_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0989_ net150 net160 net167 VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__nand3_4
Xfanout112 net113 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_2
Xfanout167 net168 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_4
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout134 net135 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
Xfanout101 addr0_reg\[6\] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_4
Xfanout145 net152 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
Xfanout123 net124 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_4
Xfanout156 net157 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0912_ net50 _0108_ _0105_ net74 VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__o211a_1
X_0843_ net139 net167 VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__and2b_4
XFILLER_0_45_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1326_ net120 net64 net46 _0442_ _0500_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_3_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1188_ net90 _0375_ _0377_ net170 VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__a31o_1
X_1257_ net115 _0063_ _0242_ _0438_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1111_ net171 net201 _0289_ _0303_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1042_ net79 _0231_ _0234_ _0235_ net83 VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0826_ net148 net165 VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__nand2_4
X_1309_ _0176_ _0491_ net173 VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1591_ net174 _0772_ _0773_ _0758_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1025_ net80 _0214_ _0215_ _0216_ net86 VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__a221o_1
X_0809_ net94 VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_16_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1 _0044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1643_ clknet_2_0__leaf_clk0 _0025_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfxtp_1
X_1574_ net104 _0431_ _0744_ _0755_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1008_ net128 _0202_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1290_ _0473_ _0474_ net120 VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_18_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1626_ clknet_2_3__leaf_clk0 _0008_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1488_ net72 net66 _0798_ _0801_ _0046_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__o32a_1
X_1557_ _0240_ _0349_ _0556_ _0226_ net74 VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__a32o_1
XFILLER_0_17_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1411_ _0587_ _0589_ _0590_ _0584_ _0582_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__o32a_1
X_1273_ _0457_ _0458_ _0126_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__o21a_1
X_1342_ _0075_ _0239_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0988_ net149 net158 net166 VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__and3_4
X_1609_ _0791_ net90 _0790_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__mux2_1
Xfanout113 addr0_reg\[5\] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_4
Xfanout102 addr0_reg\[6\] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout168 net169 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_4
Xfanout146 net147 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_4
Xfanout157 addr0_reg\[1\] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__buf_2
Xfanout135 addr0_reg\[3\] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_4
Xfanout124 addr0_reg\[4\] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_37_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0911_ net144 net162 net130 VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__a21o_1
X_0842_ net72 net65 VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__nand2_1
X_1325_ _0502_ _0508_ net93 VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__a21oi_1
X_1256_ _0429_ _0442_ net104 VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1187_ _0358_ _0376_ _0357_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1110_ _0298_ _0299_ _0302_ _0164_ net175 VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__o221a_1
XFILLER_0_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1041_ _0800_ _0044_ net122 VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__o21a_1
X_0825_ net160 net150 VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1308_ net104 _0492_ _0471_ net92 VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__a211oi_1
X_1239_ _0095_ _0425_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1590_ _0764_ _0768_ _0771_ _0731_ net90 VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__o32ai_1
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1024_ net80 _0210_ _0211_ _0218_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_50_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1642_ clknet_2_1__leaf_clk0 _0024_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfxtp_1
XANTENNA_2 _0065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1573_ net84 _0749_ _0176_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1007_ net137 net55 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__nand2_2
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1625_ clknet_2_1__leaf_clk0 _0007_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1556_ net170 net208 VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__and2_1
X_1487_ net85 _0664_ _0661_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1410_ _0808_ net49 _0112_ _0757_ net43 VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1341_ _0802_ _0045_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__nand2_1
X_1272_ net165 _0190_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_14_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0987_ net46 _0085_ _0178_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__or3_1
X_1539_ net175 net179 _0712_ _0719_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__o22a_1
X_1608_ net43 _0185_ net91 VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__a21oi_1
Xfanout125 net129 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__buf_2
Xfanout147 net152 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_2
Xfanout136 net143 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout114 net115 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__buf_2
Xfanout103 net106 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_4
Xfanout169 addr0_reg\[0\] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_4
Xfanout158 net159 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0910_ net146 net164 net137 VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__a21oi_2
X_0841_ _0704_ _0807_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1186_ net67 _0128_ _0295_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__a21oi_1
X_1255_ net114 net70 _0271_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__and3_1
X_1324_ net109 _0506_ _0507_ _0505_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1040_ net66 _0036_ _0129_ net67 VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__o22a_2
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0824_ net153 net144 VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__and2b_2
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1169_ net136 _0796_ _0059_ _0068_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__and4_1
X_1307_ net120 _0452_ _0476_ _0475_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__a31o_1
X_1238_ net75 net155 net53 _0404_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__o31a_1
XFILLER_0_34_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1023_ _0084_ _0097_ net110 VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1641_ clknet_2_3__leaf_clk0 _0023_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1572_ _0741_ _0753_ net92 _0739_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__a211o_1
XANTENNA_3 _0183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1006_ _0767_ net54 net140 VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput40 net40 VGND VGND VPWR VPWR dout0[8] sky130_fd_sc_hd__buf_2
XFILLER_0_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1555_ _0735_ _0734_ net196 net170 VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__a2bb2o_1
X_1624_ clknet_2_3__leaf_clk0 _0006_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dfxtp_1
X_1486_ _0106_ _0453_ _0663_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1340_ _0050_ _0522_ net75 VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1271_ net166 _0069_ _0158_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__a21oi_1
X_0986_ net131 _0802_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1538_ net94 _0716_ _0718_ net172 VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__a31o_1
X_1607_ _0786_ _0788_ _0789_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__or3_1
Xfanout137 net138 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_4
Xfanout126 net129 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__buf_2
Xfanout159 net161 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1469_ net123 _0290_ _0387_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__a31o_1
Xfanout104 net106 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_2
Xfanout148 net149 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__buf_4
Xfanout115 net116 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_2
XFILLER_0_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_19_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0840_ net147 _0808_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__nor2_2
X_1323_ net66 _0224_ _0215_ net79 VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__o211ai_2
X_1185_ _0366_ _0374_ _0364_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__a21bo_1
X_1254_ _0428_ _0432_ _0435_ _0440_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0969_ net71 _0757_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_2_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0823_ net158 net165 VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_43_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1306_ net105 _0481_ _0490_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__o21ba_1
X_1237_ net175 _0418_ _0424_ _0402_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_46_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1099_ net47 _0291_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__nor2_1
X_1168_ net76 _0048_ _0143_ _0227_ net85 VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__a41o_1
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_0__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1022_ _0182_ _0187_ net110 VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 _0658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1571_ net60 _0087_ _0658_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1640_ clknet_2_2__leaf_clk0 _0022_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1005_ _0198_ _0199_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput41 net41 VGND VGND VPWR VPWR dout0[9] sky130_fd_sc_hd__buf_2
Xoutput30 net30 VGND VGND VPWR VPWR dout0[28] sky130_fd_sc_hd__buf_2
XFILLER_0_50_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1554_ _0652_ _0724_ _0730_ net170 VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__a31o_1
X_1485_ _0806_ _0038_ _0137_ net127 VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__a31o_1
X_1623_ clknet_2_2__leaf_clk0 _0005_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dfxtp_1
.ends

