magic
tech sky130A
magscale 1 2
timestamp 1727228154
<< viali >>
rect 22109 37417 22143 37451
rect 22753 37417 22787 37451
rect 23397 37417 23431 37451
rect 25329 37417 25363 37451
rect 25973 37417 26007 37451
rect 27905 37417 27939 37451
rect 30205 37417 30239 37451
rect 32321 37417 32355 37451
rect 29837 37349 29871 37383
rect 22385 37145 22419 37179
rect 23029 37145 23063 37179
rect 23673 37145 23707 37179
rect 25605 37145 25639 37179
rect 26249 37145 26283 37179
rect 28181 37145 28215 37179
rect 29653 37145 29687 37179
rect 30481 37145 30515 37179
rect 32229 37145 32263 37179
rect 22385 35649 22419 35683
rect 22937 35445 22971 35479
rect 21833 35241 21867 35275
rect 24961 35105 24995 35139
rect 23213 35037 23247 35071
rect 22968 34969 23002 35003
rect 24409 34901 24443 34935
rect 23673 34697 23707 34731
rect 25421 34697 25455 34731
rect 28365 34697 28399 34731
rect 22293 34561 22327 34595
rect 22560 34561 22594 34595
rect 24041 34561 24075 34595
rect 24308 34561 24342 34595
rect 26065 34561 26099 34595
rect 26985 34561 27019 34595
rect 27252 34561 27286 34595
rect 29009 34561 29043 34595
rect 25513 34357 25547 34391
rect 28457 34357 28491 34391
rect 23581 34153 23615 34187
rect 23673 34153 23707 34187
rect 24133 34153 24167 34187
rect 24409 34153 24443 34187
rect 27077 34153 27111 34187
rect 24685 34085 24719 34119
rect 28917 34085 28951 34119
rect 21741 34017 21775 34051
rect 21833 34017 21867 34051
rect 22201 34017 22235 34051
rect 30113 34017 30147 34051
rect 21649 33949 21683 33983
rect 21925 33949 21959 33983
rect 22109 33949 22143 33983
rect 23857 33949 23891 33983
rect 23949 33949 23983 33983
rect 24225 33949 24259 33983
rect 24593 33949 24627 33983
rect 24777 33949 24811 33983
rect 24869 33949 24903 33983
rect 25053 33949 25087 33983
rect 25697 33949 25731 33983
rect 27537 33949 27571 33983
rect 22446 33881 22480 33915
rect 25964 33881 25998 33915
rect 27804 33881 27838 33915
rect 21465 33813 21499 33847
rect 29561 33813 29595 33847
rect 23305 33609 23339 33643
rect 23397 33609 23431 33643
rect 26157 33609 26191 33643
rect 27721 33609 27755 33643
rect 28825 33609 28859 33643
rect 22661 33473 22695 33507
rect 23121 33473 23155 33507
rect 23949 33473 23983 33507
rect 26341 33473 26375 33507
rect 26801 33473 26835 33507
rect 26985 33473 27019 33507
rect 27537 33473 27571 33507
rect 27905 33473 27939 33507
rect 27997 33473 28031 33507
rect 28273 33473 28307 33507
rect 29938 33473 29972 33507
rect 30849 33473 30883 33507
rect 22845 33405 22879 33439
rect 22937 33405 22971 33439
rect 26525 33405 26559 33439
rect 26617 33405 26651 33439
rect 28181 33405 28215 33439
rect 30205 33405 30239 33439
rect 23029 33337 23063 33371
rect 26433 33337 26467 33371
rect 30297 33269 30331 33303
rect 27721 33065 27755 33099
rect 28181 33065 28215 33099
rect 29561 33065 29595 33099
rect 32045 33065 32079 33099
rect 30021 32929 30055 32963
rect 32689 32929 32723 32963
rect 27905 32861 27939 32895
rect 27997 32861 28031 32895
rect 28273 32861 28307 32895
rect 29745 32861 29779 32895
rect 29837 32861 29871 32895
rect 29929 32861 29963 32895
rect 30205 32861 30239 32895
rect 30665 32861 30699 32895
rect 30932 32793 30966 32827
rect 32137 32725 32171 32759
rect 23489 32521 23523 32555
rect 23581 32521 23615 32555
rect 28825 32521 28859 32555
rect 31033 32521 31067 32555
rect 16129 32453 16163 32487
rect 29285 32453 29319 32487
rect 13185 32385 13219 32419
rect 13461 32385 13495 32419
rect 15853 32385 15887 32419
rect 19349 32385 19383 32419
rect 19441 32385 19475 32419
rect 21833 32385 21867 32419
rect 22017 32385 22051 32419
rect 23121 32385 23155 32419
rect 23305 32385 23339 32419
rect 23949 32385 23983 32419
rect 26157 32385 26191 32419
rect 26433 32385 26467 32419
rect 28365 32385 28399 32419
rect 28641 32385 28675 32419
rect 29101 32385 29135 32419
rect 29377 32385 29411 32419
rect 31217 32385 31251 32419
rect 31677 32385 31711 32419
rect 13369 32317 13403 32351
rect 16037 32317 16071 32351
rect 23857 32317 23891 32351
rect 25789 32317 25823 32351
rect 26249 32317 26283 32351
rect 28457 32317 28491 32351
rect 29469 32317 29503 32351
rect 31401 32317 31435 32351
rect 31493 32317 31527 32351
rect 15669 32249 15703 32283
rect 28917 32249 28951 32283
rect 31309 32249 31343 32283
rect 13185 32181 13219 32215
rect 13645 32181 13679 32215
rect 15945 32181 15979 32215
rect 19349 32181 19383 32215
rect 19717 32181 19751 32215
rect 22201 32181 22235 32215
rect 23213 32181 23247 32215
rect 23949 32181 23983 32215
rect 25973 32181 26007 32215
rect 26433 32181 26467 32215
rect 26525 32181 26559 32215
rect 28365 32181 28399 32215
rect 29377 32181 29411 32215
rect 29745 32181 29779 32215
rect 11069 31977 11103 32011
rect 11437 31977 11471 32011
rect 13553 31977 13587 32011
rect 17233 31977 17267 32011
rect 17693 31977 17727 32011
rect 19257 31977 19291 32011
rect 19809 31977 19843 32011
rect 23029 31977 23063 32011
rect 23213 31977 23247 32011
rect 23765 31977 23799 32011
rect 24225 31977 24259 32011
rect 26065 31977 26099 32011
rect 26525 31977 26559 32011
rect 26617 31977 26651 32011
rect 20177 31909 20211 31943
rect 11069 31841 11103 31875
rect 26157 31841 26191 31875
rect 31125 31841 31159 31875
rect 10977 31773 11011 31807
rect 11253 31773 11287 31807
rect 13185 31773 13219 31807
rect 13369 31773 13403 31807
rect 17233 31773 17267 31807
rect 17417 31773 17451 31807
rect 17509 31773 17543 31807
rect 19257 31773 19291 31807
rect 19349 31773 19383 31807
rect 19809 31773 19843 31807
rect 19993 31773 20027 31807
rect 21925 31773 21959 31807
rect 22109 31773 22143 31807
rect 22845 31773 22879 31807
rect 23029 31773 23063 31807
rect 23949 31773 23983 31807
rect 24041 31773 24075 31807
rect 26341 31773 26375 31807
rect 26801 31773 26835 31807
rect 26985 31773 27019 31807
rect 29377 31773 29411 31807
rect 31309 31773 31343 31807
rect 31493 31773 31527 31807
rect 22293 31705 22327 31739
rect 24225 31705 24259 31739
rect 26065 31705 26099 31739
rect 19625 31637 19659 31671
rect 28089 31637 28123 31671
rect 33609 31433 33643 31467
rect 11161 31365 11195 31399
rect 20729 31365 20763 31399
rect 28549 31365 28583 31399
rect 31309 31365 31343 31399
rect 33977 31365 34011 31399
rect 35633 31365 35667 31399
rect 11345 31297 11379 31331
rect 14565 31297 14599 31331
rect 14749 31297 14783 31331
rect 14841 31297 14875 31331
rect 15301 31297 15335 31331
rect 15485 31297 15519 31331
rect 19625 31297 19659 31331
rect 20085 31297 20119 31331
rect 20269 31297 20303 31331
rect 20545 31297 20579 31331
rect 22293 31297 22327 31331
rect 22569 31297 22603 31331
rect 24409 31297 24443 31331
rect 24593 31297 24627 31331
rect 26249 31297 26283 31331
rect 26525 31297 26559 31331
rect 28181 31297 28215 31331
rect 28733 31297 28767 31331
rect 31125 31297 31159 31331
rect 32873 31297 32907 31331
rect 33149 31297 33183 31331
rect 33793 31297 33827 31331
rect 35817 31297 35851 31331
rect 19717 31229 19751 31263
rect 20453 31229 20487 31263
rect 22477 31229 22511 31263
rect 26433 31229 26467 31263
rect 33057 31229 33091 31263
rect 15117 31161 15151 31195
rect 30941 31161 30975 31195
rect 33333 31161 33367 31195
rect 35449 31161 35483 31195
rect 10977 31093 11011 31127
rect 14841 31093 14875 31127
rect 15025 31093 15059 31127
rect 19625 31093 19659 31127
rect 19993 31093 20027 31127
rect 20821 31093 20855 31127
rect 22109 31093 22143 31127
rect 22385 31093 22419 31127
rect 24777 31093 24811 31127
rect 26065 31093 26099 31127
rect 26433 31093 26467 31127
rect 28917 31093 28951 31127
rect 33149 31093 33183 31127
rect 33425 31093 33459 31127
rect 12173 30889 12207 30923
rect 14841 30889 14875 30923
rect 22569 30889 22603 30923
rect 23489 30889 23523 30923
rect 23673 30889 23707 30923
rect 26065 30889 26099 30923
rect 26617 30889 26651 30923
rect 27353 30889 27387 30923
rect 27721 30889 27755 30923
rect 28733 30889 28767 30923
rect 33701 30889 33735 30923
rect 35725 30889 35759 30923
rect 36185 30889 36219 30923
rect 28549 30821 28583 30855
rect 12357 30753 12391 30787
rect 22385 30753 22419 30787
rect 33793 30753 33827 30787
rect 12449 30685 12483 30719
rect 22293 30685 22327 30719
rect 22569 30685 22603 30719
rect 23673 30685 23707 30719
rect 23765 30685 23799 30719
rect 26249 30685 26283 30719
rect 26341 30685 26375 30719
rect 27353 30685 27387 30719
rect 27445 30685 27479 30719
rect 28733 30685 28767 30719
rect 28917 30685 28951 30719
rect 33977 30685 34011 30719
rect 35909 30685 35943 30719
rect 36001 30685 36035 30719
rect 36185 30685 36219 30719
rect 12173 30617 12207 30651
rect 14381 30617 14415 30651
rect 14473 30617 14507 30651
rect 14657 30617 14691 30651
rect 20637 30617 20671 30651
rect 20821 30617 20855 30651
rect 23949 30617 23983 30651
rect 26065 30617 26099 30651
rect 26801 30617 26835 30651
rect 26985 30617 27019 30651
rect 33701 30617 33735 30651
rect 12633 30549 12667 30583
rect 20453 30549 20487 30583
rect 21005 30549 21039 30583
rect 22753 30549 22787 30583
rect 26525 30549 26559 30583
rect 33517 30549 33551 30583
rect 34161 30549 34195 30583
rect 18521 30345 18555 30379
rect 24501 30345 24535 30379
rect 10057 30277 10091 30311
rect 15945 30277 15979 30311
rect 18613 30277 18647 30311
rect 18981 30277 19015 30311
rect 23581 30277 23615 30311
rect 23949 30277 23983 30311
rect 35173 30277 35207 30311
rect 35357 30277 35391 30311
rect 9781 30209 9815 30243
rect 13093 30209 13127 30243
rect 15761 30209 15795 30243
rect 16129 30209 16163 30243
rect 17233 30209 17267 30243
rect 17509 30209 17543 30243
rect 18061 30209 18095 30243
rect 18353 30209 18387 30243
rect 18797 30209 18831 30243
rect 22661 30209 22695 30243
rect 22845 30209 22879 30243
rect 23397 30209 23431 30243
rect 24041 30209 24075 30243
rect 24317 30209 24351 30243
rect 29101 30209 29135 30243
rect 29377 30209 29411 30243
rect 29929 30209 29963 30243
rect 30205 30209 30239 30243
rect 30481 30209 30515 30243
rect 30757 30209 30791 30243
rect 31217 30209 31251 30243
rect 31493 30209 31527 30243
rect 32321 30209 32355 30243
rect 32597 30209 32631 30243
rect 34989 30209 35023 30243
rect 9873 30141 9907 30175
rect 13185 30141 13219 30175
rect 17325 30141 17359 30175
rect 18153 30141 18187 30175
rect 24225 30141 24259 30175
rect 29285 30141 29319 30175
rect 30113 30141 30147 30175
rect 30573 30141 30607 30175
rect 31309 30141 31343 30175
rect 32505 30141 32539 30175
rect 17693 30073 17727 30107
rect 23765 30073 23799 30107
rect 30389 30073 30423 30107
rect 30941 30073 30975 30107
rect 31033 30073 31067 30107
rect 32137 30073 32171 30107
rect 9413 30005 9447 30039
rect 9597 30005 9631 30039
rect 10057 30005 10091 30039
rect 13277 30005 13311 30039
rect 13461 30005 13495 30039
rect 17233 30005 17267 30039
rect 18061 30005 18095 30039
rect 22477 30005 22511 30039
rect 24041 30005 24075 30039
rect 29377 30005 29411 30039
rect 29561 30005 29595 30039
rect 29929 30005 29963 30039
rect 30481 30005 30515 30039
rect 31217 30005 31251 30039
rect 32321 30005 32355 30039
rect 9137 29801 9171 29835
rect 11621 29801 11655 29835
rect 13737 29801 13771 29835
rect 14289 29801 14323 29835
rect 16221 29801 16255 29835
rect 16773 29801 16807 29835
rect 18797 29801 18831 29835
rect 19073 29801 19107 29835
rect 19257 29801 19291 29835
rect 21005 29801 21039 29835
rect 26157 29801 26191 29835
rect 26893 29801 26927 29835
rect 27077 29801 27111 29835
rect 28733 29801 28767 29835
rect 30021 29801 30055 29835
rect 30389 29801 30423 29835
rect 31769 29801 31803 29835
rect 32137 29801 32171 29835
rect 35173 29801 35207 29835
rect 13921 29733 13955 29767
rect 16589 29733 16623 29767
rect 19717 29733 19751 29767
rect 29101 29733 29135 29767
rect 32689 29733 32723 29767
rect 11713 29665 11747 29699
rect 14473 29665 14507 29699
rect 16313 29665 16347 29699
rect 18797 29665 18831 29699
rect 19441 29665 19475 29699
rect 20913 29665 20947 29699
rect 26801 29665 26835 29699
rect 28733 29665 28767 29699
rect 31769 29665 31803 29699
rect 8953 29597 8987 29631
rect 9137 29597 9171 29631
rect 11621 29597 11655 29631
rect 11897 29597 11931 29631
rect 13553 29597 13587 29631
rect 13645 29597 13679 29631
rect 14289 29597 14323 29631
rect 14565 29597 14599 29631
rect 16129 29597 16163 29631
rect 16405 29597 16439 29631
rect 18710 29597 18744 29631
rect 19533 29597 19567 29631
rect 19991 29597 20025 29631
rect 21097 29597 21131 29631
rect 26157 29597 26191 29631
rect 26249 29597 26283 29631
rect 26709 29597 26743 29631
rect 28917 29597 28951 29631
rect 30021 29597 30055 29631
rect 30205 29597 30239 29631
rect 31684 29597 31718 29631
rect 31993 29597 32027 29631
rect 32321 29597 32355 29631
rect 35173 29597 35207 29631
rect 35265 29597 35299 29631
rect 36093 29597 36127 29631
rect 44557 29597 44591 29631
rect 16949 29529 16983 29563
rect 17141 29529 17175 29563
rect 17785 29529 17819 29563
rect 17969 29529 18003 29563
rect 19282 29529 19316 29563
rect 19809 29529 19843 29563
rect 20821 29529 20855 29563
rect 28641 29529 28675 29563
rect 32505 29529 32539 29563
rect 9321 29461 9355 29495
rect 11437 29461 11471 29495
rect 14105 29461 14139 29495
rect 18153 29461 18187 29495
rect 20177 29461 20211 29495
rect 21281 29461 21315 29495
rect 25881 29461 25915 29495
rect 35541 29461 35575 29495
rect 44373 29461 44407 29495
rect 7665 29257 7699 29291
rect 11989 29257 12023 29291
rect 12909 29257 12943 29291
rect 17601 29257 17635 29291
rect 29377 29257 29411 29291
rect 37749 29257 37783 29291
rect 7205 29189 7239 29223
rect 10517 29189 10551 29223
rect 17417 29189 17451 29223
rect 21833 29189 21867 29223
rect 22385 29189 22419 29223
rect 24593 29189 24627 29223
rect 28089 29189 28123 29223
rect 28273 29189 28307 29223
rect 34989 29189 35023 29223
rect 35081 29189 35115 29223
rect 37289 29189 37323 29223
rect 37473 29189 37507 29223
rect 7481 29121 7515 29155
rect 10793 29121 10827 29155
rect 11529 29121 11563 29155
rect 11805 29121 11839 29155
rect 13093 29121 13127 29155
rect 13369 29121 13403 29155
rect 17233 29121 17267 29155
rect 19073 29121 19107 29155
rect 19257 29121 19291 29155
rect 19349 29121 19383 29155
rect 22109 29121 22143 29155
rect 22569 29121 22603 29155
rect 24869 29121 24903 29155
rect 26341 29121 26375 29155
rect 26525 29121 26559 29155
rect 28906 29121 28940 29155
rect 29193 29121 29227 29155
rect 31125 29121 31159 29155
rect 31401 29121 31435 29155
rect 33701 29121 33735 29155
rect 33885 29121 33919 29155
rect 34069 29121 34103 29155
rect 34713 29121 34747 29155
rect 35350 29121 35384 29155
rect 35633 29121 35667 29155
rect 35909 29121 35943 29155
rect 38752 29121 38786 29155
rect 40601 29121 40635 29155
rect 44281 29121 44315 29155
rect 7389 29053 7423 29087
rect 10701 29053 10735 29087
rect 11621 29053 11655 29087
rect 13277 29053 13311 29087
rect 21925 29053 21959 29087
rect 24685 29053 24719 29087
rect 29101 29053 29135 29087
rect 31217 29053 31251 29087
rect 34805 29053 34839 29087
rect 35265 29053 35299 29087
rect 35725 29053 35759 29087
rect 38485 29053 38519 29087
rect 10977 28985 11011 29019
rect 19533 28985 19567 29019
rect 22293 28985 22327 29019
rect 28457 28985 28491 29019
rect 31585 28985 31619 29019
rect 34529 28985 34563 29019
rect 35541 28985 35575 29019
rect 36093 28985 36127 29019
rect 37657 28985 37691 29019
rect 39865 28985 39899 29019
rect 44465 28985 44499 29019
rect 7205 28917 7239 28951
rect 10701 28917 10735 28951
rect 11621 28917 11655 28951
rect 13093 28917 13127 28951
rect 19257 28917 19291 28951
rect 21833 28917 21867 28951
rect 22661 28917 22695 28951
rect 24869 28917 24903 28951
rect 25053 28917 25087 28951
rect 26341 28917 26375 28951
rect 26709 28917 26743 28951
rect 29101 28917 29135 28951
rect 31125 28917 31159 28951
rect 34713 28917 34747 28951
rect 35081 28917 35115 28951
rect 35817 28917 35851 28951
rect 39957 28917 39991 28951
rect 8953 28713 8987 28747
rect 9321 28713 9355 28747
rect 10885 28713 10919 28747
rect 11345 28713 11379 28747
rect 22937 28713 22971 28747
rect 23305 28713 23339 28747
rect 26985 28713 27019 28747
rect 27537 28713 27571 28747
rect 28825 28713 28859 28747
rect 29285 28713 29319 28747
rect 31585 28713 31619 28747
rect 37381 28713 37415 28747
rect 38209 28713 38243 28747
rect 38485 28713 38519 28747
rect 33241 28645 33275 28679
rect 36001 28645 36035 28679
rect 11069 28577 11103 28611
rect 23305 28577 23339 28611
rect 27077 28577 27111 28611
rect 27721 28577 27755 28611
rect 29193 28577 29227 28611
rect 38025 28577 38059 28611
rect 38761 28577 38795 28611
rect 38945 28577 38979 28611
rect 9137 28509 9171 28543
rect 9321 28509 9355 28543
rect 11161 28509 11195 28543
rect 18153 28509 18187 28543
rect 23121 28509 23155 28543
rect 26985 28509 27019 28543
rect 27261 28509 27295 28543
rect 27813 28509 27847 28543
rect 28969 28509 29003 28543
rect 31217 28509 31251 28543
rect 35817 28509 35851 28543
rect 38209 28509 38243 28543
rect 38669 28509 38703 28543
rect 38853 28509 38887 28543
rect 39129 28509 39163 28543
rect 41245 28509 41279 28543
rect 10425 28441 10459 28475
rect 10609 28441 10643 28475
rect 10793 28441 10827 28475
rect 10885 28441 10919 28475
rect 17969 28441 18003 28475
rect 18245 28441 18279 28475
rect 18429 28441 18463 28475
rect 23397 28441 23431 28475
rect 27537 28441 27571 28475
rect 28365 28441 28399 28475
rect 28549 28441 28583 28475
rect 29285 28441 29319 28475
rect 31401 28441 31435 28475
rect 32873 28441 32907 28475
rect 33057 28441 33091 28475
rect 34989 28441 35023 28475
rect 35173 28441 35207 28475
rect 35633 28441 35667 28475
rect 36093 28441 36127 28475
rect 37933 28441 37967 28475
rect 41512 28441 41546 28475
rect 17785 28373 17819 28407
rect 18613 28373 18647 28407
rect 27445 28373 27479 28407
rect 27997 28373 28031 28407
rect 28733 28373 28767 28407
rect 32689 28373 32723 28407
rect 35357 28373 35391 28407
rect 38393 28373 38427 28407
rect 42625 28373 42659 28407
rect 8401 28169 8435 28203
rect 10885 28169 10919 28203
rect 16313 28169 16347 28203
rect 23673 28169 23707 28203
rect 26801 28169 26835 28203
rect 27445 28169 27479 28203
rect 27537 28169 27571 28203
rect 29561 28169 29595 28203
rect 37657 28169 37691 28203
rect 8217 28101 8251 28135
rect 10425 28101 10459 28135
rect 14657 28101 14691 28135
rect 18613 28101 18647 28135
rect 19533 28101 19567 28135
rect 20453 28101 20487 28135
rect 26985 28101 27019 28135
rect 28825 28101 28859 28135
rect 29193 28101 29227 28135
rect 29745 28101 29779 28135
rect 36553 28101 36587 28135
rect 36737 28101 36771 28135
rect 37289 28101 37323 28135
rect 42165 28101 42199 28135
rect 6377 28033 6411 28067
rect 6653 28033 6687 28067
rect 8033 28033 8067 28067
rect 10701 28033 10735 28067
rect 13185 28033 13219 28067
rect 13461 28033 13495 28067
rect 14841 28033 14875 28067
rect 14933 28033 14967 28067
rect 15209 28033 15243 28067
rect 15485 28033 15519 28067
rect 15853 28033 15887 28067
rect 16129 28033 16163 28067
rect 18797 28033 18831 28067
rect 18889 28033 18923 28067
rect 19165 28033 19199 28067
rect 19349 28033 19383 28067
rect 20637 28033 20671 28067
rect 23305 28033 23339 28067
rect 24409 28033 24443 28067
rect 24685 28033 24719 28067
rect 26341 28033 26375 28067
rect 26617 28033 26651 28067
rect 27261 28033 27295 28067
rect 27721 28033 27755 28067
rect 27905 28033 27939 28067
rect 29009 28033 29043 28067
rect 29929 28033 29963 28067
rect 32689 28033 32723 28067
rect 37473 28033 37507 28067
rect 42993 28033 43027 28067
rect 43269 28033 43303 28067
rect 44281 28033 44315 28067
rect 6561 27965 6595 27999
rect 10609 27965 10643 27999
rect 13277 27965 13311 27999
rect 15301 27965 15335 27999
rect 16037 27965 16071 27999
rect 23397 27965 23431 27999
rect 24501 27965 24535 27999
rect 26525 27965 26559 27999
rect 27077 27965 27111 27999
rect 32781 27965 32815 27999
rect 41889 27965 41923 27999
rect 6837 27897 6871 27931
rect 15117 27897 15151 27931
rect 44465 27897 44499 27931
rect 6653 27829 6687 27863
rect 10425 27829 10459 27863
rect 13461 27829 13495 27863
rect 13645 27829 13679 27863
rect 14933 27829 14967 27863
rect 15209 27829 15243 27863
rect 15669 27829 15703 27863
rect 16129 27829 16163 27863
rect 18613 27829 18647 27863
rect 19073 27829 19107 27863
rect 20821 27829 20855 27863
rect 23305 27829 23339 27863
rect 24409 27829 24443 27863
rect 24869 27829 24903 27863
rect 26341 27829 26375 27863
rect 26985 27829 27019 27863
rect 27721 27829 27755 27863
rect 32689 27829 32723 27863
rect 33057 27829 33091 27863
rect 36921 27829 36955 27863
rect 42441 27829 42475 27863
rect 43361 27829 43395 27863
rect 6009 27625 6043 27659
rect 6561 27625 6595 27659
rect 6745 27625 6779 27659
rect 10149 27625 10183 27659
rect 13369 27625 13403 27659
rect 19809 27625 19843 27659
rect 21925 27625 21959 27659
rect 26709 27625 26743 27659
rect 26893 27625 26927 27659
rect 26985 27625 27019 27659
rect 29837 27625 29871 27659
rect 31953 27625 31987 27659
rect 33149 27625 33183 27659
rect 34713 27625 34747 27659
rect 35173 27625 35207 27659
rect 35541 27625 35575 27659
rect 37381 27625 37415 27659
rect 42073 27625 42107 27659
rect 42533 27625 42567 27659
rect 10333 27557 10367 27591
rect 13553 27557 13587 27591
rect 22385 27557 22419 27591
rect 27353 27557 27387 27591
rect 35265 27557 35299 27591
rect 9965 27489 9999 27523
rect 13277 27489 13311 27523
rect 17417 27489 17451 27523
rect 19993 27489 20027 27523
rect 22017 27489 22051 27523
rect 29653 27489 29687 27523
rect 33333 27489 33367 27523
rect 34805 27489 34839 27523
rect 35541 27489 35575 27523
rect 39865 27489 39899 27523
rect 41981 27489 42015 27523
rect 5825 27421 5859 27455
rect 6009 27421 6043 27455
rect 6377 27421 6411 27455
rect 6561 27421 6595 27455
rect 10149 27421 10183 27455
rect 13369 27421 13403 27455
rect 19809 27421 19843 27455
rect 20078 27421 20112 27455
rect 22201 27421 22235 27455
rect 26525 27421 26559 27455
rect 26709 27421 26743 27455
rect 26985 27421 27019 27455
rect 27169 27421 27203 27455
rect 29837 27421 29871 27455
rect 31125 27421 31159 27455
rect 31309 27421 31343 27455
rect 31769 27421 31803 27455
rect 31953 27421 31987 27455
rect 33149 27421 33183 27455
rect 33425 27421 33459 27455
rect 34989 27421 35023 27455
rect 35449 27421 35483 27455
rect 37381 27421 37415 27455
rect 37565 27421 37599 27455
rect 41337 27421 41371 27455
rect 42257 27421 42291 27455
rect 42349 27421 42383 27455
rect 42625 27421 42659 27455
rect 44281 27421 44315 27455
rect 9873 27353 9907 27387
rect 13093 27353 13127 27387
rect 15761 27353 15795 27387
rect 15945 27353 15979 27387
rect 16129 27353 16163 27387
rect 17049 27353 17083 27387
rect 17233 27353 17267 27387
rect 21925 27353 21959 27387
rect 24593 27353 24627 27387
rect 24777 27353 24811 27387
rect 29561 27353 29595 27387
rect 30941 27353 30975 27387
rect 34713 27353 34747 27387
rect 35725 27353 35759 27387
rect 40110 27353 40144 27387
rect 6193 27285 6227 27319
rect 20269 27285 20303 27319
rect 24409 27285 24443 27319
rect 30021 27285 30055 27319
rect 32137 27285 32171 27319
rect 32965 27285 32999 27319
rect 37197 27285 37231 27319
rect 41245 27285 41279 27319
rect 44465 27285 44499 27319
rect 13093 27081 13127 27115
rect 19717 27081 19751 27115
rect 22017 27081 22051 27115
rect 25237 27081 25271 27115
rect 26709 27081 26743 27115
rect 27445 27081 27479 27115
rect 35357 27081 35391 27115
rect 37749 27081 37783 27115
rect 39589 27081 39623 27115
rect 43177 27081 43211 27115
rect 20913 27013 20947 27047
rect 25329 27013 25363 27047
rect 26985 27013 27019 27047
rect 28549 27013 28583 27047
rect 42441 27013 42475 27047
rect 8033 26945 8067 26979
rect 8217 26945 8251 26979
rect 13260 26945 13294 26979
rect 13369 26945 13403 26979
rect 13553 26945 13587 26979
rect 15393 26945 15427 26979
rect 15577 26945 15611 26979
rect 19349 26945 19383 26979
rect 19533 26945 19567 26979
rect 20637 26945 20671 26979
rect 22201 26945 22235 26979
rect 22477 26945 22511 26979
rect 24777 26945 24811 26979
rect 25053 26945 25087 26979
rect 25605 26945 25639 26979
rect 26341 26945 26375 26979
rect 26525 26945 26559 26979
rect 27169 26945 27203 26979
rect 27261 26945 27295 26979
rect 28825 26945 28859 26979
rect 32137 26945 32171 26979
rect 32413 26945 32447 26979
rect 34437 26945 34471 26979
rect 34713 26945 34747 26979
rect 34989 26945 35023 26979
rect 35173 26945 35207 26979
rect 37289 26945 37323 26979
rect 37565 26945 37599 26979
rect 39773 26945 39807 26979
rect 39865 26945 39899 26979
rect 40049 26945 40083 26979
rect 40233 26945 40267 26979
rect 40509 26945 40543 26979
rect 40785 26945 40819 26979
rect 40969 26945 41003 26979
rect 41059 26945 41093 26979
rect 41521 26945 41555 26979
rect 44281 26945 44315 26979
rect 8401 26877 8435 26911
rect 20821 26877 20855 26911
rect 22385 26877 22419 26911
rect 24961 26877 24995 26911
rect 25513 26877 25547 26911
rect 28641 26877 28675 26911
rect 32229 26877 32263 26911
rect 34529 26877 34563 26911
rect 37381 26877 37415 26911
rect 39957 26877 39991 26911
rect 40601 26877 40635 26911
rect 40693 26877 40727 26911
rect 41245 26877 41279 26911
rect 41337 26877 41371 26911
rect 42993 26877 43027 26911
rect 43821 26877 43855 26911
rect 26157 26809 26191 26843
rect 28365 26809 28399 26843
rect 29009 26809 29043 26843
rect 34897 26809 34931 26843
rect 41429 26809 41463 26843
rect 13553 26741 13587 26775
rect 15761 26741 15795 26775
rect 19349 26741 19383 26775
rect 20453 26741 20487 26775
rect 20913 26741 20947 26775
rect 22477 26741 22511 26775
rect 25053 26741 25087 26775
rect 25605 26741 25639 26775
rect 25789 26741 25823 26775
rect 27261 26741 27295 26775
rect 28549 26741 28583 26775
rect 32137 26741 32171 26775
rect 32597 26741 32631 26775
rect 34437 26741 34471 26775
rect 35173 26741 35207 26775
rect 37289 26741 37323 26775
rect 40325 26741 40359 26775
rect 41705 26741 41739 26775
rect 44465 26741 44499 26775
rect 10793 26537 10827 26571
rect 10977 26537 11011 26571
rect 11161 26537 11195 26571
rect 12173 26537 12207 26571
rect 12633 26537 12667 26571
rect 14841 26537 14875 26571
rect 15485 26537 15519 26571
rect 15669 26537 15703 26571
rect 17049 26537 17083 26571
rect 18153 26537 18187 26571
rect 18889 26537 18923 26571
rect 20453 26537 20487 26571
rect 20913 26537 20947 26571
rect 22017 26537 22051 26571
rect 22201 26537 22235 26571
rect 25329 26537 25363 26571
rect 26525 26537 26559 26571
rect 29837 26537 29871 26571
rect 31585 26537 31619 26571
rect 32045 26537 32079 26571
rect 33149 26537 33183 26571
rect 33425 26537 33459 26571
rect 37197 26537 37231 26571
rect 42073 26537 42107 26571
rect 43545 26537 43579 26571
rect 10314 26469 10348 26503
rect 10425 26469 10459 26503
rect 15117 26469 15151 26503
rect 17325 26469 17359 26503
rect 18429 26469 18463 26503
rect 26341 26469 26375 26503
rect 37657 26469 37691 26503
rect 44465 26469 44499 26503
rect 10517 26401 10551 26435
rect 11345 26401 11379 26435
rect 12357 26401 12391 26435
rect 14749 26401 14783 26435
rect 15301 26401 15335 26435
rect 17049 26401 17083 26435
rect 17969 26401 18003 26435
rect 18797 26401 18831 26435
rect 21833 26401 21867 26435
rect 29653 26401 29687 26435
rect 31493 26401 31527 26435
rect 31769 26401 31803 26435
rect 40693 26401 40727 26435
rect 8033 26333 8067 26367
rect 8217 26333 8251 26367
rect 11161 26333 11195 26367
rect 11529 26333 11563 26367
rect 12449 26333 12483 26367
rect 14933 26333 14967 26367
rect 15209 26333 15243 26367
rect 15485 26333 15519 26367
rect 16957 26333 16991 26367
rect 18153 26333 18187 26367
rect 18613 26333 18647 26367
rect 20453 26333 20487 26367
rect 20637 26333 20671 26367
rect 20729 26333 20763 26367
rect 22017 26333 22051 26367
rect 25513 26333 25547 26367
rect 25697 26333 25731 26367
rect 26525 26333 26559 26367
rect 26709 26333 26743 26367
rect 29837 26333 29871 26367
rect 31125 26333 31159 26367
rect 31309 26333 31343 26367
rect 31861 26333 31895 26367
rect 33057 26333 33091 26367
rect 33241 26333 33275 26367
rect 37381 26333 37415 26367
rect 37473 26333 37507 26367
rect 40949 26333 40983 26367
rect 42165 26333 42199 26367
rect 42421 26333 42455 26367
rect 44281 26333 44315 26367
rect 7849 26265 7883 26299
rect 10149 26265 10183 26299
rect 11437 26265 11471 26299
rect 11713 26265 11747 26299
rect 11897 26265 11931 26299
rect 12173 26265 12207 26299
rect 14657 26265 14691 26299
rect 17877 26265 17911 26299
rect 18889 26265 18923 26299
rect 21741 26265 21775 26299
rect 29561 26265 29595 26299
rect 31585 26265 31619 26299
rect 37197 26265 37231 26299
rect 18337 26197 18371 26231
rect 30021 26197 30055 26231
rect 8217 25993 8251 26027
rect 9413 25993 9447 26027
rect 12449 25993 12483 26027
rect 16497 25993 16531 26027
rect 21833 25993 21867 26027
rect 24961 25993 24995 26027
rect 34805 25993 34839 26027
rect 5089 25925 5123 25959
rect 8953 25925 8987 25959
rect 10517 25925 10551 25959
rect 23213 25925 23247 25959
rect 23765 25925 23799 25959
rect 24501 25925 24535 25959
rect 28457 25925 28491 25959
rect 38945 25925 38979 25959
rect 39129 25925 39163 25959
rect 5273 25857 5307 25891
rect 5457 25857 5491 25891
rect 7757 25857 7791 25891
rect 8033 25857 8067 25891
rect 9229 25857 9263 25891
rect 10149 25857 10183 25891
rect 10333 25857 10367 25891
rect 10609 25857 10643 25891
rect 10885 25857 10919 25891
rect 11989 25857 12023 25891
rect 12265 25857 12299 25891
rect 12909 25857 12943 25891
rect 14749 25857 14783 25891
rect 14933 25857 14967 25891
rect 16129 25857 16163 25891
rect 16313 25857 16347 25891
rect 22201 25857 22235 25891
rect 22845 25857 22879 25891
rect 23029 25857 23063 25891
rect 23489 25857 23523 25891
rect 23581 25857 23615 25891
rect 23857 25857 23891 25891
rect 24133 25857 24167 25891
rect 24777 25857 24811 25891
rect 26433 25857 26467 25891
rect 26617 25857 26651 25891
rect 26801 25857 26835 25891
rect 28641 25857 28675 25891
rect 28733 25857 28767 25891
rect 32873 25857 32907 25891
rect 33793 25857 33827 25891
rect 34437 25857 34471 25891
rect 35357 25857 35391 25891
rect 37289 25857 37323 25891
rect 37473 25857 37507 25891
rect 38393 25857 38427 25891
rect 38669 25857 38703 25891
rect 39405 25857 39439 25891
rect 40509 25857 40543 25891
rect 40765 25857 40799 25891
rect 7941 25789 7975 25823
rect 9045 25789 9079 25823
rect 10701 25789 10735 25823
rect 12081 25789 12115 25823
rect 13001 25789 13035 25823
rect 22109 25789 22143 25823
rect 24041 25789 24075 25823
rect 24593 25789 24627 25823
rect 32965 25789 32999 25823
rect 33885 25789 33919 25823
rect 34529 25789 34563 25823
rect 35449 25789 35483 25823
rect 38485 25789 38519 25823
rect 39221 25789 39255 25823
rect 43085 25789 43119 25823
rect 11069 25721 11103 25755
rect 23305 25721 23339 25755
rect 24317 25721 24351 25755
rect 37657 25721 37691 25755
rect 38853 25721 38887 25755
rect 42441 25721 42475 25755
rect 8033 25653 8067 25687
rect 9229 25653 9263 25687
rect 10609 25653 10643 25687
rect 11989 25653 12023 25687
rect 13093 25653 13127 25687
rect 13277 25653 13311 25687
rect 15025 25653 15059 25687
rect 22201 25653 22235 25687
rect 23673 25653 23707 25687
rect 23857 25653 23891 25687
rect 24501 25653 24535 25687
rect 28457 25653 28491 25687
rect 28917 25653 28951 25687
rect 32873 25653 32907 25687
rect 33241 25653 33275 25687
rect 33793 25653 33827 25687
rect 34161 25653 34195 25687
rect 34437 25653 34471 25687
rect 35357 25653 35391 25687
rect 35725 25653 35759 25687
rect 37749 25653 37783 25687
rect 38393 25653 38427 25687
rect 39129 25653 39163 25687
rect 39589 25653 39623 25687
rect 41889 25653 41923 25687
rect 5273 25449 5307 25483
rect 5733 25449 5767 25483
rect 10241 25449 10275 25483
rect 19533 25449 19567 25483
rect 19717 25449 19751 25483
rect 20361 25449 20395 25483
rect 20821 25449 20855 25483
rect 23581 25449 23615 25483
rect 23765 25449 23799 25483
rect 25053 25449 25087 25483
rect 25513 25449 25547 25483
rect 28733 25449 28767 25483
rect 29837 25449 29871 25483
rect 30665 25449 30699 25483
rect 31033 25449 31067 25483
rect 31585 25449 31619 25483
rect 32045 25449 32079 25483
rect 34805 25449 34839 25483
rect 35173 25449 35207 25483
rect 36553 25449 36587 25483
rect 36921 25449 36955 25483
rect 40417 25449 40451 25483
rect 28641 25381 28675 25415
rect 32873 25381 32907 25415
rect 40693 25381 40727 25415
rect 5641 25313 5675 25347
rect 19349 25313 19383 25347
rect 20453 25313 20487 25347
rect 23397 25313 23431 25347
rect 25145 25313 25179 25347
rect 26249 25313 26283 25347
rect 30757 25313 30791 25347
rect 31769 25313 31803 25347
rect 40785 25313 40819 25347
rect 40877 25313 40911 25347
rect 43729 25313 43763 25347
rect 5457 25245 5491 25279
rect 10425 25245 10459 25279
rect 10609 25245 10643 25279
rect 19533 25245 19567 25279
rect 20637 25245 20671 25279
rect 23581 25245 23615 25279
rect 25329 25245 25363 25279
rect 26065 25245 26099 25279
rect 28273 25245 28307 25279
rect 29561 25245 29595 25279
rect 29745 25245 29779 25279
rect 29837 25245 29871 25279
rect 30665 25245 30699 25279
rect 31861 25245 31895 25279
rect 34805 25245 34839 25279
rect 34989 25245 35023 25279
rect 36461 25245 36495 25279
rect 36645 25245 36679 25279
rect 36737 25245 36771 25279
rect 40601 25245 40635 25279
rect 41061 25245 41095 25279
rect 41613 25245 41647 25279
rect 44005 25245 44039 25279
rect 44281 25245 44315 25279
rect 5733 25177 5767 25211
rect 16129 25177 16163 25211
rect 16313 25177 16347 25211
rect 19257 25177 19291 25211
rect 20361 25177 20395 25211
rect 23305 25177 23339 25211
rect 25053 25177 25087 25211
rect 25881 25177 25915 25211
rect 28457 25177 28491 25211
rect 28917 25177 28951 25211
rect 29101 25177 29135 25211
rect 31585 25177 31619 25211
rect 34161 25177 34195 25211
rect 41880 25177 41914 25211
rect 43821 25177 43855 25211
rect 16497 25109 16531 25143
rect 24961 25109 24995 25143
rect 30021 25109 30055 25143
rect 42993 25109 43027 25143
rect 43085 25109 43119 25143
rect 44465 25109 44499 25143
rect 5825 24905 5859 24939
rect 20637 24905 20671 24939
rect 23029 24905 23063 24939
rect 32137 24905 32171 24939
rect 43821 24905 43855 24939
rect 6009 24769 6043 24803
rect 6193 24769 6227 24803
rect 8401 24769 8435 24803
rect 10057 24769 10091 24803
rect 10333 24769 10367 24803
rect 11897 24769 11931 24803
rect 12173 24769 12207 24803
rect 14013 24769 14047 24803
rect 14197 24769 14231 24803
rect 17325 24769 17359 24803
rect 17601 24769 17635 24803
rect 17877 24769 17911 24803
rect 19625 24769 19659 24803
rect 19717 24769 19751 24803
rect 20269 24769 20303 24803
rect 20453 24769 20487 24803
rect 20729 24769 20763 24803
rect 20913 24769 20947 24803
rect 22569 24769 22603 24803
rect 22845 24769 22879 24803
rect 26433 24769 26467 24803
rect 32321 24769 32355 24803
rect 32505 24769 32539 24803
rect 32770 24769 32804 24803
rect 33057 24769 33091 24803
rect 38577 24769 38611 24803
rect 38853 24769 38887 24803
rect 41705 24769 41739 24803
rect 41981 24769 42015 24803
rect 42073 24769 42107 24803
rect 42257 24769 42291 24803
rect 42697 24769 42731 24803
rect 44281 24769 44315 24803
rect 8548 24701 8582 24735
rect 8769 24701 8803 24735
rect 10149 24701 10183 24735
rect 11989 24701 12023 24735
rect 17417 24701 17451 24735
rect 17969 24701 18003 24735
rect 22753 24701 22787 24735
rect 26341 24701 26375 24735
rect 32873 24701 32907 24735
rect 38761 24701 38795 24735
rect 42441 24701 42475 24735
rect 10517 24633 10551 24667
rect 17785 24633 17819 24667
rect 18245 24633 18279 24667
rect 19993 24633 20027 24667
rect 26065 24633 26099 24667
rect 8677 24565 8711 24599
rect 9045 24565 9079 24599
rect 10057 24565 10091 24599
rect 11713 24565 11747 24599
rect 11897 24565 11931 24599
rect 14381 24565 14415 24599
rect 17325 24565 17359 24599
rect 17877 24565 17911 24599
rect 19809 24565 19843 24599
rect 21097 24565 21131 24599
rect 22753 24565 22787 24599
rect 26433 24565 26467 24599
rect 32965 24565 32999 24599
rect 33241 24565 33275 24599
rect 38669 24565 38703 24599
rect 39037 24565 39071 24599
rect 41797 24565 41831 24599
rect 44465 24565 44499 24599
rect 7849 24361 7883 24395
rect 9965 24361 9999 24395
rect 10793 24361 10827 24395
rect 12817 24361 12851 24395
rect 13369 24361 13403 24395
rect 15117 24361 15151 24395
rect 15393 24361 15427 24395
rect 16313 24361 16347 24395
rect 16497 24361 16531 24395
rect 16957 24361 16991 24395
rect 17233 24361 17267 24395
rect 17877 24361 17911 24395
rect 18245 24361 18279 24395
rect 22845 24361 22879 24395
rect 23765 24361 23799 24395
rect 27997 24361 28031 24395
rect 28273 24361 28307 24395
rect 29745 24361 29779 24395
rect 31033 24361 31067 24395
rect 31585 24361 31619 24395
rect 31769 24361 31803 24395
rect 34069 24361 34103 24395
rect 34713 24361 34747 24395
rect 35265 24361 35299 24395
rect 35725 24361 35759 24395
rect 36277 24361 36311 24395
rect 18153 24293 18187 24327
rect 23029 24293 23063 24327
rect 23305 24293 23339 24327
rect 31493 24293 31527 24327
rect 35173 24293 35207 24327
rect 7757 24225 7791 24259
rect 10057 24225 10091 24259
rect 10701 24225 10735 24259
rect 13553 24225 13587 24259
rect 16129 24225 16163 24259
rect 16865 24225 16899 24259
rect 17785 24225 17819 24259
rect 22661 24225 22695 24259
rect 23673 24225 23707 24259
rect 31217 24225 31251 24259
rect 31861 24225 31895 24259
rect 34161 24225 34195 24259
rect 34897 24225 34931 24259
rect 36369 24225 36403 24259
rect 42993 24225 43027 24259
rect 7665 24157 7699 24191
rect 10241 24157 10275 24191
rect 10786 24157 10820 24191
rect 12725 24157 12759 24191
rect 12909 24157 12943 24191
rect 13645 24157 13679 24191
rect 15117 24157 15151 24191
rect 15209 24157 15243 24191
rect 16313 24157 16347 24191
rect 17049 24157 17083 24191
rect 17969 24157 18003 24191
rect 22845 24157 22879 24191
rect 23489 24157 23523 24191
rect 27997 24157 28031 24191
rect 28089 24157 28123 24191
rect 28365 24157 28399 24191
rect 28549 24157 28583 24191
rect 29561 24157 29595 24191
rect 29745 24157 29779 24191
rect 31309 24157 31343 24191
rect 31953 24157 31987 24191
rect 34345 24157 34379 24191
rect 34989 24157 35023 24191
rect 35265 24157 35299 24191
rect 35449 24157 35483 24191
rect 35541 24157 35575 24191
rect 35817 24157 35851 24191
rect 36001 24157 36035 24191
rect 36277 24157 36311 24191
rect 40601 24157 40635 24191
rect 44281 24157 44315 24191
rect 9965 24089 9999 24123
rect 10517 24089 10551 24123
rect 13369 24089 13403 24123
rect 14381 24089 14415 24123
rect 14565 24089 14599 24123
rect 14749 24089 14783 24123
rect 14933 24089 14967 24123
rect 16037 24089 16071 24123
rect 16773 24089 16807 24123
rect 17693 24089 17727 24123
rect 18429 24089 18463 24123
rect 18613 24089 18647 24123
rect 22569 24089 22603 24123
rect 23765 24089 23799 24123
rect 27813 24089 27847 24123
rect 28733 24089 28767 24123
rect 31033 24089 31067 24123
rect 34069 24089 34103 24123
rect 34713 24089 34747 24123
rect 40868 24089 40902 24123
rect 8033 24021 8067 24055
rect 10425 24021 10459 24055
rect 10977 24021 11011 24055
rect 13093 24021 13127 24055
rect 13829 24021 13863 24055
rect 29929 24021 29963 24055
rect 34529 24021 34563 24055
rect 36185 24021 36219 24055
rect 36645 24021 36679 24055
rect 41981 24021 42015 24055
rect 43637 24021 43671 24055
rect 44465 24021 44499 24055
rect 7389 23817 7423 23851
rect 7481 23817 7515 23851
rect 10425 23817 10459 23851
rect 15669 23817 15703 23851
rect 20637 23817 20671 23851
rect 26249 23817 26283 23851
rect 30205 23817 30239 23851
rect 32781 23817 32815 23851
rect 34989 23817 35023 23851
rect 41797 23817 41831 23851
rect 43177 23817 43211 23851
rect 6929 23749 6963 23783
rect 9505 23749 9539 23783
rect 20453 23749 20487 23783
rect 23581 23749 23615 23783
rect 24869 23749 24903 23783
rect 25053 23749 25087 23783
rect 26341 23749 26375 23783
rect 26525 23749 26559 23783
rect 34437 23749 34471 23783
rect 40325 23749 40359 23783
rect 4169 23681 4203 23715
rect 4353 23681 4387 23715
rect 4445 23681 4479 23715
rect 4542 23681 4576 23715
rect 7205 23681 7239 23715
rect 7665 23681 7699 23715
rect 7941 23681 7975 23715
rect 9229 23681 9263 23715
rect 9413 23681 9447 23715
rect 9597 23681 9631 23715
rect 9873 23681 9907 23715
rect 10057 23681 10091 23715
rect 10149 23681 10183 23715
rect 10241 23681 10275 23715
rect 13461 23681 13495 23715
rect 13645 23681 13679 23715
rect 13829 23681 13863 23715
rect 15209 23681 15243 23715
rect 15485 23681 15519 23715
rect 20269 23681 20303 23715
rect 22845 23681 22879 23715
rect 23397 23681 23431 23715
rect 25789 23681 25823 23715
rect 25973 23681 26007 23715
rect 26065 23681 26099 23715
rect 27261 23681 27295 23715
rect 27445 23681 27479 23715
rect 27997 23681 28031 23715
rect 29745 23681 29779 23715
rect 30021 23681 30055 23715
rect 30849 23681 30883 23715
rect 31493 23681 31527 23715
rect 31769 23681 31803 23715
rect 32321 23681 32355 23715
rect 32597 23681 32631 23715
rect 34253 23681 34287 23715
rect 34529 23681 34563 23715
rect 34713 23681 34747 23715
rect 34805 23681 34839 23715
rect 36277 23681 36311 23715
rect 36461 23681 36495 23715
rect 36737 23681 36771 23715
rect 38945 23681 38979 23715
rect 39129 23681 39163 23715
rect 39405 23681 39439 23715
rect 40509 23681 40543 23715
rect 43361 23681 43395 23715
rect 43453 23681 43487 23715
rect 43729 23681 43763 23715
rect 44281 23681 44315 23715
rect 7113 23613 7147 23647
rect 7757 23613 7791 23647
rect 15301 23613 15335 23647
rect 22937 23613 22971 23647
rect 28089 23613 28123 23647
rect 29837 23613 29871 23647
rect 30941 23613 30975 23647
rect 31585 23613 31619 23647
rect 32413 23613 32447 23647
rect 36553 23613 36587 23647
rect 39221 23613 39255 23647
rect 42993 23613 43027 23647
rect 43637 23613 43671 23647
rect 9781 23545 9815 23579
rect 23213 23545 23247 23579
rect 25237 23545 25271 23579
rect 26709 23545 26743 23579
rect 31217 23545 31251 23579
rect 4721 23477 4755 23511
rect 7205 23477 7239 23511
rect 7849 23477 7883 23511
rect 15209 23477 15243 23511
rect 22845 23477 22879 23511
rect 23673 23477 23707 23511
rect 25789 23477 25823 23511
rect 27077 23477 27111 23511
rect 27629 23477 27663 23511
rect 27905 23477 27939 23511
rect 28181 23477 28215 23511
rect 28365 23477 28399 23511
rect 29837 23477 29871 23511
rect 30941 23477 30975 23511
rect 31585 23477 31619 23511
rect 31953 23477 31987 23511
rect 32597 23477 32631 23511
rect 34069 23477 34103 23511
rect 34529 23477 34563 23511
rect 36461 23477 36495 23511
rect 36921 23477 36955 23511
rect 39129 23477 39163 23511
rect 39589 23477 39623 23511
rect 42441 23477 42475 23511
rect 44465 23477 44499 23511
rect 3157 23273 3191 23307
rect 5733 23273 5767 23307
rect 10885 23273 10919 23307
rect 12817 23273 12851 23307
rect 14657 23273 14691 23307
rect 15025 23273 15059 23307
rect 15209 23273 15243 23307
rect 18613 23273 18647 23307
rect 23581 23273 23615 23307
rect 23949 23273 23983 23307
rect 29745 23273 29779 23307
rect 33701 23273 33735 23307
rect 34161 23273 34195 23307
rect 34713 23273 34747 23307
rect 37105 23273 37139 23307
rect 37381 23273 37415 23307
rect 38209 23273 38243 23307
rect 38669 23273 38703 23307
rect 39865 23273 39899 23307
rect 5089 23205 5123 23239
rect 7849 23205 7883 23239
rect 18797 23205 18831 23239
rect 27353 23205 27387 23239
rect 29561 23205 29595 23239
rect 35173 23205 35207 23239
rect 40233 23205 40267 23239
rect 40601 23205 40635 23239
rect 41061 23205 41095 23239
rect 41337 23205 41371 23239
rect 20453 23137 20487 23171
rect 29929 23137 29963 23171
rect 33793 23137 33827 23171
rect 34805 23137 34839 23171
rect 39957 23137 39991 23171
rect 40693 23137 40727 23171
rect 40785 23137 40819 23171
rect 41429 23137 41463 23171
rect 41521 23137 41555 23171
rect 2605 23069 2639 23103
rect 2789 23069 2823 23103
rect 3025 23069 3059 23103
rect 4445 23069 4479 23103
rect 4629 23069 4663 23103
rect 4905 23069 4939 23103
rect 5181 23069 5215 23103
rect 5549 23069 5583 23103
rect 7297 23069 7331 23103
rect 7573 23069 7607 23103
rect 7717 23069 7751 23103
rect 9505 23069 9539 23103
rect 9689 23069 9723 23103
rect 10057 23069 10091 23103
rect 10333 23069 10367 23103
rect 10609 23069 10643 23103
rect 10706 23069 10740 23103
rect 12265 23069 12299 23103
rect 12633 23069 12667 23103
rect 14105 23069 14139 23103
rect 14289 23069 14323 23103
rect 14478 23069 14512 23103
rect 14841 23069 14875 23103
rect 15025 23069 15059 23103
rect 18429 23069 18463 23103
rect 18521 23069 18555 23103
rect 20085 23069 20119 23103
rect 20729 23069 20763 23103
rect 23581 23069 23615 23103
rect 23673 23069 23707 23103
rect 26433 23069 26467 23103
rect 29745 23069 29779 23103
rect 32597 23069 32631 23103
rect 33701 23069 33735 23103
rect 33977 23069 34011 23103
rect 34989 23069 35023 23103
rect 37013 23069 37047 23103
rect 37197 23069 37231 23103
rect 37381 23069 37415 23103
rect 37473 23069 37507 23103
rect 38393 23069 38427 23103
rect 38485 23069 38519 23103
rect 39865 23069 39899 23103
rect 40509 23069 40543 23103
rect 40969 23069 41003 23103
rect 41245 23069 41279 23103
rect 41705 23069 41739 23103
rect 42441 23069 42475 23103
rect 2881 23001 2915 23035
rect 5365 23001 5399 23035
rect 5457 23001 5491 23035
rect 7481 23001 7515 23035
rect 10517 23001 10551 23035
rect 12449 23001 12483 23035
rect 12541 23001 12575 23035
rect 14381 23001 14415 23035
rect 20269 23001 20303 23035
rect 20545 23001 20579 23035
rect 26065 23001 26099 23035
rect 26249 23001 26283 23035
rect 27537 23001 27571 23035
rect 27721 23001 27755 23035
rect 30021 23001 30055 23035
rect 32781 23001 32815 23035
rect 32965 23001 32999 23035
rect 34713 23001 34747 23035
rect 38209 23001 38243 23035
rect 9965 22933 9999 22967
rect 20913 22933 20947 22967
rect 36829 22933 36863 22967
rect 37749 22933 37783 22967
rect 40325 22933 40359 22967
rect 41797 22933 41831 22967
rect 8953 22729 8987 22763
rect 13369 22729 13403 22763
rect 14473 22729 14507 22763
rect 21097 22729 21131 22763
rect 26709 22729 26743 22763
rect 29469 22729 29503 22763
rect 41705 22729 41739 22763
rect 4997 22661 5031 22695
rect 5641 22661 5675 22695
rect 5733 22661 5767 22695
rect 9413 22661 9447 22695
rect 9505 22661 9539 22695
rect 10333 22661 10367 22695
rect 14013 22661 14047 22695
rect 16313 22661 16347 22695
rect 21189 22661 21223 22695
rect 21925 22661 21959 22695
rect 24501 22661 24535 22695
rect 29009 22661 29043 22695
rect 4721 22593 4755 22627
rect 4905 22593 4939 22627
rect 5135 22593 5169 22627
rect 5457 22593 5491 22627
rect 5825 22593 5859 22627
rect 8493 22593 8527 22627
rect 8769 22593 8803 22627
rect 9229 22593 9263 22627
rect 9602 22593 9636 22627
rect 10057 22593 10091 22627
rect 10241 22593 10275 22627
rect 10430 22593 10464 22627
rect 11805 22593 11839 22627
rect 11989 22593 12023 22627
rect 12265 22593 12299 22627
rect 12725 22593 12759 22627
rect 14289 22593 14323 22627
rect 16497 22593 16531 22627
rect 20637 22593 20671 22627
rect 20821 22593 20855 22627
rect 20913 22593 20947 22627
rect 21373 22593 21407 22627
rect 21465 22593 21499 22627
rect 22201 22593 22235 22627
rect 24317 22593 24351 22627
rect 26249 22593 26283 22627
rect 26525 22593 26559 22627
rect 29285 22593 29319 22627
rect 31033 22593 31067 22627
rect 31217 22593 31251 22627
rect 31769 22593 31803 22627
rect 31953 22593 31987 22627
rect 40325 22593 40359 22627
rect 40581 22593 40615 22627
rect 44281 22593 44315 22627
rect 8677 22525 8711 22559
rect 13093 22525 13127 22559
rect 14197 22525 14231 22559
rect 22017 22525 22051 22559
rect 26341 22525 26375 22559
rect 29101 22525 29135 22559
rect 6009 22457 6043 22491
rect 13001 22457 13035 22491
rect 21649 22457 21683 22491
rect 44465 22457 44499 22491
rect 5273 22389 5307 22423
rect 8677 22389 8711 22423
rect 9781 22389 9815 22423
rect 10609 22389 10643 22423
rect 12449 22389 12483 22423
rect 12890 22389 12924 22423
rect 14105 22389 14139 22423
rect 16221 22389 16255 22423
rect 20821 22389 20855 22423
rect 21465 22389 21499 22423
rect 22201 22389 22235 22423
rect 22385 22389 22419 22423
rect 24685 22389 24719 22423
rect 26525 22389 26559 22423
rect 29193 22389 29227 22423
rect 31033 22389 31067 22423
rect 31401 22389 31435 22423
rect 31585 22389 31619 22423
rect 31769 22389 31803 22423
rect 5365 22185 5399 22219
rect 7297 22185 7331 22219
rect 14933 22185 14967 22219
rect 15209 22185 15243 22219
rect 15853 22185 15887 22219
rect 17785 22185 17819 22219
rect 19349 22185 19383 22219
rect 25145 22185 25179 22219
rect 25697 22185 25731 22219
rect 26065 22185 26099 22219
rect 26801 22185 26835 22219
rect 27813 22185 27847 22219
rect 28365 22185 28399 22219
rect 32689 22185 32723 22219
rect 33149 22185 33183 22219
rect 33241 22185 33275 22219
rect 34713 22185 34747 22219
rect 35817 22185 35851 22219
rect 12173 22117 12207 22151
rect 12817 22117 12851 22151
rect 7205 22049 7239 22083
rect 7941 22049 7975 22083
rect 15853 22049 15887 22083
rect 18705 22049 18739 22083
rect 19441 22049 19475 22083
rect 24777 22049 24811 22083
rect 25605 22049 25639 22083
rect 26157 22049 26191 22083
rect 27997 22049 28031 22083
rect 35633 22049 35667 22083
rect 41521 22049 41555 22083
rect 5089 21981 5123 22015
rect 5273 21981 5307 22015
rect 5365 21981 5399 22015
rect 7113 21981 7147 22015
rect 7757 21981 7791 22015
rect 11621 21981 11655 22015
rect 11989 21981 12023 22015
rect 12265 21981 12299 22015
rect 12449 21981 12483 22015
rect 12633 21981 12667 22015
rect 14933 21981 14967 22015
rect 15025 21981 15059 22015
rect 15945 21981 15979 22015
rect 16773 21981 16807 22015
rect 17785 21981 17819 22015
rect 17877 21981 17911 22015
rect 19257 21981 19291 22015
rect 19533 21981 19567 22015
rect 25053 21981 25087 22015
rect 25145 21981 25179 22015
rect 25697 21981 25731 22015
rect 26341 21981 26375 22015
rect 26617 21981 26651 22015
rect 26801 21981 26835 22015
rect 28089 21981 28123 22015
rect 28365 21981 28399 22015
rect 28457 21981 28491 22015
rect 32873 21981 32907 22015
rect 32965 21981 32999 22015
rect 33241 21981 33275 22015
rect 33333 21981 33367 22015
rect 34897 21981 34931 22015
rect 34989 21981 35023 22015
rect 35817 21981 35851 22015
rect 40325 21981 40359 22015
rect 40417 21981 40451 22015
rect 40509 21981 40543 22015
rect 40601 21981 40635 22015
rect 40785 21981 40819 22015
rect 42993 21981 43027 22015
rect 43545 21981 43579 22015
rect 44281 21981 44315 22015
rect 6653 21913 6687 21947
rect 6837 21913 6871 21947
rect 7021 21913 7055 21947
rect 7573 21913 7607 21947
rect 11805 21913 11839 21947
rect 11897 21913 11931 21947
rect 12541 21913 12575 21947
rect 14749 21913 14783 21947
rect 15669 21913 15703 21947
rect 16589 21913 16623 21947
rect 16957 21913 16991 21947
rect 18337 21913 18371 21947
rect 18521 21913 18555 21947
rect 24409 21913 24443 21947
rect 24593 21913 24627 21947
rect 24869 21913 24903 21947
rect 25421 21913 25455 21947
rect 26065 21913 26099 21947
rect 27813 21913 27847 21947
rect 32689 21913 32723 21947
rect 34713 21913 34747 21947
rect 35541 21913 35575 21947
rect 41788 21913 41822 21947
rect 5549 21845 5583 21879
rect 7481 21845 7515 21879
rect 16129 21845 16163 21879
rect 18153 21845 18187 21879
rect 19717 21845 19751 21879
rect 25329 21845 25363 21879
rect 25881 21845 25915 21879
rect 26525 21845 26559 21879
rect 26985 21845 27019 21879
rect 28273 21845 28307 21879
rect 28733 21845 28767 21879
rect 33609 21845 33643 21879
rect 35173 21845 35207 21879
rect 36001 21845 36035 21879
rect 40141 21845 40175 21879
rect 42901 21845 42935 21879
rect 44465 21845 44499 21879
rect 6193 21641 6227 21675
rect 9873 21641 9907 21675
rect 12909 21641 12943 21675
rect 20821 21641 20855 21675
rect 33241 21641 33275 21675
rect 34713 21641 34747 21675
rect 38945 21641 38979 21675
rect 41705 21641 41739 21675
rect 2881 21573 2915 21607
rect 10241 21573 10275 21607
rect 12633 21573 12667 21607
rect 23949 21573 23983 21607
rect 24501 21573 24535 21607
rect 37289 21573 37323 21607
rect 37933 21573 37967 21607
rect 38485 21573 38519 21607
rect 40570 21573 40604 21607
rect 2697 21505 2731 21539
rect 2973 21505 3007 21539
rect 3065 21505 3099 21539
rect 5641 21505 5675 21539
rect 5825 21505 5859 21539
rect 5917 21505 5951 21539
rect 6009 21505 6043 21539
rect 9689 21505 9723 21539
rect 9965 21505 9999 21539
rect 10149 21505 10183 21539
rect 10333 21505 10367 21539
rect 12357 21505 12391 21539
rect 12541 21505 12575 21539
rect 12725 21505 12759 21539
rect 20453 21505 20487 21539
rect 20637 21505 20671 21539
rect 21189 21505 21223 21539
rect 21373 21505 21407 21539
rect 24225 21505 24259 21539
rect 24777 21505 24811 21539
rect 29825 21505 29859 21539
rect 30481 21505 30515 21539
rect 30757 21505 30791 21539
rect 31217 21505 31251 21539
rect 31493 21505 31527 21539
rect 32505 21505 32539 21539
rect 33517 21505 33551 21539
rect 33701 21505 33735 21539
rect 34345 21505 34379 21539
rect 34529 21505 34563 21539
rect 37565 21505 37599 21539
rect 38209 21505 38243 21539
rect 38761 21505 38795 21539
rect 39037 21505 39071 21539
rect 42809 21505 42843 21539
rect 43085 21505 43119 21539
rect 44281 21505 44315 21539
rect 24041 21437 24075 21471
rect 24593 21437 24627 21471
rect 29929 21437 29963 21471
rect 30665 21437 30699 21471
rect 31309 21437 31343 21471
rect 32413 21437 32447 21471
rect 37381 21437 37415 21471
rect 38025 21437 38059 21471
rect 38577 21437 38611 21471
rect 39129 21437 39163 21471
rect 40325 21437 40359 21471
rect 3249 21369 3283 21403
rect 24409 21369 24443 21403
rect 24961 21369 24995 21403
rect 31677 21369 31711 21403
rect 42625 21369 42659 21403
rect 10517 21301 10551 21335
rect 21557 21301 21591 21335
rect 23949 21301 23983 21335
rect 24501 21301 24535 21335
rect 30021 21301 30055 21335
rect 30205 21301 30239 21335
rect 30297 21301 30331 21335
rect 30481 21301 30515 21335
rect 31217 21301 31251 21335
rect 32137 21301 32171 21335
rect 32321 21301 32355 21335
rect 33333 21301 33367 21335
rect 37565 21301 37599 21335
rect 37749 21301 37783 21335
rect 38209 21301 38243 21335
rect 38393 21301 38427 21335
rect 38485 21301 38519 21335
rect 39037 21301 39071 21335
rect 39405 21301 39439 21335
rect 43637 21301 43671 21335
rect 44465 21301 44499 21335
rect 7389 21097 7423 21131
rect 8769 21097 8803 21131
rect 9781 21097 9815 21131
rect 11437 21097 11471 21131
rect 13093 21097 13127 21131
rect 13645 21097 13679 21131
rect 14749 21097 14783 21131
rect 17417 21097 17451 21131
rect 18153 21097 18187 21131
rect 19257 21097 19291 21131
rect 19717 21097 19751 21131
rect 20913 21097 20947 21131
rect 21465 21097 21499 21131
rect 21833 21097 21867 21131
rect 24777 21097 24811 21131
rect 26985 21097 27019 21131
rect 34989 21097 35023 21131
rect 36001 21097 36035 21131
rect 36461 21097 36495 21131
rect 38393 21097 38427 21131
rect 38577 21097 38611 21131
rect 43821 21097 43855 21131
rect 4353 21029 4387 21063
rect 12357 21029 12391 21063
rect 15393 21029 15427 21063
rect 42533 21029 42567 21063
rect 43361 21029 43395 21063
rect 7297 20961 7331 20995
rect 9965 20961 9999 20995
rect 10241 20961 10275 20995
rect 19349 20961 19383 20995
rect 21005 20961 21039 20995
rect 23121 20961 23155 20995
rect 24593 20961 24627 20995
rect 35173 20961 35207 20995
rect 41153 20961 41187 20995
rect 2145 20893 2179 20927
rect 2421 20893 2455 20927
rect 2513 20893 2547 20927
rect 3801 20893 3835 20927
rect 4221 20893 4255 20927
rect 7389 20893 7423 20927
rect 8217 20893 8251 20927
rect 8401 20893 8435 20927
rect 8585 20893 8619 20927
rect 9229 20893 9263 20927
rect 9505 20893 9539 20927
rect 9649 20893 9683 20927
rect 10885 20893 10919 20927
rect 11069 20893 11103 20927
rect 11161 20893 11195 20927
rect 11305 20893 11339 20927
rect 11805 20893 11839 20927
rect 11989 20893 12023 20927
rect 12225 20893 12259 20927
rect 12541 20893 12575 20927
rect 12817 20893 12851 20927
rect 12961 20893 12995 20927
rect 14105 20893 14139 20927
rect 14289 20893 14323 20927
rect 14565 20893 14599 20927
rect 14841 20893 14875 20927
rect 15209 20893 15243 20927
rect 17417 20893 17451 20927
rect 17601 20893 17635 20927
rect 17693 20893 17727 20927
rect 18245 20893 18279 20927
rect 18337 20893 18371 20927
rect 19533 20893 19567 20927
rect 21189 20893 21223 20927
rect 21465 20893 21499 20927
rect 21557 20893 21591 20927
rect 23305 20893 23339 20927
rect 24501 20893 24535 20927
rect 24777 20893 24811 20927
rect 26341 20893 26375 20927
rect 26801 20893 26835 20927
rect 26985 20893 27019 20927
rect 35265 20893 35299 20927
rect 36185 20893 36219 20927
rect 36277 20893 36311 20927
rect 38209 20893 38243 20927
rect 38301 20893 38335 20927
rect 43269 20893 43303 20927
rect 43545 20893 43579 20927
rect 43637 20893 43671 20927
rect 43913 20893 43947 20927
rect 44281 20893 44315 20927
rect 2329 20825 2363 20859
rect 3985 20825 4019 20859
rect 4077 20825 4111 20859
rect 7113 20825 7147 20859
rect 8493 20825 8527 20859
rect 9413 20825 9447 20859
rect 12081 20825 12115 20859
rect 12725 20825 12759 20859
rect 13277 20825 13311 20859
rect 13461 20825 13495 20859
rect 15025 20825 15059 20859
rect 15117 20825 15151 20859
rect 18061 20825 18095 20859
rect 19257 20825 19291 20859
rect 20913 20825 20947 20859
rect 23489 20825 23523 20859
rect 26525 20825 26559 20859
rect 26709 20825 26743 20859
rect 34989 20825 35023 20859
rect 36001 20825 36035 20859
rect 41420 20825 41454 20859
rect 2697 20757 2731 20791
rect 7573 20757 7607 20791
rect 17877 20757 17911 20791
rect 18521 20757 18555 20791
rect 21373 20757 21407 20791
rect 24961 20757 24995 20791
rect 27169 20757 27203 20791
rect 35449 20757 35483 20791
rect 42625 20757 42659 20791
rect 44465 20757 44499 20791
rect 6101 20553 6135 20587
rect 12926 20553 12960 20587
rect 19993 20553 20027 20587
rect 23305 20553 23339 20587
rect 24225 20553 24259 20587
rect 27445 20553 27479 20587
rect 27997 20553 28031 20587
rect 29377 20553 29411 20587
rect 29469 20553 29503 20587
rect 36553 20553 36587 20587
rect 38853 20553 38887 20587
rect 41613 20553 41647 20587
rect 9505 20485 9539 20519
rect 10149 20485 10183 20519
rect 12541 20485 12575 20519
rect 12633 20485 12667 20519
rect 15393 20485 15427 20519
rect 18153 20485 18187 20519
rect 26985 20485 27019 20519
rect 27537 20485 27571 20519
rect 29837 20485 29871 20519
rect 29929 20485 29963 20519
rect 38393 20485 38427 20519
rect 3709 20417 3743 20451
rect 5733 20417 5767 20451
rect 5917 20417 5951 20451
rect 9321 20417 9355 20451
rect 9597 20417 9631 20451
rect 9689 20417 9723 20451
rect 9965 20417 9999 20451
rect 10241 20417 10275 20451
rect 10338 20417 10372 20451
rect 12357 20417 12391 20451
rect 12730 20417 12764 20451
rect 13553 20417 13587 20451
rect 14473 20417 14507 20451
rect 14749 20417 14783 20451
rect 15669 20417 15703 20451
rect 16129 20417 16163 20451
rect 16221 20417 16255 20451
rect 18429 20417 18463 20451
rect 19533 20417 19567 20451
rect 19809 20417 19843 20451
rect 21005 20417 21039 20451
rect 21189 20417 21223 20451
rect 22937 20417 22971 20451
rect 23121 20417 23155 20451
rect 23765 20417 23799 20451
rect 24041 20417 24075 20451
rect 25789 20417 25823 20451
rect 26065 20417 26099 20451
rect 26341 20417 26375 20451
rect 26617 20417 26651 20451
rect 27261 20417 27295 20451
rect 27813 20417 27847 20451
rect 28089 20417 28123 20451
rect 28273 20417 28307 20451
rect 29009 20417 29043 20451
rect 29653 20417 29687 20451
rect 30113 20417 30147 20451
rect 34713 20417 34747 20451
rect 36737 20417 36771 20451
rect 37013 20417 37047 20451
rect 38669 20417 38703 20451
rect 41797 20417 41831 20451
rect 41889 20417 41923 20451
rect 42165 20417 42199 20451
rect 3433 20349 3467 20383
rect 13277 20349 13311 20383
rect 14565 20349 14599 20383
rect 15485 20349 15519 20383
rect 18245 20349 18279 20383
rect 19625 20349 19659 20383
rect 23949 20349 23983 20383
rect 25881 20349 25915 20383
rect 26433 20349 26467 20383
rect 27077 20349 27111 20383
rect 27629 20349 27663 20383
rect 29101 20349 29135 20383
rect 34805 20349 34839 20383
rect 36921 20349 36955 20383
rect 38485 20349 38519 20383
rect 42073 20349 42107 20383
rect 10517 20281 10551 20315
rect 15853 20281 15887 20315
rect 16497 20281 16531 20315
rect 18613 20281 18647 20315
rect 26249 20281 26283 20315
rect 26801 20281 26835 20315
rect 28457 20281 28491 20315
rect 5917 20213 5951 20247
rect 9873 20213 9907 20247
rect 14657 20213 14691 20247
rect 14933 20213 14967 20247
rect 15393 20213 15427 20247
rect 16313 20213 16347 20247
rect 18429 20213 18463 20247
rect 19809 20213 19843 20247
rect 21005 20213 21039 20247
rect 21373 20213 21407 20247
rect 22753 20213 22787 20247
rect 23765 20213 23799 20247
rect 25789 20213 25823 20247
rect 26341 20213 26375 20247
rect 26985 20213 27019 20247
rect 27629 20213 27663 20247
rect 29009 20213 29043 20247
rect 30297 20213 30331 20247
rect 34713 20213 34747 20247
rect 35081 20213 35115 20247
rect 36737 20213 36771 20247
rect 38393 20213 38427 20247
rect 5365 20009 5399 20043
rect 9505 20009 9539 20043
rect 13461 20009 13495 20043
rect 14565 20009 14599 20043
rect 15669 20009 15703 20043
rect 16037 20009 16071 20043
rect 18337 20009 18371 20043
rect 23581 20009 23615 20043
rect 25513 20009 25547 20043
rect 25973 20009 26007 20043
rect 26525 20009 26559 20043
rect 30021 20009 30055 20043
rect 31309 20009 31343 20043
rect 32321 20009 32355 20043
rect 33609 20009 33643 20043
rect 33977 20009 34011 20043
rect 35541 20009 35575 20043
rect 37105 20009 37139 20043
rect 3525 19941 3559 19975
rect 14381 19941 14415 19975
rect 24777 19941 24811 19975
rect 29561 19941 29595 19975
rect 6561 19873 6595 19907
rect 6745 19873 6779 19907
rect 7481 19873 7515 19907
rect 23397 19873 23431 19907
rect 25697 19873 25731 19907
rect 26617 19873 26651 19907
rect 29377 19873 29411 19907
rect 29837 19873 29871 19907
rect 32413 19873 32447 19907
rect 34069 19873 34103 19907
rect 35541 19873 35575 19907
rect 37197 19873 37231 19907
rect 2973 19805 3007 19839
rect 3341 19805 3375 19839
rect 4813 19805 4847 19839
rect 5233 19805 5267 19839
rect 6469 19805 6503 19839
rect 6837 19805 6871 19839
rect 8217 19805 8251 19839
rect 8585 19805 8619 19839
rect 8769 19805 8803 19839
rect 8953 19805 8987 19839
rect 9137 19805 9171 19839
rect 9326 19805 9360 19839
rect 12909 19805 12943 19839
rect 13093 19805 13127 19839
rect 13329 19805 13363 19839
rect 15945 19805 15979 19839
rect 16037 19805 16071 19839
rect 18061 19805 18095 19839
rect 18245 19805 18279 19839
rect 18337 19805 18371 19839
rect 23213 19805 23247 19839
rect 23581 19805 23615 19839
rect 24409 19805 24443 19839
rect 25513 19805 25547 19839
rect 25789 19805 25823 19839
rect 26525 19805 26559 19839
rect 26801 19805 26835 19839
rect 29745 19805 29779 19839
rect 31309 19805 31343 19839
rect 31401 19805 31435 19839
rect 32321 19805 32355 19839
rect 32597 19805 32631 19839
rect 33517 19805 33551 19839
rect 33609 19805 33643 19839
rect 34253 19805 34287 19839
rect 35449 19805 35483 19839
rect 37105 19805 37139 19839
rect 39681 19805 39715 19839
rect 40785 19805 40819 19839
rect 44281 19805 44315 19839
rect 3157 19737 3191 19771
rect 3249 19737 3283 19771
rect 4997 19737 5031 19771
rect 5089 19737 5123 19771
rect 9229 19737 9263 19771
rect 13185 19737 13219 19771
rect 14105 19737 14139 19771
rect 22845 19737 22879 19771
rect 23029 19737 23063 19771
rect 23305 19737 23339 19771
rect 24593 19737 24627 19771
rect 29009 19737 29043 19771
rect 29193 19737 29227 19771
rect 30021 19737 30055 19771
rect 33333 19737 33367 19771
rect 33977 19737 34011 19771
rect 8309 19669 8343 19703
rect 18521 19669 18555 19703
rect 23765 19669 23799 19703
rect 26341 19669 26375 19703
rect 31677 19669 31711 19703
rect 32781 19669 32815 19703
rect 33793 19669 33827 19703
rect 34437 19669 34471 19703
rect 35817 19669 35851 19703
rect 37473 19669 37507 19703
rect 38393 19669 38427 19703
rect 40233 19669 40267 19703
rect 44465 19669 44499 19703
rect 6929 19465 6963 19499
rect 8769 19465 8803 19499
rect 12633 19465 12667 19499
rect 19073 19465 19107 19499
rect 19165 19465 19199 19499
rect 20177 19465 20211 19499
rect 32505 19465 32539 19499
rect 34529 19465 34563 19499
rect 39957 19465 39991 19499
rect 44465 19465 44499 19499
rect 2421 19397 2455 19431
rect 2513 19397 2547 19431
rect 2973 19397 3007 19431
rect 6653 19397 6687 19431
rect 12541 19397 12575 19431
rect 13277 19397 13311 19431
rect 13662 19397 13696 19431
rect 15025 19397 15059 19431
rect 15318 19397 15352 19431
rect 15669 19397 15703 19431
rect 18613 19397 18647 19431
rect 22293 19397 22327 19431
rect 34069 19397 34103 19431
rect 2237 19329 2271 19363
rect 2610 19329 2644 19363
rect 2806 19329 2840 19363
rect 3341 19329 3375 19363
rect 6377 19329 6411 19363
rect 6561 19329 6595 19363
rect 6745 19329 6779 19363
rect 8585 19329 8619 19363
rect 10241 19329 10275 19363
rect 10425 19329 10459 19363
rect 10517 19329 10551 19363
rect 10661 19329 10695 19363
rect 13093 19329 13127 19363
rect 13369 19329 13403 19363
rect 13513 19329 13547 19363
rect 14749 19329 14783 19363
rect 14933 19329 14967 19363
rect 15169 19329 15203 19363
rect 15485 19329 15519 19363
rect 15853 19329 15887 19363
rect 18797 19329 18831 19363
rect 18889 19329 18923 19363
rect 19349 19329 19383 19363
rect 19441 19329 19475 19363
rect 19625 19329 19659 19363
rect 19717 19329 19751 19363
rect 19901 19329 19935 19363
rect 19993 19329 20027 19363
rect 20913 19329 20947 19363
rect 21097 19329 21131 19363
rect 22017 19329 22051 19363
rect 22109 19329 22143 19363
rect 31401 19329 31435 19363
rect 32137 19329 32171 19363
rect 34253 19329 34287 19363
rect 34345 19329 34379 19363
rect 38577 19329 38611 19363
rect 38833 19329 38867 19363
rect 40233 19329 40267 19363
rect 40417 19329 40451 19363
rect 42441 19329 42475 19363
rect 42708 19329 42742 19363
rect 44281 19329 44315 19363
rect 31493 19261 31527 19295
rect 32229 19261 32263 19295
rect 10793 19193 10827 19227
rect 31769 19193 31803 19227
rect 43821 19193 43855 19227
rect 18613 19125 18647 19159
rect 19349 19125 19383 19159
rect 19993 19125 20027 19159
rect 21281 19125 21315 19159
rect 21833 19125 21867 19159
rect 22109 19125 22143 19159
rect 31493 19125 31527 19159
rect 32137 19125 32171 19159
rect 34069 19125 34103 19159
rect 40049 19125 40083 19159
rect 2513 18921 2547 18955
rect 3433 18921 3467 18955
rect 4445 18921 4479 18955
rect 5733 18921 5767 18955
rect 9781 18921 9815 18955
rect 10517 18921 10551 18955
rect 11253 18921 11287 18955
rect 17049 18921 17083 18955
rect 21741 18921 21775 18955
rect 25145 18921 25179 18955
rect 27997 18921 28031 18955
rect 28917 18921 28951 18955
rect 29377 18921 29411 18955
rect 31677 18921 31711 18955
rect 37473 18921 37507 18955
rect 38485 18921 38519 18955
rect 3065 18853 3099 18887
rect 4813 18853 4847 18887
rect 7849 18853 7883 18887
rect 8677 18853 8711 18887
rect 12817 18853 12851 18887
rect 13553 18853 13587 18887
rect 15025 18853 15059 18887
rect 28457 18853 28491 18887
rect 38209 18853 38243 18887
rect 40141 18853 40175 18887
rect 42441 18853 42475 18887
rect 6193 18785 6227 18819
rect 7113 18785 7147 18819
rect 25053 18785 25087 18819
rect 28181 18785 28215 18819
rect 31493 18785 31527 18819
rect 37565 18785 37599 18819
rect 41061 18785 41095 18819
rect 43821 18785 43855 18819
rect 3249 18717 3283 18751
rect 3617 18717 3651 18751
rect 3893 18717 3927 18751
rect 4077 18717 4111 18751
rect 4313 18717 4347 18751
rect 5181 18717 5215 18751
rect 5601 18717 5635 18751
rect 6101 18717 6135 18751
rect 6469 18717 6503 18751
rect 6653 18717 6687 18751
rect 8033 18717 8067 18751
rect 8125 18717 8159 18751
rect 8309 18717 8343 18751
rect 8401 18717 8435 18751
rect 8545 18717 8579 18751
rect 9229 18717 9263 18751
rect 9505 18717 9539 18751
rect 9649 18717 9683 18751
rect 9965 18717 9999 18751
rect 10338 18717 10372 18751
rect 10701 18717 10735 18751
rect 11069 18717 11103 18751
rect 12265 18717 12299 18751
rect 12541 18717 12575 18751
rect 12638 18717 12672 18751
rect 13001 18717 13035 18751
rect 13369 18717 13403 18751
rect 14473 18717 14507 18751
rect 14657 18717 14691 18751
rect 14841 18717 14875 18751
rect 16773 18717 16807 18751
rect 16865 18717 16899 18751
rect 17049 18717 17083 18751
rect 19257 18717 19291 18751
rect 19441 18717 19475 18751
rect 21557 18717 21591 18751
rect 21741 18717 21775 18751
rect 21833 18717 21867 18751
rect 24961 18717 24995 18751
rect 27997 18717 28031 18751
rect 28273 18717 28307 18751
rect 29101 18717 29135 18751
rect 29193 18717 29227 18751
rect 31401 18717 31435 18751
rect 31677 18717 31711 18751
rect 37473 18717 37507 18751
rect 38025 18717 38059 18751
rect 38117 18717 38151 18751
rect 38301 18717 38335 18751
rect 40049 18717 40083 18751
rect 40233 18717 40267 18751
rect 40325 18717 40359 18751
rect 40509 18717 40543 18751
rect 43177 18717 43211 18751
rect 44281 18717 44315 18751
rect 2421 18649 2455 18683
rect 4169 18649 4203 18683
rect 4997 18649 5031 18683
rect 5365 18649 5399 18683
rect 5457 18649 5491 18683
rect 9413 18649 9447 18683
rect 10149 18649 10183 18683
rect 10241 18649 10275 18683
rect 10885 18649 10919 18683
rect 10977 18649 11011 18683
rect 12449 18649 12483 18683
rect 13185 18649 13219 18683
rect 13277 18649 13311 18683
rect 14749 18649 14783 18683
rect 29377 18649 29411 18683
rect 41328 18649 41362 18683
rect 16589 18581 16623 18615
rect 19625 18581 19659 18615
rect 22017 18581 22051 18615
rect 25329 18581 25363 18615
rect 28733 18581 28767 18615
rect 31861 18581 31895 18615
rect 37841 18581 37875 18615
rect 39865 18581 39899 18615
rect 42533 18581 42567 18615
rect 43269 18581 43303 18615
rect 44465 18581 44499 18615
rect 3433 18377 3467 18411
rect 15301 18377 15335 18411
rect 18153 18377 18187 18411
rect 19809 18377 19843 18411
rect 23305 18377 23339 18411
rect 24041 18377 24075 18411
rect 29745 18377 29779 18411
rect 31677 18377 31711 18411
rect 32597 18377 32631 18411
rect 37105 18377 37139 18411
rect 40877 18377 40911 18411
rect 41613 18377 41647 18411
rect 4077 18309 4111 18343
rect 5273 18309 5307 18343
rect 5365 18309 5399 18343
rect 6653 18309 6687 18343
rect 8309 18309 8343 18343
rect 8401 18309 8435 18343
rect 9137 18309 9171 18343
rect 12466 18309 12500 18343
rect 13921 18309 13955 18343
rect 15025 18309 15059 18343
rect 26985 18309 27019 18343
rect 29292 18309 29326 18343
rect 32137 18309 32171 18343
rect 36645 18309 36679 18343
rect 2513 18241 2547 18275
rect 2881 18241 2915 18275
rect 3709 18241 3743 18275
rect 4261 18241 4295 18275
rect 5176 18241 5210 18275
rect 5549 18241 5583 18275
rect 5733 18241 5767 18275
rect 6101 18241 6135 18275
rect 6469 18241 6503 18275
rect 6745 18241 6779 18275
rect 6842 18241 6876 18275
rect 8125 18241 8159 18275
rect 8498 18241 8532 18275
rect 8861 18241 8895 18275
rect 9045 18241 9079 18275
rect 9234 18241 9268 18275
rect 11897 18241 11931 18275
rect 12081 18241 12115 18275
rect 12173 18241 12207 18275
rect 12270 18241 12304 18275
rect 13737 18241 13771 18275
rect 14013 18241 14047 18275
rect 14105 18241 14139 18275
rect 14749 18241 14783 18275
rect 14933 18241 14967 18275
rect 15117 18241 15151 18275
rect 17049 18241 17083 18275
rect 17233 18241 17267 18275
rect 17325 18241 17359 18275
rect 17693 18241 17727 18275
rect 17969 18241 18003 18275
rect 19349 18241 19383 18275
rect 19625 18241 19659 18275
rect 22201 18241 22235 18275
rect 22385 18241 22419 18275
rect 22477 18241 22511 18275
rect 22845 18241 22879 18275
rect 23121 18241 23155 18275
rect 23581 18241 23615 18275
rect 23857 18241 23891 18275
rect 25329 18241 25363 18275
rect 25421 18241 25455 18275
rect 27261 18241 27295 18275
rect 29561 18241 29595 18275
rect 31217 18241 31251 18275
rect 31493 18241 31527 18275
rect 32321 18241 32355 18275
rect 32413 18241 32447 18275
rect 34161 18241 34195 18275
rect 34253 18241 34287 18275
rect 34437 18241 34471 18275
rect 34529 18263 34563 18297
rect 34713 18241 34747 18275
rect 36921 18241 36955 18275
rect 37381 18241 37415 18275
rect 37657 18241 37691 18275
rect 41521 18241 41555 18275
rect 41797 18241 41831 18275
rect 41889 18241 41923 18275
rect 42165 18241 42199 18275
rect 44281 18241 44315 18275
rect 2605 18173 2639 18207
rect 3065 18173 3099 18207
rect 8694 18173 8728 18207
rect 9430 18173 9464 18207
rect 12817 18173 12851 18207
rect 13093 18173 13127 18207
rect 17785 18173 17819 18207
rect 19165 18173 19199 18207
rect 19441 18173 19475 18207
rect 22937 18173 22971 18207
rect 23673 18173 23707 18207
rect 27077 18173 27111 18207
rect 29377 18173 29411 18207
rect 31309 18173 31343 18207
rect 36737 18173 36771 18207
rect 37749 18173 37783 18207
rect 40325 18173 40359 18207
rect 42073 18173 42107 18207
rect 4997 18105 5031 18139
rect 7021 18105 7055 18139
rect 14289 18105 14323 18139
rect 22661 18105 22695 18139
rect 29101 18105 29135 18139
rect 37381 18105 37415 18139
rect 4537 18037 4571 18071
rect 17049 18037 17083 18071
rect 17509 18037 17543 18071
rect 17693 18037 17727 18071
rect 19349 18037 19383 18071
rect 22385 18037 22419 18071
rect 23121 18037 23155 18071
rect 23765 18037 23799 18071
rect 25421 18037 25455 18071
rect 25697 18037 25731 18071
rect 26985 18037 27019 18071
rect 27445 18037 27479 18071
rect 29285 18037 29319 18071
rect 31309 18037 31343 18071
rect 32137 18037 32171 18071
rect 33977 18037 34011 18071
rect 34161 18037 34195 18071
rect 34529 18037 34563 18071
rect 34897 18037 34931 18071
rect 36645 18037 36679 18071
rect 37565 18037 37599 18071
rect 39681 18037 39715 18071
rect 44465 18037 44499 18071
rect 2421 17833 2455 17867
rect 3157 17833 3191 17867
rect 5365 17833 5399 17867
rect 8125 17833 8159 17867
rect 9965 17833 9999 17867
rect 15209 17833 15243 17867
rect 16681 17833 16715 17867
rect 17141 17833 17175 17867
rect 22937 17833 22971 17867
rect 23397 17833 23431 17867
rect 25973 17833 26007 17867
rect 26249 17833 26283 17867
rect 26985 17833 27019 17867
rect 27721 17833 27755 17867
rect 29837 17833 29871 17867
rect 31401 17833 31435 17867
rect 31953 17833 31987 17867
rect 32505 17833 32539 17867
rect 33241 17833 33275 17867
rect 33885 17833 33919 17867
rect 34069 17833 34103 17867
rect 35357 17833 35391 17867
rect 35725 17833 35759 17867
rect 36185 17833 36219 17867
rect 37289 17833 37323 17867
rect 37749 17833 37783 17867
rect 41521 17833 41555 17867
rect 4445 17765 4479 17799
rect 6745 17765 6779 17799
rect 12265 17765 12299 17799
rect 34345 17765 34379 17799
rect 35265 17765 35299 17799
rect 38393 17765 38427 17799
rect 41245 17765 41279 17799
rect 41981 17765 42015 17799
rect 16773 17697 16807 17731
rect 19809 17697 19843 17731
rect 23029 17697 23063 17731
rect 27905 17697 27939 17731
rect 31217 17697 31251 17731
rect 31769 17697 31803 17731
rect 32413 17697 32447 17731
rect 33149 17697 33183 17731
rect 35449 17697 35483 17731
rect 36369 17697 36403 17731
rect 42165 17697 42199 17731
rect 43085 17697 43119 17731
rect 2605 17629 2639 17663
rect 2973 17629 3007 17663
rect 3341 17629 3375 17663
rect 4261 17629 4295 17663
rect 5549 17629 5583 17663
rect 6193 17629 6227 17663
rect 6469 17629 6503 17663
rect 6613 17629 6647 17663
rect 7481 17629 7515 17663
rect 7757 17629 7791 17663
rect 9413 17629 9447 17663
rect 9786 17629 9820 17663
rect 11713 17629 11747 17663
rect 11989 17629 12023 17663
rect 12086 17629 12120 17663
rect 12449 17629 12483 17663
rect 12725 17629 12759 17663
rect 16681 17629 16715 17663
rect 16957 17629 16991 17663
rect 19625 17629 19659 17663
rect 23213 17629 23247 17663
rect 25605 17629 25639 17663
rect 26249 17629 26283 17663
rect 26433 17629 26467 17663
rect 26525 17629 26559 17663
rect 27169 17629 27203 17663
rect 27261 17629 27295 17663
rect 27997 17629 28031 17663
rect 29745 17629 29779 17663
rect 29837 17629 29871 17663
rect 31125 17629 31159 17663
rect 31401 17629 31435 17663
rect 31953 17629 31987 17663
rect 32505 17629 32539 17663
rect 33241 17629 33275 17663
rect 33517 17629 33551 17663
rect 33977 17629 34011 17663
rect 34069 17629 34103 17663
rect 35357 17629 35391 17663
rect 36461 17629 36495 17663
rect 37105 17629 37139 17663
rect 37473 17629 37507 17663
rect 37565 17629 37599 17663
rect 38209 17629 38243 17663
rect 38853 17629 38887 17663
rect 39865 17629 39899 17663
rect 40132 17629 40166 17663
rect 41429 17629 41463 17663
rect 41705 17629 41739 17663
rect 41797 17629 41831 17663
rect 42073 17629 42107 17663
rect 42289 17629 42323 17663
rect 42441 17629 42475 17663
rect 43729 17629 43763 17663
rect 5733 17561 5767 17595
rect 5917 17561 5951 17595
rect 6377 17561 6411 17595
rect 7849 17561 7883 17595
rect 7966 17561 8000 17595
rect 9597 17561 9631 17595
rect 9689 17561 9723 17595
rect 11897 17561 11931 17595
rect 14933 17561 14967 17595
rect 15117 17561 15151 17595
rect 19441 17561 19475 17595
rect 22937 17561 22971 17595
rect 25789 17561 25823 17595
rect 26985 17561 27019 17595
rect 27721 17561 27755 17595
rect 29567 17561 29601 17595
rect 31677 17561 31711 17595
rect 32229 17561 32263 17595
rect 32965 17561 32999 17595
rect 33701 17561 33735 17595
rect 34897 17561 34931 17595
rect 35081 17561 35115 17595
rect 36185 17561 36219 17595
rect 37289 17561 37323 17595
rect 38669 17561 38703 17595
rect 39037 17561 39071 17595
rect 3525 17493 3559 17527
rect 26709 17493 26743 17527
rect 26893 17493 26927 17527
rect 27445 17493 27479 17527
rect 28181 17493 28215 17527
rect 30021 17493 30055 17527
rect 31585 17493 31619 17527
rect 32137 17493 32171 17527
rect 32689 17493 32723 17527
rect 33425 17493 33459 17527
rect 36645 17493 36679 17527
rect 42625 17493 42659 17527
rect 3801 17289 3835 17323
rect 8401 17289 8435 17323
rect 8953 17289 8987 17323
rect 9321 17289 9355 17323
rect 10701 17289 10735 17323
rect 11713 17289 11747 17323
rect 14933 17289 14967 17323
rect 19090 17289 19124 17323
rect 23397 17289 23431 17323
rect 27353 17289 27387 17323
rect 36093 17289 36127 17323
rect 36829 17289 36863 17323
rect 38301 17289 38335 17323
rect 40693 17289 40727 17323
rect 43821 17289 43855 17323
rect 7113 17221 7147 17255
rect 7665 17221 7699 17255
rect 8125 17221 8159 17255
rect 12541 17221 12575 17255
rect 14013 17221 14047 17255
rect 23213 17221 23247 17255
rect 27721 17221 27755 17255
rect 32137 17221 32171 17255
rect 32321 17221 32355 17255
rect 35633 17221 35667 17255
rect 36369 17221 36403 17255
rect 2237 17153 2271 17187
rect 3617 17153 3651 17187
rect 4261 17153 4295 17187
rect 4445 17153 4479 17187
rect 6101 17153 6135 17187
rect 6929 17153 6963 17187
rect 7297 17153 7331 17187
rect 8769 17153 8803 17187
rect 9137 17153 9171 17187
rect 9505 17153 9539 17187
rect 9689 17153 9723 17187
rect 9781 17153 9815 17187
rect 9878 17153 9912 17187
rect 10793 17153 10827 17187
rect 11989 17153 12023 17187
rect 12173 17153 12207 17187
rect 12357 17153 12391 17187
rect 13001 17153 13035 17187
rect 13185 17153 13219 17187
rect 13277 17153 13311 17187
rect 13374 17153 13408 17187
rect 13737 17153 13771 17187
rect 13921 17153 13955 17187
rect 14110 17153 14144 17187
rect 14657 17153 14691 17187
rect 15025 17153 15059 17187
rect 18521 17153 18555 17187
rect 18705 17153 18739 17187
rect 18797 17153 18831 17187
rect 18894 17153 18928 17187
rect 19257 17153 19291 17187
rect 19441 17153 19475 17187
rect 23029 17153 23063 17187
rect 24777 17153 24811 17187
rect 25053 17153 25087 17187
rect 26985 17153 27019 17187
rect 27905 17153 27939 17187
rect 27997 17153 28031 17187
rect 29469 17153 29503 17187
rect 31573 17159 31607 17193
rect 31769 17153 31803 17187
rect 35909 17153 35943 17187
rect 36645 17153 36679 17187
rect 37657 17153 37691 17187
rect 37841 17153 37875 17187
rect 38393 17153 38427 17187
rect 38577 17153 38611 17187
rect 38761 17153 38795 17187
rect 39037 17153 39071 17187
rect 39313 17153 39347 17187
rect 39569 17153 39603 17187
rect 42441 17153 42475 17187
rect 42708 17153 42742 17187
rect 44281 17153 44315 17187
rect 8217 17085 8251 17119
rect 11621 17085 11655 17119
rect 14473 17085 14507 17119
rect 24869 17085 24903 17119
rect 27077 17085 27111 17119
rect 29561 17085 29595 17119
rect 35725 17085 35759 17119
rect 36461 17085 36495 17119
rect 38853 17085 38887 17119
rect 39221 17085 39255 17119
rect 5917 17017 5951 17051
rect 7481 17017 7515 17051
rect 7665 17017 7699 17051
rect 10057 17017 10091 17051
rect 13553 17017 13587 17051
rect 14289 17017 14323 17051
rect 29837 17017 29871 17051
rect 31953 17017 31987 17051
rect 32505 17017 32539 17051
rect 38025 17017 38059 17051
rect 38945 17017 38979 17051
rect 44465 17017 44499 17051
rect 2329 16949 2363 16983
rect 4077 16949 4111 16983
rect 4721 16949 4755 16983
rect 19349 16949 19383 16983
rect 19625 16949 19659 16983
rect 24961 16949 24995 16983
rect 25237 16949 25271 16983
rect 27169 16949 27203 16983
rect 27813 16949 27847 16983
rect 28181 16949 28215 16983
rect 29469 16949 29503 16983
rect 31677 16949 31711 16983
rect 35633 16949 35667 16983
rect 36369 16949 36403 16983
rect 37381 16949 37415 16983
rect 2513 16745 2547 16779
rect 3617 16745 3651 16779
rect 4353 16745 4387 16779
rect 8769 16745 8803 16779
rect 21097 16745 21131 16779
rect 21833 16745 21867 16779
rect 22477 16745 22511 16779
rect 22845 16745 22879 16779
rect 24685 16745 24719 16779
rect 24869 16745 24903 16779
rect 25513 16745 25547 16779
rect 28457 16745 28491 16779
rect 31677 16745 31711 16779
rect 32137 16745 32171 16779
rect 32505 16745 32539 16779
rect 38577 16745 38611 16779
rect 1777 16677 1811 16711
rect 2881 16677 2915 16711
rect 3065 16677 3099 16711
rect 8033 16677 8067 16711
rect 17417 16677 17451 16711
rect 17877 16677 17911 16711
rect 21373 16677 21407 16711
rect 25881 16677 25915 16711
rect 32045 16677 32079 16711
rect 37657 16677 37691 16711
rect 38393 16677 38427 16711
rect 2329 16609 2363 16643
rect 4077 16609 4111 16643
rect 4721 16609 4755 16643
rect 7113 16609 7147 16643
rect 10609 16609 10643 16643
rect 10977 16609 11011 16643
rect 21005 16609 21039 16643
rect 25053 16609 25087 16643
rect 25513 16609 25547 16643
rect 26341 16609 26375 16643
rect 28549 16609 28583 16643
rect 31769 16609 31803 16643
rect 32229 16609 32263 16643
rect 37749 16609 37783 16643
rect 37841 16609 37875 16643
rect 1409 16541 1443 16575
rect 2697 16541 2731 16575
rect 3249 16541 3283 16575
rect 3893 16541 3927 16575
rect 3985 16541 4019 16575
rect 4169 16541 4203 16575
rect 4905 16541 4939 16575
rect 5273 16541 5307 16575
rect 5457 16541 5491 16575
rect 5825 16541 5859 16575
rect 6101 16541 6135 16575
rect 6469 16541 6503 16575
rect 7021 16541 7055 16575
rect 7665 16541 7699 16575
rect 8585 16541 8619 16575
rect 9137 16541 9171 16575
rect 9510 16541 9544 16575
rect 9965 16541 9999 16575
rect 10057 16541 10091 16575
rect 10425 16541 10459 16575
rect 11253 16541 11287 16575
rect 11626 16541 11660 16575
rect 15761 16541 15795 16575
rect 16129 16541 16163 16575
rect 21189 16541 21223 16575
rect 22661 16541 22695 16575
rect 22845 16541 22879 16575
rect 24869 16541 24903 16575
rect 25145 16541 25179 16575
rect 25697 16541 25731 16575
rect 28773 16541 28807 16575
rect 31677 16541 31711 16575
rect 32137 16541 32171 16575
rect 37565 16541 37599 16575
rect 38025 16541 38059 16575
rect 38669 16541 38703 16575
rect 44281 16541 44315 16575
rect 1777 16473 1811 16507
rect 2237 16473 2271 16507
rect 3433 16473 3467 16507
rect 5641 16473 5675 16507
rect 5733 16473 5767 16507
rect 8033 16473 8067 16507
rect 9321 16473 9355 16507
rect 9413 16473 9447 16507
rect 11437 16473 11471 16507
rect 11529 16473 11563 16507
rect 15945 16473 15979 16507
rect 16037 16473 16071 16507
rect 17049 16473 17083 16507
rect 17233 16473 17267 16507
rect 17509 16473 17543 16507
rect 17693 16473 17727 16507
rect 20913 16473 20947 16507
rect 21465 16473 21499 16507
rect 21649 16473 21683 16507
rect 25421 16473 25455 16507
rect 25973 16473 26007 16507
rect 26157 16473 26191 16507
rect 28457 16473 28491 16507
rect 38209 16473 38243 16507
rect 1593 16405 1627 16439
rect 3341 16405 3375 16439
rect 5181 16405 5215 16439
rect 6009 16405 6043 16439
rect 7389 16405 7423 16439
rect 8493 16405 8527 16439
rect 9706 16405 9740 16439
rect 11813 16405 11847 16439
rect 16313 16405 16347 16439
rect 25329 16405 25363 16439
rect 28917 16405 28951 16439
rect 37381 16405 37415 16439
rect 44465 16405 44499 16439
rect 1593 16201 1627 16235
rect 5457 16201 5491 16235
rect 6653 16201 6687 16235
rect 8585 16201 8619 16235
rect 10885 16201 10919 16235
rect 15301 16201 15335 16235
rect 17509 16201 17543 16235
rect 20545 16201 20579 16235
rect 22201 16201 22235 16235
rect 25421 16201 25455 16235
rect 26157 16201 26191 16235
rect 29009 16201 29043 16235
rect 32413 16201 32447 16235
rect 32965 16201 32999 16235
rect 38761 16201 38795 16235
rect 4537 16133 4571 16167
rect 5549 16133 5583 16167
rect 6193 16133 6227 16167
rect 10517 16133 10551 16167
rect 11805 16133 11839 16167
rect 15209 16133 15243 16167
rect 18613 16133 18647 16167
rect 25053 16133 25087 16167
rect 25789 16133 25823 16167
rect 25973 16133 26007 16167
rect 37289 16133 37323 16167
rect 1409 16065 1443 16099
rect 1961 16065 1995 16099
rect 2053 16065 2087 16099
rect 2145 16065 2179 16099
rect 2789 16065 2823 16099
rect 3525 16065 3559 16099
rect 3893 16065 3927 16099
rect 4629 16065 4663 16099
rect 5825 16065 5859 16099
rect 7021 16065 7055 16099
rect 7389 16065 7423 16099
rect 7573 16065 7607 16099
rect 7941 16065 7975 16099
rect 8769 16065 8803 16099
rect 9229 16065 9263 16099
rect 9597 16065 9631 16099
rect 10333 16065 10367 16099
rect 10609 16065 10643 16099
rect 10701 16065 10735 16099
rect 11621 16065 11655 16099
rect 11897 16065 11931 16099
rect 12041 16065 12075 16099
rect 12357 16065 12391 16099
rect 12725 16065 12759 16099
rect 13001 16065 13035 16099
rect 15669 16065 15703 16099
rect 15853 16065 15887 16099
rect 15945 16065 15979 16099
rect 16089 16065 16123 16099
rect 17049 16065 17083 16099
rect 17325 16065 17359 16099
rect 18889 16065 18923 16099
rect 20085 16065 20119 16099
rect 20361 16065 20395 16099
rect 22385 16065 22419 16099
rect 22661 16065 22695 16099
rect 22753 16065 22787 16099
rect 22937 16065 22971 16099
rect 23029 16065 23063 16099
rect 25237 16065 25271 16099
rect 29193 16065 29227 16099
rect 29469 16065 29503 16099
rect 29561 16065 29595 16099
rect 29745 16065 29779 16099
rect 32597 16065 32631 16099
rect 33057 16065 33091 16099
rect 35081 16065 35115 16099
rect 35357 16065 35391 16099
rect 35817 16065 35851 16099
rect 36001 16065 36035 16099
rect 36277 16065 36311 16099
rect 36369 16065 36403 16099
rect 36829 16065 36863 16099
rect 39405 16065 39439 16099
rect 44281 16065 44315 16099
rect 2237 15997 2271 16031
rect 2421 15997 2455 16031
rect 3617 15997 3651 16031
rect 4077 15997 4111 16031
rect 6929 15997 6963 16031
rect 8217 15997 8251 16031
rect 8309 15997 8343 16031
rect 8426 15997 8460 16031
rect 9321 15997 9355 16031
rect 9505 15997 9539 16031
rect 13093 15997 13127 16031
rect 17141 15997 17175 16031
rect 18705 15997 18739 16031
rect 20177 15997 20211 16031
rect 22477 15997 22511 16031
rect 29377 15997 29411 16031
rect 32689 15997 32723 16031
rect 35173 15997 35207 16031
rect 36093 15997 36127 16031
rect 36553 15997 36587 16031
rect 36645 15997 36679 16031
rect 37933 15997 37967 16031
rect 38669 15997 38703 16031
rect 8953 15929 8987 15963
rect 12173 15929 12207 15963
rect 16221 15929 16255 15963
rect 35541 15929 35575 15963
rect 35909 15929 35943 15963
rect 36737 15929 36771 15963
rect 38025 15929 38059 15963
rect 2881 15861 2915 15895
rect 4813 15861 4847 15895
rect 9965 15861 9999 15895
rect 13185 15861 13219 15895
rect 13369 15861 13403 15895
rect 17233 15861 17267 15895
rect 18797 15861 18831 15895
rect 19073 15861 19107 15895
rect 20085 15861 20119 15895
rect 22385 15861 22419 15895
rect 23029 15861 23063 15895
rect 23213 15861 23247 15895
rect 29193 15861 29227 15895
rect 29745 15861 29779 15895
rect 29929 15861 29963 15895
rect 32597 15861 32631 15895
rect 35081 15861 35115 15895
rect 35633 15861 35667 15895
rect 37013 15861 37047 15895
rect 44465 15861 44499 15895
rect 1593 15657 1627 15691
rect 5365 15657 5399 15691
rect 5917 15657 5951 15691
rect 6653 15657 6687 15691
rect 8493 15657 8527 15691
rect 14657 15657 14691 15691
rect 16497 15657 16531 15691
rect 22293 15657 22327 15691
rect 22753 15657 22787 15691
rect 23857 15657 23891 15691
rect 25605 15657 25639 15691
rect 28089 15657 28123 15691
rect 28273 15657 28307 15691
rect 29561 15657 29595 15691
rect 29929 15657 29963 15691
rect 32413 15657 32447 15691
rect 32597 15657 32631 15691
rect 32873 15657 32907 15691
rect 33333 15657 33367 15691
rect 33517 15657 33551 15691
rect 34253 15657 34287 15691
rect 34437 15657 34471 15691
rect 34805 15657 34839 15691
rect 35173 15657 35207 15691
rect 37013 15657 37047 15691
rect 2881 15589 2915 15623
rect 5641 15589 5675 15623
rect 7389 15589 7423 15623
rect 13093 15589 13127 15623
rect 13921 15589 13955 15623
rect 3617 15521 3651 15555
rect 9505 15521 9539 15555
rect 9965 15521 9999 15555
rect 10425 15521 10459 15555
rect 11069 15521 11103 15555
rect 14841 15521 14875 15555
rect 15117 15521 15151 15555
rect 22477 15521 22511 15555
rect 27905 15521 27939 15555
rect 32873 15521 32907 15555
rect 33149 15521 33183 15555
rect 34805 15521 34839 15555
rect 40969 15521 41003 15555
rect 1409 15453 1443 15487
rect 2421 15453 2455 15487
rect 3433 15453 3467 15487
rect 5181 15453 5215 15487
rect 5457 15453 5491 15487
rect 5733 15453 5767 15487
rect 6101 15453 6135 15487
rect 6377 15453 6411 15487
rect 6521 15453 6555 15487
rect 6837 15453 6871 15487
rect 7257 15453 7291 15487
rect 7573 15453 7607 15487
rect 8033 15453 8067 15487
rect 8125 15453 8159 15487
rect 8217 15453 8251 15487
rect 8401 15453 8435 15487
rect 8493 15453 8527 15487
rect 8677 15453 8711 15487
rect 8953 15453 8987 15487
rect 9413 15453 9447 15487
rect 9781 15453 9815 15487
rect 11161 15453 11195 15487
rect 11529 15453 11563 15487
rect 11713 15453 11747 15487
rect 12541 15453 12575 15487
rect 12725 15453 12759 15487
rect 12914 15453 12948 15487
rect 14105 15453 14139 15487
rect 14473 15453 14507 15487
rect 15945 15453 15979 15487
rect 16365 15453 16399 15487
rect 17693 15453 17727 15487
rect 17969 15453 18003 15487
rect 18066 15453 18100 15487
rect 18262 15453 18296 15487
rect 18429 15453 18463 15487
rect 18705 15453 18739 15487
rect 18849 15453 18883 15487
rect 22569 15453 22603 15487
rect 23857 15453 23891 15487
rect 23949 15453 23983 15487
rect 25421 15453 25455 15487
rect 25513 15453 25547 15487
rect 25697 15453 25731 15487
rect 26709 15453 26743 15487
rect 28089 15453 28123 15487
rect 29561 15453 29595 15487
rect 29653 15453 29687 15487
rect 32965 15453 32999 15487
rect 33057 15453 33091 15487
rect 33333 15453 33367 15487
rect 33609 15453 33643 15487
rect 34069 15453 34103 15487
rect 34253 15453 34287 15487
rect 34989 15453 35023 15487
rect 35633 15453 35667 15487
rect 35900 15453 35934 15487
rect 37105 15453 37139 15487
rect 40877 15453 40911 15487
rect 41153 15453 41187 15487
rect 41245 15453 41279 15487
rect 41521 15453 41555 15487
rect 44281 15453 44315 15487
rect 2881 15385 2915 15419
rect 6285 15385 6319 15419
rect 7021 15385 7055 15419
rect 7113 15385 7147 15419
rect 12173 15385 12207 15419
rect 12817 15385 12851 15419
rect 13737 15385 13771 15419
rect 14289 15385 14323 15419
rect 14381 15385 14415 15419
rect 16129 15385 16163 15419
rect 16221 15385 16255 15419
rect 17877 15385 17911 15419
rect 18613 15385 18647 15419
rect 22293 15385 22327 15419
rect 26893 15385 26927 15419
rect 27813 15385 27847 15419
rect 33793 15385 33827 15419
rect 33977 15385 34011 15419
rect 34713 15385 34747 15419
rect 37350 15385 37384 15419
rect 41429 15385 41463 15419
rect 41766 15385 41800 15419
rect 2605 15317 2639 15351
rect 3341 15317 3375 15351
rect 7757 15317 7791 15351
rect 9137 15317 9171 15351
rect 10793 15317 10827 15351
rect 12081 15317 12115 15351
rect 18998 15317 19032 15351
rect 24225 15317 24259 15351
rect 25237 15317 25271 15351
rect 27077 15317 27111 15351
rect 38485 15317 38519 15351
rect 42901 15317 42935 15351
rect 44465 15317 44499 15351
rect 3157 15113 3191 15147
rect 8861 15113 8895 15147
rect 9045 15113 9079 15147
rect 11069 15113 11103 15147
rect 12173 15113 12207 15147
rect 12541 15113 12575 15147
rect 23857 15113 23891 15147
rect 26617 15113 26651 15147
rect 27353 15113 27387 15147
rect 27905 15113 27939 15147
rect 31953 15113 31987 15147
rect 33977 15113 34011 15147
rect 39037 15113 39071 15147
rect 42441 15113 42475 15147
rect 3065 15045 3099 15079
rect 6469 15045 6503 15079
rect 8309 15045 8343 15079
rect 8769 15045 8803 15079
rect 9505 15045 9539 15079
rect 14841 15045 14875 15079
rect 18889 15045 18923 15079
rect 18981 15045 19015 15079
rect 30665 15045 30699 15079
rect 33517 15045 33551 15079
rect 37902 15045 37936 15079
rect 3341 14977 3375 15011
rect 6009 14977 6043 15011
rect 7113 14977 7147 15011
rect 7297 14977 7331 15011
rect 9137 14977 9171 15011
rect 10333 14977 10367 15011
rect 10701 14977 10735 15011
rect 11713 14977 11747 15011
rect 12081 14977 12115 15011
rect 12357 14977 12391 15011
rect 14657 14977 14691 15011
rect 14933 14977 14967 15011
rect 15077 14977 15111 15011
rect 18705 14977 18739 15011
rect 19078 14977 19112 15011
rect 24041 14977 24075 15011
rect 24317 14977 24351 15011
rect 26157 14977 26191 15011
rect 26433 14977 26467 15011
rect 26985 14977 27019 15011
rect 27537 14977 27571 15011
rect 30849 14977 30883 15011
rect 30941 14977 30975 15011
rect 31217 14977 31251 15011
rect 31493 14977 31527 15011
rect 31677 14977 31711 15011
rect 31769 14977 31803 15011
rect 33701 14977 33735 15011
rect 33793 14977 33827 15011
rect 37657 14977 37691 15011
rect 2605 14909 2639 14943
rect 2697 14909 2731 14943
rect 2789 14909 2823 14943
rect 2881 14909 2915 14943
rect 9413 14909 9447 14943
rect 9622 14909 9656 14943
rect 10425 14909 10459 14943
rect 10609 14909 10643 14943
rect 24133 14909 24167 14943
rect 26249 14909 26283 14943
rect 27077 14909 27111 14943
rect 27629 14909 27663 14943
rect 31033 14909 31067 14943
rect 43085 14909 43119 14943
rect 6653 14841 6687 14875
rect 8309 14841 8343 14875
rect 11897 14841 11931 14875
rect 15209 14841 15243 14875
rect 19257 14841 19291 14875
rect 30481 14841 30515 14875
rect 6101 14773 6135 14807
rect 7021 14773 7055 14807
rect 7481 14773 7515 14807
rect 9781 14773 9815 14807
rect 24317 14773 24351 14807
rect 26341 14773 26375 14807
rect 27077 14773 27111 14807
rect 27721 14773 27755 14807
rect 30941 14773 30975 14807
rect 31401 14773 31435 14807
rect 31769 14773 31803 14807
rect 33517 14773 33551 14807
rect 1593 14569 1627 14603
rect 6101 14569 6135 14603
rect 7941 14569 7975 14603
rect 8585 14569 8619 14603
rect 20085 14569 20119 14603
rect 21833 14569 21867 14603
rect 22753 14569 22787 14603
rect 22937 14569 22971 14603
rect 23581 14569 23615 14603
rect 24041 14569 24075 14603
rect 30941 14569 30975 14603
rect 31125 14569 31159 14603
rect 6285 14501 6319 14535
rect 8769 14501 8803 14535
rect 9597 14501 9631 14535
rect 16497 14501 16531 14535
rect 19901 14501 19935 14535
rect 5641 14433 5675 14467
rect 5917 14433 5951 14467
rect 6745 14433 6779 14467
rect 7849 14433 7883 14467
rect 8033 14433 8067 14467
rect 8953 14433 8987 14467
rect 9438 14433 9472 14467
rect 14657 14433 14691 14467
rect 22569 14433 22603 14467
rect 23765 14433 23799 14467
rect 1409 14365 1443 14399
rect 5089 14365 5123 14399
rect 5733 14365 5767 14399
rect 5825 14365 5859 14399
rect 8493 14365 8527 14399
rect 8585 14365 8619 14399
rect 9321 14365 9355 14399
rect 9689 14365 9723 14399
rect 14105 14365 14139 14399
rect 14289 14365 14323 14399
rect 15577 14365 15611 14399
rect 15945 14365 15979 14399
rect 16129 14365 16163 14399
rect 16318 14365 16352 14399
rect 20085 14365 20119 14399
rect 20177 14365 20211 14399
rect 21373 14365 21407 14399
rect 21741 14365 21775 14399
rect 21833 14365 21867 14399
rect 22753 14365 22787 14399
rect 23581 14365 23615 14399
rect 23857 14365 23891 14399
rect 30757 14365 30791 14399
rect 30849 14365 30883 14399
rect 44281 14365 44315 14399
rect 2329 14297 2363 14331
rect 6285 14297 6319 14331
rect 8217 14297 8251 14331
rect 8309 14297 8343 14331
rect 9229 14297 9263 14331
rect 15209 14297 15243 14331
rect 16221 14297 16255 14331
rect 20361 14297 20395 14331
rect 22477 14297 22511 14331
rect 2237 14229 2271 14263
rect 5273 14229 5307 14263
rect 6837 14229 6871 14263
rect 7021 14229 7055 14263
rect 8125 14229 8159 14263
rect 9873 14229 9907 14263
rect 14565 14229 14599 14263
rect 15301 14229 15335 14263
rect 15669 14229 15703 14263
rect 22017 14229 22051 14263
rect 44465 14229 44499 14263
rect 1593 14025 1627 14059
rect 2513 14025 2547 14059
rect 3249 14025 3283 14059
rect 5733 14025 5767 14059
rect 5917 14025 5951 14059
rect 12089 14025 12123 14059
rect 15577 14025 15611 14059
rect 16313 14025 16347 14059
rect 17141 14025 17175 14059
rect 23029 14025 23063 14059
rect 28089 14025 28123 14059
rect 28365 14025 28399 14059
rect 29009 14025 29043 14059
rect 32505 14025 32539 14059
rect 44465 14025 44499 14059
rect 2973 13957 3007 13991
rect 3090 13957 3124 13991
rect 5181 13957 5215 13991
rect 17049 13957 17083 13991
rect 21097 13957 21131 13991
rect 22017 13957 22051 13991
rect 22201 13957 22235 13991
rect 22845 13957 22879 13991
rect 27629 13957 27663 13991
rect 32137 13957 32171 13991
rect 32321 13957 32355 13991
rect 1409 13889 1443 13923
rect 1685 13889 1719 13923
rect 2329 13889 2363 13923
rect 4169 13889 4203 13923
rect 4445 13889 4479 13923
rect 8217 13889 8251 13923
rect 8309 13889 8343 13923
rect 8585 13889 8619 13923
rect 9045 13889 9079 13923
rect 9413 13889 9447 13923
rect 10425 13889 10459 13923
rect 11161 13889 11195 13923
rect 11529 13889 11563 13923
rect 11713 13889 11747 13923
rect 11805 13889 11839 13923
rect 11949 13889 11983 13923
rect 14565 13889 14599 13923
rect 14657 13889 14691 13923
rect 15025 13889 15059 13923
rect 15761 13889 15795 13923
rect 15945 13889 15979 13923
rect 16037 13889 16071 13923
rect 16129 13889 16163 13923
rect 17417 13889 17451 13923
rect 17601 13889 17635 13923
rect 17693 13889 17727 13923
rect 17785 13889 17819 13923
rect 18705 13889 18739 13923
rect 18889 13889 18923 13923
rect 18981 13889 19015 13923
rect 19125 13889 19159 13923
rect 19274 13889 19308 13923
rect 20913 13889 20947 13923
rect 21833 13889 21867 13923
rect 22661 13889 22695 13923
rect 25881 13889 25915 13923
rect 26065 13889 26099 13923
rect 26433 13889 26467 13923
rect 26617 13889 26651 13923
rect 26801 13889 26835 13923
rect 26985 13889 27019 13923
rect 27169 13889 27203 13923
rect 27537 13889 27571 13923
rect 27905 13889 27939 13923
rect 28181 13889 28215 13923
rect 28825 13889 28859 13923
rect 44281 13889 44315 13923
rect 1869 13821 1903 13855
rect 1961 13821 1995 13855
rect 2053 13821 2087 13855
rect 2145 13821 2179 13855
rect 2605 13821 2639 13855
rect 2881 13821 2915 13855
rect 4629 13821 4663 13855
rect 4721 13821 4755 13855
rect 4813 13821 4847 13855
rect 4905 13821 4939 13855
rect 5641 13821 5675 13855
rect 8769 13821 8803 13855
rect 15117 13821 15151 13855
rect 21281 13821 21315 13855
rect 27721 13821 27755 13855
rect 4353 13753 4387 13787
rect 5181 13753 5215 13787
rect 17969 13753 18003 13787
rect 9229 13685 9263 13719
rect 10609 13685 10643 13719
rect 10977 13685 11011 13719
rect 25881 13685 25915 13719
rect 26249 13685 26283 13719
rect 27905 13685 27939 13719
rect 2237 13481 2271 13515
rect 4629 13481 4663 13515
rect 4905 13481 4939 13515
rect 5549 13481 5583 13515
rect 7389 13481 7423 13515
rect 7665 13481 7699 13515
rect 11253 13481 11287 13515
rect 11897 13481 11931 13515
rect 13093 13481 13127 13515
rect 17417 13481 17451 13515
rect 22293 13481 22327 13515
rect 22477 13481 22511 13515
rect 25329 13481 25363 13515
rect 26709 13481 26743 13515
rect 28917 13481 28951 13515
rect 29285 13481 29319 13515
rect 31401 13481 31435 13515
rect 2421 13413 2455 13447
rect 3893 13413 3927 13447
rect 5181 13413 5215 13447
rect 8677 13413 8711 13447
rect 9137 13413 9171 13447
rect 11529 13413 11563 13447
rect 27077 13413 27111 13447
rect 1593 13345 1627 13379
rect 2078 13345 2112 13379
rect 3525 13345 3559 13379
rect 5641 13345 5675 13379
rect 6009 13345 6043 13379
rect 6377 13345 6411 13379
rect 6469 13345 6503 13379
rect 22201 13345 22235 13379
rect 26801 13345 26835 13379
rect 28917 13345 28951 13379
rect 1961 13277 1995 13311
rect 2973 13277 3007 13311
rect 4721 13277 4755 13311
rect 4997 13277 5031 13311
rect 5420 13277 5454 13311
rect 6745 13277 6779 13311
rect 7205 13277 7239 13311
rect 7481 13277 7515 13311
rect 7849 13277 7883 13311
rect 8401 13277 8435 13311
rect 9269 13277 9303 13311
rect 9400 13277 9434 13311
rect 9505 13277 9539 13311
rect 9689 13277 9723 13311
rect 9965 13277 9999 13311
rect 10333 13277 10367 13311
rect 10701 13277 10735 13311
rect 10977 13277 11011 13311
rect 11121 13277 11155 13311
rect 11713 13277 11747 13311
rect 12029 13277 12063 13311
rect 12176 13277 12210 13311
rect 12449 13277 12483 13311
rect 12541 13277 12575 13311
rect 12725 13277 12759 13311
rect 12914 13277 12948 13311
rect 13277 13277 13311 13311
rect 13645 13277 13679 13311
rect 14657 13277 14691 13311
rect 15025 13277 15059 13311
rect 15209 13277 15243 13311
rect 16865 13277 16899 13311
rect 17238 13277 17272 13311
rect 22109 13277 22143 13311
rect 26709 13277 26743 13311
rect 28549 13277 28583 13311
rect 28733 13277 28767 13311
rect 29101 13277 29135 13311
rect 2421 13209 2455 13243
rect 3341 13209 3375 13243
rect 3893 13209 3927 13243
rect 4353 13209 4387 13243
rect 5273 13209 5307 13243
rect 6260 13209 6294 13243
rect 6837 13209 6871 13243
rect 7113 13209 7147 13243
rect 10885 13209 10919 13243
rect 12265 13209 12299 13243
rect 12817 13209 12851 13243
rect 13461 13209 13495 13243
rect 13553 13209 13587 13243
rect 17049 13209 17083 13243
rect 17141 13209 17175 13243
rect 25513 13209 25547 13243
rect 25697 13209 25731 13243
rect 28365 13209 28399 13243
rect 28825 13209 28859 13243
rect 30757 13209 30791 13243
rect 30941 13209 30975 13243
rect 31125 13209 31159 13243
rect 31493 13209 31527 13243
rect 31677 13209 31711 13243
rect 1869 13141 1903 13175
rect 2881 13141 2915 13175
rect 3157 13141 3191 13175
rect 4445 13141 4479 13175
rect 6101 13141 6135 13175
rect 7021 13141 7055 13175
rect 8125 13141 8159 13175
rect 10149 13141 10183 13175
rect 10517 13141 10551 13175
rect 13829 13141 13863 13175
rect 14749 13141 14783 13175
rect 1685 12937 1719 12971
rect 2605 12937 2639 12971
rect 2789 12937 2823 12971
rect 3433 12937 3467 12971
rect 5089 12937 5123 12971
rect 6101 12937 6135 12971
rect 11621 12937 11655 12971
rect 13369 12937 13403 12971
rect 15485 12937 15519 12971
rect 20085 12937 20119 12971
rect 23029 12937 23063 12971
rect 23581 12937 23615 12971
rect 26065 12937 26099 12971
rect 31493 12937 31527 12971
rect 2053 12869 2087 12903
rect 5365 12869 5399 12903
rect 10241 12869 10275 12903
rect 10333 12869 10367 12903
rect 12909 12869 12943 12903
rect 13277 12869 13311 12903
rect 14013 12869 14047 12903
rect 14105 12869 14139 12903
rect 17325 12869 17359 12903
rect 17417 12869 17451 12903
rect 18337 12869 18371 12903
rect 19809 12869 19843 12903
rect 31033 12869 31067 12903
rect 1777 12801 1811 12835
rect 2973 12801 3007 12835
rect 3249 12801 3283 12835
rect 3985 12801 4019 12835
rect 4261 12801 4295 12835
rect 5825 12801 5859 12835
rect 6745 12801 6779 12835
rect 8401 12801 8435 12835
rect 8769 12801 8803 12835
rect 8953 12801 8987 12835
rect 9689 12801 9723 12835
rect 10057 12801 10091 12835
rect 10430 12801 10464 12835
rect 10793 12801 10827 12835
rect 11161 12801 11195 12835
rect 12173 12801 12207 12835
rect 12541 12801 12575 12835
rect 12725 12801 12759 12835
rect 13093 12801 13127 12835
rect 13829 12801 13863 12835
rect 14249 12801 14283 12835
rect 14565 12801 14599 12835
rect 14749 12801 14783 12835
rect 14841 12801 14875 12835
rect 14938 12801 14972 12835
rect 15301 12801 15335 12835
rect 17141 12801 17175 12835
rect 17514 12801 17548 12835
rect 18061 12801 18095 12835
rect 18245 12801 18279 12835
rect 18481 12801 18515 12835
rect 18797 12801 18831 12835
rect 18981 12801 19015 12835
rect 19073 12801 19107 12835
rect 19217 12801 19251 12835
rect 19533 12801 19567 12835
rect 19717 12801 19751 12835
rect 19901 12801 19935 12835
rect 23213 12801 23247 12835
rect 23305 12801 23339 12835
rect 23489 12801 23523 12835
rect 23857 12801 23891 12835
rect 23949 12801 23983 12835
rect 25697 12801 25731 12835
rect 25881 12801 25915 12835
rect 31309 12801 31343 12835
rect 2513 12733 2547 12767
rect 3157 12733 3191 12767
rect 4813 12733 4847 12767
rect 5917 12733 5951 12767
rect 6469 12733 6503 12767
rect 6561 12733 6595 12767
rect 6653 12733 6687 12767
rect 7941 12733 7975 12767
rect 8217 12733 8251 12767
rect 12265 12733 12299 12767
rect 31125 12733 31159 12767
rect 2053 12665 2087 12699
rect 4169 12665 4203 12699
rect 4629 12665 4663 12699
rect 4721 12665 4755 12699
rect 5365 12665 5399 12699
rect 6929 12665 6963 12699
rect 9505 12665 9539 12699
rect 15117 12665 15151 12699
rect 17693 12665 17727 12699
rect 10609 12597 10643 12631
rect 14381 12597 14415 12631
rect 18613 12597 18647 12631
rect 19349 12597 19383 12631
rect 23213 12597 23247 12631
rect 23949 12597 23983 12631
rect 25697 12597 25731 12631
rect 31033 12597 31067 12631
rect 1593 12393 1627 12427
rect 1869 12393 1903 12427
rect 5549 12393 5583 12427
rect 10241 12393 10275 12427
rect 12449 12393 12483 12427
rect 14381 12393 14415 12427
rect 17693 12393 17727 12427
rect 4721 12325 4755 12359
rect 19809 12325 19843 12359
rect 6193 12257 6227 12291
rect 7757 12257 7791 12291
rect 8677 12257 8711 12291
rect 14749 12257 14783 12291
rect 1409 12189 1443 12223
rect 1685 12189 1719 12223
rect 5181 12189 5215 12223
rect 5825 12189 5859 12223
rect 5917 12189 5951 12223
rect 7665 12189 7699 12223
rect 8033 12189 8067 12223
rect 8217 12189 8251 12223
rect 12357 12189 12391 12223
rect 14197 12189 14231 12223
rect 15117 12189 15151 12223
rect 15301 12189 15335 12223
rect 17141 12189 17175 12223
rect 17325 12189 17359 12223
rect 17514 12189 17548 12223
rect 19257 12189 19291 12223
rect 19533 12189 19567 12223
rect 19630 12189 19664 12223
rect 4721 12121 4755 12155
rect 5273 12121 5307 12155
rect 5708 12121 5742 12155
rect 10517 12121 10551 12155
rect 12725 12121 12759 12155
rect 12909 12121 12943 12155
rect 17417 12121 17451 12155
rect 19441 12121 19475 12155
rect 5457 12053 5491 12087
rect 14841 12053 14875 12087
rect 1593 11849 1627 11883
rect 1409 11713 1443 11747
<< metal1 >>
rect 1104 37562 44896 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 44896 37562
rect 1104 37488 44896 37510
rect 21910 37408 21916 37460
rect 21968 37448 21974 37460
rect 22097 37451 22155 37457
rect 22097 37448 22109 37451
rect 21968 37420 22109 37448
rect 21968 37408 21974 37420
rect 22097 37417 22109 37420
rect 22143 37417 22155 37451
rect 22097 37411 22155 37417
rect 22554 37408 22560 37460
rect 22612 37448 22618 37460
rect 22741 37451 22799 37457
rect 22741 37448 22753 37451
rect 22612 37420 22753 37448
rect 22612 37408 22618 37420
rect 22741 37417 22753 37420
rect 22787 37417 22799 37451
rect 22741 37411 22799 37417
rect 23198 37408 23204 37460
rect 23256 37448 23262 37460
rect 23385 37451 23443 37457
rect 23385 37448 23397 37451
rect 23256 37420 23397 37448
rect 23256 37408 23262 37420
rect 23385 37417 23397 37420
rect 23431 37417 23443 37451
rect 23385 37411 23443 37417
rect 25130 37408 25136 37460
rect 25188 37448 25194 37460
rect 25317 37451 25375 37457
rect 25317 37448 25329 37451
rect 25188 37420 25329 37448
rect 25188 37408 25194 37420
rect 25317 37417 25329 37420
rect 25363 37417 25375 37451
rect 25317 37411 25375 37417
rect 25774 37408 25780 37460
rect 25832 37448 25838 37460
rect 25961 37451 26019 37457
rect 25961 37448 25973 37451
rect 25832 37420 25973 37448
rect 25832 37408 25838 37420
rect 25961 37417 25973 37420
rect 26007 37417 26019 37451
rect 25961 37411 26019 37417
rect 27706 37408 27712 37460
rect 27764 37448 27770 37460
rect 27893 37451 27951 37457
rect 27893 37448 27905 37451
rect 27764 37420 27905 37448
rect 27764 37408 27770 37420
rect 27893 37417 27905 37420
rect 27939 37417 27951 37451
rect 27893 37411 27951 37417
rect 29638 37408 29644 37460
rect 29696 37448 29702 37460
rect 30193 37451 30251 37457
rect 30193 37448 30205 37451
rect 29696 37420 30205 37448
rect 29696 37408 29702 37420
rect 30193 37417 30205 37420
rect 30239 37417 30251 37451
rect 30193 37411 30251 37417
rect 31570 37408 31576 37460
rect 31628 37448 31634 37460
rect 32309 37451 32367 37457
rect 32309 37448 32321 37451
rect 31628 37420 32321 37448
rect 31628 37408 31634 37420
rect 32309 37417 32321 37420
rect 32355 37417 32367 37451
rect 32309 37411 32367 37417
rect 28994 37340 29000 37392
rect 29052 37380 29058 37392
rect 29825 37383 29883 37389
rect 29825 37380 29837 37383
rect 29052 37352 29837 37380
rect 29052 37340 29058 37352
rect 29825 37349 29837 37352
rect 29871 37349 29883 37383
rect 29825 37343 29883 37349
rect 22370 37136 22376 37188
rect 22428 37136 22434 37188
rect 23017 37179 23075 37185
rect 23017 37145 23029 37179
rect 23063 37176 23075 37179
rect 23382 37176 23388 37188
rect 23063 37148 23388 37176
rect 23063 37145 23075 37148
rect 23017 37139 23075 37145
rect 23382 37136 23388 37148
rect 23440 37136 23446 37188
rect 23658 37136 23664 37188
rect 23716 37136 23722 37188
rect 25590 37136 25596 37188
rect 25648 37136 25654 37188
rect 26237 37179 26295 37185
rect 26237 37145 26249 37179
rect 26283 37176 26295 37179
rect 27062 37176 27068 37188
rect 26283 37148 27068 37176
rect 26283 37145 26295 37148
rect 26237 37139 26295 37145
rect 27062 37136 27068 37148
rect 27120 37136 27126 37188
rect 28166 37136 28172 37188
rect 28224 37136 28230 37188
rect 29638 37136 29644 37188
rect 29696 37136 29702 37188
rect 30466 37136 30472 37188
rect 30524 37136 30530 37188
rect 32214 37136 32220 37188
rect 32272 37136 32278 37188
rect 1104 37018 44896 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 44896 37018
rect 1104 36944 44896 36966
rect 1104 36474 44896 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 44896 36474
rect 1104 36400 44896 36422
rect 1104 35930 44896 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 44896 35930
rect 1104 35856 44896 35878
rect 22370 35640 22376 35692
rect 22428 35640 22434 35692
rect 22646 35436 22652 35488
rect 22704 35476 22710 35488
rect 22925 35479 22983 35485
rect 22925 35476 22937 35479
rect 22704 35448 22937 35476
rect 22704 35436 22710 35448
rect 22925 35445 22937 35448
rect 22971 35445 22983 35479
rect 22925 35439 22983 35445
rect 1104 35386 44896 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 44896 35386
rect 1104 35312 44896 35334
rect 21821 35275 21879 35281
rect 21821 35241 21833 35275
rect 21867 35272 21879 35275
rect 22278 35272 22284 35284
rect 21867 35244 22284 35272
rect 21867 35241 21879 35244
rect 21821 35235 21879 35241
rect 22278 35232 22284 35244
rect 22336 35232 22342 35284
rect 23658 35096 23664 35148
rect 23716 35136 23722 35148
rect 24949 35139 25007 35145
rect 24949 35136 24961 35139
rect 23716 35108 24961 35136
rect 23716 35096 23722 35108
rect 24949 35105 24961 35108
rect 24995 35105 25007 35139
rect 24949 35099 25007 35105
rect 23198 35028 23204 35080
rect 23256 35028 23262 35080
rect 22956 35003 23014 35009
rect 22956 34969 22968 35003
rect 23002 35000 23014 35003
rect 23290 35000 23296 35012
rect 23002 34972 23296 35000
rect 23002 34969 23014 34972
rect 22956 34963 23014 34969
rect 23290 34960 23296 34972
rect 23348 34960 23354 35012
rect 23566 34960 23572 35012
rect 23624 35000 23630 35012
rect 26970 35000 26976 35012
rect 23624 34972 26976 35000
rect 23624 34960 23630 34972
rect 26970 34960 26976 34972
rect 27028 34960 27034 35012
rect 24118 34892 24124 34944
rect 24176 34932 24182 34944
rect 24397 34935 24455 34941
rect 24397 34932 24409 34935
rect 24176 34904 24409 34932
rect 24176 34892 24182 34904
rect 24397 34901 24409 34904
rect 24443 34901 24455 34935
rect 24397 34895 24455 34901
rect 1104 34842 44896 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 44896 34842
rect 1104 34768 44896 34790
rect 14366 34688 14372 34740
rect 14424 34728 14430 34740
rect 23566 34728 23572 34740
rect 14424 34700 23572 34728
rect 14424 34688 14430 34700
rect 23566 34688 23572 34700
rect 23624 34688 23630 34740
rect 23658 34688 23664 34740
rect 23716 34688 23722 34740
rect 25409 34731 25467 34737
rect 25409 34697 25421 34731
rect 25455 34728 25467 34731
rect 25590 34728 25596 34740
rect 25455 34700 25596 34728
rect 25455 34697 25467 34700
rect 25409 34691 25467 34697
rect 25590 34688 25596 34700
rect 25648 34688 25654 34740
rect 28166 34688 28172 34740
rect 28224 34728 28230 34740
rect 28353 34731 28411 34737
rect 28353 34728 28365 34731
rect 28224 34700 28365 34728
rect 28224 34688 28230 34700
rect 28353 34697 28365 34700
rect 28399 34728 28411 34731
rect 28399 34700 29040 34728
rect 28399 34697 28411 34700
rect 28353 34691 28411 34697
rect 23198 34660 23204 34672
rect 22296 34632 23204 34660
rect 22186 34552 22192 34604
rect 22244 34592 22250 34604
rect 22296 34601 22324 34632
rect 23198 34620 23204 34632
rect 23256 34660 23262 34672
rect 27522 34660 27528 34672
rect 23256 34632 27528 34660
rect 23256 34620 23262 34632
rect 22281 34595 22339 34601
rect 22281 34592 22293 34595
rect 22244 34564 22293 34592
rect 22244 34552 22250 34564
rect 22281 34561 22293 34564
rect 22327 34561 22339 34595
rect 22281 34555 22339 34561
rect 22548 34595 22606 34601
rect 22548 34561 22560 34595
rect 22594 34592 22606 34595
rect 23658 34592 23664 34604
rect 22594 34564 23664 34592
rect 22594 34561 22606 34564
rect 22548 34555 22606 34561
rect 23658 34552 23664 34564
rect 23716 34552 23722 34604
rect 24044 34601 24072 34632
rect 24302 34601 24308 34604
rect 24029 34595 24087 34601
rect 24029 34561 24041 34595
rect 24075 34561 24087 34595
rect 24029 34555 24087 34561
rect 24296 34555 24308 34601
rect 24302 34552 24308 34555
rect 24360 34552 24366 34604
rect 25590 34552 25596 34604
rect 25648 34592 25654 34604
rect 26988 34601 27016 34632
rect 27522 34620 27528 34632
rect 27580 34620 27586 34672
rect 26053 34595 26111 34601
rect 26053 34592 26065 34595
rect 25648 34564 26065 34592
rect 25648 34552 25654 34564
rect 26053 34561 26065 34564
rect 26099 34561 26111 34595
rect 26053 34555 26111 34561
rect 26973 34595 27031 34601
rect 26973 34561 26985 34595
rect 27019 34561 27031 34595
rect 26973 34555 27031 34561
rect 27240 34595 27298 34601
rect 27240 34561 27252 34595
rect 27286 34592 27298 34595
rect 27706 34592 27712 34604
rect 27286 34564 27712 34592
rect 27286 34561 27298 34564
rect 27240 34555 27298 34561
rect 27706 34552 27712 34564
rect 27764 34552 27770 34604
rect 29012 34601 29040 34700
rect 28997 34595 29055 34601
rect 28997 34561 29009 34595
rect 29043 34561 29055 34595
rect 28997 34555 29055 34561
rect 25498 34348 25504 34400
rect 25556 34348 25562 34400
rect 28442 34348 28448 34400
rect 28500 34348 28506 34400
rect 1104 34298 44896 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 44896 34298
rect 1104 34224 44896 34246
rect 22830 34184 22836 34196
rect 22066 34156 22836 34184
rect 16298 34008 16304 34060
rect 16356 34048 16362 34060
rect 21729 34051 21787 34057
rect 21729 34048 21741 34051
rect 16356 34020 21741 34048
rect 16356 34008 16362 34020
rect 21729 34017 21741 34020
rect 21775 34017 21787 34051
rect 21729 34011 21787 34017
rect 21821 34051 21879 34057
rect 21821 34017 21833 34051
rect 21867 34048 21879 34051
rect 22066 34048 22094 34156
rect 22830 34144 22836 34156
rect 22888 34144 22894 34196
rect 23106 34144 23112 34196
rect 23164 34144 23170 34196
rect 23198 34144 23204 34196
rect 23256 34184 23262 34196
rect 23382 34184 23388 34196
rect 23256 34156 23388 34184
rect 23256 34144 23262 34156
rect 23382 34144 23388 34156
rect 23440 34184 23446 34196
rect 23569 34187 23627 34193
rect 23569 34184 23581 34187
rect 23440 34156 23581 34184
rect 23440 34144 23446 34156
rect 23569 34153 23581 34156
rect 23615 34153 23627 34187
rect 23569 34147 23627 34153
rect 23658 34144 23664 34196
rect 23716 34144 23722 34196
rect 24118 34144 24124 34196
rect 24176 34144 24182 34196
rect 24302 34144 24308 34196
rect 24360 34184 24366 34196
rect 24397 34187 24455 34193
rect 24397 34184 24409 34187
rect 24360 34156 24409 34184
rect 24360 34144 24366 34156
rect 24397 34153 24409 34156
rect 24443 34153 24455 34187
rect 24397 34147 24455 34153
rect 27062 34144 27068 34196
rect 27120 34144 27126 34196
rect 23124 34116 23152 34144
rect 24673 34119 24731 34125
rect 24673 34116 24685 34119
rect 23124 34088 24685 34116
rect 24673 34085 24685 34088
rect 24719 34085 24731 34119
rect 24673 34079 24731 34085
rect 28905 34119 28963 34125
rect 28905 34085 28917 34119
rect 28951 34085 28963 34119
rect 28905 34079 28963 34085
rect 21867 34020 22094 34048
rect 21867 34017 21879 34020
rect 21821 34011 21879 34017
rect 22186 34008 22192 34060
rect 22244 34008 22250 34060
rect 28920 34048 28948 34079
rect 29638 34048 29644 34060
rect 23860 34020 24624 34048
rect 28920 34020 29644 34048
rect 21634 33940 21640 33992
rect 21692 33940 21698 33992
rect 21910 33940 21916 33992
rect 21968 33940 21974 33992
rect 22097 33983 22155 33989
rect 22097 33949 22109 33983
rect 22143 33980 22155 33983
rect 23382 33980 23388 33992
rect 22143 33952 23388 33980
rect 22143 33949 22155 33952
rect 22097 33943 22155 33949
rect 23382 33940 23388 33952
rect 23440 33940 23446 33992
rect 23860 33989 23888 34020
rect 24596 33992 24624 34020
rect 29638 34008 29644 34020
rect 29696 34048 29702 34060
rect 30101 34051 30159 34057
rect 30101 34048 30113 34051
rect 29696 34020 30113 34048
rect 29696 34008 29702 34020
rect 30101 34017 30113 34020
rect 30147 34017 30159 34051
rect 30101 34011 30159 34017
rect 23845 33983 23903 33989
rect 23845 33949 23857 33983
rect 23891 33949 23903 33983
rect 23845 33943 23903 33949
rect 23937 33983 23995 33989
rect 23937 33949 23949 33983
rect 23983 33949 23995 33983
rect 23937 33943 23995 33949
rect 24213 33983 24271 33989
rect 24213 33949 24225 33983
rect 24259 33982 24271 33983
rect 24259 33980 24348 33982
rect 24259 33954 24532 33980
rect 24259 33949 24271 33954
rect 24320 33952 24532 33954
rect 24213 33943 24271 33949
rect 22434 33915 22492 33921
rect 22434 33912 22446 33915
rect 22066 33884 22446 33912
rect 21453 33847 21511 33853
rect 21453 33813 21465 33847
rect 21499 33844 21511 33847
rect 22066 33844 22094 33884
rect 22434 33881 22446 33884
rect 22480 33881 22492 33915
rect 22434 33875 22492 33881
rect 23474 33872 23480 33924
rect 23532 33912 23538 33924
rect 23952 33912 23980 33943
rect 23532 33884 23980 33912
rect 23532 33872 23538 33884
rect 21499 33816 22094 33844
rect 21499 33813 21511 33816
rect 21453 33807 21511 33813
rect 22738 33804 22744 33856
rect 22796 33844 22802 33856
rect 24504 33844 24532 33952
rect 24578 33940 24584 33992
rect 24636 33940 24642 33992
rect 24762 33940 24768 33992
rect 24820 33940 24826 33992
rect 24857 33983 24915 33989
rect 24857 33949 24869 33983
rect 24903 33949 24915 33983
rect 24857 33943 24915 33949
rect 25041 33983 25099 33989
rect 25041 33949 25053 33983
rect 25087 33980 25099 33983
rect 25498 33980 25504 33992
rect 25087 33952 25504 33980
rect 25087 33949 25099 33952
rect 25041 33943 25099 33949
rect 24872 33844 24900 33943
rect 25498 33940 25504 33952
rect 25556 33940 25562 33992
rect 25685 33983 25743 33989
rect 25685 33949 25697 33983
rect 25731 33980 25743 33983
rect 27522 33980 27528 33992
rect 25731 33952 27528 33980
rect 25731 33949 25743 33952
rect 25685 33943 25743 33949
rect 27522 33940 27528 33952
rect 27580 33940 27586 33992
rect 25952 33915 26010 33921
rect 25952 33881 25964 33915
rect 25998 33912 26010 33915
rect 26142 33912 26148 33924
rect 25998 33884 26148 33912
rect 25998 33881 26010 33884
rect 25952 33875 26010 33881
rect 26142 33872 26148 33884
rect 26200 33872 26206 33924
rect 27798 33921 27804 33924
rect 27792 33875 27804 33921
rect 27798 33872 27804 33875
rect 27856 33872 27862 33924
rect 26602 33844 26608 33856
rect 22796 33816 26608 33844
rect 22796 33804 22802 33816
rect 26602 33804 26608 33816
rect 26660 33804 26666 33856
rect 28994 33804 29000 33856
rect 29052 33844 29058 33856
rect 29549 33847 29607 33853
rect 29549 33844 29561 33847
rect 29052 33816 29561 33844
rect 29052 33804 29058 33816
rect 29549 33813 29561 33816
rect 29595 33813 29607 33847
rect 29549 33807 29607 33813
rect 1104 33754 44896 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 44896 33754
rect 1104 33680 44896 33702
rect 17770 33600 17776 33652
rect 17828 33640 17834 33652
rect 23106 33640 23112 33652
rect 17828 33612 23112 33640
rect 17828 33600 17834 33612
rect 23106 33600 23112 33612
rect 23164 33600 23170 33652
rect 23290 33600 23296 33652
rect 23348 33600 23354 33652
rect 23382 33600 23388 33652
rect 23440 33600 23446 33652
rect 26142 33600 26148 33652
rect 26200 33600 26206 33652
rect 27706 33600 27712 33652
rect 27764 33600 27770 33652
rect 28813 33643 28871 33649
rect 28813 33609 28825 33643
rect 28859 33640 28871 33643
rect 30466 33640 30472 33652
rect 28859 33612 30472 33640
rect 28859 33609 28871 33612
rect 28813 33603 28871 33609
rect 30466 33600 30472 33612
rect 30524 33600 30530 33652
rect 24578 33572 24584 33584
rect 23124 33544 24584 33572
rect 22646 33464 22652 33516
rect 22704 33464 22710 33516
rect 23124 33513 23152 33544
rect 24578 33532 24584 33544
rect 24636 33572 24642 33584
rect 24636 33544 27936 33572
rect 24636 33532 24642 33544
rect 23109 33507 23167 33513
rect 23109 33504 23121 33507
rect 22756 33476 23121 33504
rect 21634 33396 21640 33448
rect 21692 33436 21698 33448
rect 22756 33436 22784 33476
rect 23109 33473 23121 33476
rect 23155 33473 23167 33507
rect 23109 33467 23167 33473
rect 23198 33464 23204 33516
rect 23256 33504 23262 33516
rect 26344 33513 26372 33544
rect 27908 33516 27936 33544
rect 23937 33507 23995 33513
rect 23937 33504 23949 33507
rect 23256 33476 23949 33504
rect 23256 33464 23262 33476
rect 23937 33473 23949 33476
rect 23983 33473 23995 33507
rect 23937 33467 23995 33473
rect 26329 33507 26387 33513
rect 26329 33473 26341 33507
rect 26375 33473 26387 33507
rect 26329 33467 26387 33473
rect 26789 33507 26847 33513
rect 26789 33473 26801 33507
rect 26835 33504 26847 33507
rect 26973 33507 27031 33513
rect 26973 33504 26985 33507
rect 26835 33476 26985 33504
rect 26835 33473 26847 33476
rect 26789 33467 26847 33473
rect 26973 33473 26985 33476
rect 27019 33473 27031 33507
rect 26973 33467 27031 33473
rect 27062 33464 27068 33516
rect 27120 33504 27126 33516
rect 27525 33507 27583 33513
rect 27525 33504 27537 33507
rect 27120 33476 27537 33504
rect 27120 33464 27126 33476
rect 27525 33473 27537 33476
rect 27571 33473 27583 33507
rect 27525 33467 27583 33473
rect 27890 33464 27896 33516
rect 27948 33464 27954 33516
rect 27982 33464 27988 33516
rect 28040 33464 28046 33516
rect 28258 33504 28264 33516
rect 28092 33476 28264 33504
rect 21692 33408 22784 33436
rect 22833 33439 22891 33445
rect 21692 33396 21698 33408
rect 22833 33405 22845 33439
rect 22879 33405 22891 33439
rect 22833 33399 22891 33405
rect 21910 33328 21916 33380
rect 21968 33368 21974 33380
rect 22738 33368 22744 33380
rect 21968 33340 22744 33368
rect 21968 33328 21974 33340
rect 22738 33328 22744 33340
rect 22796 33368 22802 33380
rect 22848 33368 22876 33399
rect 22922 33396 22928 33448
rect 22980 33396 22986 33448
rect 26510 33396 26516 33448
rect 26568 33396 26574 33448
rect 26602 33396 26608 33448
rect 26660 33436 26666 33448
rect 28092 33436 28120 33476
rect 28258 33464 28264 33476
rect 28316 33464 28322 33516
rect 29546 33464 29552 33516
rect 29604 33504 29610 33516
rect 29926 33507 29984 33513
rect 29926 33504 29938 33507
rect 29604 33476 29938 33504
rect 29604 33464 29610 33476
rect 29926 33473 29938 33476
rect 29972 33473 29984 33507
rect 29926 33467 29984 33473
rect 30466 33464 30472 33516
rect 30524 33504 30530 33516
rect 30837 33507 30895 33513
rect 30837 33504 30849 33507
rect 30524 33476 30849 33504
rect 30524 33464 30530 33476
rect 30837 33473 30849 33476
rect 30883 33473 30895 33507
rect 30837 33467 30895 33473
rect 26660 33408 28120 33436
rect 28169 33439 28227 33445
rect 26660 33396 26666 33408
rect 28169 33405 28181 33439
rect 28215 33436 28227 33439
rect 28442 33436 28448 33448
rect 28215 33408 28448 33436
rect 28215 33405 28227 33408
rect 28169 33399 28227 33405
rect 28442 33396 28448 33408
rect 28500 33396 28506 33448
rect 30193 33439 30251 33445
rect 30193 33405 30205 33439
rect 30239 33436 30251 33439
rect 30650 33436 30656 33448
rect 30239 33408 30656 33436
rect 30239 33405 30251 33408
rect 30193 33399 30251 33405
rect 30650 33396 30656 33408
rect 30708 33396 30714 33448
rect 22796 33340 22876 33368
rect 23017 33371 23075 33377
rect 22796 33328 22802 33340
rect 23017 33337 23029 33371
rect 23063 33368 23075 33371
rect 23566 33368 23572 33380
rect 23063 33340 23572 33368
rect 23063 33337 23075 33340
rect 23017 33331 23075 33337
rect 23566 33328 23572 33340
rect 23624 33328 23630 33380
rect 26421 33371 26479 33377
rect 26421 33337 26433 33371
rect 26467 33368 26479 33371
rect 27430 33368 27436 33380
rect 26467 33340 27436 33368
rect 26467 33337 26479 33340
rect 26421 33331 26479 33337
rect 27430 33328 27436 33340
rect 27488 33328 27494 33380
rect 30190 33260 30196 33312
rect 30248 33300 30254 33312
rect 30285 33303 30343 33309
rect 30285 33300 30297 33303
rect 30248 33272 30297 33300
rect 30248 33260 30254 33272
rect 30285 33269 30297 33272
rect 30331 33269 30343 33303
rect 30285 33263 30343 33269
rect 1104 33210 44896 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 44896 33210
rect 1104 33136 44896 33158
rect 27709 33099 27767 33105
rect 27709 33065 27721 33099
rect 27755 33096 27767 33099
rect 27798 33096 27804 33108
rect 27755 33068 27804 33096
rect 27755 33065 27767 33068
rect 27709 33059 27767 33065
rect 27798 33056 27804 33068
rect 27856 33056 27862 33108
rect 28169 33099 28227 33105
rect 28169 33065 28181 33099
rect 28215 33096 28227 33099
rect 28994 33096 29000 33108
rect 28215 33068 29000 33096
rect 28215 33065 28227 33068
rect 28169 33059 28227 33065
rect 28994 33056 29000 33068
rect 29052 33056 29058 33108
rect 29546 33056 29552 33108
rect 29604 33056 29610 33108
rect 31570 33096 31576 33108
rect 30024 33068 31576 33096
rect 21818 32988 21824 33040
rect 21876 33028 21882 33040
rect 21876 33000 28120 33028
rect 21876 32988 21882 33000
rect 20714 32920 20720 32972
rect 20772 32960 20778 32972
rect 23382 32960 23388 32972
rect 20772 32932 23388 32960
rect 20772 32920 20778 32932
rect 23382 32920 23388 32932
rect 23440 32920 23446 32972
rect 18414 32852 18420 32904
rect 18472 32892 18478 32904
rect 21910 32892 21916 32904
rect 18472 32864 21916 32892
rect 18472 32852 18478 32864
rect 21910 32852 21916 32864
rect 21968 32892 21974 32904
rect 27798 32892 27804 32904
rect 21968 32864 27804 32892
rect 21968 32852 21974 32864
rect 27798 32852 27804 32864
rect 27856 32852 27862 32904
rect 27890 32852 27896 32904
rect 27948 32852 27954 32904
rect 27985 32895 28043 32901
rect 27985 32861 27997 32895
rect 28031 32861 28043 32895
rect 27985 32855 28043 32861
rect 27614 32784 27620 32836
rect 27672 32824 27678 32836
rect 28000 32824 28028 32855
rect 27672 32796 28028 32824
rect 28092 32824 28120 33000
rect 28258 32988 28264 33040
rect 28316 33028 28322 33040
rect 30024 33028 30052 33068
rect 31570 33056 31576 33068
rect 31628 33056 31634 33108
rect 32033 33099 32091 33105
rect 32033 33065 32045 33099
rect 32079 33096 32091 33099
rect 32214 33096 32220 33108
rect 32079 33068 32220 33096
rect 32079 33065 32091 33068
rect 32033 33059 32091 33065
rect 32214 33056 32220 33068
rect 32272 33056 32278 33108
rect 28316 33000 30052 33028
rect 28316 32988 28322 33000
rect 30024 32969 30052 33000
rect 30009 32963 30067 32969
rect 30009 32929 30021 32963
rect 30055 32929 30067 32963
rect 32232 32960 32260 33056
rect 32677 32963 32735 32969
rect 32677 32960 32689 32963
rect 32232 32932 32689 32960
rect 30009 32923 30067 32929
rect 32677 32929 32689 32932
rect 32723 32929 32735 32963
rect 32677 32923 32735 32929
rect 28258 32852 28264 32904
rect 28316 32852 28322 32904
rect 29730 32852 29736 32904
rect 29788 32852 29794 32904
rect 29822 32852 29828 32904
rect 29880 32852 29886 32904
rect 29914 32852 29920 32904
rect 29972 32852 29978 32904
rect 30190 32852 30196 32904
rect 30248 32852 30254 32904
rect 30650 32852 30656 32904
rect 30708 32892 30714 32904
rect 30708 32864 32260 32892
rect 30708 32852 30714 32864
rect 30282 32824 30288 32836
rect 28092 32796 30288 32824
rect 27672 32784 27678 32796
rect 30282 32784 30288 32796
rect 30340 32784 30346 32836
rect 30920 32827 30978 32833
rect 30920 32793 30932 32827
rect 30966 32824 30978 32827
rect 31018 32824 31024 32836
rect 30966 32796 31024 32824
rect 30966 32793 30978 32796
rect 30920 32787 30978 32793
rect 31018 32784 31024 32796
rect 31076 32784 31082 32836
rect 32232 32824 32260 32864
rect 36078 32824 36084 32836
rect 32232 32796 36084 32824
rect 36078 32784 36084 32796
rect 36136 32784 36142 32836
rect 13722 32716 13728 32768
rect 13780 32756 13786 32768
rect 22002 32756 22008 32768
rect 13780 32728 22008 32756
rect 13780 32716 13786 32728
rect 22002 32716 22008 32728
rect 22060 32756 22066 32768
rect 26142 32756 26148 32768
rect 22060 32728 26148 32756
rect 22060 32716 22066 32728
rect 26142 32716 26148 32728
rect 26200 32716 26206 32768
rect 27890 32716 27896 32768
rect 27948 32756 27954 32768
rect 29730 32756 29736 32768
rect 27948 32728 29736 32756
rect 27948 32716 27954 32728
rect 29730 32716 29736 32728
rect 29788 32716 29794 32768
rect 32122 32716 32128 32768
rect 32180 32716 32186 32768
rect 1104 32666 44896 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 44896 32666
rect 1104 32592 44896 32614
rect 14826 32512 14832 32564
rect 14884 32552 14890 32564
rect 14884 32524 16252 32552
rect 14884 32512 14890 32524
rect 12342 32444 12348 32496
rect 12400 32484 12406 32496
rect 16117 32487 16175 32493
rect 16117 32484 16129 32487
rect 12400 32456 16129 32484
rect 12400 32444 12406 32456
rect 16117 32453 16129 32456
rect 16163 32453 16175 32487
rect 16224 32484 16252 32524
rect 19334 32512 19340 32564
rect 19392 32552 19398 32564
rect 23106 32552 23112 32564
rect 19392 32524 23112 32552
rect 19392 32512 19398 32524
rect 23106 32512 23112 32524
rect 23164 32512 23170 32564
rect 23474 32512 23480 32564
rect 23532 32512 23538 32564
rect 23566 32512 23572 32564
rect 23624 32512 23630 32564
rect 28813 32555 28871 32561
rect 28813 32521 28825 32555
rect 28859 32552 28871 32555
rect 29822 32552 29828 32564
rect 28859 32524 29828 32552
rect 28859 32521 28871 32524
rect 28813 32515 28871 32521
rect 29822 32512 29828 32524
rect 29880 32512 29886 32564
rect 31018 32512 31024 32564
rect 31076 32512 31082 32564
rect 37458 32552 37464 32564
rect 35866 32524 37464 32552
rect 16224 32456 20852 32484
rect 16117 32447 16175 32453
rect 11422 32376 11428 32428
rect 11480 32416 11486 32428
rect 13173 32419 13231 32425
rect 13173 32416 13185 32419
rect 11480 32388 13185 32416
rect 11480 32376 11486 32388
rect 13173 32385 13185 32388
rect 13219 32385 13231 32419
rect 13173 32379 13231 32385
rect 13449 32419 13507 32425
rect 13449 32385 13461 32419
rect 13495 32385 13507 32419
rect 13449 32379 13507 32385
rect 13357 32351 13415 32357
rect 13357 32317 13369 32351
rect 13403 32317 13415 32351
rect 13464 32348 13492 32379
rect 15838 32376 15844 32428
rect 15896 32376 15902 32428
rect 19058 32376 19064 32428
rect 19116 32416 19122 32428
rect 19337 32419 19395 32425
rect 19337 32416 19349 32419
rect 19116 32388 19349 32416
rect 19116 32376 19122 32388
rect 19337 32385 19349 32388
rect 19383 32385 19395 32419
rect 19337 32379 19395 32385
rect 19426 32376 19432 32428
rect 19484 32376 19490 32428
rect 13538 32348 13544 32360
rect 13464 32320 13544 32348
rect 13357 32311 13415 32317
rect 13372 32280 13400 32311
rect 13538 32308 13544 32320
rect 13596 32348 13602 32360
rect 13596 32320 15792 32348
rect 13596 32308 13602 32320
rect 15657 32283 15715 32289
rect 15657 32280 15669 32283
rect 13372 32252 15669 32280
rect 15657 32249 15669 32252
rect 15703 32249 15715 32283
rect 15764 32280 15792 32320
rect 16022 32308 16028 32360
rect 16080 32308 16086 32360
rect 16114 32308 16120 32360
rect 16172 32348 16178 32360
rect 20714 32348 20720 32360
rect 16172 32320 20720 32348
rect 16172 32308 16178 32320
rect 20714 32308 20720 32320
rect 20772 32308 20778 32360
rect 20824 32348 20852 32456
rect 21928 32456 22968 32484
rect 21818 32376 21824 32428
rect 21876 32376 21882 32428
rect 21928 32348 21956 32456
rect 22005 32419 22063 32425
rect 22005 32385 22017 32419
rect 22051 32385 22063 32419
rect 22005 32379 22063 32385
rect 20824 32320 21956 32348
rect 15764 32252 19380 32280
rect 15657 32243 15715 32249
rect 13170 32172 13176 32224
rect 13228 32172 13234 32224
rect 13630 32172 13636 32224
rect 13688 32172 13694 32224
rect 15930 32172 15936 32224
rect 15988 32172 15994 32224
rect 19352 32221 19380 32252
rect 19518 32240 19524 32292
rect 19576 32280 19582 32292
rect 22020 32280 22048 32379
rect 22940 32348 22968 32456
rect 23014 32444 23020 32496
rect 23072 32484 23078 32496
rect 29273 32487 29331 32493
rect 23072 32456 23980 32484
rect 23072 32444 23078 32456
rect 23109 32419 23167 32425
rect 23109 32385 23121 32419
rect 23155 32416 23167 32419
rect 23155 32388 23244 32416
rect 23155 32385 23167 32388
rect 23109 32379 23167 32385
rect 23216 32348 23244 32388
rect 23290 32376 23296 32428
rect 23348 32376 23354 32428
rect 23952 32425 23980 32456
rect 29273 32453 29285 32487
rect 29319 32484 29331 32487
rect 31386 32484 31392 32496
rect 29319 32456 31392 32484
rect 29319 32453 29331 32456
rect 29273 32447 29331 32453
rect 31386 32444 31392 32456
rect 31444 32444 31450 32496
rect 35866 32484 35894 32524
rect 37458 32512 37464 32524
rect 37516 32512 37522 32564
rect 31496 32456 35894 32484
rect 23937 32419 23995 32425
rect 23937 32385 23949 32419
rect 23983 32385 23995 32419
rect 26145 32419 26203 32425
rect 26145 32416 26157 32419
rect 23937 32379 23995 32385
rect 25792 32388 26157 32416
rect 23750 32348 23756 32360
rect 22940 32320 23152 32348
rect 23216 32320 23756 32348
rect 23014 32280 23020 32292
rect 19576 32252 22048 32280
rect 22112 32252 23020 32280
rect 19576 32240 19582 32252
rect 19337 32215 19395 32221
rect 19337 32181 19349 32215
rect 19383 32181 19395 32215
rect 19337 32175 19395 32181
rect 19705 32215 19763 32221
rect 19705 32181 19717 32215
rect 19751 32212 19763 32215
rect 22112 32212 22140 32252
rect 23014 32240 23020 32252
rect 23072 32240 23078 32292
rect 23124 32280 23152 32320
rect 23750 32308 23756 32320
rect 23808 32308 23814 32360
rect 23845 32351 23903 32357
rect 23845 32317 23857 32351
rect 23891 32348 23903 32351
rect 24026 32348 24032 32360
rect 23891 32320 24032 32348
rect 23891 32317 23903 32320
rect 23845 32311 23903 32317
rect 24026 32308 24032 32320
rect 24084 32308 24090 32360
rect 25792 32357 25820 32388
rect 26145 32385 26157 32388
rect 26191 32385 26203 32419
rect 26145 32379 26203 32385
rect 26421 32419 26479 32425
rect 26421 32385 26433 32419
rect 26467 32416 26479 32419
rect 26602 32416 26608 32428
rect 26467 32388 26608 32416
rect 26467 32385 26479 32388
rect 26421 32379 26479 32385
rect 26602 32376 26608 32388
rect 26660 32376 26666 32428
rect 28350 32376 28356 32428
rect 28408 32376 28414 32428
rect 28534 32376 28540 32428
rect 28592 32416 28598 32428
rect 28629 32419 28687 32425
rect 28629 32416 28641 32419
rect 28592 32388 28641 32416
rect 28592 32376 28598 32388
rect 28629 32385 28641 32388
rect 28675 32385 28687 32419
rect 28629 32379 28687 32385
rect 25777 32351 25835 32357
rect 25777 32348 25789 32351
rect 24688 32320 25789 32348
rect 24688 32280 24716 32320
rect 25777 32317 25789 32320
rect 25823 32317 25835 32351
rect 25777 32311 25835 32317
rect 26234 32308 26240 32360
rect 26292 32308 26298 32360
rect 27246 32308 27252 32360
rect 27304 32348 27310 32360
rect 28445 32351 28503 32357
rect 28445 32348 28457 32351
rect 27304 32320 28457 32348
rect 27304 32308 27310 32320
rect 28445 32317 28457 32320
rect 28491 32317 28503 32351
rect 28644 32348 28672 32379
rect 28994 32376 29000 32428
rect 29052 32416 29058 32428
rect 29089 32419 29147 32425
rect 29089 32416 29101 32419
rect 29052 32388 29101 32416
rect 29052 32376 29058 32388
rect 29089 32385 29101 32388
rect 29135 32385 29147 32419
rect 29089 32379 29147 32385
rect 29365 32419 29423 32425
rect 29365 32385 29377 32419
rect 29411 32416 29423 32419
rect 29638 32416 29644 32428
rect 29411 32388 29644 32416
rect 29411 32385 29423 32388
rect 29365 32379 29423 32385
rect 29638 32376 29644 32388
rect 29696 32376 29702 32428
rect 31205 32419 31263 32425
rect 31205 32416 31217 32419
rect 29932 32388 31217 32416
rect 29457 32351 29515 32357
rect 29457 32348 29469 32351
rect 28644 32320 29469 32348
rect 28445 32311 28503 32317
rect 29457 32317 29469 32320
rect 29503 32317 29515 32351
rect 29457 32311 29515 32317
rect 23124 32252 24716 32280
rect 25682 32240 25688 32292
rect 25740 32280 25746 32292
rect 28460 32280 28488 32311
rect 29730 32308 29736 32360
rect 29788 32348 29794 32360
rect 29932 32348 29960 32388
rect 31205 32385 31217 32388
rect 31251 32416 31263 32419
rect 31496 32416 31524 32456
rect 31251 32388 31524 32416
rect 31665 32419 31723 32425
rect 31251 32385 31263 32388
rect 31205 32379 31263 32385
rect 31665 32385 31677 32419
rect 31711 32416 31723 32419
rect 32122 32416 32128 32428
rect 31711 32388 32128 32416
rect 31711 32385 31723 32388
rect 31665 32379 31723 32385
rect 32122 32376 32128 32388
rect 32180 32376 32186 32428
rect 29788 32320 29960 32348
rect 29788 32308 29794 32320
rect 30374 32308 30380 32360
rect 30432 32348 30438 32360
rect 31389 32351 31447 32357
rect 31389 32348 31401 32351
rect 30432 32320 31401 32348
rect 30432 32308 30438 32320
rect 31389 32317 31401 32320
rect 31435 32317 31447 32351
rect 31389 32311 31447 32317
rect 31481 32351 31539 32357
rect 31481 32317 31493 32351
rect 31527 32348 31539 32351
rect 31570 32348 31576 32360
rect 31527 32320 31576 32348
rect 31527 32317 31539 32320
rect 31481 32311 31539 32317
rect 31570 32308 31576 32320
rect 31628 32348 31634 32360
rect 37090 32348 37096 32360
rect 31628 32320 37096 32348
rect 31628 32308 31634 32320
rect 37090 32308 37096 32320
rect 37148 32308 37154 32360
rect 28905 32283 28963 32289
rect 28905 32280 28917 32283
rect 25740 32252 26464 32280
rect 28460 32252 28917 32280
rect 25740 32240 25746 32252
rect 19751 32184 22140 32212
rect 22189 32215 22247 32221
rect 19751 32181 19763 32184
rect 19705 32175 19763 32181
rect 22189 32181 22201 32215
rect 22235 32212 22247 32215
rect 22278 32212 22284 32224
rect 22235 32184 22284 32212
rect 22235 32181 22247 32184
rect 22189 32175 22247 32181
rect 22278 32172 22284 32184
rect 22336 32172 22342 32224
rect 23198 32172 23204 32224
rect 23256 32172 23262 32224
rect 23934 32172 23940 32224
rect 23992 32172 23998 32224
rect 25961 32215 26019 32221
rect 25961 32181 25973 32215
rect 26007 32212 26019 32215
rect 26050 32212 26056 32224
rect 26007 32184 26056 32212
rect 26007 32181 26019 32184
rect 25961 32175 26019 32181
rect 26050 32172 26056 32184
rect 26108 32172 26114 32224
rect 26436 32221 26464 32252
rect 28905 32249 28917 32252
rect 28951 32249 28963 32283
rect 31297 32283 31355 32289
rect 28905 32243 28963 32249
rect 29380 32252 30880 32280
rect 26421 32215 26479 32221
rect 26421 32181 26433 32215
rect 26467 32212 26479 32215
rect 26513 32215 26571 32221
rect 26513 32212 26525 32215
rect 26467 32184 26525 32212
rect 26467 32181 26479 32184
rect 26421 32175 26479 32181
rect 26513 32181 26525 32184
rect 26559 32181 26571 32215
rect 26513 32175 26571 32181
rect 27798 32172 27804 32224
rect 27856 32212 27862 32224
rect 29380 32221 29408 32252
rect 28353 32215 28411 32221
rect 28353 32212 28365 32215
rect 27856 32184 28365 32212
rect 27856 32172 27862 32184
rect 28353 32181 28365 32184
rect 28399 32212 28411 32215
rect 29365 32215 29423 32221
rect 29365 32212 29377 32215
rect 28399 32184 29377 32212
rect 28399 32181 28411 32184
rect 28353 32175 28411 32181
rect 29365 32181 29377 32184
rect 29411 32181 29423 32215
rect 29365 32175 29423 32181
rect 29730 32172 29736 32224
rect 29788 32172 29794 32224
rect 30852 32212 30880 32252
rect 31297 32249 31309 32283
rect 31343 32280 31355 32283
rect 32122 32280 32128 32292
rect 31343 32252 32128 32280
rect 31343 32249 31355 32252
rect 31297 32243 31355 32249
rect 32122 32240 32128 32252
rect 32180 32240 32186 32292
rect 36354 32212 36360 32224
rect 30852 32184 36360 32212
rect 36354 32172 36360 32184
rect 36412 32172 36418 32224
rect 1104 32122 44896 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 44896 32122
rect 1104 32048 44896 32070
rect 11054 31968 11060 32020
rect 11112 31968 11118 32020
rect 11422 31968 11428 32020
rect 11480 31968 11486 32020
rect 13538 31968 13544 32020
rect 13596 31968 13602 32020
rect 17218 31968 17224 32020
rect 17276 31968 17282 32020
rect 17678 31968 17684 32020
rect 17736 31968 17742 32020
rect 19245 32011 19303 32017
rect 19245 31977 19257 32011
rect 19291 31977 19303 32011
rect 19797 32011 19855 32017
rect 19797 32008 19809 32011
rect 19245 31971 19303 31977
rect 19352 31980 19809 32008
rect 9122 31900 9128 31952
rect 9180 31940 9186 31952
rect 9180 31912 16252 31940
rect 9180 31900 9186 31912
rect 11057 31875 11115 31881
rect 11057 31841 11069 31875
rect 11103 31872 11115 31875
rect 13630 31872 13636 31884
rect 11103 31844 13636 31872
rect 11103 31841 11115 31844
rect 11057 31835 11115 31841
rect 13630 31832 13636 31844
rect 13688 31832 13694 31884
rect 7926 31764 7932 31816
rect 7984 31804 7990 31816
rect 7984 31776 10916 31804
rect 7984 31764 7990 31776
rect 10888 31736 10916 31776
rect 10962 31764 10968 31816
rect 11020 31764 11026 31816
rect 11146 31764 11152 31816
rect 11204 31804 11210 31816
rect 11241 31807 11299 31813
rect 11241 31804 11253 31807
rect 11204 31776 11253 31804
rect 11204 31764 11210 31776
rect 11241 31773 11253 31776
rect 11287 31773 11299 31807
rect 13173 31807 13231 31813
rect 13173 31804 13185 31807
rect 11241 31767 11299 31773
rect 11348 31776 13185 31804
rect 11348 31736 11376 31776
rect 13173 31773 13185 31776
rect 13219 31773 13231 31807
rect 13173 31767 13231 31773
rect 13357 31807 13415 31813
rect 13357 31773 13369 31807
rect 13403 31804 13415 31807
rect 16114 31804 16120 31816
rect 13403 31776 16120 31804
rect 13403 31773 13415 31776
rect 13357 31767 13415 31773
rect 16114 31764 16120 31776
rect 16172 31764 16178 31816
rect 16224 31804 16252 31912
rect 17034 31900 17040 31952
rect 17092 31940 17098 31952
rect 19260 31940 19288 31971
rect 17092 31912 19288 31940
rect 17092 31900 17098 31912
rect 19352 31872 19380 31980
rect 19797 31977 19809 31980
rect 19843 31977 19855 32011
rect 19797 31971 19855 31977
rect 23014 31968 23020 32020
rect 23072 31968 23078 32020
rect 23198 31968 23204 32020
rect 23256 31968 23262 32020
rect 23750 31968 23756 32020
rect 23808 31968 23814 32020
rect 23934 31968 23940 32020
rect 23992 32008 23998 32020
rect 24213 32011 24271 32017
rect 24213 32008 24225 32011
rect 23992 31980 24225 32008
rect 23992 31968 23998 31980
rect 24213 31977 24225 31980
rect 24259 31977 24271 32011
rect 24213 31971 24271 31977
rect 20165 31943 20223 31949
rect 20165 31909 20177 31943
rect 20211 31940 20223 31943
rect 24228 31940 24256 31971
rect 26050 31968 26056 32020
rect 26108 31968 26114 32020
rect 26252 31980 26464 32008
rect 26252 31940 26280 31980
rect 20211 31912 21312 31940
rect 24228 31912 26280 31940
rect 26436 31940 26464 31980
rect 26510 31968 26516 32020
rect 26568 31968 26574 32020
rect 26602 31968 26608 32020
rect 26660 31968 26666 32020
rect 34422 32008 34428 32020
rect 29840 31980 34428 32008
rect 29730 31940 29736 31952
rect 26436 31912 29736 31940
rect 20211 31909 20223 31912
rect 20165 31903 20223 31909
rect 20806 31872 20812 31884
rect 17236 31844 18920 31872
rect 17236 31813 17264 31844
rect 17221 31807 17279 31813
rect 17221 31804 17233 31807
rect 16224 31776 17233 31804
rect 17221 31773 17233 31776
rect 17267 31773 17279 31807
rect 17221 31767 17279 31773
rect 17405 31807 17463 31813
rect 17405 31773 17417 31807
rect 17451 31773 17463 31807
rect 17405 31767 17463 31773
rect 17497 31807 17555 31813
rect 17497 31773 17509 31807
rect 17543 31804 17555 31807
rect 17862 31804 17868 31816
rect 17543 31776 17868 31804
rect 17543 31773 17555 31776
rect 17497 31767 17555 31773
rect 10888 31708 11376 31736
rect 17420 31736 17448 31767
rect 17862 31764 17868 31776
rect 17920 31764 17926 31816
rect 18892 31736 18920 31844
rect 19260 31844 19380 31872
rect 19812 31844 20812 31872
rect 18966 31764 18972 31816
rect 19024 31804 19030 31816
rect 19260 31813 19288 31844
rect 19245 31807 19303 31813
rect 19245 31804 19257 31807
rect 19024 31776 19257 31804
rect 19024 31764 19030 31776
rect 19245 31773 19257 31776
rect 19291 31773 19303 31807
rect 19245 31767 19303 31773
rect 19334 31764 19340 31816
rect 19392 31804 19398 31816
rect 19812 31813 19840 31844
rect 20806 31832 20812 31844
rect 20864 31832 20870 31884
rect 21284 31872 21312 31912
rect 29730 31900 29736 31912
rect 29788 31900 29794 31952
rect 26145 31875 26203 31881
rect 26145 31872 26157 31875
rect 21284 31844 26157 31872
rect 26145 31841 26157 31844
rect 26191 31841 26203 31875
rect 26145 31835 26203 31841
rect 26418 31832 26424 31884
rect 26476 31872 26482 31884
rect 29840 31872 29868 31980
rect 34422 31968 34428 31980
rect 34480 31968 34486 32020
rect 26476 31844 29868 31872
rect 26476 31832 26482 31844
rect 30926 31832 30932 31884
rect 30984 31872 30990 31884
rect 31113 31875 31171 31881
rect 31113 31872 31125 31875
rect 30984 31844 31125 31872
rect 30984 31832 30990 31844
rect 31113 31841 31125 31844
rect 31159 31841 31171 31875
rect 31113 31835 31171 31841
rect 31386 31832 31392 31884
rect 31444 31872 31450 31884
rect 32766 31872 32772 31884
rect 31444 31844 32772 31872
rect 31444 31832 31450 31844
rect 32766 31832 32772 31844
rect 32824 31832 32830 31884
rect 19797 31807 19855 31813
rect 19392 31776 19437 31804
rect 19392 31764 19398 31776
rect 19797 31773 19809 31807
rect 19843 31773 19855 31807
rect 19797 31767 19855 31773
rect 19978 31764 19984 31816
rect 20036 31764 20042 31816
rect 21910 31764 21916 31816
rect 21968 31764 21974 31816
rect 22002 31764 22008 31816
rect 22060 31804 22066 31816
rect 22097 31807 22155 31813
rect 22097 31804 22109 31807
rect 22060 31776 22109 31804
rect 22060 31764 22066 31776
rect 22097 31773 22109 31776
rect 22143 31773 22155 31807
rect 22097 31767 22155 31773
rect 22738 31764 22744 31816
rect 22796 31804 22802 31816
rect 22833 31807 22891 31813
rect 22833 31804 22845 31807
rect 22796 31776 22845 31804
rect 22796 31764 22802 31776
rect 22833 31773 22845 31776
rect 22879 31773 22891 31807
rect 22833 31767 22891 31773
rect 23014 31764 23020 31816
rect 23072 31764 23078 31816
rect 23934 31764 23940 31816
rect 23992 31764 23998 31816
rect 24029 31807 24087 31813
rect 24029 31773 24041 31807
rect 24075 31804 24087 31807
rect 24118 31804 24124 31816
rect 24075 31776 24124 31804
rect 24075 31773 24087 31776
rect 24029 31767 24087 31773
rect 24118 31764 24124 31776
rect 24176 31764 24182 31816
rect 26329 31807 26387 31813
rect 26329 31804 26341 31807
rect 24320 31776 26341 31804
rect 19352 31736 19380 31764
rect 17420 31708 17540 31736
rect 18892 31708 19380 31736
rect 22281 31739 22339 31745
rect 17512 31680 17540 31708
rect 22281 31705 22293 31739
rect 22327 31736 22339 31739
rect 22462 31736 22468 31748
rect 22327 31708 22468 31736
rect 22327 31705 22339 31708
rect 22281 31699 22339 31705
rect 22462 31696 22468 31708
rect 22520 31696 22526 31748
rect 23474 31696 23480 31748
rect 23532 31736 23538 31748
rect 24213 31739 24271 31745
rect 24213 31736 24225 31739
rect 23532 31708 24225 31736
rect 23532 31696 23538 31708
rect 24213 31705 24225 31708
rect 24259 31705 24271 31739
rect 24213 31699 24271 31705
rect 17494 31628 17500 31680
rect 17552 31628 17558 31680
rect 19610 31628 19616 31680
rect 19668 31628 19674 31680
rect 22370 31628 22376 31680
rect 22428 31668 22434 31680
rect 24320 31668 24348 31776
rect 26329 31773 26341 31776
rect 26375 31773 26387 31807
rect 26789 31807 26847 31813
rect 26789 31804 26801 31807
rect 26329 31767 26387 31773
rect 26620 31776 26801 31804
rect 26053 31739 26111 31745
rect 26053 31705 26065 31739
rect 26099 31705 26111 31739
rect 26053 31699 26111 31705
rect 22428 31640 24348 31668
rect 26068 31668 26096 31699
rect 26142 31696 26148 31748
rect 26200 31736 26206 31748
rect 26620 31736 26648 31776
rect 26789 31773 26801 31776
rect 26835 31773 26847 31807
rect 26789 31767 26847 31773
rect 26970 31764 26976 31816
rect 27028 31764 27034 31816
rect 28810 31804 28816 31816
rect 27080 31776 28816 31804
rect 26200 31708 26648 31736
rect 26200 31696 26206 31708
rect 27080 31668 27108 31776
rect 28810 31764 28816 31776
rect 28868 31764 28874 31816
rect 29365 31807 29423 31813
rect 29365 31773 29377 31807
rect 29411 31804 29423 31807
rect 31018 31804 31024 31816
rect 29411 31776 31024 31804
rect 29411 31773 29423 31776
rect 29365 31767 29423 31773
rect 31018 31764 31024 31776
rect 31076 31764 31082 31816
rect 31297 31807 31355 31813
rect 31297 31804 31309 31807
rect 31275 31776 31309 31804
rect 31297 31773 31309 31776
rect 31343 31773 31355 31807
rect 31297 31767 31355 31773
rect 28350 31696 28356 31748
rect 28408 31736 28414 31748
rect 31312 31736 31340 31767
rect 31478 31764 31484 31816
rect 31536 31764 31542 31816
rect 33318 31736 33324 31748
rect 28408 31708 33324 31736
rect 28408 31696 28414 31708
rect 33318 31696 33324 31708
rect 33376 31696 33382 31748
rect 26068 31640 27108 31668
rect 22428 31628 22434 31640
rect 27522 31628 27528 31680
rect 27580 31668 27586 31680
rect 28074 31668 28080 31680
rect 27580 31640 28080 31668
rect 27580 31628 27586 31640
rect 28074 31628 28080 31640
rect 28132 31628 28138 31680
rect 1104 31578 44896 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 44896 31578
rect 1104 31504 44896 31526
rect 12066 31424 12072 31476
rect 12124 31464 12130 31476
rect 22186 31464 22192 31476
rect 12124 31436 14872 31464
rect 12124 31424 12130 31436
rect 11146 31356 11152 31408
rect 11204 31356 11210 31408
rect 11333 31331 11391 31337
rect 11333 31297 11345 31331
rect 11379 31328 11391 31331
rect 11379 31300 12434 31328
rect 11379 31297 11391 31300
rect 11333 31291 11391 31297
rect 12406 31260 12434 31300
rect 14550 31288 14556 31340
rect 14608 31288 14614 31340
rect 14734 31328 14740 31340
rect 14660 31300 14740 31328
rect 14660 31260 14688 31300
rect 14734 31288 14740 31300
rect 14792 31288 14798 31340
rect 14844 31337 14872 31436
rect 19628 31436 22192 31464
rect 14829 31331 14887 31337
rect 14829 31297 14841 31331
rect 14875 31297 14887 31331
rect 14829 31291 14887 31297
rect 15194 31288 15200 31340
rect 15252 31328 15258 31340
rect 15289 31331 15347 31337
rect 15289 31328 15301 31331
rect 15252 31300 15301 31328
rect 15252 31288 15258 31300
rect 15289 31297 15301 31300
rect 15335 31297 15347 31331
rect 15289 31291 15347 31297
rect 15470 31288 15476 31340
rect 15528 31288 15534 31340
rect 19628 31337 19656 31436
rect 22186 31424 22192 31436
rect 22244 31464 22250 31476
rect 22738 31464 22744 31476
rect 22244 31436 22744 31464
rect 22244 31424 22250 31436
rect 22738 31424 22744 31436
rect 22796 31424 22802 31476
rect 33597 31467 33655 31473
rect 33597 31464 33609 31467
rect 26252 31436 33609 31464
rect 20714 31356 20720 31408
rect 20772 31356 20778 31408
rect 19613 31331 19671 31337
rect 19613 31297 19625 31331
rect 19659 31297 19671 31331
rect 19613 31291 19671 31297
rect 20070 31288 20076 31340
rect 20128 31288 20134 31340
rect 20257 31331 20315 31337
rect 20257 31297 20269 31331
rect 20303 31328 20315 31331
rect 20533 31331 20591 31337
rect 20533 31328 20545 31331
rect 20303 31300 20545 31328
rect 20303 31297 20315 31300
rect 20257 31291 20315 31297
rect 20533 31297 20545 31300
rect 20579 31297 20591 31331
rect 20533 31291 20591 31297
rect 12406 31232 14688 31260
rect 16022 31220 16028 31272
rect 16080 31260 16086 31272
rect 16482 31260 16488 31272
rect 16080 31232 16488 31260
rect 16080 31220 16086 31232
rect 16482 31220 16488 31232
rect 16540 31260 16546 31272
rect 19705 31263 19763 31269
rect 19705 31260 19717 31263
rect 16540 31232 19717 31260
rect 16540 31220 16546 31232
rect 19705 31229 19717 31232
rect 19751 31229 19763 31263
rect 19705 31223 19763 31229
rect 19886 31220 19892 31272
rect 19944 31260 19950 31272
rect 20272 31260 20300 31291
rect 22278 31288 22284 31340
rect 22336 31288 22342 31340
rect 22557 31331 22615 31337
rect 22557 31297 22569 31331
rect 22603 31328 22615 31331
rect 23382 31328 23388 31340
rect 22603 31300 23388 31328
rect 22603 31297 22615 31300
rect 22557 31291 22615 31297
rect 23382 31288 23388 31300
rect 23440 31288 23446 31340
rect 23566 31288 23572 31340
rect 23624 31328 23630 31340
rect 26252 31337 26280 31436
rect 33597 31433 33609 31436
rect 33643 31464 33655 31467
rect 33778 31464 33784 31476
rect 33643 31436 33784 31464
rect 33643 31433 33655 31436
rect 33597 31427 33655 31433
rect 33778 31424 33784 31436
rect 33836 31424 33842 31476
rect 28534 31356 28540 31408
rect 28592 31356 28598 31408
rect 30282 31356 30288 31408
rect 30340 31396 30346 31408
rect 31297 31399 31355 31405
rect 31297 31396 31309 31399
rect 30340 31368 31309 31396
rect 30340 31356 30346 31368
rect 31297 31365 31309 31368
rect 31343 31365 31355 31399
rect 33965 31399 34023 31405
rect 33965 31396 33977 31399
rect 31297 31359 31355 31365
rect 32784 31368 33977 31396
rect 24397 31331 24455 31337
rect 24397 31328 24409 31331
rect 23624 31300 24409 31328
rect 23624 31288 23630 31300
rect 24397 31297 24409 31300
rect 24443 31297 24455 31331
rect 24397 31291 24455 31297
rect 24581 31331 24639 31337
rect 24581 31297 24593 31331
rect 24627 31297 24639 31331
rect 24581 31291 24639 31297
rect 26237 31331 26295 31337
rect 26237 31297 26249 31331
rect 26283 31297 26295 31331
rect 26513 31331 26571 31337
rect 26513 31328 26525 31331
rect 26237 31291 26295 31297
rect 26344 31300 26525 31328
rect 19944 31232 20300 31260
rect 20441 31263 20499 31269
rect 19944 31220 19950 31232
rect 20441 31229 20453 31263
rect 20487 31260 20499 31263
rect 20487 31232 22416 31260
rect 20487 31229 20499 31232
rect 20441 31223 20499 31229
rect 15105 31195 15163 31201
rect 15105 31192 15117 31195
rect 14844 31164 15117 31192
rect 10318 31084 10324 31136
rect 10376 31124 10382 31136
rect 14844 31133 14872 31164
rect 15105 31161 15117 31164
rect 15151 31161 15163 31195
rect 22388 31192 22416 31232
rect 22462 31220 22468 31272
rect 22520 31220 22526 31272
rect 23290 31220 23296 31272
rect 23348 31260 23354 31272
rect 24596 31260 24624 31291
rect 25958 31260 25964 31272
rect 23348 31232 25964 31260
rect 23348 31220 23354 31232
rect 25958 31220 25964 31232
rect 26016 31220 26022 31272
rect 26142 31220 26148 31272
rect 26200 31260 26206 31272
rect 26344 31260 26372 31300
rect 26513 31297 26525 31300
rect 26559 31297 26571 31331
rect 26513 31291 26571 31297
rect 28074 31288 28080 31340
rect 28132 31328 28138 31340
rect 28169 31331 28227 31337
rect 28169 31328 28181 31331
rect 28132 31300 28181 31328
rect 28132 31288 28138 31300
rect 28169 31297 28181 31300
rect 28215 31297 28227 31331
rect 28169 31291 28227 31297
rect 28350 31288 28356 31340
rect 28408 31328 28414 31340
rect 28721 31331 28779 31337
rect 28721 31328 28733 31331
rect 28408 31300 28733 31328
rect 28408 31288 28414 31300
rect 28721 31297 28733 31300
rect 28767 31297 28779 31331
rect 28721 31291 28779 31297
rect 31110 31288 31116 31340
rect 31168 31288 31174 31340
rect 31478 31288 31484 31340
rect 31536 31328 31542 31340
rect 32784 31328 32812 31368
rect 33965 31365 33977 31368
rect 34011 31396 34023 31399
rect 35621 31399 35679 31405
rect 35621 31396 35633 31399
rect 34011 31368 35633 31396
rect 34011 31365 34023 31368
rect 33965 31359 34023 31365
rect 35621 31365 35633 31368
rect 35667 31365 35679 31399
rect 35621 31359 35679 31365
rect 31536 31300 32812 31328
rect 31536 31288 31542 31300
rect 32858 31288 32864 31340
rect 32916 31288 32922 31340
rect 33134 31288 33140 31340
rect 33192 31288 33198 31340
rect 33410 31288 33416 31340
rect 33468 31328 33474 31340
rect 33781 31331 33839 31337
rect 33781 31328 33793 31331
rect 33468 31300 33793 31328
rect 33468 31288 33474 31300
rect 33781 31297 33793 31300
rect 33827 31297 33839 31331
rect 33781 31291 33839 31297
rect 34606 31288 34612 31340
rect 34664 31328 34670 31340
rect 35805 31331 35863 31337
rect 35805 31328 35817 31331
rect 34664 31300 35817 31328
rect 34664 31288 34670 31300
rect 35805 31297 35817 31300
rect 35851 31297 35863 31331
rect 35805 31291 35863 31297
rect 26200 31232 26372 31260
rect 26421 31263 26479 31269
rect 26200 31220 26206 31232
rect 26421 31229 26433 31263
rect 26467 31260 26479 31263
rect 26602 31260 26608 31272
rect 26467 31232 26608 31260
rect 26467 31229 26479 31232
rect 26421 31223 26479 31229
rect 26602 31220 26608 31232
rect 26660 31220 26666 31272
rect 26694 31220 26700 31272
rect 26752 31260 26758 31272
rect 29362 31260 29368 31272
rect 26752 31232 29368 31260
rect 26752 31220 26758 31232
rect 29362 31220 29368 31232
rect 29420 31220 29426 31272
rect 33045 31263 33103 31269
rect 33045 31229 33057 31263
rect 33091 31229 33103 31263
rect 36538 31260 36544 31272
rect 33045 31223 33103 31229
rect 33244 31232 36544 31260
rect 22388 31164 22508 31192
rect 15105 31155 15163 31161
rect 10965 31127 11023 31133
rect 10965 31124 10977 31127
rect 10376 31096 10977 31124
rect 10376 31084 10382 31096
rect 10965 31093 10977 31096
rect 11011 31093 11023 31127
rect 10965 31087 11023 31093
rect 14829 31127 14887 31133
rect 14829 31093 14841 31127
rect 14875 31093 14887 31127
rect 14829 31087 14887 31093
rect 15013 31127 15071 31133
rect 15013 31093 15025 31127
rect 15059 31124 15071 31127
rect 15286 31124 15292 31136
rect 15059 31096 15292 31124
rect 15059 31093 15071 31096
rect 15013 31087 15071 31093
rect 15286 31084 15292 31096
rect 15344 31084 15350 31136
rect 19610 31084 19616 31136
rect 19668 31084 19674 31136
rect 19978 31084 19984 31136
rect 20036 31084 20042 31136
rect 20714 31084 20720 31136
rect 20772 31124 20778 31136
rect 20809 31127 20867 31133
rect 20809 31124 20821 31127
rect 20772 31096 20821 31124
rect 20772 31084 20778 31096
rect 20809 31093 20821 31096
rect 20855 31093 20867 31127
rect 20809 31087 20867 31093
rect 22094 31084 22100 31136
rect 22152 31084 22158 31136
rect 22370 31084 22376 31136
rect 22428 31084 22434 31136
rect 22480 31124 22508 31164
rect 24688 31164 26188 31192
rect 24688 31124 24716 31164
rect 22480 31096 24716 31124
rect 24765 31127 24823 31133
rect 24765 31093 24777 31127
rect 24811 31124 24823 31127
rect 25866 31124 25872 31136
rect 24811 31096 25872 31124
rect 24811 31093 24823 31096
rect 24765 31087 24823 31093
rect 25866 31084 25872 31096
rect 25924 31084 25930 31136
rect 26050 31084 26056 31136
rect 26108 31084 26114 31136
rect 26160 31124 26188 31164
rect 26326 31152 26332 31204
rect 26384 31192 26390 31204
rect 30929 31195 30987 31201
rect 30929 31192 30941 31195
rect 26384 31164 30941 31192
rect 26384 31152 26390 31164
rect 30929 31161 30941 31164
rect 30975 31161 30987 31195
rect 30929 31155 30987 31161
rect 32950 31152 32956 31204
rect 33008 31192 33014 31204
rect 33060 31192 33088 31223
rect 33008 31164 33088 31192
rect 33008 31152 33014 31164
rect 26234 31124 26240 31136
rect 26160 31096 26240 31124
rect 26234 31084 26240 31096
rect 26292 31124 26298 31136
rect 26421 31127 26479 31133
rect 26421 31124 26433 31127
rect 26292 31096 26433 31124
rect 26292 31084 26298 31096
rect 26421 31093 26433 31096
rect 26467 31093 26479 31127
rect 26421 31087 26479 31093
rect 28902 31084 28908 31136
rect 28960 31084 28966 31136
rect 32858 31084 32864 31136
rect 32916 31124 32922 31136
rect 33137 31127 33195 31133
rect 33137 31124 33149 31127
rect 32916 31096 33149 31124
rect 32916 31084 32922 31096
rect 33137 31093 33149 31096
rect 33183 31124 33195 31127
rect 33244 31124 33272 31232
rect 36538 31220 36544 31232
rect 36596 31220 36602 31272
rect 33321 31195 33379 31201
rect 33321 31161 33333 31195
rect 33367 31192 33379 31195
rect 33594 31192 33600 31204
rect 33367 31164 33600 31192
rect 33367 31161 33379 31164
rect 33321 31155 33379 31161
rect 33594 31152 33600 31164
rect 33652 31152 33658 31204
rect 33686 31152 33692 31204
rect 33744 31192 33750 31204
rect 35437 31195 35495 31201
rect 35437 31192 35449 31195
rect 33744 31164 35449 31192
rect 33744 31152 33750 31164
rect 35437 31161 35449 31164
rect 35483 31192 35495 31195
rect 36262 31192 36268 31204
rect 35483 31164 36268 31192
rect 35483 31161 35495 31164
rect 35437 31155 35495 31161
rect 36262 31152 36268 31164
rect 36320 31152 36326 31204
rect 33183 31096 33272 31124
rect 33183 31093 33195 31096
rect 33137 31087 33195 31093
rect 33410 31084 33416 31136
rect 33468 31084 33474 31136
rect 1104 31034 44896 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 44896 31034
rect 1104 30960 44896 30982
rect 11882 30880 11888 30932
rect 11940 30920 11946 30932
rect 12161 30923 12219 30929
rect 12161 30920 12173 30923
rect 11940 30892 12173 30920
rect 11940 30880 11946 30892
rect 12161 30889 12173 30892
rect 12207 30920 12219 30923
rect 12342 30920 12348 30932
rect 12207 30892 12348 30920
rect 12207 30889 12219 30892
rect 12161 30883 12219 30889
rect 12342 30880 12348 30892
rect 12400 30880 12406 30932
rect 14550 30880 14556 30932
rect 14608 30920 14614 30932
rect 14829 30923 14887 30929
rect 14829 30920 14841 30923
rect 14608 30892 14841 30920
rect 14608 30880 14614 30892
rect 14829 30889 14841 30892
rect 14875 30889 14887 30923
rect 19518 30920 19524 30932
rect 14829 30883 14887 30889
rect 14936 30892 19524 30920
rect 12345 30787 12403 30793
rect 12345 30753 12357 30787
rect 12391 30784 12403 30787
rect 12802 30784 12808 30796
rect 12391 30756 12808 30784
rect 12391 30753 12403 30756
rect 12345 30747 12403 30753
rect 12802 30744 12808 30756
rect 12860 30784 12866 30796
rect 14936 30784 14964 30892
rect 19518 30880 19524 30892
rect 19576 30880 19582 30932
rect 22554 30880 22560 30932
rect 22612 30880 22618 30932
rect 23474 30880 23480 30932
rect 23532 30880 23538 30932
rect 23566 30880 23572 30932
rect 23624 30920 23630 30932
rect 23661 30923 23719 30929
rect 23661 30920 23673 30923
rect 23624 30892 23673 30920
rect 23624 30880 23630 30892
rect 23661 30889 23673 30892
rect 23707 30889 23719 30923
rect 23661 30883 23719 30889
rect 24486 30880 24492 30932
rect 24544 30920 24550 30932
rect 26053 30923 26111 30929
rect 26053 30920 26065 30923
rect 24544 30892 26065 30920
rect 24544 30880 24550 30892
rect 26053 30889 26065 30892
rect 26099 30889 26111 30923
rect 26053 30883 26111 30889
rect 26142 30880 26148 30932
rect 26200 30920 26206 30932
rect 26605 30923 26663 30929
rect 26605 30920 26617 30923
rect 26200 30892 26617 30920
rect 26200 30880 26206 30892
rect 26605 30889 26617 30892
rect 26651 30889 26663 30923
rect 26605 30883 26663 30889
rect 27338 30880 27344 30932
rect 27396 30880 27402 30932
rect 27709 30923 27767 30929
rect 27709 30889 27721 30923
rect 27755 30920 27767 30923
rect 27982 30920 27988 30932
rect 27755 30892 27988 30920
rect 27755 30889 27767 30892
rect 27709 30883 27767 30889
rect 27982 30880 27988 30892
rect 28040 30880 28046 30932
rect 28718 30880 28724 30932
rect 28776 30920 28782 30932
rect 32214 30920 32220 30932
rect 28776 30892 32220 30920
rect 28776 30880 28782 30892
rect 32214 30880 32220 30892
rect 32272 30920 32278 30932
rect 33042 30920 33048 30932
rect 32272 30892 33048 30920
rect 32272 30880 32278 30892
rect 33042 30880 33048 30892
rect 33100 30880 33106 30932
rect 33502 30880 33508 30932
rect 33560 30920 33566 30932
rect 33689 30923 33747 30929
rect 33689 30920 33701 30923
rect 33560 30892 33701 30920
rect 33560 30880 33566 30892
rect 33689 30889 33701 30892
rect 33735 30889 33747 30923
rect 33689 30883 33747 30889
rect 34422 30880 34428 30932
rect 34480 30920 34486 30932
rect 35713 30923 35771 30929
rect 35713 30920 35725 30923
rect 34480 30892 35725 30920
rect 34480 30880 34486 30892
rect 35713 30889 35725 30892
rect 35759 30889 35771 30923
rect 35713 30883 35771 30889
rect 36173 30923 36231 30929
rect 36173 30889 36185 30923
rect 36219 30920 36231 30923
rect 38010 30920 38016 30932
rect 36219 30892 38016 30920
rect 36219 30889 36231 30892
rect 36173 30883 36231 30889
rect 38010 30880 38016 30892
rect 38068 30880 38074 30932
rect 17678 30812 17684 30864
rect 17736 30852 17742 30864
rect 17736 30824 25636 30852
rect 17736 30812 17742 30824
rect 12860 30756 14964 30784
rect 12860 30744 12866 30756
rect 18506 30744 18512 30796
rect 18564 30784 18570 30796
rect 22373 30787 22431 30793
rect 22373 30784 22385 30787
rect 18564 30756 22385 30784
rect 18564 30744 18570 30756
rect 22373 30753 22385 30756
rect 22419 30753 22431 30787
rect 23014 30784 23020 30796
rect 22373 30747 22431 30753
rect 22572 30756 23020 30784
rect 12437 30719 12495 30725
rect 12437 30685 12449 30719
rect 12483 30716 12495 30719
rect 13354 30716 13360 30728
rect 12483 30688 13360 30716
rect 12483 30685 12495 30688
rect 12437 30679 12495 30685
rect 13354 30676 13360 30688
rect 13412 30676 13418 30728
rect 15654 30676 15660 30728
rect 15712 30716 15718 30728
rect 22572 30725 22600 30756
rect 23014 30744 23020 30756
rect 23072 30784 23078 30796
rect 23072 30756 25544 30784
rect 23072 30744 23078 30756
rect 22281 30719 22339 30725
rect 22281 30716 22293 30719
rect 15712 30688 22293 30716
rect 15712 30676 15718 30688
rect 22281 30685 22293 30688
rect 22327 30685 22339 30719
rect 22281 30679 22339 30685
rect 22557 30719 22615 30725
rect 22557 30685 22569 30719
rect 22603 30685 22615 30719
rect 22557 30679 22615 30685
rect 22738 30676 22744 30728
rect 22796 30716 22802 30728
rect 23661 30719 23719 30725
rect 23661 30716 23673 30719
rect 22796 30688 23673 30716
rect 22796 30676 22802 30688
rect 23661 30685 23673 30688
rect 23707 30685 23719 30719
rect 23661 30679 23719 30685
rect 23750 30676 23756 30728
rect 23808 30716 23814 30728
rect 24762 30716 24768 30728
rect 23808 30688 24768 30716
rect 23808 30676 23814 30688
rect 24762 30676 24768 30688
rect 24820 30676 24826 30728
rect 12066 30608 12072 30660
rect 12124 30648 12130 30660
rect 12161 30651 12219 30657
rect 12161 30648 12173 30651
rect 12124 30620 12173 30648
rect 12124 30608 12130 30620
rect 12161 30617 12173 30620
rect 12207 30617 12219 30651
rect 12161 30611 12219 30617
rect 14369 30651 14427 30657
rect 14369 30617 14381 30651
rect 14415 30648 14427 30651
rect 14458 30648 14464 30660
rect 14415 30620 14464 30648
rect 14415 30617 14427 30620
rect 14369 30611 14427 30617
rect 14458 30608 14464 30620
rect 14516 30608 14522 30660
rect 14645 30651 14703 30657
rect 14645 30617 14657 30651
rect 14691 30617 14703 30651
rect 14645 30611 14703 30617
rect 12621 30583 12679 30589
rect 12621 30549 12633 30583
rect 12667 30580 12679 30583
rect 12894 30580 12900 30592
rect 12667 30552 12900 30580
rect 12667 30549 12679 30552
rect 12621 30543 12679 30549
rect 12894 30540 12900 30552
rect 12952 30540 12958 30592
rect 13630 30540 13636 30592
rect 13688 30580 13694 30592
rect 14660 30580 14688 30611
rect 14734 30608 14740 30660
rect 14792 30648 14798 30660
rect 19794 30648 19800 30660
rect 14792 30620 19800 30648
rect 14792 30608 14798 30620
rect 19794 30608 19800 30620
rect 19852 30648 19858 30660
rect 20625 30651 20683 30657
rect 20625 30648 20637 30651
rect 19852 30620 20637 30648
rect 19852 30608 19858 30620
rect 20625 30617 20637 30620
rect 20671 30617 20683 30651
rect 20625 30611 20683 30617
rect 20809 30651 20867 30657
rect 20809 30617 20821 30651
rect 20855 30617 20867 30651
rect 20809 30611 20867 30617
rect 18230 30580 18236 30592
rect 13688 30552 18236 30580
rect 13688 30540 13694 30552
rect 18230 30540 18236 30552
rect 18288 30580 18294 30592
rect 19150 30580 19156 30592
rect 18288 30552 19156 30580
rect 18288 30540 18294 30552
rect 19150 30540 19156 30552
rect 19208 30540 19214 30592
rect 20438 30540 20444 30592
rect 20496 30580 20502 30592
rect 20824 30580 20852 30611
rect 23934 30608 23940 30660
rect 23992 30608 23998 30660
rect 25516 30648 25544 30756
rect 25608 30716 25636 30824
rect 25958 30812 25964 30864
rect 26016 30852 26022 30864
rect 28258 30852 28264 30864
rect 26016 30824 28264 30852
rect 26016 30812 26022 30824
rect 28258 30812 28264 30824
rect 28316 30812 28322 30864
rect 28537 30855 28595 30861
rect 28537 30821 28549 30855
rect 28583 30821 28595 30855
rect 28537 30815 28595 30821
rect 26602 30784 26608 30796
rect 26344 30756 26608 30784
rect 26344 30725 26372 30756
rect 26602 30744 26608 30756
rect 26660 30784 26666 30796
rect 28552 30784 28580 30815
rect 31110 30812 31116 30864
rect 31168 30852 31174 30864
rect 33134 30852 33140 30864
rect 31168 30824 33140 30852
rect 31168 30812 31174 30824
rect 33134 30812 33140 30824
rect 33192 30812 33198 30864
rect 33686 30784 33692 30796
rect 26660 30756 28580 30784
rect 28828 30756 33692 30784
rect 26660 30744 26666 30756
rect 26237 30719 26295 30725
rect 26237 30716 26249 30719
rect 25608 30688 26249 30716
rect 26237 30685 26249 30688
rect 26283 30685 26295 30719
rect 26237 30679 26295 30685
rect 26329 30719 26387 30725
rect 26329 30685 26341 30719
rect 26375 30685 26387 30719
rect 27341 30719 27399 30725
rect 27341 30716 27353 30719
rect 26329 30679 26387 30685
rect 26528 30688 27353 30716
rect 25516 30620 26004 30648
rect 20496 30552 20852 30580
rect 20993 30583 21051 30589
rect 20496 30540 20502 30552
rect 20993 30549 21005 30583
rect 21039 30580 21051 30583
rect 21818 30580 21824 30592
rect 21039 30552 21824 30580
rect 21039 30549 21051 30552
rect 20993 30543 21051 30549
rect 21818 30540 21824 30552
rect 21876 30540 21882 30592
rect 22741 30583 22799 30589
rect 22741 30549 22753 30583
rect 22787 30580 22799 30583
rect 25498 30580 25504 30592
rect 22787 30552 25504 30580
rect 22787 30549 22799 30552
rect 22741 30543 22799 30549
rect 25498 30540 25504 30552
rect 25556 30540 25562 30592
rect 25976 30580 26004 30620
rect 26050 30608 26056 30660
rect 26108 30608 26114 30660
rect 26326 30580 26332 30592
rect 25976 30552 26332 30580
rect 26326 30540 26332 30552
rect 26384 30540 26390 30592
rect 26528 30589 26556 30688
rect 27341 30685 27353 30688
rect 27387 30685 27399 30719
rect 27341 30679 27399 30685
rect 27430 30676 27436 30728
rect 27488 30676 27494 30728
rect 27982 30676 27988 30728
rect 28040 30716 28046 30728
rect 28721 30719 28779 30725
rect 28721 30716 28733 30719
rect 28040 30688 28733 30716
rect 28040 30676 28046 30688
rect 28721 30685 28733 30688
rect 28767 30685 28779 30719
rect 28721 30679 28779 30685
rect 26789 30651 26847 30657
rect 26789 30617 26801 30651
rect 26835 30617 26847 30651
rect 26789 30611 26847 30617
rect 26513 30583 26571 30589
rect 26513 30549 26525 30583
rect 26559 30549 26571 30583
rect 26804 30580 26832 30611
rect 26970 30608 26976 30660
rect 27028 30608 27034 30660
rect 27062 30608 27068 30660
rect 27120 30648 27126 30660
rect 28828 30648 28856 30756
rect 33686 30744 33692 30756
rect 33744 30744 33750 30796
rect 33778 30744 33784 30796
rect 33836 30744 33842 30796
rect 28902 30676 28908 30728
rect 28960 30716 28966 30728
rect 33226 30716 33232 30728
rect 28960 30688 33232 30716
rect 28960 30676 28966 30688
rect 33226 30676 33232 30688
rect 33284 30676 33290 30728
rect 33318 30676 33324 30728
rect 33376 30716 33382 30728
rect 33965 30719 34023 30725
rect 33965 30716 33977 30719
rect 33376 30688 33977 30716
rect 33376 30676 33382 30688
rect 33796 30660 33824 30688
rect 33965 30685 33977 30688
rect 34011 30685 34023 30719
rect 33965 30679 34023 30685
rect 34514 30676 34520 30728
rect 34572 30716 34578 30728
rect 35897 30719 35955 30725
rect 35897 30716 35909 30719
rect 34572 30688 35909 30716
rect 34572 30676 34578 30688
rect 35897 30685 35909 30688
rect 35943 30685 35955 30719
rect 35897 30679 35955 30685
rect 35986 30676 35992 30728
rect 36044 30676 36050 30728
rect 36170 30676 36176 30728
rect 36228 30676 36234 30728
rect 27120 30620 28856 30648
rect 27120 30608 27126 30620
rect 33134 30608 33140 30660
rect 33192 30648 33198 30660
rect 33192 30620 33640 30648
rect 33192 30608 33198 30620
rect 28442 30580 28448 30592
rect 26804 30552 28448 30580
rect 26513 30543 26571 30549
rect 28442 30540 28448 30552
rect 28500 30540 28506 30592
rect 29914 30540 29920 30592
rect 29972 30580 29978 30592
rect 31110 30580 31116 30592
rect 29972 30552 31116 30580
rect 29972 30540 29978 30552
rect 31110 30540 31116 30552
rect 31168 30540 31174 30592
rect 32306 30540 32312 30592
rect 32364 30580 32370 30592
rect 32766 30580 32772 30592
rect 32364 30552 32772 30580
rect 32364 30540 32370 30552
rect 32766 30540 32772 30552
rect 32824 30540 32830 30592
rect 33502 30540 33508 30592
rect 33560 30540 33566 30592
rect 33612 30580 33640 30620
rect 33686 30608 33692 30660
rect 33744 30608 33750 30660
rect 33778 30608 33784 30660
rect 33836 30608 33842 30660
rect 34790 30648 34796 30660
rect 34072 30620 34796 30648
rect 34072 30580 34100 30620
rect 34790 30608 34796 30620
rect 34848 30608 34854 30660
rect 33612 30552 34100 30580
rect 34149 30583 34207 30589
rect 34149 30549 34161 30583
rect 34195 30580 34207 30583
rect 35342 30580 35348 30592
rect 34195 30552 35348 30580
rect 34195 30549 34207 30552
rect 34149 30543 34207 30549
rect 35342 30540 35348 30552
rect 35400 30540 35406 30592
rect 1104 30490 44896 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 44896 30490
rect 1104 30416 44896 30438
rect 14458 30376 14464 30388
rect 10060 30348 14464 30376
rect 7834 30268 7840 30320
rect 7892 30308 7898 30320
rect 10060 30317 10088 30348
rect 14458 30336 14464 30348
rect 14516 30336 14522 30388
rect 18506 30336 18512 30388
rect 18564 30336 18570 30388
rect 18782 30336 18788 30388
rect 18840 30376 18846 30388
rect 22462 30376 22468 30388
rect 18840 30348 22468 30376
rect 18840 30336 18846 30348
rect 22462 30336 22468 30348
rect 22520 30336 22526 30388
rect 22554 30336 22560 30388
rect 22612 30376 22618 30388
rect 24302 30376 24308 30388
rect 22612 30348 24308 30376
rect 22612 30336 22618 30348
rect 24302 30336 24308 30348
rect 24360 30336 24366 30388
rect 24486 30336 24492 30388
rect 24544 30336 24550 30388
rect 25958 30336 25964 30388
rect 26016 30376 26022 30388
rect 33686 30376 33692 30388
rect 26016 30348 33692 30376
rect 26016 30336 26022 30348
rect 33686 30336 33692 30348
rect 33744 30336 33750 30388
rect 10045 30311 10103 30317
rect 7892 30280 9996 30308
rect 7892 30268 7898 30280
rect 9766 30200 9772 30252
rect 9824 30200 9830 30252
rect 9861 30175 9919 30181
rect 9861 30172 9873 30175
rect 9416 30144 9873 30172
rect 6546 29996 6552 30048
rect 6604 30036 6610 30048
rect 9416 30045 9444 30144
rect 9861 30141 9873 30144
rect 9907 30141 9919 30175
rect 9968 30172 9996 30280
rect 10045 30277 10057 30311
rect 10091 30277 10103 30311
rect 10045 30271 10103 30277
rect 10870 30268 10876 30320
rect 10928 30308 10934 30320
rect 15933 30311 15991 30317
rect 15933 30308 15945 30311
rect 10928 30280 15945 30308
rect 10928 30268 10934 30280
rect 15933 30277 15945 30280
rect 15979 30277 15991 30311
rect 18601 30311 18659 30317
rect 18601 30308 18613 30311
rect 15933 30271 15991 30277
rect 18524 30280 18613 30308
rect 13081 30243 13139 30249
rect 13081 30209 13093 30243
rect 13127 30240 13139 30243
rect 13127 30212 13584 30240
rect 13127 30209 13139 30212
rect 13081 30203 13139 30209
rect 11054 30172 11060 30184
rect 9968 30144 11060 30172
rect 9861 30135 9919 30141
rect 11054 30132 11060 30144
rect 11112 30172 11118 30184
rect 13173 30175 13231 30181
rect 13173 30172 13185 30175
rect 11112 30144 13185 30172
rect 11112 30132 11118 30144
rect 13173 30141 13185 30144
rect 13219 30172 13231 30175
rect 13446 30172 13452 30184
rect 13219 30144 13452 30172
rect 13219 30141 13231 30144
rect 13173 30135 13231 30141
rect 13446 30132 13452 30144
rect 13504 30132 13510 30184
rect 13556 30172 13584 30212
rect 15746 30200 15752 30252
rect 15804 30200 15810 30252
rect 15838 30200 15844 30252
rect 15896 30240 15902 30252
rect 16117 30243 16175 30249
rect 16117 30240 16129 30243
rect 15896 30212 16129 30240
rect 15896 30200 15902 30212
rect 16117 30209 16129 30212
rect 16163 30209 16175 30243
rect 16117 30203 16175 30209
rect 17221 30243 17279 30249
rect 17221 30209 17233 30243
rect 17267 30240 17279 30243
rect 17402 30240 17408 30252
rect 17267 30212 17408 30240
rect 17267 30209 17279 30212
rect 17221 30203 17279 30209
rect 13814 30172 13820 30184
rect 13556 30144 13820 30172
rect 13814 30132 13820 30144
rect 13872 30132 13878 30184
rect 17236 30172 17264 30203
rect 17402 30200 17408 30212
rect 17460 30200 17466 30252
rect 17497 30243 17555 30249
rect 17497 30209 17509 30243
rect 17543 30240 17555 30243
rect 17586 30240 17592 30252
rect 17543 30212 17592 30240
rect 17543 30209 17555 30212
rect 17497 30203 17555 30209
rect 17586 30200 17592 30212
rect 17644 30200 17650 30252
rect 18046 30200 18052 30252
rect 18104 30200 18110 30252
rect 18230 30200 18236 30252
rect 18288 30240 18294 30252
rect 18341 30243 18399 30249
rect 18341 30240 18353 30243
rect 18288 30212 18353 30240
rect 18288 30200 18294 30212
rect 18341 30209 18353 30212
rect 18387 30209 18399 30243
rect 18341 30203 18399 30209
rect 15764 30144 17264 30172
rect 15764 30116 15792 30144
rect 17310 30132 17316 30184
rect 17368 30132 17374 30184
rect 18141 30175 18199 30181
rect 18141 30172 18153 30175
rect 17604 30144 18153 30172
rect 9766 30064 9772 30116
rect 9824 30104 9830 30116
rect 10870 30104 10876 30116
rect 9824 30076 10876 30104
rect 9824 30064 9830 30076
rect 10870 30064 10876 30076
rect 10928 30064 10934 30116
rect 13722 30104 13728 30116
rect 13280 30076 13728 30104
rect 9401 30039 9459 30045
rect 9401 30036 9413 30039
rect 6604 30008 9413 30036
rect 6604 29996 6610 30008
rect 9401 30005 9413 30008
rect 9447 30005 9459 30039
rect 9401 29999 9459 30005
rect 9585 30039 9643 30045
rect 9585 30005 9597 30039
rect 9631 30036 9643 30039
rect 9674 30036 9680 30048
rect 9631 30008 9680 30036
rect 9631 30005 9643 30008
rect 9585 29999 9643 30005
rect 9674 29996 9680 30008
rect 9732 29996 9738 30048
rect 10042 29996 10048 30048
rect 10100 29996 10106 30048
rect 13280 30045 13308 30076
rect 13722 30064 13728 30076
rect 13780 30064 13786 30116
rect 15746 30064 15752 30116
rect 15804 30064 15810 30116
rect 16850 30064 16856 30116
rect 16908 30104 16914 30116
rect 17604 30104 17632 30144
rect 18141 30141 18153 30144
rect 18187 30141 18199 30175
rect 18141 30135 18199 30141
rect 16908 30076 17632 30104
rect 16908 30064 16914 30076
rect 17678 30064 17684 30116
rect 17736 30064 17742 30116
rect 18156 30104 18184 30135
rect 18524 30104 18552 30280
rect 18601 30277 18613 30280
rect 18647 30277 18659 30311
rect 18601 30271 18659 30277
rect 18690 30268 18696 30320
rect 18748 30308 18754 30320
rect 18748 30280 18920 30308
rect 18748 30268 18754 30280
rect 18782 30200 18788 30252
rect 18840 30200 18846 30252
rect 18892 30240 18920 30280
rect 18966 30268 18972 30320
rect 19024 30268 19030 30320
rect 21634 30268 21640 30320
rect 21692 30308 21698 30320
rect 23569 30311 23627 30317
rect 23569 30308 23581 30311
rect 21692 30280 23581 30308
rect 21692 30268 21698 30280
rect 23569 30277 23581 30280
rect 23615 30308 23627 30311
rect 23842 30308 23848 30320
rect 23615 30280 23848 30308
rect 23615 30277 23627 30280
rect 23569 30271 23627 30277
rect 23842 30268 23848 30280
rect 23900 30268 23906 30320
rect 23937 30311 23995 30317
rect 23937 30277 23949 30311
rect 23983 30308 23995 30311
rect 23983 30280 24164 30308
rect 23983 30277 23995 30280
rect 23937 30271 23995 30277
rect 19426 30240 19432 30252
rect 18892 30212 19432 30240
rect 19426 30200 19432 30212
rect 19484 30200 19490 30252
rect 19518 30200 19524 30252
rect 19576 30240 19582 30252
rect 19886 30240 19892 30252
rect 19576 30212 19892 30240
rect 19576 30200 19582 30212
rect 19886 30200 19892 30212
rect 19944 30200 19950 30252
rect 22646 30200 22652 30252
rect 22704 30200 22710 30252
rect 22833 30243 22891 30249
rect 22833 30209 22845 30243
rect 22879 30240 22891 30243
rect 23014 30240 23020 30252
rect 22879 30212 23020 30240
rect 22879 30209 22891 30212
rect 22833 30203 22891 30209
rect 23014 30200 23020 30212
rect 23072 30200 23078 30252
rect 23385 30243 23443 30249
rect 23385 30209 23397 30243
rect 23431 30240 23443 30243
rect 23474 30240 23480 30252
rect 23431 30212 23480 30240
rect 23431 30209 23443 30212
rect 23385 30203 23443 30209
rect 23474 30200 23480 30212
rect 23532 30200 23538 30252
rect 18874 30132 18880 30184
rect 18932 30172 18938 30184
rect 21910 30172 21916 30184
rect 18932 30144 21916 30172
rect 18932 30132 18938 30144
rect 21910 30132 21916 30144
rect 21968 30132 21974 30184
rect 23952 30172 23980 30271
rect 24026 30200 24032 30252
rect 24084 30200 24090 30252
rect 24136 30240 24164 30280
rect 24210 30268 24216 30320
rect 24268 30308 24274 30320
rect 31662 30308 31668 30320
rect 24268 30280 29500 30308
rect 24268 30268 24274 30280
rect 24305 30243 24363 30249
rect 24305 30240 24317 30243
rect 24136 30212 24317 30240
rect 24305 30209 24317 30212
rect 24351 30240 24363 30243
rect 24351 30212 26832 30240
rect 24351 30209 24363 30212
rect 24305 30203 24363 30209
rect 22204 30144 23980 30172
rect 18156 30076 18552 30104
rect 18598 30064 18604 30116
rect 18656 30104 18662 30116
rect 22204 30104 22232 30144
rect 24210 30132 24216 30184
rect 24268 30132 24274 30184
rect 23474 30104 23480 30116
rect 18656 30076 22232 30104
rect 22296 30076 23480 30104
rect 18656 30064 18662 30076
rect 13265 30039 13323 30045
rect 13265 30005 13277 30039
rect 13311 30005 13323 30039
rect 13265 29999 13323 30005
rect 13449 30039 13507 30045
rect 13449 30005 13461 30039
rect 13495 30036 13507 30039
rect 14550 30036 14556 30048
rect 13495 30008 14556 30036
rect 13495 30005 13507 30008
rect 13449 29999 13507 30005
rect 14550 29996 14556 30008
rect 14608 29996 14614 30048
rect 16022 29996 16028 30048
rect 16080 30036 16086 30048
rect 17218 30036 17224 30048
rect 16080 30008 17224 30036
rect 16080 29996 16086 30008
rect 17218 29996 17224 30008
rect 17276 29996 17282 30048
rect 17862 29996 17868 30048
rect 17920 30036 17926 30048
rect 18049 30039 18107 30045
rect 18049 30036 18061 30039
rect 17920 30008 18061 30036
rect 17920 29996 17926 30008
rect 18049 30005 18061 30008
rect 18095 30005 18107 30039
rect 18049 29999 18107 30005
rect 18138 29996 18144 30048
rect 18196 30036 18202 30048
rect 18782 30036 18788 30048
rect 18196 30008 18788 30036
rect 18196 29996 18202 30008
rect 18782 29996 18788 30008
rect 18840 29996 18846 30048
rect 19150 29996 19156 30048
rect 19208 30036 19214 30048
rect 19518 30036 19524 30048
rect 19208 30008 19524 30036
rect 19208 29996 19214 30008
rect 19518 29996 19524 30008
rect 19576 29996 19582 30048
rect 19610 29996 19616 30048
rect 19668 30036 19674 30048
rect 22296 30036 22324 30076
rect 23474 30064 23480 30076
rect 23532 30064 23538 30116
rect 23753 30107 23811 30113
rect 23753 30073 23765 30107
rect 23799 30104 23811 30107
rect 23934 30104 23940 30116
rect 23799 30076 23940 30104
rect 23799 30073 23811 30076
rect 23753 30067 23811 30073
rect 23934 30064 23940 30076
rect 23992 30104 23998 30116
rect 23992 30076 24072 30104
rect 23992 30064 23998 30076
rect 19668 30008 22324 30036
rect 19668 29996 19674 30008
rect 22370 29996 22376 30048
rect 22428 30036 22434 30048
rect 22465 30039 22523 30045
rect 22465 30036 22477 30039
rect 22428 30008 22477 30036
rect 22428 29996 22434 30008
rect 22465 30005 22477 30008
rect 22511 30036 22523 30039
rect 23382 30036 23388 30048
rect 22511 30008 23388 30036
rect 22511 30005 22523 30008
rect 22465 29999 22523 30005
rect 23382 29996 23388 30008
rect 23440 29996 23446 30048
rect 24044 30045 24072 30076
rect 24486 30064 24492 30116
rect 24544 30104 24550 30116
rect 26804 30104 26832 30212
rect 29086 30200 29092 30252
rect 29144 30200 29150 30252
rect 29362 30200 29368 30252
rect 29420 30200 29426 30252
rect 29472 30240 29500 30280
rect 31227 30280 31668 30308
rect 29917 30243 29975 30249
rect 29917 30240 29929 30243
rect 29472 30212 29929 30240
rect 29917 30209 29929 30212
rect 29963 30209 29975 30243
rect 29917 30203 29975 30209
rect 30190 30200 30196 30252
rect 30248 30200 30254 30252
rect 30374 30200 30380 30252
rect 30432 30240 30438 30252
rect 30469 30243 30527 30249
rect 30469 30240 30481 30243
rect 30432 30212 30481 30240
rect 30432 30200 30438 30212
rect 30469 30209 30481 30212
rect 30515 30209 30527 30243
rect 30469 30203 30527 30209
rect 30742 30200 30748 30252
rect 30800 30200 30806 30252
rect 31227 30249 31255 30280
rect 31662 30268 31668 30280
rect 31720 30268 31726 30320
rect 31846 30268 31852 30320
rect 31904 30308 31910 30320
rect 31904 30280 32628 30308
rect 31904 30268 31910 30280
rect 31205 30243 31263 30249
rect 31205 30209 31217 30243
rect 31251 30209 31263 30243
rect 31205 30203 31263 30209
rect 31478 30200 31484 30252
rect 31536 30200 31542 30252
rect 31754 30200 31760 30252
rect 31812 30240 31818 30252
rect 32309 30243 32367 30249
rect 32309 30240 32321 30243
rect 31812 30212 32321 30240
rect 31812 30200 31818 30212
rect 32309 30209 32321 30212
rect 32355 30240 32367 30243
rect 32398 30240 32404 30252
rect 32355 30212 32404 30240
rect 32355 30209 32367 30212
rect 32309 30203 32367 30209
rect 32398 30200 32404 30212
rect 32456 30200 32462 30252
rect 32600 30249 32628 30280
rect 33410 30268 33416 30320
rect 33468 30308 33474 30320
rect 35161 30311 35219 30317
rect 35161 30308 35173 30311
rect 33468 30280 35173 30308
rect 33468 30268 33474 30280
rect 35161 30277 35173 30280
rect 35207 30277 35219 30311
rect 35161 30271 35219 30277
rect 35345 30311 35403 30317
rect 35345 30277 35357 30311
rect 35391 30308 35403 30311
rect 35986 30308 35992 30320
rect 35391 30280 35992 30308
rect 35391 30277 35403 30280
rect 35345 30271 35403 30277
rect 35986 30268 35992 30280
rect 36044 30268 36050 30320
rect 32585 30243 32643 30249
rect 32585 30209 32597 30243
rect 32631 30209 32643 30243
rect 32585 30203 32643 30209
rect 32674 30200 32680 30252
rect 32732 30240 32738 30252
rect 34977 30243 35035 30249
rect 34977 30240 34989 30243
rect 32732 30212 34989 30240
rect 32732 30200 32738 30212
rect 34977 30209 34989 30212
rect 35023 30209 35035 30243
rect 34977 30203 35035 30209
rect 27706 30132 27712 30184
rect 27764 30172 27770 30184
rect 29270 30172 29276 30184
rect 27764 30144 29276 30172
rect 27764 30132 27770 30144
rect 29270 30132 29276 30144
rect 29328 30132 29334 30184
rect 29822 30132 29828 30184
rect 29880 30172 29886 30184
rect 30098 30172 30104 30184
rect 29880 30144 30104 30172
rect 29880 30132 29886 30144
rect 30098 30132 30104 30144
rect 30156 30132 30162 30184
rect 30558 30132 30564 30184
rect 30616 30132 30622 30184
rect 31297 30175 31355 30181
rect 31297 30172 31309 30175
rect 30944 30144 31309 30172
rect 30282 30104 30288 30116
rect 24544 30076 26372 30104
rect 26804 30076 30288 30104
rect 24544 30064 24550 30076
rect 24029 30039 24087 30045
rect 24029 30005 24041 30039
rect 24075 30005 24087 30039
rect 24029 29999 24087 30005
rect 25866 29996 25872 30048
rect 25924 30036 25930 30048
rect 26234 30036 26240 30048
rect 25924 30008 26240 30036
rect 25924 29996 25930 30008
rect 26234 29996 26240 30008
rect 26292 29996 26298 30048
rect 26344 30036 26372 30076
rect 30282 30064 30288 30076
rect 30340 30064 30346 30116
rect 30944 30113 30972 30144
rect 31297 30141 31309 30144
rect 31343 30141 31355 30175
rect 31297 30135 31355 30141
rect 32493 30175 32551 30181
rect 32493 30141 32505 30175
rect 32539 30172 32551 30175
rect 33778 30172 33784 30184
rect 32539 30144 33784 30172
rect 32539 30141 32551 30144
rect 32493 30135 32551 30141
rect 33778 30132 33784 30144
rect 33836 30132 33842 30184
rect 30377 30107 30435 30113
rect 30377 30073 30389 30107
rect 30423 30104 30435 30107
rect 30929 30107 30987 30113
rect 30423 30076 30880 30104
rect 30423 30073 30435 30076
rect 30377 30067 30435 30073
rect 29365 30039 29423 30045
rect 29365 30036 29377 30039
rect 26344 30008 29377 30036
rect 29365 30005 29377 30008
rect 29411 30036 29423 30039
rect 29454 30036 29460 30048
rect 29411 30008 29460 30036
rect 29411 30005 29423 30008
rect 29365 29999 29423 30005
rect 29454 29996 29460 30008
rect 29512 29996 29518 30048
rect 29546 29996 29552 30048
rect 29604 29996 29610 30048
rect 29914 29996 29920 30048
rect 29972 29996 29978 30048
rect 30466 29996 30472 30048
rect 30524 29996 30530 30048
rect 30852 30036 30880 30076
rect 30929 30073 30941 30107
rect 30975 30073 30987 30107
rect 30929 30067 30987 30073
rect 31021 30107 31079 30113
rect 31021 30073 31033 30107
rect 31067 30104 31079 30107
rect 31110 30104 31116 30116
rect 31067 30076 31116 30104
rect 31067 30073 31079 30076
rect 31021 30067 31079 30073
rect 31110 30064 31116 30076
rect 31168 30064 31174 30116
rect 32122 30064 32128 30116
rect 32180 30064 32186 30116
rect 31205 30039 31263 30045
rect 31205 30036 31217 30039
rect 30852 30008 31217 30036
rect 31205 30005 31217 30008
rect 31251 30005 31263 30039
rect 31205 29999 31263 30005
rect 31938 29996 31944 30048
rect 31996 30036 32002 30048
rect 32309 30039 32367 30045
rect 32309 30036 32321 30039
rect 31996 30008 32321 30036
rect 31996 29996 32002 30008
rect 32309 30005 32321 30008
rect 32355 30005 32367 30039
rect 32309 29999 32367 30005
rect 34790 29996 34796 30048
rect 34848 30036 34854 30048
rect 36998 30036 37004 30048
rect 34848 30008 37004 30036
rect 34848 29996 34854 30008
rect 36998 29996 37004 30008
rect 37056 29996 37062 30048
rect 1104 29946 44896 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 44896 29946
rect 1104 29872 44896 29894
rect 9122 29792 9128 29844
rect 9180 29792 9186 29844
rect 9950 29792 9956 29844
rect 10008 29832 10014 29844
rect 11609 29835 11667 29841
rect 11609 29832 11621 29835
rect 10008 29804 11621 29832
rect 10008 29792 10014 29804
rect 11609 29801 11621 29804
rect 11655 29801 11667 29835
rect 13630 29832 13636 29844
rect 11609 29795 11667 29801
rect 11716 29804 13636 29832
rect 9306 29696 9312 29708
rect 8956 29668 9312 29696
rect 8956 29637 8984 29668
rect 9306 29656 9312 29668
rect 9364 29656 9370 29708
rect 11146 29656 11152 29708
rect 11204 29696 11210 29708
rect 11716 29705 11744 29804
rect 13630 29792 13636 29804
rect 13688 29792 13694 29844
rect 13722 29792 13728 29844
rect 13780 29792 13786 29844
rect 14277 29835 14335 29841
rect 14277 29832 14289 29835
rect 13832 29804 14289 29832
rect 13446 29724 13452 29776
rect 13504 29764 13510 29776
rect 13832 29764 13860 29804
rect 14277 29801 14289 29804
rect 14323 29832 14335 29835
rect 16022 29832 16028 29844
rect 14323 29804 16028 29832
rect 14323 29801 14335 29804
rect 14277 29795 14335 29801
rect 16022 29792 16028 29804
rect 16080 29792 16086 29844
rect 16209 29835 16267 29841
rect 16209 29801 16221 29835
rect 16255 29801 16267 29835
rect 16758 29832 16764 29844
rect 16209 29795 16267 29801
rect 16316 29804 16764 29832
rect 13504 29736 13860 29764
rect 13909 29767 13967 29773
rect 13504 29724 13510 29736
rect 13909 29733 13921 29767
rect 13955 29733 13967 29767
rect 13909 29727 13967 29733
rect 11701 29699 11759 29705
rect 11701 29696 11713 29699
rect 11204 29668 11713 29696
rect 11204 29656 11210 29668
rect 11701 29665 11713 29668
rect 11747 29665 11759 29699
rect 13722 29696 13728 29708
rect 11701 29659 11759 29665
rect 11900 29668 13728 29696
rect 8941 29631 8999 29637
rect 8941 29597 8953 29631
rect 8987 29597 8999 29631
rect 8941 29591 8999 29597
rect 9125 29631 9183 29637
rect 9125 29597 9137 29631
rect 9171 29628 9183 29631
rect 11054 29628 11060 29640
rect 9171 29600 11060 29628
rect 9171 29597 9183 29600
rect 9125 29591 9183 29597
rect 11054 29588 11060 29600
rect 11112 29588 11118 29640
rect 11238 29588 11244 29640
rect 11296 29628 11302 29640
rect 11900 29637 11928 29668
rect 13722 29656 13728 29668
rect 13780 29656 13786 29708
rect 13924 29696 13952 29727
rect 14458 29696 14464 29708
rect 13924 29668 14464 29696
rect 14458 29656 14464 29668
rect 14516 29656 14522 29708
rect 11609 29631 11667 29637
rect 11609 29628 11621 29631
rect 11296 29600 11621 29628
rect 11296 29588 11302 29600
rect 11609 29597 11621 29600
rect 11655 29597 11667 29631
rect 11609 29591 11667 29597
rect 11885 29631 11943 29637
rect 11885 29597 11897 29631
rect 11931 29597 11943 29631
rect 11885 29591 11943 29597
rect 13541 29631 13599 29637
rect 13541 29597 13553 29631
rect 13587 29597 13599 29631
rect 13541 29591 13599 29597
rect 10686 29520 10692 29572
rect 10744 29560 10750 29572
rect 13556 29560 13584 29591
rect 13630 29588 13636 29640
rect 13688 29588 13694 29640
rect 14274 29588 14280 29640
rect 14332 29588 14338 29640
rect 14550 29588 14556 29640
rect 14608 29628 14614 29640
rect 16117 29631 16175 29637
rect 16117 29628 16129 29631
rect 14608 29600 16129 29628
rect 14608 29588 14614 29600
rect 16117 29597 16129 29600
rect 16163 29597 16175 29631
rect 16117 29591 16175 29597
rect 15194 29560 15200 29572
rect 10744 29532 15200 29560
rect 10744 29520 10750 29532
rect 15194 29520 15200 29532
rect 15252 29520 15258 29572
rect 16224 29560 16252 29795
rect 16316 29705 16344 29804
rect 16758 29792 16764 29804
rect 16816 29792 16822 29844
rect 18782 29792 18788 29844
rect 18840 29792 18846 29844
rect 19058 29792 19064 29844
rect 19116 29792 19122 29844
rect 19150 29792 19156 29844
rect 19208 29832 19214 29844
rect 19245 29835 19303 29841
rect 19245 29832 19257 29835
rect 19208 29804 19257 29832
rect 19208 29792 19214 29804
rect 19245 29801 19257 29804
rect 19291 29801 19303 29835
rect 20898 29832 20904 29844
rect 19245 29795 19303 29801
rect 19628 29804 20904 29832
rect 16577 29767 16635 29773
rect 16577 29733 16589 29767
rect 16623 29764 16635 29767
rect 19628 29764 19656 29804
rect 20898 29792 20904 29804
rect 20956 29792 20962 29844
rect 20993 29835 21051 29841
rect 20993 29801 21005 29835
rect 21039 29832 21051 29835
rect 21818 29832 21824 29844
rect 21039 29804 21824 29832
rect 21039 29801 21051 29804
rect 20993 29795 21051 29801
rect 21818 29792 21824 29804
rect 21876 29792 21882 29844
rect 21910 29792 21916 29844
rect 21968 29832 21974 29844
rect 21968 29804 26096 29832
rect 21968 29792 21974 29804
rect 16623 29736 19656 29764
rect 19705 29767 19763 29773
rect 16623 29733 16635 29736
rect 16577 29727 16635 29733
rect 19705 29733 19717 29767
rect 19751 29764 19763 29767
rect 19751 29736 20852 29764
rect 19751 29733 19763 29736
rect 19705 29727 19763 29733
rect 16301 29699 16359 29705
rect 16301 29665 16313 29699
rect 16347 29665 16359 29699
rect 16301 29659 16359 29665
rect 16758 29656 16764 29708
rect 16816 29696 16822 29708
rect 18785 29699 18843 29705
rect 18785 29696 18797 29699
rect 16816 29668 18797 29696
rect 16816 29656 16822 29668
rect 18785 29665 18797 29668
rect 18831 29696 18843 29699
rect 18831 29668 19334 29696
rect 18831 29665 18843 29668
rect 18785 29659 18843 29665
rect 16390 29588 16396 29640
rect 16448 29628 16454 29640
rect 18138 29628 18144 29640
rect 16448 29600 18144 29628
rect 16448 29588 16454 29600
rect 16574 29560 16580 29572
rect 16224 29532 16580 29560
rect 16574 29520 16580 29532
rect 16632 29520 16638 29572
rect 16758 29520 16764 29572
rect 16816 29560 16822 29572
rect 16937 29563 16995 29569
rect 16937 29560 16949 29563
rect 16816 29532 16949 29560
rect 16816 29520 16822 29532
rect 16937 29529 16949 29532
rect 16983 29529 16995 29563
rect 16937 29523 16995 29529
rect 17034 29520 17040 29572
rect 17092 29560 17098 29572
rect 17129 29563 17187 29569
rect 17129 29560 17141 29563
rect 17092 29532 17141 29560
rect 17092 29520 17098 29532
rect 17129 29529 17141 29532
rect 17175 29529 17187 29563
rect 17129 29523 17187 29529
rect 17402 29520 17408 29572
rect 17460 29560 17466 29572
rect 17972 29569 18000 29600
rect 18138 29588 18144 29600
rect 18196 29588 18202 29640
rect 18690 29628 18696 29640
rect 18748 29637 18754 29640
rect 18656 29600 18696 29628
rect 18690 29588 18696 29600
rect 18748 29591 18756 29637
rect 19306 29628 19334 29668
rect 19426 29656 19432 29708
rect 19484 29656 19490 29708
rect 20530 29696 20536 29708
rect 19536 29668 20536 29696
rect 19536 29637 19564 29668
rect 20530 29656 20536 29668
rect 20588 29656 20594 29708
rect 19521 29631 19579 29637
rect 19521 29628 19533 29631
rect 19306 29600 19533 29628
rect 19521 29597 19533 29600
rect 19567 29597 19579 29631
rect 19521 29591 19579 29597
rect 18748 29588 18754 29591
rect 19978 29588 19984 29640
rect 20036 29628 20042 29640
rect 20824 29628 20852 29736
rect 21082 29724 21088 29776
rect 21140 29764 21146 29776
rect 24486 29764 24492 29776
rect 21140 29736 24492 29764
rect 21140 29724 21146 29736
rect 24486 29724 24492 29736
rect 24544 29724 24550 29776
rect 26068 29764 26096 29804
rect 26142 29792 26148 29844
rect 26200 29792 26206 29844
rect 26878 29792 26884 29844
rect 26936 29792 26942 29844
rect 27065 29835 27123 29841
rect 27065 29801 27077 29835
rect 27111 29832 27123 29835
rect 27430 29832 27436 29844
rect 27111 29804 27436 29832
rect 27111 29801 27123 29804
rect 27065 29795 27123 29801
rect 27430 29792 27436 29804
rect 27488 29792 27494 29844
rect 28718 29792 28724 29844
rect 28776 29792 28782 29844
rect 28966 29804 29960 29832
rect 26068 29736 27936 29764
rect 20898 29656 20904 29708
rect 20956 29656 20962 29708
rect 21450 29656 21456 29708
rect 21508 29696 21514 29708
rect 24210 29696 24216 29708
rect 21508 29668 24216 29696
rect 21508 29656 21514 29668
rect 24210 29656 24216 29668
rect 24268 29656 24274 29708
rect 24394 29656 24400 29708
rect 24452 29696 24458 29708
rect 26789 29699 26847 29705
rect 24452 29668 26648 29696
rect 24452 29656 24458 29668
rect 20036 29600 20079 29628
rect 20824 29600 21036 29628
rect 20036 29588 20042 29600
rect 17773 29563 17831 29569
rect 17773 29560 17785 29563
rect 17460 29532 17785 29560
rect 17460 29520 17466 29532
rect 17773 29529 17785 29532
rect 17819 29529 17831 29563
rect 17773 29523 17831 29529
rect 17957 29563 18015 29569
rect 17957 29529 17969 29563
rect 18003 29529 18015 29563
rect 18598 29560 18604 29572
rect 17957 29523 18015 29529
rect 18064 29532 18604 29560
rect 9309 29495 9367 29501
rect 9309 29461 9321 29495
rect 9355 29492 9367 29495
rect 10778 29492 10784 29504
rect 9355 29464 10784 29492
rect 9355 29461 9367 29464
rect 9309 29455 9367 29461
rect 10778 29452 10784 29464
rect 10836 29452 10842 29504
rect 11425 29495 11483 29501
rect 11425 29461 11437 29495
rect 11471 29492 11483 29495
rect 11790 29492 11796 29504
rect 11471 29464 11796 29492
rect 11471 29461 11483 29464
rect 11425 29455 11483 29461
rect 11790 29452 11796 29464
rect 11848 29452 11854 29504
rect 14090 29452 14096 29504
rect 14148 29452 14154 29504
rect 14734 29452 14740 29504
rect 14792 29492 14798 29504
rect 18064 29492 18092 29532
rect 18598 29520 18604 29532
rect 18656 29520 18662 29572
rect 19288 29569 19294 29572
rect 19270 29563 19294 29569
rect 19270 29529 19282 29563
rect 19270 29523 19294 29529
rect 19288 29520 19294 29523
rect 19346 29520 19352 29572
rect 19794 29520 19800 29572
rect 19852 29520 19858 29572
rect 20622 29520 20628 29572
rect 20680 29560 20686 29572
rect 20809 29563 20867 29569
rect 20809 29560 20821 29563
rect 20680 29532 20821 29560
rect 20680 29520 20686 29532
rect 20809 29529 20821 29532
rect 20855 29529 20867 29563
rect 21008 29560 21036 29600
rect 21082 29588 21088 29640
rect 21140 29588 21146 29640
rect 26145 29631 26203 29637
rect 26145 29597 26157 29631
rect 26191 29597 26203 29631
rect 26145 29591 26203 29597
rect 26160 29560 26188 29591
rect 26234 29588 26240 29640
rect 26292 29588 26298 29640
rect 26510 29560 26516 29572
rect 21008 29532 25995 29560
rect 26160 29532 26516 29560
rect 20809 29523 20867 29529
rect 14792 29464 18092 29492
rect 18141 29495 18199 29501
rect 14792 29452 14798 29464
rect 18141 29461 18153 29495
rect 18187 29492 18199 29495
rect 19150 29492 19156 29504
rect 18187 29464 19156 29492
rect 18187 29461 18199 29464
rect 18141 29455 18199 29461
rect 19150 29452 19156 29464
rect 19208 29492 19214 29504
rect 19702 29492 19708 29504
rect 19208 29464 19708 29492
rect 19208 29452 19214 29464
rect 19702 29452 19708 29464
rect 19760 29452 19766 29504
rect 20162 29452 20168 29504
rect 20220 29452 20226 29504
rect 21269 29495 21327 29501
rect 21269 29461 21281 29495
rect 21315 29492 21327 29495
rect 22002 29492 22008 29504
rect 21315 29464 22008 29492
rect 21315 29461 21327 29464
rect 21269 29455 21327 29461
rect 22002 29452 22008 29464
rect 22060 29452 22066 29504
rect 22646 29452 22652 29504
rect 22704 29492 22710 29504
rect 23014 29492 23020 29504
rect 22704 29464 23020 29492
rect 22704 29452 22710 29464
rect 23014 29452 23020 29464
rect 23072 29452 23078 29504
rect 23198 29452 23204 29504
rect 23256 29492 23262 29504
rect 24394 29492 24400 29504
rect 23256 29464 24400 29492
rect 23256 29452 23262 29464
rect 24394 29452 24400 29464
rect 24452 29452 24458 29504
rect 25866 29452 25872 29504
rect 25924 29452 25930 29504
rect 25967 29492 25995 29532
rect 26510 29520 26516 29532
rect 26568 29520 26574 29572
rect 26620 29560 26648 29668
rect 26789 29665 26801 29699
rect 26835 29696 26847 29699
rect 27706 29696 27712 29708
rect 26835 29668 27712 29696
rect 26835 29665 26847 29668
rect 26789 29659 26847 29665
rect 27706 29656 27712 29668
rect 27764 29656 27770 29708
rect 27908 29696 27936 29736
rect 27982 29724 27988 29776
rect 28040 29764 28046 29776
rect 28966 29764 28994 29804
rect 28040 29736 28994 29764
rect 28040 29724 28046 29736
rect 29086 29724 29092 29776
rect 29144 29724 29150 29776
rect 29178 29724 29184 29776
rect 29236 29764 29242 29776
rect 29730 29764 29736 29776
rect 29236 29736 29736 29764
rect 29236 29724 29242 29736
rect 29730 29724 29736 29736
rect 29788 29724 29794 29776
rect 29932 29764 29960 29804
rect 30006 29792 30012 29844
rect 30064 29792 30070 29844
rect 30374 29792 30380 29844
rect 30432 29792 30438 29844
rect 31662 29832 31668 29844
rect 30484 29804 31668 29832
rect 30484 29764 30512 29804
rect 31662 29792 31668 29804
rect 31720 29792 31726 29844
rect 31757 29835 31815 29841
rect 31757 29801 31769 29835
rect 31803 29801 31815 29835
rect 31757 29795 31815 29801
rect 29932 29736 30512 29764
rect 30558 29724 30564 29776
rect 30616 29764 30622 29776
rect 31772 29764 31800 29795
rect 31846 29792 31852 29844
rect 31904 29832 31910 29844
rect 32125 29835 32183 29841
rect 32125 29832 32137 29835
rect 31904 29804 32137 29832
rect 31904 29792 31910 29804
rect 32125 29801 32137 29804
rect 32171 29801 32183 29835
rect 32125 29795 32183 29801
rect 33962 29792 33968 29844
rect 34020 29832 34026 29844
rect 35161 29835 35219 29841
rect 35161 29832 35173 29835
rect 34020 29804 35173 29832
rect 34020 29792 34026 29804
rect 35161 29801 35173 29804
rect 35207 29801 35219 29835
rect 35161 29795 35219 29801
rect 32030 29764 32036 29776
rect 30616 29736 31800 29764
rect 31864 29736 32036 29764
rect 30616 29724 30622 29736
rect 28721 29699 28779 29705
rect 28721 29696 28733 29699
rect 27908 29668 28733 29696
rect 28721 29665 28733 29668
rect 28767 29696 28779 29699
rect 29822 29696 29828 29708
rect 28767 29668 29828 29696
rect 28767 29665 28779 29668
rect 28721 29659 28779 29665
rect 29822 29656 29828 29668
rect 29880 29656 29886 29708
rect 30374 29696 30380 29708
rect 29932 29668 30380 29696
rect 26694 29588 26700 29640
rect 26752 29588 26758 29640
rect 28905 29631 28963 29637
rect 28905 29597 28917 29631
rect 28951 29628 28963 29631
rect 29932 29628 29960 29668
rect 30374 29656 30380 29668
rect 30432 29696 30438 29708
rect 31386 29696 31392 29708
rect 30432 29668 31392 29696
rect 30432 29656 30438 29668
rect 31386 29656 31392 29668
rect 31444 29656 31450 29708
rect 31757 29699 31815 29705
rect 31757 29665 31769 29699
rect 31803 29696 31815 29699
rect 31864 29696 31892 29736
rect 32030 29724 32036 29736
rect 32088 29724 32094 29776
rect 32398 29724 32404 29776
rect 32456 29764 32462 29776
rect 32677 29767 32735 29773
rect 32677 29764 32689 29767
rect 32456 29736 32689 29764
rect 32456 29724 32462 29736
rect 32677 29733 32689 29736
rect 32723 29764 32735 29767
rect 38378 29764 38384 29776
rect 32723 29736 38384 29764
rect 32723 29733 32735 29736
rect 32677 29727 32735 29733
rect 38378 29724 38384 29736
rect 38436 29724 38442 29776
rect 35986 29696 35992 29708
rect 31803 29668 31892 29696
rect 35176 29668 35992 29696
rect 31803 29665 31815 29668
rect 31757 29659 31815 29665
rect 28951 29600 29960 29628
rect 30009 29631 30067 29637
rect 28951 29597 28963 29600
rect 28905 29591 28963 29597
rect 30009 29597 30021 29631
rect 30055 29628 30067 29631
rect 30193 29631 30251 29637
rect 30055 29600 30144 29628
rect 30055 29597 30067 29600
rect 30009 29591 30067 29597
rect 28350 29560 28356 29572
rect 26620 29532 28356 29560
rect 28350 29520 28356 29532
rect 28408 29520 28414 29572
rect 28626 29520 28632 29572
rect 28684 29560 28690 29572
rect 29546 29560 29552 29572
rect 28684 29532 29552 29560
rect 28684 29520 28690 29532
rect 29546 29520 29552 29532
rect 29604 29520 29610 29572
rect 30116 29560 30144 29600
rect 30193 29597 30205 29631
rect 30239 29628 30251 29631
rect 31110 29628 31116 29640
rect 30239 29600 31116 29628
rect 30239 29597 30251 29600
rect 30193 29591 30251 29597
rect 31110 29588 31116 29600
rect 31168 29588 31174 29640
rect 31662 29588 31668 29640
rect 31720 29637 31726 29640
rect 31720 29628 31730 29637
rect 31981 29631 32039 29637
rect 31720 29600 31765 29628
rect 31720 29591 31730 29600
rect 31981 29597 31993 29631
rect 32027 29628 32039 29631
rect 32122 29628 32128 29640
rect 32027 29600 32128 29628
rect 32027 29597 32039 29600
rect 31981 29591 32039 29597
rect 31720 29588 31726 29591
rect 32122 29588 32128 29600
rect 32180 29588 32186 29640
rect 32309 29631 32367 29637
rect 32309 29597 32321 29631
rect 32355 29628 32367 29631
rect 32674 29628 32680 29640
rect 32355 29600 32680 29628
rect 32355 29597 32367 29600
rect 32309 29591 32367 29597
rect 32324 29560 32352 29591
rect 32674 29588 32680 29600
rect 32732 29588 32738 29640
rect 35176 29637 35204 29668
rect 35986 29656 35992 29668
rect 36044 29656 36050 29708
rect 35161 29631 35219 29637
rect 35161 29597 35173 29631
rect 35207 29597 35219 29631
rect 35161 29591 35219 29597
rect 35253 29631 35311 29637
rect 35253 29597 35265 29631
rect 35299 29597 35311 29631
rect 35253 29591 35311 29597
rect 29656 29532 30144 29560
rect 31588 29532 32352 29560
rect 29656 29492 29684 29532
rect 25967 29464 29684 29492
rect 30098 29452 30104 29504
rect 30156 29492 30162 29504
rect 30558 29492 30564 29504
rect 30156 29464 30564 29492
rect 30156 29452 30162 29464
rect 30558 29452 30564 29464
rect 30616 29452 30622 29504
rect 30650 29452 30656 29504
rect 30708 29492 30714 29504
rect 31588 29492 31616 29532
rect 32490 29520 32496 29572
rect 32548 29520 32554 29572
rect 34698 29520 34704 29572
rect 34756 29560 34762 29572
rect 35268 29560 35296 29591
rect 36078 29588 36084 29640
rect 36136 29588 36142 29640
rect 44542 29588 44548 29640
rect 44600 29588 44606 29640
rect 37642 29560 37648 29572
rect 34756 29532 35296 29560
rect 35360 29532 37648 29560
rect 34756 29520 34762 29532
rect 30708 29464 31616 29492
rect 30708 29452 30714 29464
rect 32030 29452 32036 29504
rect 32088 29492 32094 29504
rect 35360 29492 35388 29532
rect 37642 29520 37648 29532
rect 37700 29520 37706 29572
rect 32088 29464 35388 29492
rect 32088 29452 32094 29464
rect 35434 29452 35440 29504
rect 35492 29492 35498 29504
rect 35529 29495 35587 29501
rect 35529 29492 35541 29495
rect 35492 29464 35541 29492
rect 35492 29452 35498 29464
rect 35529 29461 35541 29464
rect 35575 29461 35587 29495
rect 35529 29455 35587 29461
rect 42794 29452 42800 29504
rect 42852 29492 42858 29504
rect 44361 29495 44419 29501
rect 44361 29492 44373 29495
rect 42852 29464 44373 29492
rect 42852 29452 42858 29464
rect 44361 29461 44373 29464
rect 44407 29461 44419 29495
rect 44361 29455 44419 29461
rect 1104 29402 44896 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 44896 29402
rect 1104 29328 44896 29350
rect 7650 29248 7656 29300
rect 7708 29248 7714 29300
rect 9306 29248 9312 29300
rect 9364 29288 9370 29300
rect 9364 29260 11836 29288
rect 9364 29248 9370 29260
rect 7193 29223 7251 29229
rect 7193 29189 7205 29223
rect 7239 29220 7251 29223
rect 8938 29220 8944 29232
rect 7239 29192 8944 29220
rect 7239 29189 7251 29192
rect 7193 29183 7251 29189
rect 8938 29180 8944 29192
rect 8996 29180 9002 29232
rect 10502 29180 10508 29232
rect 10560 29180 10566 29232
rect 11808 29220 11836 29260
rect 11974 29248 11980 29300
rect 12032 29248 12038 29300
rect 12897 29291 12955 29297
rect 12897 29257 12909 29291
rect 12943 29288 12955 29291
rect 12986 29288 12992 29300
rect 12943 29260 12992 29288
rect 12943 29257 12955 29260
rect 12897 29251 12955 29257
rect 12986 29248 12992 29260
rect 13044 29248 13050 29300
rect 17586 29248 17592 29300
rect 17644 29248 17650 29300
rect 19426 29248 19432 29300
rect 19484 29288 19490 29300
rect 19978 29288 19984 29300
rect 19484 29260 19984 29288
rect 19484 29248 19490 29260
rect 19978 29248 19984 29260
rect 20036 29248 20042 29300
rect 21744 29260 22094 29288
rect 17034 29220 17040 29232
rect 11808 29192 17040 29220
rect 17034 29180 17040 29192
rect 17092 29180 17098 29232
rect 17126 29180 17132 29232
rect 17184 29220 17190 29232
rect 17402 29220 17408 29232
rect 17184 29192 17408 29220
rect 17184 29180 17190 29192
rect 17402 29180 17408 29192
rect 17460 29180 17466 29232
rect 18046 29180 18052 29232
rect 18104 29220 18110 29232
rect 21744 29220 21772 29260
rect 18104 29192 21772 29220
rect 18104 29180 18110 29192
rect 21818 29180 21824 29232
rect 21876 29180 21882 29232
rect 22066 29220 22094 29260
rect 23842 29248 23848 29300
rect 23900 29288 23906 29300
rect 23900 29260 28120 29288
rect 23900 29248 23906 29260
rect 22373 29223 22431 29229
rect 22373 29220 22385 29223
rect 22066 29192 22385 29220
rect 22373 29189 22385 29192
rect 22419 29220 22431 29223
rect 22738 29220 22744 29232
rect 22419 29192 22744 29220
rect 22419 29189 22431 29192
rect 22373 29183 22431 29189
rect 22738 29180 22744 29192
rect 22796 29180 22802 29232
rect 24581 29223 24639 29229
rect 24581 29189 24593 29223
rect 24627 29220 24639 29223
rect 25866 29220 25872 29232
rect 24627 29192 25872 29220
rect 24627 29189 24639 29192
rect 24581 29183 24639 29189
rect 25866 29180 25872 29192
rect 25924 29180 25930 29232
rect 27982 29220 27988 29232
rect 26436 29192 27988 29220
rect 6914 29112 6920 29164
rect 6972 29152 6978 29164
rect 7469 29155 7527 29161
rect 7469 29152 7481 29155
rect 6972 29124 7481 29152
rect 6972 29112 6978 29124
rect 7469 29121 7481 29124
rect 7515 29121 7527 29155
rect 7469 29115 7527 29121
rect 10226 29112 10232 29164
rect 10284 29152 10290 29164
rect 10781 29155 10839 29161
rect 10781 29152 10793 29155
rect 10284 29124 10793 29152
rect 10284 29112 10290 29124
rect 10781 29121 10793 29124
rect 10827 29121 10839 29155
rect 10781 29115 10839 29121
rect 11422 29112 11428 29164
rect 11480 29152 11486 29164
rect 11517 29155 11575 29161
rect 11517 29152 11529 29155
rect 11480 29124 11529 29152
rect 11480 29112 11486 29124
rect 11517 29121 11529 29124
rect 11563 29121 11575 29155
rect 11517 29115 11575 29121
rect 11790 29112 11796 29164
rect 11848 29112 11854 29164
rect 12986 29112 12992 29164
rect 13044 29152 13050 29164
rect 13081 29155 13139 29161
rect 13081 29152 13093 29155
rect 13044 29124 13093 29152
rect 13044 29112 13050 29124
rect 13081 29121 13093 29124
rect 13127 29121 13139 29155
rect 13081 29115 13139 29121
rect 13357 29155 13415 29161
rect 13357 29121 13369 29155
rect 13403 29152 13415 29155
rect 13538 29152 13544 29164
rect 13403 29124 13544 29152
rect 13403 29121 13415 29124
rect 13357 29115 13415 29121
rect 13538 29112 13544 29124
rect 13596 29112 13602 29164
rect 13630 29112 13636 29164
rect 13688 29152 13694 29164
rect 13688 29124 16712 29152
rect 13688 29112 13694 29124
rect 7374 29044 7380 29096
rect 7432 29044 7438 29096
rect 10686 29044 10692 29096
rect 10744 29044 10750 29096
rect 11054 29044 11060 29096
rect 11112 29084 11118 29096
rect 11609 29087 11667 29093
rect 11609 29084 11621 29087
rect 11112 29056 11621 29084
rect 11112 29044 11118 29056
rect 11609 29053 11621 29056
rect 11655 29053 11667 29087
rect 11609 29047 11667 29053
rect 13262 29044 13268 29096
rect 13320 29044 13326 29096
rect 13722 29044 13728 29096
rect 13780 29084 13786 29096
rect 16684 29084 16712 29124
rect 16942 29112 16948 29164
rect 17000 29152 17006 29164
rect 17221 29155 17279 29161
rect 17221 29152 17233 29155
rect 17000 29124 17233 29152
rect 17000 29112 17006 29124
rect 17221 29121 17233 29124
rect 17267 29121 17279 29155
rect 17221 29115 17279 29121
rect 18138 29112 18144 29164
rect 18196 29152 18202 29164
rect 19061 29155 19119 29161
rect 19061 29152 19073 29155
rect 18196 29124 19073 29152
rect 18196 29112 18202 29124
rect 19061 29121 19073 29124
rect 19107 29121 19119 29155
rect 19061 29115 19119 29121
rect 19242 29112 19248 29164
rect 19300 29112 19306 29164
rect 19337 29155 19395 29161
rect 19337 29121 19349 29155
rect 19383 29152 19395 29155
rect 19426 29152 19432 29164
rect 19383 29124 19432 29152
rect 19383 29121 19395 29124
rect 19337 29115 19395 29121
rect 19426 29112 19432 29124
rect 19484 29112 19490 29164
rect 22097 29155 22155 29161
rect 22097 29121 22109 29155
rect 22143 29152 22155 29155
rect 22186 29152 22192 29164
rect 22143 29124 22192 29152
rect 22143 29121 22155 29124
rect 22097 29115 22155 29121
rect 22186 29112 22192 29124
rect 22244 29112 22250 29164
rect 22557 29155 22615 29161
rect 22557 29121 22569 29155
rect 22603 29152 22615 29155
rect 23290 29152 23296 29164
rect 22603 29124 23296 29152
rect 22603 29121 22615 29124
rect 22557 29115 22615 29121
rect 23290 29112 23296 29124
rect 23348 29112 23354 29164
rect 23474 29112 23480 29164
rect 23532 29152 23538 29164
rect 23532 29124 24808 29152
rect 23532 29112 23538 29124
rect 21634 29084 21640 29096
rect 13780 29056 16528 29084
rect 16684 29056 21640 29084
rect 13780 29044 13786 29056
rect 10965 29019 11023 29025
rect 10965 28985 10977 29019
rect 11011 29016 11023 29019
rect 11011 28988 11652 29016
rect 11011 28985 11023 28988
rect 10965 28979 11023 28985
rect 7190 28908 7196 28960
rect 7248 28948 7254 28960
rect 9674 28948 9680 28960
rect 7248 28920 9680 28948
rect 7248 28908 7254 28920
rect 9674 28908 9680 28920
rect 9732 28908 9738 28960
rect 10686 28908 10692 28960
rect 10744 28908 10750 28960
rect 11624 28957 11652 28988
rect 11698 28976 11704 29028
rect 11756 29016 11762 29028
rect 16390 29016 16396 29028
rect 11756 28988 16396 29016
rect 11756 28976 11762 28988
rect 16390 28976 16396 28988
rect 16448 28976 16454 29028
rect 16500 29016 16528 29056
rect 21634 29044 21640 29056
rect 21692 29044 21698 29096
rect 21910 29044 21916 29096
rect 21968 29044 21974 29096
rect 24673 29087 24731 29093
rect 24673 29084 24685 29087
rect 22066 29056 24685 29084
rect 19334 29016 19340 29028
rect 16500 28988 19340 29016
rect 19334 28976 19340 28988
rect 19392 28976 19398 29028
rect 19521 29019 19579 29025
rect 19521 28985 19533 29019
rect 19567 29016 19579 29019
rect 22066 29016 22094 29056
rect 24673 29053 24685 29056
rect 24719 29053 24731 29087
rect 24780 29084 24808 29124
rect 24854 29112 24860 29164
rect 24912 29112 24918 29164
rect 26329 29155 26387 29161
rect 26329 29121 26341 29155
rect 26375 29152 26387 29155
rect 26436 29152 26464 29192
rect 27982 29180 27988 29192
rect 28040 29180 28046 29232
rect 28092 29229 28120 29260
rect 28350 29248 28356 29300
rect 28408 29288 28414 29300
rect 29178 29288 29184 29300
rect 28408 29260 29184 29288
rect 28408 29248 28414 29260
rect 29178 29248 29184 29260
rect 29236 29248 29242 29300
rect 29270 29248 29276 29300
rect 29328 29288 29334 29300
rect 29365 29291 29423 29297
rect 29365 29288 29377 29291
rect 29328 29260 29377 29288
rect 29328 29248 29334 29260
rect 29365 29257 29377 29260
rect 29411 29257 29423 29291
rect 29365 29251 29423 29257
rect 29546 29248 29552 29300
rect 29604 29288 29610 29300
rect 31938 29288 31944 29300
rect 29604 29260 31944 29288
rect 29604 29248 29610 29260
rect 31938 29248 31944 29260
rect 31996 29248 32002 29300
rect 34790 29248 34796 29300
rect 34848 29288 34854 29300
rect 34848 29260 35388 29288
rect 34848 29248 34854 29260
rect 28077 29223 28135 29229
rect 28077 29189 28089 29223
rect 28123 29189 28135 29223
rect 28077 29183 28135 29189
rect 28258 29180 28264 29232
rect 28316 29180 28322 29232
rect 28994 29180 29000 29232
rect 29052 29220 29058 29232
rect 29052 29192 29592 29220
rect 29052 29180 29058 29192
rect 29564 29164 29592 29192
rect 29730 29180 29736 29232
rect 29788 29220 29794 29232
rect 29788 29192 31248 29220
rect 29788 29180 29794 29192
rect 26375 29124 26464 29152
rect 26513 29155 26571 29161
rect 26375 29121 26387 29124
rect 26329 29115 26387 29121
rect 26513 29121 26525 29155
rect 26559 29152 26571 29155
rect 26786 29152 26792 29164
rect 26559 29124 26792 29152
rect 26559 29121 26571 29124
rect 26513 29115 26571 29121
rect 26786 29112 26792 29124
rect 26844 29112 26850 29164
rect 28350 29112 28356 29164
rect 28408 29152 28414 29164
rect 28894 29155 28952 29161
rect 28894 29152 28906 29155
rect 28408 29124 28906 29152
rect 28408 29112 28414 29124
rect 28894 29121 28906 29124
rect 28940 29121 28952 29155
rect 28894 29115 28952 29121
rect 29181 29155 29239 29161
rect 29181 29121 29193 29155
rect 29227 29152 29239 29155
rect 29270 29152 29276 29164
rect 29227 29124 29276 29152
rect 29227 29121 29239 29124
rect 29181 29115 29239 29121
rect 29270 29112 29276 29124
rect 29328 29112 29334 29164
rect 29546 29112 29552 29164
rect 29604 29112 29610 29164
rect 30558 29112 30564 29164
rect 30616 29152 30622 29164
rect 30926 29152 30932 29164
rect 30616 29124 30932 29152
rect 30616 29112 30622 29124
rect 30926 29112 30932 29124
rect 30984 29112 30990 29164
rect 31110 29112 31116 29164
rect 31168 29112 31174 29164
rect 31220 29152 31248 29192
rect 31294 29180 31300 29232
rect 31352 29220 31358 29232
rect 34977 29223 35035 29229
rect 34977 29220 34989 29223
rect 31352 29192 34989 29220
rect 31352 29180 31358 29192
rect 34977 29189 34989 29192
rect 35023 29189 35035 29223
rect 34977 29183 35035 29189
rect 35066 29180 35072 29232
rect 35124 29180 35130 29232
rect 31389 29155 31447 29161
rect 31389 29152 31401 29155
rect 31220 29124 31401 29152
rect 31389 29121 31401 29124
rect 31435 29121 31447 29155
rect 33689 29155 33747 29161
rect 33689 29152 33701 29155
rect 31389 29115 31447 29121
rect 33612 29124 33701 29152
rect 28534 29084 28540 29096
rect 24780 29056 28540 29084
rect 24673 29047 24731 29053
rect 28534 29044 28540 29056
rect 28592 29044 28598 29096
rect 29089 29087 29147 29093
rect 29089 29053 29101 29087
rect 29135 29084 29147 29087
rect 29454 29084 29460 29096
rect 29135 29056 29460 29084
rect 29135 29053 29147 29056
rect 29089 29047 29147 29053
rect 29454 29044 29460 29056
rect 29512 29084 29518 29096
rect 29512 29056 29592 29084
rect 29512 29044 29518 29056
rect 19567 28988 22094 29016
rect 22281 29019 22339 29025
rect 19567 28985 19579 28988
rect 19521 28979 19579 28985
rect 22281 28985 22293 29019
rect 22327 29016 22339 29019
rect 23290 29016 23296 29028
rect 22327 28988 23296 29016
rect 22327 28985 22339 28988
rect 22281 28979 22339 28985
rect 23290 28976 23296 28988
rect 23348 28976 23354 29028
rect 23382 28976 23388 29028
rect 23440 29016 23446 29028
rect 28074 29016 28080 29028
rect 23440 28988 28080 29016
rect 23440 28976 23446 28988
rect 28074 28976 28080 28988
rect 28132 28976 28138 29028
rect 28445 29019 28503 29025
rect 28445 28985 28457 29019
rect 28491 29016 28503 29019
rect 28902 29016 28908 29028
rect 28491 28988 28908 29016
rect 28491 28985 28503 28988
rect 28445 28979 28503 28985
rect 28902 28976 28908 28988
rect 28960 28976 28966 29028
rect 29564 29016 29592 29056
rect 31202 29044 31208 29096
rect 31260 29044 31266 29096
rect 29914 29016 29920 29028
rect 29564 28988 29920 29016
rect 29914 28976 29920 28988
rect 29972 28976 29978 29028
rect 31570 28976 31576 29028
rect 31628 28976 31634 29028
rect 33612 28994 33640 29124
rect 33689 29121 33701 29124
rect 33735 29121 33747 29155
rect 33689 29115 33747 29121
rect 33870 29112 33876 29164
rect 33928 29112 33934 29164
rect 34057 29155 34115 29161
rect 34057 29121 34069 29155
rect 34103 29152 34115 29155
rect 34514 29152 34520 29164
rect 34103 29124 34520 29152
rect 34103 29121 34115 29124
rect 34057 29115 34115 29121
rect 34514 29112 34520 29124
rect 34572 29112 34578 29164
rect 34698 29112 34704 29164
rect 34756 29112 34762 29164
rect 35360 29161 35388 29260
rect 35710 29248 35716 29300
rect 35768 29288 35774 29300
rect 37737 29291 37795 29297
rect 37737 29288 37749 29291
rect 35768 29260 37749 29288
rect 35768 29248 35774 29260
rect 35434 29180 35440 29232
rect 35492 29220 35498 29232
rect 35802 29220 35808 29232
rect 35492 29192 35808 29220
rect 35492 29180 35498 29192
rect 35802 29180 35808 29192
rect 35860 29220 35866 29232
rect 37292 29229 37320 29260
rect 37737 29257 37749 29260
rect 37783 29257 37795 29291
rect 37737 29251 37795 29257
rect 37277 29223 37335 29229
rect 35860 29192 35940 29220
rect 35860 29180 35866 29192
rect 35912 29161 35940 29192
rect 37277 29189 37289 29223
rect 37323 29189 37335 29223
rect 37277 29183 37335 29189
rect 37366 29180 37372 29232
rect 37424 29220 37430 29232
rect 37461 29223 37519 29229
rect 37461 29220 37473 29223
rect 37424 29192 37473 29220
rect 37424 29180 37430 29192
rect 37461 29189 37473 29192
rect 37507 29189 37519 29223
rect 37461 29183 37519 29189
rect 38746 29161 38752 29164
rect 35338 29155 35396 29161
rect 35338 29121 35350 29155
rect 35384 29121 35396 29155
rect 35621 29155 35679 29161
rect 35621 29152 35633 29155
rect 35338 29115 35396 29121
rect 35452 29124 35633 29152
rect 35452 29096 35480 29124
rect 35621 29121 35633 29124
rect 35667 29121 35679 29155
rect 35621 29115 35679 29121
rect 35897 29155 35955 29161
rect 35897 29121 35909 29155
rect 35943 29121 35955 29155
rect 35897 29115 35955 29121
rect 38740 29115 38752 29161
rect 38746 29112 38752 29115
rect 38804 29112 38810 29164
rect 40589 29155 40647 29161
rect 40589 29121 40601 29155
rect 40635 29152 40647 29155
rect 44269 29155 44327 29161
rect 44269 29152 44281 29155
rect 40635 29124 44281 29152
rect 40635 29121 40647 29124
rect 40589 29115 40647 29121
rect 44269 29121 44281 29124
rect 44315 29121 44327 29155
rect 44269 29115 44327 29121
rect 34790 29044 34796 29096
rect 34848 29044 34854 29096
rect 35250 29044 35256 29096
rect 35308 29044 35314 29096
rect 35434 29044 35440 29096
rect 35492 29044 35498 29096
rect 35713 29087 35771 29093
rect 35713 29084 35725 29087
rect 35544 29056 35725 29084
rect 33612 28966 33732 28994
rect 34146 28976 34152 29028
rect 34204 29016 34210 29028
rect 35544 29025 35572 29056
rect 35713 29053 35725 29056
rect 35759 29053 35771 29087
rect 36262 29084 36268 29096
rect 35713 29047 35771 29053
rect 35820 29056 36268 29084
rect 34517 29019 34575 29025
rect 34517 29016 34529 29019
rect 34204 28988 34529 29016
rect 34204 28976 34210 28988
rect 34517 28985 34529 28988
rect 34563 28985 34575 29019
rect 34517 28979 34575 28985
rect 35529 29019 35587 29025
rect 35529 28985 35541 29019
rect 35575 28985 35587 29019
rect 35529 28979 35587 28985
rect 35618 28976 35624 29028
rect 35676 29016 35682 29028
rect 35820 29016 35848 29056
rect 36262 29044 36268 29056
rect 36320 29044 36326 29096
rect 37182 29044 37188 29096
rect 37240 29084 37246 29096
rect 38473 29087 38531 29093
rect 38473 29084 38485 29087
rect 37240 29056 38485 29084
rect 37240 29044 37246 29056
rect 38473 29053 38485 29056
rect 38519 29053 38531 29087
rect 38473 29047 38531 29053
rect 35676 28988 35848 29016
rect 36081 29019 36139 29025
rect 35676 28976 35682 28988
rect 36081 28985 36093 29019
rect 36127 29016 36139 29019
rect 36170 29016 36176 29028
rect 36127 28988 36176 29016
rect 36127 28985 36139 28988
rect 36081 28979 36139 28985
rect 36170 28976 36176 28988
rect 36228 28976 36234 29028
rect 37642 28976 37648 29028
rect 37700 29016 37706 29028
rect 38286 29016 38292 29028
rect 37700 28988 38292 29016
rect 37700 28976 37706 28988
rect 38286 28976 38292 28988
rect 38344 28976 38350 29028
rect 39853 29019 39911 29025
rect 39853 28985 39865 29019
rect 39899 29016 39911 29019
rect 40604 29016 40632 29115
rect 39899 28988 40632 29016
rect 39899 28985 39911 28988
rect 39853 28979 39911 28985
rect 44082 28976 44088 29028
rect 44140 29016 44146 29028
rect 44453 29019 44511 29025
rect 44453 29016 44465 29019
rect 44140 28988 44465 29016
rect 44140 28976 44146 28988
rect 44453 28985 44465 28988
rect 44499 28985 44511 29019
rect 44453 28979 44511 28985
rect 11609 28951 11667 28957
rect 11609 28948 11621 28951
rect 11587 28920 11621 28948
rect 11609 28917 11621 28920
rect 11655 28917 11667 28951
rect 11609 28911 11667 28917
rect 13078 28908 13084 28960
rect 13136 28948 13142 28960
rect 17954 28948 17960 28960
rect 13136 28920 17960 28948
rect 13136 28908 13142 28920
rect 17954 28908 17960 28920
rect 18012 28908 18018 28960
rect 19245 28951 19303 28957
rect 19245 28917 19257 28951
rect 19291 28948 19303 28951
rect 20162 28948 20168 28960
rect 19291 28920 20168 28948
rect 19291 28917 19303 28920
rect 19245 28911 19303 28917
rect 20162 28908 20168 28920
rect 20220 28908 20226 28960
rect 21818 28908 21824 28960
rect 21876 28908 21882 28960
rect 22462 28908 22468 28960
rect 22520 28948 22526 28960
rect 22649 28951 22707 28957
rect 22649 28948 22661 28951
rect 22520 28920 22661 28948
rect 22520 28908 22526 28920
rect 22649 28917 22661 28920
rect 22695 28948 22707 28951
rect 23198 28948 23204 28960
rect 22695 28920 23204 28948
rect 22695 28917 22707 28920
rect 22649 28911 22707 28917
rect 23198 28908 23204 28920
rect 23256 28908 23262 28960
rect 24857 28951 24915 28957
rect 24857 28917 24869 28951
rect 24903 28948 24915 28951
rect 24946 28948 24952 28960
rect 24903 28920 24952 28948
rect 24903 28917 24915 28920
rect 24857 28911 24915 28917
rect 24946 28908 24952 28920
rect 25004 28908 25010 28960
rect 25038 28908 25044 28960
rect 25096 28908 25102 28960
rect 26326 28908 26332 28960
rect 26384 28908 26390 28960
rect 26694 28908 26700 28960
rect 26752 28908 26758 28960
rect 26786 28908 26792 28960
rect 26844 28948 26850 28960
rect 28626 28948 28632 28960
rect 26844 28920 28632 28948
rect 26844 28908 26850 28920
rect 28626 28908 28632 28920
rect 28684 28908 28690 28960
rect 29089 28951 29147 28957
rect 29089 28917 29101 28951
rect 29135 28948 29147 28951
rect 29362 28948 29368 28960
rect 29135 28920 29368 28948
rect 29135 28917 29147 28920
rect 29089 28911 29147 28917
rect 29362 28908 29368 28920
rect 29420 28908 29426 28960
rect 29822 28908 29828 28960
rect 29880 28948 29886 28960
rect 31113 28951 31171 28957
rect 31113 28948 31125 28951
rect 29880 28920 31125 28948
rect 29880 28908 29886 28920
rect 31113 28917 31125 28920
rect 31159 28917 31171 28951
rect 33704 28948 33732 28966
rect 33870 28948 33876 28960
rect 33704 28920 33876 28948
rect 31113 28911 31171 28917
rect 33870 28908 33876 28920
rect 33928 28908 33934 28960
rect 34330 28908 34336 28960
rect 34388 28948 34394 28960
rect 34701 28951 34759 28957
rect 34701 28948 34713 28951
rect 34388 28920 34713 28948
rect 34388 28908 34394 28920
rect 34701 28917 34713 28920
rect 34747 28917 34759 28951
rect 34701 28911 34759 28917
rect 34882 28908 34888 28960
rect 34940 28948 34946 28960
rect 35069 28951 35127 28957
rect 35069 28948 35081 28951
rect 34940 28920 35081 28948
rect 34940 28908 34946 28920
rect 35069 28917 35081 28920
rect 35115 28917 35127 28951
rect 35069 28911 35127 28917
rect 35805 28951 35863 28957
rect 35805 28917 35817 28951
rect 35851 28948 35863 28951
rect 36262 28948 36268 28960
rect 35851 28920 36268 28948
rect 35851 28917 35863 28920
rect 35805 28911 35863 28917
rect 36262 28908 36268 28920
rect 36320 28908 36326 28960
rect 39942 28908 39948 28960
rect 40000 28908 40006 28960
rect 1104 28858 44896 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 44896 28858
rect 1104 28784 44896 28806
rect 8938 28704 8944 28756
rect 8996 28704 9002 28756
rect 9306 28704 9312 28756
rect 9364 28704 9370 28756
rect 9674 28704 9680 28756
rect 9732 28744 9738 28756
rect 10873 28747 10931 28753
rect 10873 28744 10885 28747
rect 9732 28716 10885 28744
rect 9732 28704 9738 28716
rect 10873 28713 10885 28716
rect 10919 28744 10931 28747
rect 11054 28744 11060 28756
rect 10919 28716 11060 28744
rect 10919 28713 10931 28716
rect 10873 28707 10931 28713
rect 11054 28704 11060 28716
rect 11112 28704 11118 28756
rect 11330 28704 11336 28756
rect 11388 28704 11394 28756
rect 21818 28744 21824 28756
rect 11440 28716 21824 28744
rect 8018 28636 8024 28688
rect 8076 28676 8082 28688
rect 11440 28676 11468 28716
rect 21818 28704 21824 28716
rect 21876 28704 21882 28756
rect 22830 28704 22836 28756
rect 22888 28744 22894 28756
rect 22925 28747 22983 28753
rect 22925 28744 22937 28747
rect 22888 28716 22937 28744
rect 22888 28704 22894 28716
rect 22925 28713 22937 28716
rect 22971 28713 22983 28747
rect 22925 28707 22983 28713
rect 23290 28704 23296 28756
rect 23348 28704 23354 28756
rect 26973 28747 27031 28753
rect 26973 28713 26985 28747
rect 27019 28713 27031 28747
rect 26973 28707 27031 28713
rect 8076 28648 11468 28676
rect 8076 28636 8082 28648
rect 11514 28636 11520 28688
rect 11572 28676 11578 28688
rect 13170 28676 13176 28688
rect 11572 28648 13176 28676
rect 11572 28636 11578 28648
rect 13170 28636 13176 28648
rect 13228 28676 13234 28688
rect 13722 28676 13728 28688
rect 13228 28648 13728 28676
rect 13228 28636 13234 28648
rect 13722 28636 13728 28648
rect 13780 28636 13786 28688
rect 16114 28636 16120 28688
rect 16172 28676 16178 28688
rect 26988 28676 27016 28707
rect 27430 28704 27436 28756
rect 27488 28744 27494 28756
rect 27525 28747 27583 28753
rect 27525 28744 27537 28747
rect 27488 28716 27537 28744
rect 27488 28704 27494 28716
rect 27525 28713 27537 28716
rect 27571 28713 27583 28747
rect 27525 28707 27583 28713
rect 28810 28704 28816 28756
rect 28868 28704 28874 28756
rect 29273 28747 29331 28753
rect 29273 28713 29285 28747
rect 29319 28744 29331 28747
rect 29730 28744 29736 28756
rect 29319 28716 29736 28744
rect 29319 28713 29331 28716
rect 29273 28707 29331 28713
rect 29730 28704 29736 28716
rect 29788 28704 29794 28756
rect 31110 28704 31116 28756
rect 31168 28744 31174 28756
rect 31573 28747 31631 28753
rect 31573 28744 31585 28747
rect 31168 28716 31585 28744
rect 31168 28704 31174 28716
rect 31573 28713 31585 28716
rect 31619 28744 31631 28747
rect 31662 28744 31668 28756
rect 31619 28716 31668 28744
rect 31619 28713 31631 28716
rect 31573 28707 31631 28713
rect 31662 28704 31668 28716
rect 31720 28704 31726 28756
rect 34330 28704 34336 28756
rect 34388 28744 34394 28756
rect 35342 28744 35348 28756
rect 34388 28716 35348 28744
rect 34388 28704 34394 28716
rect 35342 28704 35348 28716
rect 35400 28704 35406 28756
rect 36078 28704 36084 28756
rect 36136 28744 36142 28756
rect 37182 28744 37188 28756
rect 36136 28716 37188 28744
rect 36136 28704 36142 28716
rect 37182 28704 37188 28716
rect 37240 28744 37246 28756
rect 37369 28747 37427 28753
rect 37369 28744 37381 28747
rect 37240 28716 37381 28744
rect 37240 28704 37246 28716
rect 37369 28713 37381 28716
rect 37415 28713 37427 28747
rect 37369 28707 37427 28713
rect 38197 28747 38255 28753
rect 38197 28713 38209 28747
rect 38243 28744 38255 28747
rect 38378 28744 38384 28756
rect 38243 28716 38384 28744
rect 38243 28713 38255 28716
rect 38197 28707 38255 28713
rect 38378 28704 38384 28716
rect 38436 28704 38442 28756
rect 38473 28747 38531 28753
rect 38473 28713 38485 28747
rect 38519 28744 38531 28747
rect 38746 28744 38752 28756
rect 38519 28716 38752 28744
rect 38519 28713 38531 28716
rect 38473 28707 38531 28713
rect 38746 28704 38752 28716
rect 38804 28704 38810 28756
rect 28902 28676 28908 28688
rect 16172 28648 27016 28676
rect 27080 28648 28908 28676
rect 16172 28636 16178 28648
rect 11057 28611 11115 28617
rect 11057 28577 11069 28611
rect 11103 28608 11115 28611
rect 11422 28608 11428 28620
rect 11103 28580 11428 28608
rect 11103 28577 11115 28580
rect 11057 28571 11115 28577
rect 11422 28568 11428 28580
rect 11480 28568 11486 28620
rect 23198 28608 23204 28620
rect 11624 28580 23204 28608
rect 9122 28500 9128 28552
rect 9180 28500 9186 28552
rect 9309 28543 9367 28549
rect 9309 28509 9321 28543
rect 9355 28540 9367 28543
rect 9582 28540 9588 28552
rect 9355 28512 9588 28540
rect 9355 28509 9367 28512
rect 9309 28503 9367 28509
rect 9582 28500 9588 28512
rect 9640 28500 9646 28552
rect 9950 28500 9956 28552
rect 10008 28540 10014 28552
rect 10008 28512 10640 28540
rect 10008 28500 10014 28512
rect 10612 28484 10640 28512
rect 10686 28500 10692 28552
rect 10744 28540 10750 28552
rect 11149 28543 11207 28549
rect 11149 28540 11161 28543
rect 10744 28512 11161 28540
rect 10744 28500 10750 28512
rect 11149 28509 11161 28512
rect 11195 28540 11207 28543
rect 11624 28540 11652 28580
rect 23198 28568 23204 28580
rect 23256 28568 23262 28620
rect 23293 28611 23351 28617
rect 23293 28577 23305 28611
rect 23339 28608 23351 28611
rect 23382 28608 23388 28620
rect 23339 28580 23388 28608
rect 23339 28577 23351 28580
rect 23293 28571 23351 28577
rect 23382 28568 23388 28580
rect 23440 28568 23446 28620
rect 25498 28568 25504 28620
rect 25556 28608 25562 28620
rect 26142 28608 26148 28620
rect 25556 28580 26148 28608
rect 25556 28568 25562 28580
rect 26142 28568 26148 28580
rect 26200 28568 26206 28620
rect 27080 28617 27108 28648
rect 28902 28636 28908 28648
rect 28960 28636 28966 28688
rect 28994 28636 29000 28688
rect 29052 28636 29058 28688
rect 31294 28676 31300 28688
rect 29288 28648 31300 28676
rect 27065 28611 27123 28617
rect 27065 28577 27077 28611
rect 27111 28577 27123 28611
rect 27065 28571 27123 28577
rect 27709 28611 27767 28617
rect 27709 28577 27721 28611
rect 27755 28608 27767 28611
rect 28810 28608 28816 28620
rect 27755 28580 28816 28608
rect 27755 28577 27767 28580
rect 27709 28571 27767 28577
rect 28810 28568 28816 28580
rect 28868 28568 28874 28620
rect 29012 28608 29040 28636
rect 29181 28611 29239 28617
rect 29181 28608 29193 28611
rect 29012 28580 29193 28608
rect 29181 28577 29193 28580
rect 29227 28608 29239 28611
rect 29288 28608 29316 28648
rect 31294 28636 31300 28648
rect 31352 28636 31358 28688
rect 33134 28636 33140 28688
rect 33192 28676 33198 28688
rect 33229 28679 33287 28685
rect 33229 28676 33241 28679
rect 33192 28648 33241 28676
rect 33192 28636 33198 28648
rect 33229 28645 33241 28648
rect 33275 28676 33287 28679
rect 33318 28676 33324 28688
rect 33275 28648 33324 28676
rect 33275 28645 33287 28648
rect 33229 28639 33287 28645
rect 33318 28636 33324 28648
rect 33376 28636 33382 28688
rect 35989 28679 36047 28685
rect 35989 28645 36001 28679
rect 36035 28676 36047 28679
rect 41138 28676 41144 28688
rect 36035 28648 41144 28676
rect 36035 28645 36047 28648
rect 35989 28639 36047 28645
rect 41138 28636 41144 28648
rect 41196 28636 41202 28688
rect 29227 28580 29316 28608
rect 29227 28577 29239 28580
rect 29181 28571 29239 28577
rect 34054 28568 34060 28620
rect 34112 28608 34118 28620
rect 34606 28608 34612 28620
rect 34112 28580 34612 28608
rect 34112 28568 34118 28580
rect 34606 28568 34612 28580
rect 34664 28608 34670 28620
rect 36722 28608 36728 28620
rect 34664 28580 36728 28608
rect 34664 28568 34670 28580
rect 36722 28568 36728 28580
rect 36780 28568 36786 28620
rect 38010 28568 38016 28620
rect 38068 28568 38074 28620
rect 38562 28568 38568 28620
rect 38620 28608 38626 28620
rect 38749 28611 38807 28617
rect 38749 28608 38761 28611
rect 38620 28580 38761 28608
rect 38620 28568 38626 28580
rect 38749 28577 38761 28580
rect 38795 28577 38807 28611
rect 38749 28571 38807 28577
rect 38933 28611 38991 28617
rect 38933 28577 38945 28611
rect 38979 28608 38991 28611
rect 40034 28608 40040 28620
rect 38979 28580 40040 28608
rect 38979 28577 38991 28580
rect 38933 28571 38991 28577
rect 40034 28568 40040 28580
rect 40092 28568 40098 28620
rect 11195 28512 11652 28540
rect 18141 28543 18199 28549
rect 11195 28509 11207 28512
rect 11149 28503 11207 28509
rect 18141 28509 18153 28543
rect 18187 28540 18199 28543
rect 18187 28512 18644 28540
rect 18187 28509 18199 28512
rect 18141 28503 18199 28509
rect 5718 28432 5724 28484
rect 5776 28472 5782 28484
rect 10413 28475 10471 28481
rect 10413 28472 10425 28475
rect 5776 28444 10425 28472
rect 5776 28432 5782 28444
rect 10413 28441 10425 28444
rect 10459 28441 10471 28475
rect 10413 28435 10471 28441
rect 10428 28404 10456 28435
rect 10594 28432 10600 28484
rect 10652 28432 10658 28484
rect 10778 28432 10784 28484
rect 10836 28432 10842 28484
rect 10870 28432 10876 28484
rect 10928 28432 10934 28484
rect 17957 28475 18015 28481
rect 17957 28441 17969 28475
rect 18003 28472 18015 28475
rect 18046 28472 18052 28484
rect 18003 28444 18052 28472
rect 18003 28441 18015 28444
rect 17957 28435 18015 28441
rect 18046 28432 18052 28444
rect 18104 28432 18110 28484
rect 18230 28432 18236 28484
rect 18288 28432 18294 28484
rect 18414 28432 18420 28484
rect 18472 28432 18478 28484
rect 18616 28416 18644 28512
rect 23106 28500 23112 28552
rect 23164 28500 23170 28552
rect 26694 28500 26700 28552
rect 26752 28540 26758 28552
rect 26973 28543 27031 28549
rect 26973 28540 26985 28543
rect 26752 28512 26985 28540
rect 26752 28500 26758 28512
rect 26973 28509 26985 28512
rect 27019 28509 27031 28543
rect 26973 28503 27031 28509
rect 27246 28500 27252 28552
rect 27304 28500 27310 28552
rect 27801 28543 27859 28549
rect 27801 28509 27813 28543
rect 27847 28540 27859 28543
rect 27890 28540 27896 28552
rect 27847 28512 27896 28540
rect 27847 28509 27859 28512
rect 27801 28503 27859 28509
rect 27890 28500 27896 28512
rect 27948 28500 27954 28552
rect 28957 28543 29015 28549
rect 28957 28509 28969 28543
rect 29003 28509 29015 28543
rect 28957 28503 29015 28509
rect 20254 28432 20260 28484
rect 20312 28472 20318 28484
rect 22186 28472 22192 28484
rect 20312 28444 22192 28472
rect 20312 28432 20318 28444
rect 22186 28432 22192 28444
rect 22244 28432 22250 28484
rect 23382 28432 23388 28484
rect 23440 28432 23446 28484
rect 24946 28432 24952 28484
rect 25004 28472 25010 28484
rect 25590 28472 25596 28484
rect 25004 28444 25596 28472
rect 25004 28432 25010 28444
rect 25590 28432 25596 28444
rect 25648 28432 25654 28484
rect 26142 28432 26148 28484
rect 26200 28472 26206 28484
rect 27525 28475 27583 28481
rect 27525 28472 27537 28475
rect 26200 28444 26924 28472
rect 26200 28432 26206 28444
rect 11514 28404 11520 28416
rect 10428 28376 11520 28404
rect 11514 28364 11520 28376
rect 11572 28364 11578 28416
rect 14918 28364 14924 28416
rect 14976 28404 14982 28416
rect 17773 28407 17831 28413
rect 17773 28404 17785 28407
rect 14976 28376 17785 28404
rect 14976 28364 14982 28376
rect 17773 28373 17785 28376
rect 17819 28404 17831 28407
rect 18506 28404 18512 28416
rect 17819 28376 18512 28404
rect 17819 28373 17831 28376
rect 17773 28367 17831 28373
rect 18506 28364 18512 28376
rect 18564 28364 18570 28416
rect 18598 28364 18604 28416
rect 18656 28364 18662 28416
rect 18782 28364 18788 28416
rect 18840 28404 18846 28416
rect 20070 28404 20076 28416
rect 18840 28376 20076 28404
rect 18840 28364 18846 28376
rect 20070 28364 20076 28376
rect 20128 28364 20134 28416
rect 20162 28364 20168 28416
rect 20220 28404 20226 28416
rect 26786 28404 26792 28416
rect 20220 28376 26792 28404
rect 20220 28364 20226 28376
rect 26786 28364 26792 28376
rect 26844 28364 26850 28416
rect 26896 28404 26924 28444
rect 27080 28444 27537 28472
rect 27080 28404 27108 28444
rect 27525 28441 27537 28444
rect 27571 28441 27583 28475
rect 27525 28435 27583 28441
rect 28258 28432 28264 28484
rect 28316 28472 28322 28484
rect 28353 28475 28411 28481
rect 28353 28472 28365 28475
rect 28316 28444 28365 28472
rect 28316 28432 28322 28444
rect 28353 28441 28365 28444
rect 28399 28441 28411 28475
rect 28353 28435 28411 28441
rect 28442 28432 28448 28484
rect 28500 28472 28506 28484
rect 28537 28475 28595 28481
rect 28537 28472 28549 28475
rect 28500 28444 28549 28472
rect 28500 28432 28506 28444
rect 28537 28441 28549 28444
rect 28583 28441 28595 28475
rect 28537 28435 28595 28441
rect 28966 28416 28994 28503
rect 30282 28500 30288 28552
rect 30340 28540 30346 28552
rect 30742 28540 30748 28552
rect 30340 28512 30748 28540
rect 30340 28500 30346 28512
rect 30742 28500 30748 28512
rect 30800 28540 30806 28552
rect 31205 28543 31263 28549
rect 31205 28540 31217 28543
rect 30800 28512 31217 28540
rect 30800 28500 30806 28512
rect 31205 28509 31217 28512
rect 31251 28509 31263 28543
rect 35710 28540 35716 28552
rect 31205 28503 31263 28509
rect 35176 28512 35716 28540
rect 29273 28475 29331 28481
rect 29273 28441 29285 28475
rect 29319 28441 29331 28475
rect 29273 28435 29331 28441
rect 26896 28376 27108 28404
rect 27433 28407 27491 28413
rect 27433 28373 27445 28407
rect 27479 28404 27491 28407
rect 27706 28404 27712 28416
rect 27479 28376 27712 28404
rect 27479 28373 27491 28376
rect 27433 28367 27491 28373
rect 27706 28364 27712 28376
rect 27764 28364 27770 28416
rect 27982 28364 27988 28416
rect 28040 28364 28046 28416
rect 28718 28364 28724 28416
rect 28776 28364 28782 28416
rect 28966 28376 29000 28416
rect 28994 28364 29000 28376
rect 29052 28364 29058 28416
rect 29288 28404 29316 28435
rect 31386 28432 31392 28484
rect 31444 28432 31450 28484
rect 32858 28432 32864 28484
rect 32916 28432 32922 28484
rect 33045 28475 33103 28481
rect 33045 28441 33057 28475
rect 33091 28472 33103 28475
rect 33502 28472 33508 28484
rect 33091 28444 33508 28472
rect 33091 28441 33103 28444
rect 33045 28435 33103 28441
rect 29362 28404 29368 28416
rect 29288 28376 29368 28404
rect 29362 28364 29368 28376
rect 29420 28364 29426 28416
rect 32674 28364 32680 28416
rect 32732 28404 32738 28416
rect 33060 28404 33088 28435
rect 33502 28432 33508 28444
rect 33560 28432 33566 28484
rect 33870 28432 33876 28484
rect 33928 28472 33934 28484
rect 34606 28472 34612 28484
rect 33928 28444 34612 28472
rect 33928 28432 33934 28444
rect 34606 28432 34612 28444
rect 34664 28472 34670 28484
rect 35176 28481 35204 28512
rect 35710 28500 35716 28512
rect 35768 28500 35774 28552
rect 35802 28500 35808 28552
rect 35860 28500 35866 28552
rect 36998 28500 37004 28552
rect 37056 28540 37062 28552
rect 38197 28543 38255 28549
rect 38197 28540 38209 28543
rect 37056 28512 38209 28540
rect 37056 28500 37062 28512
rect 38197 28509 38209 28512
rect 38243 28509 38255 28543
rect 38197 28503 38255 28509
rect 38657 28543 38715 28549
rect 38657 28509 38669 28543
rect 38703 28540 38715 28543
rect 38841 28543 38899 28549
rect 38703 28512 38792 28540
rect 38703 28509 38715 28512
rect 38657 28503 38715 28509
rect 38764 28484 38792 28512
rect 38841 28509 38853 28543
rect 38887 28509 38899 28543
rect 38841 28503 38899 28509
rect 39117 28543 39175 28549
rect 39117 28509 39129 28543
rect 39163 28540 39175 28543
rect 39942 28540 39948 28552
rect 39163 28512 39948 28540
rect 39163 28509 39175 28512
rect 39117 28503 39175 28509
rect 34977 28475 35035 28481
rect 34977 28472 34989 28475
rect 34664 28444 34989 28472
rect 34664 28432 34670 28444
rect 34977 28441 34989 28444
rect 35023 28441 35035 28475
rect 34977 28435 35035 28441
rect 35161 28475 35219 28481
rect 35161 28441 35173 28475
rect 35207 28441 35219 28475
rect 35161 28435 35219 28441
rect 32732 28376 33088 28404
rect 32732 28364 32738 28376
rect 34330 28364 34336 28416
rect 34388 28404 34394 28416
rect 35176 28404 35204 28435
rect 35618 28432 35624 28484
rect 35676 28432 35682 28484
rect 35986 28432 35992 28484
rect 36044 28472 36050 28484
rect 36081 28475 36139 28481
rect 36081 28472 36093 28475
rect 36044 28444 36093 28472
rect 36044 28432 36050 28444
rect 36081 28441 36093 28444
rect 36127 28441 36139 28475
rect 36081 28435 36139 28441
rect 37458 28432 37464 28484
rect 37516 28472 37522 28484
rect 37921 28475 37979 28481
rect 37921 28472 37933 28475
rect 37516 28444 37933 28472
rect 37516 28432 37522 28444
rect 37921 28441 37933 28444
rect 37967 28441 37979 28475
rect 37921 28435 37979 28441
rect 38746 28432 38752 28484
rect 38804 28432 38810 28484
rect 34388 28376 35204 28404
rect 34388 28364 34394 28376
rect 35342 28364 35348 28416
rect 35400 28364 35406 28416
rect 35526 28364 35532 28416
rect 35584 28404 35590 28416
rect 36446 28404 36452 28416
rect 35584 28376 36452 28404
rect 35584 28364 35590 28376
rect 36446 28364 36452 28376
rect 36504 28364 36510 28416
rect 38194 28364 38200 28416
rect 38252 28404 38258 28416
rect 38381 28407 38439 28413
rect 38381 28404 38393 28407
rect 38252 28376 38393 28404
rect 38252 28364 38258 28376
rect 38381 28373 38393 28376
rect 38427 28373 38439 28407
rect 38381 28367 38439 28373
rect 38654 28364 38660 28416
rect 38712 28404 38718 28416
rect 38856 28404 38884 28503
rect 39942 28500 39948 28512
rect 40000 28500 40006 28552
rect 41230 28500 41236 28552
rect 41288 28500 41294 28552
rect 41500 28475 41558 28481
rect 41500 28441 41512 28475
rect 41546 28472 41558 28475
rect 42058 28472 42064 28484
rect 41546 28444 42064 28472
rect 41546 28441 41558 28444
rect 41500 28435 41558 28441
rect 42058 28432 42064 28444
rect 42116 28432 42122 28484
rect 38712 28376 38884 28404
rect 42613 28407 42671 28413
rect 38712 28364 38718 28376
rect 42613 28373 42625 28407
rect 42659 28404 42671 28407
rect 42978 28404 42984 28416
rect 42659 28376 42984 28404
rect 42659 28373 42671 28376
rect 42613 28367 42671 28373
rect 42978 28364 42984 28376
rect 43036 28364 43042 28416
rect 1104 28314 44896 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 44896 28314
rect 1104 28240 44896 28262
rect 8389 28203 8447 28209
rect 8389 28169 8401 28203
rect 8435 28200 8447 28203
rect 10686 28200 10692 28212
rect 8435 28172 10692 28200
rect 8435 28169 8447 28172
rect 8389 28163 8447 28169
rect 10686 28160 10692 28172
rect 10744 28160 10750 28212
rect 10870 28160 10876 28212
rect 10928 28160 10934 28212
rect 15562 28200 15568 28212
rect 14936 28172 15568 28200
rect 7558 28092 7564 28144
rect 7616 28132 7622 28144
rect 8205 28135 8263 28141
rect 8205 28132 8217 28135
rect 7616 28104 8217 28132
rect 7616 28092 7622 28104
rect 8205 28101 8217 28104
rect 8251 28101 8263 28135
rect 8205 28095 8263 28101
rect 10413 28135 10471 28141
rect 10413 28101 10425 28135
rect 10459 28132 10471 28135
rect 11606 28132 11612 28144
rect 10459 28104 11612 28132
rect 10459 28101 10471 28104
rect 10413 28095 10471 28101
rect 11606 28092 11612 28104
rect 11664 28092 11670 28144
rect 14458 28092 14464 28144
rect 14516 28132 14522 28144
rect 14645 28135 14703 28141
rect 14645 28132 14657 28135
rect 14516 28104 14657 28132
rect 14516 28092 14522 28104
rect 14645 28101 14657 28104
rect 14691 28101 14703 28135
rect 14936 28132 14964 28172
rect 15562 28160 15568 28172
rect 15620 28160 15626 28212
rect 16298 28160 16304 28212
rect 16356 28160 16362 28212
rect 16666 28160 16672 28212
rect 16724 28200 16730 28212
rect 18782 28200 18788 28212
rect 16724 28172 18788 28200
rect 16724 28160 16730 28172
rect 18782 28160 18788 28172
rect 18840 28160 18846 28212
rect 18966 28160 18972 28212
rect 19024 28200 19030 28212
rect 21634 28200 21640 28212
rect 19024 28172 21640 28200
rect 19024 28160 19030 28172
rect 21634 28160 21640 28172
rect 21692 28160 21698 28212
rect 23661 28203 23719 28209
rect 23661 28169 23673 28203
rect 23707 28200 23719 28203
rect 23707 28172 24716 28200
rect 23707 28169 23719 28172
rect 23661 28163 23719 28169
rect 17402 28132 17408 28144
rect 14645 28095 14703 28101
rect 14844 28104 14964 28132
rect 15304 28104 17408 28132
rect 5258 28024 5264 28076
rect 5316 28064 5322 28076
rect 6365 28067 6423 28073
rect 6365 28064 6377 28067
rect 5316 28036 6377 28064
rect 5316 28024 5322 28036
rect 6365 28033 6377 28036
rect 6411 28033 6423 28067
rect 6641 28067 6699 28073
rect 6641 28064 6653 28067
rect 6365 28027 6423 28033
rect 6472 28036 6653 28064
rect 6086 27956 6092 28008
rect 6144 27996 6150 28008
rect 6472 27996 6500 28036
rect 6641 28033 6653 28036
rect 6687 28033 6699 28067
rect 6641 28027 6699 28033
rect 7006 28024 7012 28076
rect 7064 28064 7070 28076
rect 8018 28064 8024 28076
rect 7064 28036 8024 28064
rect 7064 28024 7070 28036
rect 8018 28024 8024 28036
rect 8076 28024 8082 28076
rect 10689 28067 10747 28073
rect 10689 28033 10701 28067
rect 10735 28033 10747 28067
rect 10689 28027 10747 28033
rect 6144 27968 6500 27996
rect 6549 27999 6607 28005
rect 6144 27956 6150 27968
rect 6549 27965 6561 27999
rect 6595 27996 6607 27999
rect 6730 27996 6736 28008
rect 6595 27968 6736 27996
rect 6595 27965 6607 27968
rect 6549 27959 6607 27965
rect 6730 27956 6736 27968
rect 6788 27956 6794 28008
rect 10597 27999 10655 28005
rect 10597 27965 10609 27999
rect 10643 27965 10655 27999
rect 10704 27996 10732 28027
rect 11054 28024 11060 28076
rect 11112 28064 11118 28076
rect 13173 28067 13231 28073
rect 13173 28064 13185 28067
rect 11112 28036 13185 28064
rect 11112 28024 11118 28036
rect 13173 28033 13185 28036
rect 13219 28033 13231 28067
rect 13173 28027 13231 28033
rect 13449 28067 13507 28073
rect 13449 28033 13461 28067
rect 13495 28064 13507 28067
rect 13538 28064 13544 28076
rect 13495 28036 13544 28064
rect 13495 28033 13507 28036
rect 13449 28027 13507 28033
rect 13538 28024 13544 28036
rect 13596 28064 13602 28076
rect 14274 28064 14280 28076
rect 13596 28036 14280 28064
rect 13596 28024 13602 28036
rect 14274 28024 14280 28036
rect 14332 28024 14338 28076
rect 14844 28073 14872 28104
rect 14829 28067 14887 28073
rect 14829 28033 14841 28067
rect 14875 28033 14887 28067
rect 14829 28027 14887 28033
rect 14921 28067 14979 28073
rect 14921 28033 14933 28067
rect 14967 28064 14979 28067
rect 15010 28064 15016 28076
rect 14967 28036 15016 28064
rect 14967 28033 14979 28036
rect 14921 28027 14979 28033
rect 15010 28024 15016 28036
rect 15068 28024 15074 28076
rect 15194 28024 15200 28076
rect 15252 28024 15258 28076
rect 11790 27996 11796 28008
rect 10704 27968 11796 27996
rect 10597 27959 10655 27965
rect 6822 27888 6828 27940
rect 6880 27888 6886 27940
rect 10612 27928 10640 27959
rect 11790 27956 11796 27968
rect 11848 27956 11854 28008
rect 13262 27956 13268 28008
rect 13320 27956 13326 28008
rect 15304 28005 15332 28104
rect 17402 28092 17408 28104
rect 17460 28092 17466 28144
rect 18601 28135 18659 28141
rect 18601 28101 18613 28135
rect 18647 28132 18659 28135
rect 19521 28135 19579 28141
rect 19521 28132 19533 28135
rect 18647 28104 19533 28132
rect 18647 28101 18659 28104
rect 18601 28095 18659 28101
rect 19521 28101 19533 28104
rect 19567 28132 19579 28135
rect 19794 28132 19800 28144
rect 19567 28104 19800 28132
rect 19567 28101 19579 28104
rect 19521 28095 19579 28101
rect 19794 28092 19800 28104
rect 19852 28092 19858 28144
rect 20070 28092 20076 28144
rect 20128 28132 20134 28144
rect 20441 28135 20499 28141
rect 20441 28132 20453 28135
rect 20128 28104 20453 28132
rect 20128 28092 20134 28104
rect 20441 28101 20453 28104
rect 20487 28101 20499 28135
rect 20441 28095 20499 28101
rect 15470 28024 15476 28076
rect 15528 28024 15534 28076
rect 15838 28024 15844 28076
rect 15896 28024 15902 28076
rect 16117 28067 16175 28073
rect 16117 28064 16129 28067
rect 15948 28036 16129 28064
rect 15289 27999 15347 28005
rect 15289 27996 15301 27999
rect 14844 27968 15301 27996
rect 11514 27928 11520 27940
rect 10612 27900 11520 27928
rect 11514 27888 11520 27900
rect 11572 27888 11578 27940
rect 13078 27888 13084 27940
rect 13136 27928 13142 27940
rect 14844 27928 14872 27968
rect 15289 27965 15301 27968
rect 15335 27965 15347 27999
rect 15289 27959 15347 27965
rect 15562 27956 15568 28008
rect 15620 27996 15626 28008
rect 15948 27996 15976 28036
rect 16117 28033 16129 28036
rect 16163 28033 16175 28067
rect 16117 28027 16175 28033
rect 18506 28024 18512 28076
rect 18564 28064 18570 28076
rect 18785 28067 18843 28073
rect 18785 28064 18797 28067
rect 18564 28036 18797 28064
rect 18564 28024 18570 28036
rect 18785 28033 18797 28036
rect 18831 28033 18843 28067
rect 18785 28027 18843 28033
rect 18874 28024 18880 28076
rect 18932 28024 18938 28076
rect 19150 28024 19156 28076
rect 19208 28024 19214 28076
rect 19242 28024 19248 28076
rect 19300 28064 19306 28076
rect 19337 28067 19395 28073
rect 19337 28064 19349 28067
rect 19300 28036 19349 28064
rect 19300 28024 19306 28036
rect 19337 28033 19349 28036
rect 19383 28033 19395 28067
rect 19337 28027 19395 28033
rect 20530 28024 20536 28076
rect 20588 28064 20594 28076
rect 20625 28067 20683 28073
rect 20625 28064 20637 28067
rect 20588 28036 20637 28064
rect 20588 28024 20594 28036
rect 20625 28033 20637 28036
rect 20671 28033 20683 28067
rect 20625 28027 20683 28033
rect 23293 28067 23351 28073
rect 23293 28033 23305 28067
rect 23339 28064 23351 28067
rect 24118 28064 24124 28076
rect 23339 28036 24124 28064
rect 23339 28033 23351 28036
rect 23293 28027 23351 28033
rect 24118 28024 24124 28036
rect 24176 28024 24182 28076
rect 24210 28024 24216 28076
rect 24268 28064 24274 28076
rect 24688 28073 24716 28172
rect 26786 28160 26792 28212
rect 26844 28160 26850 28212
rect 27430 28160 27436 28212
rect 27488 28160 27494 28212
rect 27522 28160 27528 28212
rect 27580 28160 27586 28212
rect 28994 28160 29000 28212
rect 29052 28200 29058 28212
rect 29454 28200 29460 28212
rect 29052 28172 29460 28200
rect 29052 28160 29058 28172
rect 29454 28160 29460 28172
rect 29512 28200 29518 28212
rect 29549 28203 29607 28209
rect 29549 28200 29561 28203
rect 29512 28172 29561 28200
rect 29512 28160 29518 28172
rect 29549 28169 29561 28172
rect 29595 28169 29607 28203
rect 30466 28200 30472 28212
rect 29549 28163 29607 28169
rect 29656 28172 30472 28200
rect 26973 28135 27031 28141
rect 26973 28132 26985 28135
rect 24964 28104 26985 28132
rect 24397 28067 24455 28073
rect 24397 28064 24409 28067
rect 24268 28036 24409 28064
rect 24268 28024 24274 28036
rect 24397 28033 24409 28036
rect 24443 28033 24455 28067
rect 24397 28027 24455 28033
rect 24673 28067 24731 28073
rect 24673 28033 24685 28067
rect 24719 28064 24731 28067
rect 24854 28064 24860 28076
rect 24719 28036 24860 28064
rect 24719 28033 24731 28036
rect 24673 28027 24731 28033
rect 24854 28024 24860 28036
rect 24912 28024 24918 28076
rect 15620 27968 15976 27996
rect 15620 27956 15626 27968
rect 16022 27956 16028 28008
rect 16080 27956 16086 28008
rect 18892 27996 18920 28024
rect 22830 27996 22836 28008
rect 18892 27968 22836 27996
rect 22830 27956 22836 27968
rect 22888 27956 22894 28008
rect 23385 27999 23443 28005
rect 23385 27965 23397 27999
rect 23431 27996 23443 27999
rect 23474 27996 23480 28008
rect 23431 27968 23480 27996
rect 23431 27965 23443 27968
rect 23385 27959 23443 27965
rect 23474 27956 23480 27968
rect 23532 27956 23538 28008
rect 24486 27956 24492 28008
rect 24544 27956 24550 28008
rect 13136 27900 14872 27928
rect 15105 27931 15163 27937
rect 13136 27888 13142 27900
rect 15105 27897 15117 27931
rect 15151 27928 15163 27931
rect 21910 27928 21916 27940
rect 15151 27900 21916 27928
rect 15151 27897 15163 27900
rect 15105 27891 15163 27897
rect 21910 27888 21916 27900
rect 21968 27888 21974 27940
rect 22002 27888 22008 27940
rect 22060 27928 22066 27940
rect 24964 27928 24992 28104
rect 26973 28101 26985 28104
rect 27019 28101 27031 28135
rect 26973 28095 27031 28101
rect 27062 28092 27068 28144
rect 27120 28132 27126 28144
rect 27120 28104 28028 28132
rect 27120 28092 27126 28104
rect 25038 28024 25044 28076
rect 25096 28064 25102 28076
rect 26329 28067 26387 28073
rect 26329 28064 26341 28067
rect 25096 28036 26341 28064
rect 25096 28024 25102 28036
rect 26329 28033 26341 28036
rect 26375 28033 26387 28067
rect 26329 28027 26387 28033
rect 26602 28024 26608 28076
rect 26660 28024 26666 28076
rect 27246 28024 27252 28076
rect 27304 28024 27310 28076
rect 27706 28024 27712 28076
rect 27764 28024 27770 28076
rect 27893 28067 27951 28073
rect 27893 28033 27905 28067
rect 27939 28033 27951 28067
rect 27893 28027 27951 28033
rect 26513 27999 26571 28005
rect 26513 27965 26525 27999
rect 26559 27965 26571 27999
rect 26513 27959 26571 27965
rect 22060 27900 24992 27928
rect 26528 27928 26556 27959
rect 26694 27956 26700 28008
rect 26752 27996 26758 28008
rect 27065 27999 27123 28005
rect 27065 27996 27077 27999
rect 26752 27968 27077 27996
rect 26752 27956 26758 27968
rect 27065 27965 27077 27968
rect 27111 27965 27123 27999
rect 27065 27959 27123 27965
rect 27430 27928 27436 27940
rect 26528 27900 27436 27928
rect 22060 27888 22066 27900
rect 27430 27888 27436 27900
rect 27488 27888 27494 27940
rect 27908 27928 27936 28027
rect 28000 27996 28028 28104
rect 28810 28092 28816 28144
rect 28868 28092 28874 28144
rect 29181 28135 29239 28141
rect 29181 28101 29193 28135
rect 29227 28132 29239 28135
rect 29656 28132 29684 28172
rect 30466 28160 30472 28172
rect 30524 28200 30530 28212
rect 33962 28200 33968 28212
rect 30524 28172 33968 28200
rect 30524 28160 30530 28172
rect 33962 28160 33968 28172
rect 34020 28160 34026 28212
rect 37645 28203 37703 28209
rect 37645 28169 37657 28203
rect 37691 28200 37703 28203
rect 38010 28200 38016 28212
rect 37691 28172 38016 28200
rect 37691 28169 37703 28172
rect 37645 28163 37703 28169
rect 38010 28160 38016 28172
rect 38068 28160 38074 28212
rect 29227 28104 29684 28132
rect 29733 28135 29791 28141
rect 29227 28101 29239 28104
rect 29181 28095 29239 28101
rect 29733 28101 29745 28135
rect 29779 28132 29791 28135
rect 30190 28132 30196 28144
rect 29779 28104 30196 28132
rect 29779 28101 29791 28104
rect 29733 28095 29791 28101
rect 30190 28092 30196 28104
rect 30248 28092 30254 28144
rect 30374 28092 30380 28144
rect 30432 28132 30438 28144
rect 34054 28132 34060 28144
rect 30432 28104 34060 28132
rect 30432 28092 30438 28104
rect 34054 28092 34060 28104
rect 34112 28092 34118 28144
rect 36538 28092 36544 28144
rect 36596 28092 36602 28144
rect 36722 28092 36728 28144
rect 36780 28092 36786 28144
rect 37277 28135 37335 28141
rect 37277 28101 37289 28135
rect 37323 28132 37335 28135
rect 37550 28132 37556 28144
rect 37323 28104 37556 28132
rect 37323 28101 37335 28104
rect 37277 28095 37335 28101
rect 37550 28092 37556 28104
rect 37608 28092 37614 28144
rect 42153 28135 42211 28141
rect 42153 28101 42165 28135
rect 42199 28132 42211 28135
rect 42794 28132 42800 28144
rect 42199 28104 42800 28132
rect 42199 28101 42211 28104
rect 42153 28095 42211 28101
rect 42794 28092 42800 28104
rect 42852 28092 42858 28144
rect 42996 28104 44312 28132
rect 42996 28076 43024 28104
rect 28718 28024 28724 28076
rect 28776 28064 28782 28076
rect 28997 28067 29055 28073
rect 28997 28064 29009 28067
rect 28776 28036 29009 28064
rect 28776 28024 28782 28036
rect 28997 28033 29009 28036
rect 29043 28033 29055 28067
rect 28997 28027 29055 28033
rect 29914 28024 29920 28076
rect 29972 28024 29978 28076
rect 32677 28067 32735 28073
rect 32677 28064 32689 28067
rect 31726 28036 32689 28064
rect 31726 27996 31754 28036
rect 32677 28033 32689 28036
rect 32723 28033 32735 28067
rect 32677 28027 32735 28033
rect 37461 28067 37519 28073
rect 37461 28033 37473 28067
rect 37507 28064 37519 28067
rect 38010 28064 38016 28076
rect 37507 28036 38016 28064
rect 37507 28033 37519 28036
rect 37461 28027 37519 28033
rect 38010 28024 38016 28036
rect 38068 28024 38074 28076
rect 42978 28024 42984 28076
rect 43036 28024 43042 28076
rect 44284 28073 44312 28104
rect 43257 28067 43315 28073
rect 43257 28033 43269 28067
rect 43303 28033 43315 28067
rect 43257 28027 43315 28033
rect 44269 28067 44327 28073
rect 44269 28033 44281 28067
rect 44315 28033 44327 28067
rect 44269 28027 44327 28033
rect 28000 27968 31754 27996
rect 32766 27956 32772 28008
rect 32824 27956 32830 28008
rect 34054 27956 34060 28008
rect 34112 27996 34118 28008
rect 36906 27996 36912 28008
rect 34112 27968 36912 27996
rect 34112 27956 34118 27968
rect 36906 27956 36912 27968
rect 36964 27956 36970 28008
rect 37090 27956 37096 28008
rect 37148 27996 37154 28008
rect 41877 27999 41935 28005
rect 41877 27996 41889 27999
rect 37148 27968 41889 27996
rect 37148 27956 37154 27968
rect 41877 27965 41889 27968
rect 41923 27996 41935 27999
rect 43272 27996 43300 28027
rect 41923 27968 43300 27996
rect 41923 27965 41935 27968
rect 41877 27959 41935 27965
rect 35802 27928 35808 27940
rect 27908 27900 35808 27928
rect 35802 27888 35808 27900
rect 35860 27888 35866 27940
rect 44450 27888 44456 27940
rect 44508 27888 44514 27940
rect 6641 27863 6699 27869
rect 6641 27829 6653 27863
rect 6687 27860 6699 27863
rect 7190 27860 7196 27872
rect 6687 27832 7196 27860
rect 6687 27829 6699 27832
rect 6641 27823 6699 27829
rect 7190 27820 7196 27832
rect 7248 27820 7254 27872
rect 9858 27820 9864 27872
rect 9916 27860 9922 27872
rect 10410 27860 10416 27872
rect 9916 27832 10416 27860
rect 9916 27820 9922 27832
rect 10410 27820 10416 27832
rect 10468 27820 10474 27872
rect 13446 27820 13452 27872
rect 13504 27820 13510 27872
rect 13630 27820 13636 27872
rect 13688 27820 13694 27872
rect 14918 27820 14924 27872
rect 14976 27820 14982 27872
rect 15010 27820 15016 27872
rect 15068 27860 15074 27872
rect 15197 27863 15255 27869
rect 15197 27860 15209 27863
rect 15068 27832 15209 27860
rect 15068 27820 15074 27832
rect 15197 27829 15209 27832
rect 15243 27829 15255 27863
rect 15197 27823 15255 27829
rect 15654 27820 15660 27872
rect 15712 27820 15718 27872
rect 16114 27820 16120 27872
rect 16172 27820 16178 27872
rect 17954 27820 17960 27872
rect 18012 27860 18018 27872
rect 18601 27863 18659 27869
rect 18601 27860 18613 27863
rect 18012 27832 18613 27860
rect 18012 27820 18018 27832
rect 18601 27829 18613 27832
rect 18647 27860 18659 27863
rect 18966 27860 18972 27872
rect 18647 27832 18972 27860
rect 18647 27829 18659 27832
rect 18601 27823 18659 27829
rect 18966 27820 18972 27832
rect 19024 27820 19030 27872
rect 19058 27820 19064 27872
rect 19116 27820 19122 27872
rect 19702 27820 19708 27872
rect 19760 27860 19766 27872
rect 20438 27860 20444 27872
rect 19760 27832 20444 27860
rect 19760 27820 19766 27832
rect 20438 27820 20444 27832
rect 20496 27820 20502 27872
rect 20809 27863 20867 27869
rect 20809 27829 20821 27863
rect 20855 27860 20867 27863
rect 21542 27860 21548 27872
rect 20855 27832 21548 27860
rect 20855 27829 20867 27832
rect 20809 27823 20867 27829
rect 21542 27820 21548 27832
rect 21600 27820 21606 27872
rect 21634 27820 21640 27872
rect 21692 27860 21698 27872
rect 23293 27863 23351 27869
rect 23293 27860 23305 27863
rect 21692 27832 23305 27860
rect 21692 27820 21698 27832
rect 23293 27829 23305 27832
rect 23339 27829 23351 27863
rect 23293 27823 23351 27829
rect 23382 27820 23388 27872
rect 23440 27860 23446 27872
rect 24397 27863 24455 27869
rect 24397 27860 24409 27863
rect 23440 27832 24409 27860
rect 23440 27820 23446 27832
rect 24397 27829 24409 27832
rect 24443 27829 24455 27863
rect 24397 27823 24455 27829
rect 24857 27863 24915 27869
rect 24857 27829 24869 27863
rect 24903 27860 24915 27863
rect 26234 27860 26240 27872
rect 24903 27832 26240 27860
rect 24903 27829 24915 27832
rect 24857 27823 24915 27829
rect 26234 27820 26240 27832
rect 26292 27820 26298 27872
rect 26326 27820 26332 27872
rect 26384 27820 26390 27872
rect 26602 27820 26608 27872
rect 26660 27860 26666 27872
rect 26973 27863 27031 27869
rect 26973 27860 26985 27863
rect 26660 27832 26985 27860
rect 26660 27820 26666 27832
rect 26973 27829 26985 27832
rect 27019 27860 27031 27863
rect 27062 27860 27068 27872
rect 27019 27832 27068 27860
rect 27019 27829 27031 27832
rect 26973 27823 27031 27829
rect 27062 27820 27068 27832
rect 27120 27820 27126 27872
rect 27154 27820 27160 27872
rect 27212 27860 27218 27872
rect 27709 27863 27767 27869
rect 27709 27860 27721 27863
rect 27212 27832 27721 27860
rect 27212 27820 27218 27832
rect 27709 27829 27721 27832
rect 27755 27829 27767 27863
rect 27709 27823 27767 27829
rect 28902 27820 28908 27872
rect 28960 27860 28966 27872
rect 32677 27863 32735 27869
rect 32677 27860 32689 27863
rect 28960 27832 32689 27860
rect 28960 27820 28966 27832
rect 32677 27829 32689 27832
rect 32723 27829 32735 27863
rect 32677 27823 32735 27829
rect 33045 27863 33103 27869
rect 33045 27829 33057 27863
rect 33091 27860 33103 27863
rect 33134 27860 33140 27872
rect 33091 27832 33140 27860
rect 33091 27829 33103 27832
rect 33045 27823 33103 27829
rect 33134 27820 33140 27832
rect 33192 27820 33198 27872
rect 34698 27820 34704 27872
rect 34756 27860 34762 27872
rect 36538 27860 36544 27872
rect 34756 27832 36544 27860
rect 34756 27820 34762 27832
rect 36538 27820 36544 27832
rect 36596 27820 36602 27872
rect 36909 27863 36967 27869
rect 36909 27829 36921 27863
rect 36955 27860 36967 27863
rect 37458 27860 37464 27872
rect 36955 27832 37464 27860
rect 36955 27829 36967 27832
rect 36909 27823 36967 27829
rect 37458 27820 37464 27832
rect 37516 27820 37522 27872
rect 40034 27820 40040 27872
rect 40092 27860 40098 27872
rect 40770 27860 40776 27872
rect 40092 27832 40776 27860
rect 40092 27820 40098 27832
rect 40770 27820 40776 27832
rect 40828 27820 40834 27872
rect 42426 27820 42432 27872
rect 42484 27820 42490 27872
rect 42610 27820 42616 27872
rect 42668 27860 42674 27872
rect 43349 27863 43407 27869
rect 43349 27860 43361 27863
rect 42668 27832 43361 27860
rect 42668 27820 42674 27832
rect 43349 27829 43361 27832
rect 43395 27829 43407 27863
rect 43349 27823 43407 27829
rect 1104 27770 44896 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 44896 27770
rect 1104 27696 44896 27718
rect 5350 27616 5356 27668
rect 5408 27656 5414 27668
rect 5997 27659 6055 27665
rect 5997 27656 6009 27659
rect 5408 27628 6009 27656
rect 5408 27616 5414 27628
rect 5997 27625 6009 27628
rect 6043 27656 6055 27659
rect 6549 27659 6607 27665
rect 6549 27656 6561 27659
rect 6043 27628 6561 27656
rect 6043 27625 6055 27628
rect 5997 27619 6055 27625
rect 6549 27625 6561 27628
rect 6595 27656 6607 27659
rect 6595 27628 6684 27656
rect 6595 27625 6607 27628
rect 6549 27619 6607 27625
rect 6656 27588 6684 27628
rect 6730 27616 6736 27668
rect 6788 27616 6794 27668
rect 7558 27616 7564 27668
rect 7616 27656 7622 27668
rect 10137 27659 10195 27665
rect 7616 27628 9674 27656
rect 7616 27616 7622 27628
rect 7926 27588 7932 27600
rect 6656 27560 7932 27588
rect 7926 27548 7932 27560
rect 7984 27548 7990 27600
rect 9646 27588 9674 27628
rect 10137 27625 10149 27659
rect 10183 27656 10195 27659
rect 10410 27656 10416 27668
rect 10183 27628 10416 27656
rect 10183 27625 10195 27628
rect 10137 27619 10195 27625
rect 10410 27616 10416 27628
rect 10468 27656 10474 27668
rect 13357 27659 13415 27665
rect 10468 27628 11192 27656
rect 10468 27616 10474 27628
rect 10321 27591 10379 27597
rect 9646 27560 10272 27588
rect 6822 27520 6828 27532
rect 5828 27492 6828 27520
rect 5828 27461 5856 27492
rect 5813 27455 5871 27461
rect 5813 27421 5825 27455
rect 5859 27421 5871 27455
rect 5813 27415 5871 27421
rect 5994 27412 6000 27464
rect 6052 27412 6058 27464
rect 6380 27461 6408 27492
rect 6822 27480 6828 27492
rect 6880 27480 6886 27532
rect 9858 27480 9864 27532
rect 9916 27520 9922 27532
rect 9953 27523 10011 27529
rect 9953 27520 9965 27523
rect 9916 27492 9965 27520
rect 9916 27480 9922 27492
rect 9953 27489 9965 27492
rect 9999 27489 10011 27523
rect 10244 27520 10272 27560
rect 10321 27557 10333 27591
rect 10367 27588 10379 27591
rect 11054 27588 11060 27600
rect 10367 27560 11060 27588
rect 10367 27557 10379 27560
rect 10321 27551 10379 27557
rect 11054 27548 11060 27560
rect 11112 27548 11118 27600
rect 11164 27588 11192 27628
rect 13357 27625 13369 27659
rect 13403 27656 13415 27659
rect 18874 27656 18880 27668
rect 13403 27628 18880 27656
rect 13403 27625 13415 27628
rect 13357 27619 13415 27625
rect 18874 27616 18880 27628
rect 18932 27616 18938 27668
rect 19334 27616 19340 27668
rect 19392 27656 19398 27668
rect 19610 27656 19616 27668
rect 19392 27628 19616 27656
rect 19392 27616 19398 27628
rect 19610 27616 19616 27628
rect 19668 27656 19674 27668
rect 19797 27659 19855 27665
rect 19797 27656 19809 27659
rect 19668 27628 19809 27656
rect 19668 27616 19674 27628
rect 19797 27625 19809 27628
rect 19843 27625 19855 27659
rect 19797 27619 19855 27625
rect 21910 27616 21916 27668
rect 21968 27616 21974 27668
rect 22554 27616 22560 27668
rect 22612 27656 22618 27668
rect 26602 27656 26608 27668
rect 22612 27628 26608 27656
rect 22612 27616 22618 27628
rect 26602 27616 26608 27628
rect 26660 27616 26666 27668
rect 26694 27616 26700 27668
rect 26752 27616 26758 27668
rect 26878 27616 26884 27668
rect 26936 27616 26942 27668
rect 26973 27659 27031 27665
rect 26973 27625 26985 27659
rect 27019 27625 27031 27659
rect 26973 27619 27031 27625
rect 29825 27659 29883 27665
rect 29825 27625 29837 27659
rect 29871 27656 29883 27659
rect 31941 27659 31999 27665
rect 29871 27628 31892 27656
rect 29871 27625 29883 27628
rect 29825 27619 29883 27625
rect 13541 27591 13599 27597
rect 11164 27560 13492 27588
rect 13078 27520 13084 27532
rect 10244 27492 13084 27520
rect 9953 27483 10011 27489
rect 13078 27480 13084 27492
rect 13136 27480 13142 27532
rect 13262 27480 13268 27532
rect 13320 27480 13326 27532
rect 6365 27455 6423 27461
rect 6365 27421 6377 27455
rect 6411 27421 6423 27455
rect 6365 27415 6423 27421
rect 6549 27455 6607 27461
rect 6549 27421 6561 27455
rect 6595 27452 6607 27455
rect 8202 27452 8208 27464
rect 6595 27424 8208 27452
rect 6595 27421 6607 27424
rect 6549 27415 6607 27421
rect 5442 27344 5448 27396
rect 5500 27384 5506 27396
rect 6564 27384 6592 27415
rect 8202 27412 8208 27424
rect 8260 27412 8266 27464
rect 8754 27412 8760 27464
rect 8812 27452 8818 27464
rect 10137 27455 10195 27461
rect 10137 27452 10149 27455
rect 8812 27424 10149 27452
rect 8812 27412 8818 27424
rect 10137 27421 10149 27424
rect 10183 27421 10195 27455
rect 10137 27415 10195 27421
rect 12986 27412 12992 27464
rect 13044 27452 13050 27464
rect 13357 27455 13415 27461
rect 13357 27452 13369 27455
rect 13044 27424 13369 27452
rect 13044 27412 13050 27424
rect 13357 27421 13369 27424
rect 13403 27421 13415 27455
rect 13464 27452 13492 27560
rect 13541 27557 13553 27591
rect 13587 27588 13599 27591
rect 19702 27588 19708 27600
rect 13587 27560 19708 27588
rect 13587 27557 13599 27560
rect 13541 27551 13599 27557
rect 19702 27548 19708 27560
rect 19760 27548 19766 27600
rect 22373 27591 22431 27597
rect 19904 27560 22140 27588
rect 14550 27480 14556 27532
rect 14608 27520 14614 27532
rect 15194 27520 15200 27532
rect 14608 27492 15200 27520
rect 14608 27480 14614 27492
rect 15194 27480 15200 27492
rect 15252 27520 15258 27532
rect 17405 27523 17463 27529
rect 15252 27492 17356 27520
rect 15252 27480 15258 27492
rect 17328 27452 17356 27492
rect 17405 27489 17417 27523
rect 17451 27520 17463 27523
rect 17494 27520 17500 27532
rect 17451 27492 17500 27520
rect 17451 27489 17463 27492
rect 17405 27483 17463 27489
rect 17494 27480 17500 27492
rect 17552 27520 17558 27532
rect 19904 27520 19932 27560
rect 17552 27492 19932 27520
rect 19981 27523 20039 27529
rect 17552 27480 17558 27492
rect 19981 27489 19993 27523
rect 20027 27520 20039 27523
rect 20027 27492 20392 27520
rect 20027 27489 20039 27492
rect 19981 27483 20039 27489
rect 19610 27452 19616 27464
rect 13464 27424 17264 27452
rect 17328 27424 19616 27452
rect 13357 27415 13415 27421
rect 17236 27396 17264 27424
rect 19610 27412 19616 27424
rect 19668 27412 19674 27464
rect 19794 27412 19800 27464
rect 19852 27412 19858 27464
rect 20066 27455 20124 27461
rect 20066 27421 20078 27455
rect 20112 27421 20124 27455
rect 20066 27415 20124 27421
rect 5500 27356 6592 27384
rect 5500 27344 5506 27356
rect 9582 27344 9588 27396
rect 9640 27384 9646 27396
rect 9861 27387 9919 27393
rect 9861 27384 9873 27387
rect 9640 27356 9873 27384
rect 9640 27344 9646 27356
rect 9861 27353 9873 27356
rect 9907 27353 9919 27387
rect 9861 27347 9919 27353
rect 13078 27344 13084 27396
rect 13136 27344 13142 27396
rect 15378 27344 15384 27396
rect 15436 27384 15442 27396
rect 15749 27387 15807 27393
rect 15749 27384 15761 27387
rect 15436 27356 15761 27384
rect 15436 27344 15442 27356
rect 15749 27353 15761 27356
rect 15795 27353 15807 27387
rect 15749 27347 15807 27353
rect 15930 27344 15936 27396
rect 15988 27344 15994 27396
rect 16114 27344 16120 27396
rect 16172 27344 16178 27396
rect 16942 27344 16948 27396
rect 17000 27384 17006 27396
rect 17037 27387 17095 27393
rect 17037 27384 17049 27387
rect 17000 27356 17049 27384
rect 17000 27344 17006 27356
rect 17037 27353 17049 27356
rect 17083 27353 17095 27387
rect 17037 27347 17095 27353
rect 17218 27344 17224 27396
rect 17276 27344 17282 27396
rect 17402 27344 17408 27396
rect 17460 27384 17466 27396
rect 19978 27384 19984 27396
rect 17460 27356 19984 27384
rect 17460 27344 17466 27356
rect 19978 27344 19984 27356
rect 20036 27344 20042 27396
rect 6181 27319 6239 27325
rect 6181 27285 6193 27319
rect 6227 27316 6239 27319
rect 6914 27316 6920 27328
rect 6227 27288 6920 27316
rect 6227 27285 6239 27288
rect 6181 27279 6239 27285
rect 6914 27276 6920 27288
rect 6972 27276 6978 27328
rect 11238 27276 11244 27328
rect 11296 27316 11302 27328
rect 15102 27316 15108 27328
rect 11296 27288 15108 27316
rect 11296 27276 11302 27288
rect 15102 27276 15108 27288
rect 15160 27276 15166 27328
rect 16390 27276 16396 27328
rect 16448 27316 16454 27328
rect 20088 27316 20116 27415
rect 20364 27384 20392 27492
rect 20438 27480 20444 27532
rect 20496 27520 20502 27532
rect 22005 27523 22063 27529
rect 22005 27520 22017 27523
rect 20496 27492 22017 27520
rect 20496 27480 20502 27492
rect 22005 27489 22017 27492
rect 22051 27489 22063 27523
rect 22112 27520 22140 27560
rect 22373 27557 22385 27591
rect 22419 27588 22431 27591
rect 22922 27588 22928 27600
rect 22419 27560 22928 27588
rect 22419 27557 22431 27560
rect 22373 27551 22431 27557
rect 22922 27548 22928 27560
rect 22980 27548 22986 27600
rect 26786 27548 26792 27600
rect 26844 27588 26850 27600
rect 26988 27588 27016 27619
rect 26844 27560 27016 27588
rect 27341 27591 27399 27597
rect 26844 27548 26850 27560
rect 27341 27557 27353 27591
rect 27387 27588 27399 27591
rect 27798 27588 27804 27600
rect 27387 27560 27804 27588
rect 27387 27557 27399 27560
rect 27341 27551 27399 27557
rect 27798 27548 27804 27560
rect 27856 27548 27862 27600
rect 30466 27588 30472 27600
rect 28966 27560 30472 27588
rect 25406 27520 25412 27532
rect 22112 27492 25412 27520
rect 22005 27483 22063 27489
rect 25406 27480 25412 27492
rect 25464 27480 25470 27532
rect 26234 27480 26240 27532
rect 26292 27520 26298 27532
rect 26292 27492 27016 27520
rect 26292 27480 26298 27492
rect 22186 27412 22192 27464
rect 22244 27412 22250 27464
rect 25314 27412 25320 27464
rect 25372 27452 25378 27464
rect 26513 27455 26571 27461
rect 26513 27452 26525 27455
rect 25372 27424 26525 27452
rect 25372 27412 25378 27424
rect 26513 27421 26525 27424
rect 26559 27421 26571 27455
rect 26513 27415 26571 27421
rect 26697 27455 26755 27461
rect 26697 27421 26709 27455
rect 26743 27452 26755 27455
rect 26786 27452 26792 27464
rect 26743 27424 26792 27452
rect 26743 27421 26755 27424
rect 26697 27415 26755 27421
rect 26786 27412 26792 27424
rect 26844 27412 26850 27464
rect 26988 27461 27016 27492
rect 27522 27480 27528 27532
rect 27580 27520 27586 27532
rect 28966 27520 28994 27560
rect 30466 27548 30472 27560
rect 30524 27548 30530 27600
rect 31662 27548 31668 27600
rect 31720 27588 31726 27600
rect 31864 27588 31892 27628
rect 31941 27625 31953 27659
rect 31987 27656 31999 27659
rect 32030 27656 32036 27668
rect 31987 27628 32036 27656
rect 31987 27625 31999 27628
rect 31941 27619 31999 27625
rect 32030 27616 32036 27628
rect 32088 27616 32094 27668
rect 32858 27616 32864 27668
rect 32916 27656 32922 27668
rect 33137 27659 33195 27665
rect 33137 27656 33149 27659
rect 32916 27628 33149 27656
rect 32916 27616 32922 27628
rect 33137 27625 33149 27628
rect 33183 27625 33195 27659
rect 34054 27656 34060 27668
rect 33137 27619 33195 27625
rect 33336 27628 34060 27656
rect 33336 27588 33364 27628
rect 34054 27616 34060 27628
rect 34112 27616 34118 27668
rect 34698 27616 34704 27668
rect 34756 27616 34762 27668
rect 35158 27616 35164 27668
rect 35216 27616 35222 27668
rect 35526 27616 35532 27668
rect 35584 27616 35590 27668
rect 37182 27616 37188 27668
rect 37240 27656 37246 27668
rect 37240 27628 37320 27656
rect 37240 27616 37246 27628
rect 35253 27591 35311 27597
rect 35253 27588 35265 27591
rect 31720 27560 31800 27588
rect 31864 27560 33364 27588
rect 33428 27560 35265 27588
rect 31720 27548 31726 27560
rect 27580 27492 28994 27520
rect 27580 27480 27586 27492
rect 29454 27480 29460 27532
rect 29512 27520 29518 27532
rect 29641 27523 29699 27529
rect 29641 27520 29653 27523
rect 29512 27492 29653 27520
rect 29512 27480 29518 27492
rect 29641 27489 29653 27492
rect 29687 27520 29699 27523
rect 29730 27520 29736 27532
rect 29687 27492 29736 27520
rect 29687 27489 29699 27492
rect 29641 27483 29699 27489
rect 29730 27480 29736 27492
rect 29788 27480 29794 27532
rect 31772 27520 31800 27560
rect 32398 27520 32404 27532
rect 29840 27492 31708 27520
rect 26973 27455 27031 27461
rect 26973 27421 26985 27455
rect 27019 27421 27031 27455
rect 26973 27415 27031 27421
rect 27157 27455 27215 27461
rect 27157 27421 27169 27455
rect 27203 27452 27215 27455
rect 27706 27452 27712 27464
rect 27203 27424 27712 27452
rect 27203 27421 27215 27424
rect 27157 27415 27215 27421
rect 27706 27412 27712 27424
rect 27764 27412 27770 27464
rect 28810 27412 28816 27464
rect 28868 27452 28874 27464
rect 29840 27461 29868 27492
rect 31680 27464 31708 27492
rect 31772 27492 32404 27520
rect 29825 27455 29883 27461
rect 29825 27452 29837 27455
rect 28868 27424 29837 27452
rect 28868 27412 28874 27424
rect 29825 27421 29837 27424
rect 29871 27421 29883 27455
rect 31113 27455 31171 27461
rect 31113 27452 31125 27455
rect 29825 27415 29883 27421
rect 29932 27424 31125 27452
rect 21726 27384 21732 27396
rect 20364 27356 21732 27384
rect 21726 27344 21732 27356
rect 21784 27344 21790 27396
rect 21910 27344 21916 27396
rect 21968 27344 21974 27396
rect 23290 27344 23296 27396
rect 23348 27384 23354 27396
rect 24581 27387 24639 27393
rect 24581 27384 24593 27387
rect 23348 27356 24593 27384
rect 23348 27344 23354 27356
rect 24581 27353 24593 27356
rect 24627 27353 24639 27387
rect 24581 27347 24639 27353
rect 24765 27387 24823 27393
rect 24765 27353 24777 27387
rect 24811 27384 24823 27387
rect 26234 27384 26240 27396
rect 24811 27356 26240 27384
rect 24811 27353 24823 27356
rect 24765 27347 24823 27353
rect 26234 27344 26240 27356
rect 26292 27344 26298 27396
rect 26418 27344 26424 27396
rect 26476 27384 26482 27396
rect 29546 27384 29552 27396
rect 26476 27356 29552 27384
rect 26476 27344 26482 27356
rect 29546 27344 29552 27356
rect 29604 27344 29610 27396
rect 29932 27384 29960 27424
rect 31113 27421 31125 27424
rect 31159 27421 31171 27455
rect 31113 27415 31171 27421
rect 31297 27455 31355 27461
rect 31297 27421 31309 27455
rect 31343 27452 31355 27455
rect 31343 27424 31524 27452
rect 31343 27421 31355 27424
rect 31297 27415 31355 27421
rect 29656 27356 29960 27384
rect 16448 27288 20116 27316
rect 20257 27319 20315 27325
rect 16448 27276 16454 27288
rect 20257 27285 20269 27319
rect 20303 27316 20315 27319
rect 20714 27316 20720 27328
rect 20303 27288 20720 27316
rect 20303 27285 20315 27288
rect 20257 27279 20315 27285
rect 20714 27276 20720 27288
rect 20772 27276 20778 27328
rect 21082 27276 21088 27328
rect 21140 27316 21146 27328
rect 22370 27316 22376 27328
rect 21140 27288 22376 27316
rect 21140 27276 21146 27288
rect 22370 27276 22376 27288
rect 22428 27276 22434 27328
rect 24394 27276 24400 27328
rect 24452 27276 24458 27328
rect 24670 27276 24676 27328
rect 24728 27316 24734 27328
rect 29086 27316 29092 27328
rect 24728 27288 29092 27316
rect 24728 27276 24734 27288
rect 29086 27276 29092 27288
rect 29144 27276 29150 27328
rect 29362 27276 29368 27328
rect 29420 27316 29426 27328
rect 29656 27316 29684 27356
rect 30926 27344 30932 27396
rect 30984 27344 30990 27396
rect 31496 27384 31524 27424
rect 31662 27412 31668 27464
rect 31720 27412 31726 27464
rect 31772 27461 31800 27492
rect 32398 27480 32404 27492
rect 32456 27480 32462 27532
rect 32582 27480 32588 27532
rect 32640 27520 32646 27532
rect 33042 27520 33048 27532
rect 32640 27492 33048 27520
rect 32640 27480 32646 27492
rect 33042 27480 33048 27492
rect 33100 27480 33106 27532
rect 33318 27480 33324 27532
rect 33376 27480 33382 27532
rect 31757 27455 31815 27461
rect 31757 27421 31769 27455
rect 31803 27452 31815 27455
rect 31941 27455 31999 27461
rect 31803 27424 31837 27452
rect 31803 27421 31815 27424
rect 31757 27415 31815 27421
rect 31941 27421 31953 27455
rect 31987 27452 31999 27455
rect 32122 27452 32128 27464
rect 31987 27424 32128 27452
rect 31987 27421 31999 27424
rect 31941 27415 31999 27421
rect 32122 27412 32128 27424
rect 32180 27412 32186 27464
rect 33137 27455 33195 27461
rect 33137 27421 33149 27455
rect 33183 27452 33195 27455
rect 33226 27452 33232 27464
rect 33183 27424 33232 27452
rect 33183 27421 33195 27424
rect 33137 27415 33195 27421
rect 33226 27412 33232 27424
rect 33284 27412 33290 27464
rect 33428 27461 33456 27560
rect 35253 27557 35265 27560
rect 35299 27557 35311 27591
rect 37292 27588 37320 27628
rect 37366 27616 37372 27668
rect 37424 27616 37430 27668
rect 40586 27656 40592 27668
rect 37476 27628 40592 27656
rect 37476 27588 37504 27628
rect 37292 27560 37504 27588
rect 35253 27551 35311 27557
rect 34330 27480 34336 27532
rect 34388 27520 34394 27532
rect 34793 27523 34851 27529
rect 34793 27520 34805 27523
rect 34388 27492 34805 27520
rect 34388 27480 34394 27492
rect 34793 27489 34805 27492
rect 34839 27489 34851 27523
rect 34793 27483 34851 27489
rect 35342 27480 35348 27532
rect 35400 27520 35406 27532
rect 39868 27529 39896 27628
rect 40586 27616 40592 27628
rect 40644 27656 40650 27668
rect 41230 27656 41236 27668
rect 40644 27628 41236 27656
rect 40644 27616 40650 27628
rect 41230 27616 41236 27628
rect 41288 27616 41294 27668
rect 42058 27616 42064 27668
rect 42116 27616 42122 27668
rect 42426 27616 42432 27668
rect 42484 27656 42490 27668
rect 42521 27659 42579 27665
rect 42521 27656 42533 27659
rect 42484 27628 42533 27656
rect 42484 27616 42490 27628
rect 42521 27625 42533 27628
rect 42567 27625 42579 27659
rect 42521 27619 42579 27625
rect 35529 27523 35587 27529
rect 35529 27520 35541 27523
rect 35400 27492 35541 27520
rect 35400 27480 35406 27492
rect 35529 27489 35541 27492
rect 35575 27489 35587 27523
rect 35529 27483 35587 27489
rect 39853 27523 39911 27529
rect 39853 27489 39865 27523
rect 39899 27489 39911 27523
rect 39853 27483 39911 27489
rect 41969 27523 42027 27529
rect 41969 27489 41981 27523
rect 42015 27520 42027 27523
rect 42015 27492 44312 27520
rect 42015 27489 42027 27492
rect 41969 27483 42027 27489
rect 33413 27455 33471 27461
rect 33413 27421 33425 27455
rect 33459 27421 33471 27455
rect 34977 27455 35035 27461
rect 34977 27452 34989 27455
rect 33413 27415 33471 27421
rect 34072 27424 34989 27452
rect 34072 27384 34100 27424
rect 34977 27421 34989 27424
rect 35023 27452 35035 27455
rect 35437 27455 35495 27461
rect 35437 27452 35449 27455
rect 35023 27424 35449 27452
rect 35023 27421 35035 27424
rect 34977 27415 35035 27421
rect 35437 27421 35449 27424
rect 35483 27421 35495 27455
rect 36722 27452 36728 27464
rect 35437 27415 35495 27421
rect 35636 27424 36728 27452
rect 31496 27356 34100 27384
rect 34422 27344 34428 27396
rect 34480 27384 34486 27396
rect 34701 27387 34759 27393
rect 34701 27384 34713 27387
rect 34480 27356 34713 27384
rect 34480 27344 34486 27356
rect 34701 27353 34713 27356
rect 34747 27384 34759 27387
rect 35636 27384 35664 27424
rect 36722 27412 36728 27424
rect 36780 27452 36786 27464
rect 37369 27455 37427 27461
rect 37369 27452 37381 27455
rect 36780 27424 37381 27452
rect 36780 27412 36786 27424
rect 37369 27421 37381 27424
rect 37415 27421 37427 27455
rect 37369 27415 37427 27421
rect 37550 27412 37556 27464
rect 37608 27412 37614 27464
rect 40402 27412 40408 27464
rect 40460 27452 40466 27464
rect 41325 27455 41383 27461
rect 41325 27452 41337 27455
rect 40460 27424 41337 27452
rect 40460 27412 40466 27424
rect 41325 27421 41337 27424
rect 41371 27421 41383 27455
rect 41325 27415 41383 27421
rect 34747 27356 35664 27384
rect 35713 27387 35771 27393
rect 34747 27353 34759 27356
rect 34701 27347 34759 27353
rect 35713 27353 35725 27387
rect 35759 27384 35771 27387
rect 36078 27384 36084 27396
rect 35759 27356 36084 27384
rect 35759 27353 35771 27356
rect 35713 27347 35771 27353
rect 36078 27344 36084 27356
rect 36136 27344 36142 27396
rect 39574 27344 39580 27396
rect 39632 27384 39638 27396
rect 40098 27387 40156 27393
rect 40098 27384 40110 27387
rect 39632 27356 40110 27384
rect 39632 27344 39638 27356
rect 40098 27353 40110 27356
rect 40144 27353 40156 27387
rect 41984 27384 42012 27483
rect 42242 27412 42248 27464
rect 42300 27412 42306 27464
rect 42334 27412 42340 27464
rect 42392 27412 42398 27464
rect 42610 27412 42616 27464
rect 42668 27412 42674 27464
rect 44284 27461 44312 27492
rect 44269 27455 44327 27461
rect 44269 27421 44281 27455
rect 44315 27421 44327 27455
rect 44269 27415 44327 27421
rect 40098 27347 40156 27353
rect 41248 27356 42012 27384
rect 29420 27288 29684 27316
rect 30009 27319 30067 27325
rect 29420 27276 29426 27288
rect 30009 27285 30021 27319
rect 30055 27316 30067 27319
rect 31478 27316 31484 27328
rect 30055 27288 31484 27316
rect 30055 27285 30067 27288
rect 30009 27279 30067 27285
rect 31478 27276 31484 27288
rect 31536 27276 31542 27328
rect 32122 27276 32128 27328
rect 32180 27316 32186 27328
rect 32582 27316 32588 27328
rect 32180 27288 32588 27316
rect 32180 27276 32186 27288
rect 32582 27276 32588 27288
rect 32640 27276 32646 27328
rect 32858 27276 32864 27328
rect 32916 27316 32922 27328
rect 32953 27319 33011 27325
rect 32953 27316 32965 27319
rect 32916 27288 32965 27316
rect 32916 27276 32922 27288
rect 32953 27285 32965 27288
rect 32999 27285 33011 27319
rect 32953 27279 33011 27285
rect 33042 27276 33048 27328
rect 33100 27316 33106 27328
rect 34330 27316 34336 27328
rect 33100 27288 34336 27316
rect 33100 27276 33106 27288
rect 34330 27276 34336 27288
rect 34388 27276 34394 27328
rect 35802 27276 35808 27328
rect 35860 27316 35866 27328
rect 41248 27325 41276 27356
rect 37185 27319 37243 27325
rect 37185 27316 37197 27319
rect 35860 27288 37197 27316
rect 35860 27276 35866 27288
rect 37185 27285 37197 27288
rect 37231 27285 37243 27319
rect 37185 27279 37243 27285
rect 41233 27319 41291 27325
rect 41233 27285 41245 27319
rect 41279 27285 41291 27319
rect 41233 27279 41291 27285
rect 41322 27276 41328 27328
rect 41380 27316 41386 27328
rect 42628 27316 42656 27412
rect 41380 27288 42656 27316
rect 41380 27276 41386 27288
rect 44450 27276 44456 27328
rect 44508 27276 44514 27328
rect 1104 27226 44896 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 44896 27226
rect 1104 27152 44896 27174
rect 5994 27072 6000 27124
rect 6052 27112 6058 27124
rect 8754 27112 8760 27124
rect 6052 27084 8760 27112
rect 6052 27072 6058 27084
rect 8754 27072 8760 27084
rect 8812 27072 8818 27124
rect 13081 27115 13139 27121
rect 13081 27081 13093 27115
rect 13127 27112 13139 27115
rect 13262 27112 13268 27124
rect 13127 27084 13268 27112
rect 13127 27081 13139 27084
rect 13081 27075 13139 27081
rect 13262 27072 13268 27084
rect 13320 27072 13326 27124
rect 13372 27084 13768 27112
rect 8478 27004 8484 27056
rect 8536 27044 8542 27056
rect 12986 27044 12992 27056
rect 8536 27016 12992 27044
rect 8536 27004 8542 27016
rect 12986 27004 12992 27016
rect 13044 27004 13050 27056
rect 13372 27044 13400 27084
rect 13630 27044 13636 27056
rect 13096 27016 13400 27044
rect 13464 27016 13636 27044
rect 6822 26936 6828 26988
rect 6880 26976 6886 26988
rect 8021 26979 8079 26985
rect 8021 26976 8033 26979
rect 6880 26948 8033 26976
rect 6880 26936 6886 26948
rect 8021 26945 8033 26948
rect 8067 26945 8079 26979
rect 8021 26939 8079 26945
rect 8202 26936 8208 26988
rect 8260 26936 8266 26988
rect 10870 26936 10876 26988
rect 10928 26976 10934 26988
rect 11422 26976 11428 26988
rect 10928 26948 11428 26976
rect 10928 26936 10934 26948
rect 11422 26936 11428 26948
rect 11480 26976 11486 26988
rect 13096 26976 13124 27016
rect 13262 26985 13268 26988
rect 13248 26979 13268 26985
rect 13248 26976 13260 26979
rect 11480 26948 13124 26976
rect 13188 26948 13260 26976
rect 11480 26936 11486 26948
rect 8386 26868 8392 26920
rect 8444 26868 8450 26920
rect 13188 26908 13216 26948
rect 13248 26945 13260 26948
rect 13248 26939 13268 26945
rect 13262 26936 13268 26939
rect 13320 26936 13326 26988
rect 13357 26979 13415 26985
rect 13357 26945 13369 26979
rect 13403 26976 13415 26979
rect 13464 26976 13492 27016
rect 13630 27004 13636 27016
rect 13688 27004 13694 27056
rect 13740 27044 13768 27084
rect 15102 27072 15108 27124
rect 15160 27112 15166 27124
rect 18046 27112 18052 27124
rect 15160 27084 18052 27112
rect 15160 27072 15166 27084
rect 18046 27072 18052 27084
rect 18104 27072 18110 27124
rect 19702 27072 19708 27124
rect 19760 27072 19766 27124
rect 22005 27115 22063 27121
rect 20824 27084 21036 27112
rect 15470 27044 15476 27056
rect 13740 27016 15476 27044
rect 15470 27004 15476 27016
rect 15528 27044 15534 27056
rect 20824 27044 20852 27084
rect 15528 27016 20852 27044
rect 15528 27004 15534 27016
rect 20898 27004 20904 27056
rect 20956 27004 20962 27056
rect 21008 27044 21036 27084
rect 22005 27081 22017 27115
rect 22051 27112 22063 27115
rect 22186 27112 22192 27124
rect 22051 27084 22192 27112
rect 22051 27081 22063 27084
rect 22005 27075 22063 27081
rect 22186 27072 22192 27084
rect 22244 27072 22250 27124
rect 24670 27112 24676 27124
rect 24136 27084 24676 27112
rect 24136 27044 24164 27084
rect 24670 27072 24676 27084
rect 24728 27072 24734 27124
rect 25225 27115 25283 27121
rect 25225 27081 25237 27115
rect 25271 27112 25283 27115
rect 25271 27084 25360 27112
rect 25271 27081 25283 27084
rect 25225 27075 25283 27081
rect 21008 27016 24164 27044
rect 24394 27004 24400 27056
rect 24452 27044 24458 27056
rect 25332 27053 25360 27084
rect 25590 27072 25596 27124
rect 25648 27112 25654 27124
rect 26050 27112 26056 27124
rect 25648 27084 26056 27112
rect 25648 27072 25654 27084
rect 26050 27072 26056 27084
rect 26108 27072 26114 27124
rect 26694 27072 26700 27124
rect 26752 27112 26758 27124
rect 26752 27084 27016 27112
rect 26752 27072 26758 27084
rect 25317 27047 25375 27053
rect 24452 27016 25176 27044
rect 24452 27004 24458 27016
rect 13403 26948 13492 26976
rect 13541 26979 13599 26985
rect 13403 26945 13415 26948
rect 13357 26939 13415 26945
rect 13541 26945 13553 26979
rect 13587 26976 13599 26979
rect 14734 26976 14740 26988
rect 13587 26948 14740 26976
rect 13587 26945 13599 26948
rect 13541 26939 13599 26945
rect 14734 26936 14740 26948
rect 14792 26976 14798 26988
rect 15010 26976 15016 26988
rect 14792 26948 15016 26976
rect 14792 26936 14798 26948
rect 15010 26936 15016 26948
rect 15068 26936 15074 26988
rect 15194 26936 15200 26988
rect 15252 26976 15258 26988
rect 15381 26979 15439 26985
rect 15381 26976 15393 26979
rect 15252 26948 15393 26976
rect 15252 26936 15258 26948
rect 15381 26945 15393 26948
rect 15427 26945 15439 26979
rect 15381 26939 15439 26945
rect 15565 26979 15623 26985
rect 15565 26945 15577 26979
rect 15611 26945 15623 26979
rect 15565 26939 15623 26945
rect 8496 26880 13216 26908
rect 15580 26908 15608 26939
rect 15654 26936 15660 26988
rect 15712 26976 15718 26988
rect 19337 26979 19395 26985
rect 19337 26976 19349 26979
rect 15712 26948 19349 26976
rect 15712 26936 15718 26948
rect 19337 26945 19349 26948
rect 19383 26945 19395 26979
rect 19337 26939 19395 26945
rect 19518 26936 19524 26988
rect 19576 26936 19582 26988
rect 20622 26936 20628 26988
rect 20680 26936 20686 26988
rect 22189 26979 22247 26985
rect 22189 26976 22201 26979
rect 20732 26948 22201 26976
rect 17218 26908 17224 26920
rect 15580 26880 17224 26908
rect 7190 26800 7196 26852
rect 7248 26840 7254 26852
rect 8496 26840 8524 26880
rect 17218 26868 17224 26880
rect 17276 26868 17282 26920
rect 19426 26908 19432 26920
rect 18524 26880 19432 26908
rect 7248 26812 8524 26840
rect 7248 26800 7254 26812
rect 11422 26800 11428 26852
rect 11480 26840 11486 26852
rect 11698 26840 11704 26852
rect 11480 26812 11704 26840
rect 11480 26800 11486 26812
rect 11698 26800 11704 26812
rect 11756 26800 11762 26852
rect 18524 26784 18552 26880
rect 19426 26868 19432 26880
rect 19484 26908 19490 26920
rect 20732 26908 20760 26948
rect 22189 26945 22201 26948
rect 22235 26945 22247 26979
rect 22189 26939 22247 26945
rect 22465 26979 22523 26985
rect 22465 26945 22477 26979
rect 22511 26976 22523 26979
rect 24670 26976 24676 26988
rect 22511 26948 24676 26976
rect 22511 26945 22523 26948
rect 22465 26939 22523 26945
rect 24670 26936 24676 26948
rect 24728 26936 24734 26988
rect 24762 26936 24768 26988
rect 24820 26936 24826 26988
rect 25041 26979 25099 26985
rect 25041 26976 25053 26979
rect 24872 26948 25053 26976
rect 19484 26880 20760 26908
rect 20809 26911 20867 26917
rect 19484 26868 19490 26880
rect 20809 26877 20821 26911
rect 20855 26908 20867 26911
rect 21174 26908 21180 26920
rect 20855 26880 21180 26908
rect 20855 26877 20867 26880
rect 20809 26871 20867 26877
rect 21174 26868 21180 26880
rect 21232 26868 21238 26920
rect 22370 26868 22376 26920
rect 22428 26868 22434 26920
rect 23198 26868 23204 26920
rect 23256 26908 23262 26920
rect 24872 26908 24900 26948
rect 25041 26945 25053 26948
rect 25087 26945 25099 26979
rect 25148 26976 25176 27016
rect 25317 27013 25329 27047
rect 25363 27013 25375 27047
rect 25317 27007 25375 27013
rect 25958 27004 25964 27056
rect 26016 27044 26022 27056
rect 26988 27053 27016 27084
rect 27430 27072 27436 27124
rect 27488 27072 27494 27124
rect 27798 27072 27804 27124
rect 27856 27112 27862 27124
rect 33410 27112 33416 27124
rect 27856 27084 33416 27112
rect 27856 27072 27862 27084
rect 33410 27072 33416 27084
rect 33468 27072 33474 27124
rect 34514 27072 34520 27124
rect 34572 27112 34578 27124
rect 35345 27115 35403 27121
rect 35345 27112 35357 27115
rect 34572 27084 35357 27112
rect 34572 27072 34578 27084
rect 35345 27081 35357 27084
rect 35391 27081 35403 27115
rect 35345 27075 35403 27081
rect 37366 27072 37372 27124
rect 37424 27112 37430 27124
rect 37737 27115 37795 27121
rect 37737 27112 37749 27115
rect 37424 27084 37749 27112
rect 37424 27072 37430 27084
rect 37737 27081 37749 27084
rect 37783 27081 37795 27115
rect 37737 27075 37795 27081
rect 39574 27072 39580 27124
rect 39632 27072 39638 27124
rect 41046 27072 41052 27124
rect 41104 27112 41110 27124
rect 43165 27115 43223 27121
rect 43165 27112 43177 27115
rect 41104 27084 43177 27112
rect 41104 27072 41110 27084
rect 43165 27081 43177 27084
rect 43211 27081 43223 27115
rect 43165 27075 43223 27081
rect 26973 27047 27031 27053
rect 26016 27016 26648 27044
rect 26016 27004 26022 27016
rect 25593 26979 25651 26985
rect 25593 26976 25605 26979
rect 25148 26948 25605 26976
rect 25041 26939 25099 26945
rect 25593 26945 25605 26948
rect 25639 26945 25651 26979
rect 26329 26979 26387 26985
rect 26329 26976 26341 26979
rect 25593 26939 25651 26945
rect 26160 26948 26341 26976
rect 23256 26880 24900 26908
rect 23256 26868 23262 26880
rect 24946 26868 24952 26920
rect 25004 26868 25010 26920
rect 25498 26868 25504 26920
rect 25556 26868 25562 26920
rect 18598 26800 18604 26852
rect 18656 26840 18662 26852
rect 23290 26840 23296 26852
rect 18656 26812 23296 26840
rect 18656 26800 18662 26812
rect 7742 26732 7748 26784
rect 7800 26772 7806 26784
rect 12250 26772 12256 26784
rect 7800 26744 12256 26772
rect 7800 26732 7806 26744
rect 12250 26732 12256 26744
rect 12308 26732 12314 26784
rect 13541 26775 13599 26781
rect 13541 26741 13553 26775
rect 13587 26772 13599 26775
rect 13722 26772 13728 26784
rect 13587 26744 13728 26772
rect 13587 26741 13599 26744
rect 13541 26735 13599 26741
rect 13722 26732 13728 26744
rect 13780 26732 13786 26784
rect 15749 26775 15807 26781
rect 15749 26741 15761 26775
rect 15795 26772 15807 26775
rect 18506 26772 18512 26784
rect 15795 26744 18512 26772
rect 15795 26741 15807 26744
rect 15749 26735 15807 26741
rect 18506 26732 18512 26744
rect 18564 26732 18570 26784
rect 19058 26732 19064 26784
rect 19116 26772 19122 26784
rect 19337 26775 19395 26781
rect 19337 26772 19349 26775
rect 19116 26744 19349 26772
rect 19116 26732 19122 26744
rect 19337 26741 19349 26744
rect 19383 26741 19395 26775
rect 19337 26735 19395 26741
rect 20438 26732 20444 26784
rect 20496 26732 20502 26784
rect 20916 26781 20944 26812
rect 23290 26800 23296 26812
rect 23348 26800 23354 26852
rect 23934 26800 23940 26852
rect 23992 26840 23998 26852
rect 25130 26840 25136 26852
rect 23992 26812 25136 26840
rect 23992 26800 23998 26812
rect 25130 26800 25136 26812
rect 25188 26840 25194 26852
rect 26160 26849 26188 26948
rect 26329 26945 26341 26948
rect 26375 26945 26387 26979
rect 26329 26939 26387 26945
rect 26418 26936 26424 26988
rect 26476 26976 26482 26988
rect 26513 26979 26571 26985
rect 26513 26976 26525 26979
rect 26476 26948 26525 26976
rect 26476 26936 26482 26948
rect 26513 26945 26525 26948
rect 26559 26945 26571 26979
rect 26620 26976 26648 27016
rect 26973 27013 26985 27047
rect 27019 27013 27031 27047
rect 26973 27007 27031 27013
rect 27062 27004 27068 27056
rect 27120 27044 27126 27056
rect 27120 27016 27292 27044
rect 27120 27004 27126 27016
rect 27264 26985 27292 27016
rect 27614 27004 27620 27056
rect 27672 27044 27678 27056
rect 28537 27047 28595 27053
rect 28537 27044 28549 27047
rect 27672 27016 28549 27044
rect 27672 27004 27678 27016
rect 28537 27013 28549 27016
rect 28583 27013 28595 27047
rect 28537 27007 28595 27013
rect 31478 27004 31484 27056
rect 31536 27044 31542 27056
rect 31536 27016 35020 27044
rect 31536 27004 31542 27016
rect 27157 26979 27215 26985
rect 27157 26976 27169 26979
rect 26620 26948 27169 26976
rect 26513 26939 26571 26945
rect 27157 26945 27169 26948
rect 27203 26945 27215 26979
rect 27157 26939 27215 26945
rect 27249 26979 27307 26985
rect 27249 26945 27261 26979
rect 27295 26945 27307 26979
rect 27249 26939 27307 26945
rect 28442 26936 28448 26988
rect 28500 26976 28506 26988
rect 28813 26979 28871 26985
rect 28813 26976 28825 26979
rect 28500 26948 28825 26976
rect 28500 26936 28506 26948
rect 28813 26945 28825 26948
rect 28859 26976 28871 26979
rect 29362 26976 29368 26988
rect 28859 26948 29368 26976
rect 28859 26945 28871 26948
rect 28813 26939 28871 26945
rect 29362 26936 29368 26948
rect 29420 26936 29426 26988
rect 32122 26936 32128 26988
rect 32180 26936 32186 26988
rect 32401 26979 32459 26985
rect 32401 26945 32413 26979
rect 32447 26976 32459 26979
rect 32490 26976 32496 26988
rect 32447 26948 32496 26976
rect 32447 26945 32459 26948
rect 32401 26939 32459 26945
rect 32490 26936 32496 26948
rect 32548 26936 32554 26988
rect 32582 26936 32588 26988
rect 32640 26976 32646 26988
rect 34238 26976 34244 26988
rect 32640 26948 34244 26976
rect 32640 26936 32646 26948
rect 34238 26936 34244 26948
rect 34296 26936 34302 26988
rect 34330 26936 34336 26988
rect 34388 26976 34394 26988
rect 34425 26979 34483 26985
rect 34425 26976 34437 26979
rect 34388 26948 34437 26976
rect 34388 26936 34394 26948
rect 34425 26945 34437 26948
rect 34471 26945 34483 26979
rect 34425 26939 34483 26945
rect 34701 26979 34759 26985
rect 34701 26945 34713 26979
rect 34747 26976 34759 26979
rect 34790 26976 34796 26988
rect 34747 26948 34796 26976
rect 34747 26945 34759 26948
rect 34701 26939 34759 26945
rect 34790 26936 34796 26948
rect 34848 26936 34854 26988
rect 34992 26985 35020 27016
rect 35250 27004 35256 27056
rect 35308 27044 35314 27056
rect 35308 27016 37596 27044
rect 35308 27004 35314 27016
rect 34977 26979 35035 26985
rect 34977 26945 34989 26979
rect 35023 26945 35035 26979
rect 34977 26939 35035 26945
rect 35158 26936 35164 26988
rect 35216 26936 35222 26988
rect 35434 26936 35440 26988
rect 35492 26976 35498 26988
rect 37568 26985 37596 27016
rect 38746 27004 38752 27056
rect 38804 27044 38810 27056
rect 38804 27016 40540 27044
rect 38804 27004 38810 27016
rect 39776 26988 39804 27016
rect 40512 26988 40540 27016
rect 42426 27004 42432 27056
rect 42484 27004 42490 27056
rect 37277 26979 37335 26985
rect 37277 26976 37289 26979
rect 35492 26948 37289 26976
rect 35492 26936 35498 26948
rect 37277 26945 37289 26948
rect 37323 26945 37335 26979
rect 37277 26939 37335 26945
rect 37553 26979 37611 26985
rect 37553 26945 37565 26979
rect 37599 26945 37611 26979
rect 37553 26939 37611 26945
rect 39758 26936 39764 26988
rect 39816 26936 39822 26988
rect 39850 26936 39856 26988
rect 39908 26936 39914 26988
rect 40034 26936 40040 26988
rect 40092 26936 40098 26988
rect 40221 26979 40279 26985
rect 40221 26945 40233 26979
rect 40267 26976 40279 26979
rect 40402 26976 40408 26988
rect 40267 26948 40408 26976
rect 40267 26945 40279 26948
rect 40221 26939 40279 26945
rect 40402 26936 40408 26948
rect 40460 26936 40466 26988
rect 40494 26936 40500 26988
rect 40552 26936 40558 26988
rect 40770 26936 40776 26988
rect 40828 26936 40834 26988
rect 40954 26936 40960 26988
rect 41012 26936 41018 26988
rect 41046 26936 41052 26988
rect 41104 26976 41110 26988
rect 41509 26979 41567 26985
rect 41104 26948 41147 26976
rect 41104 26936 41110 26948
rect 41509 26945 41521 26979
rect 41555 26976 41567 26979
rect 42242 26976 42248 26988
rect 41555 26948 42248 26976
rect 41555 26945 41567 26948
rect 41509 26939 41567 26945
rect 28629 26911 28687 26917
rect 28629 26908 28641 26911
rect 27080 26880 28641 26908
rect 26145 26843 26203 26849
rect 26145 26840 26157 26843
rect 25188 26812 26157 26840
rect 25188 26800 25194 26812
rect 26145 26809 26157 26812
rect 26191 26809 26203 26843
rect 26145 26803 26203 26809
rect 26602 26800 26608 26852
rect 26660 26840 26666 26852
rect 27080 26840 27108 26880
rect 28368 26852 28396 26880
rect 28629 26877 28641 26880
rect 28675 26877 28687 26911
rect 28629 26871 28687 26877
rect 32030 26868 32036 26920
rect 32088 26908 32094 26920
rect 32217 26911 32275 26917
rect 32217 26908 32229 26911
rect 32088 26880 32229 26908
rect 32088 26868 32094 26880
rect 32217 26877 32229 26880
rect 32263 26877 32275 26911
rect 32217 26871 32275 26877
rect 34514 26868 34520 26920
rect 34572 26868 34578 26920
rect 35176 26908 35204 26936
rect 34992 26880 35204 26908
rect 27522 26840 27528 26852
rect 26660 26812 27108 26840
rect 27172 26812 27528 26840
rect 26660 26800 26666 26812
rect 20901 26775 20959 26781
rect 20901 26741 20913 26775
rect 20947 26741 20959 26775
rect 20901 26735 20959 26741
rect 22465 26775 22523 26781
rect 22465 26741 22477 26775
rect 22511 26772 22523 26775
rect 22554 26772 22560 26784
rect 22511 26744 22560 26772
rect 22511 26741 22523 26744
rect 22465 26735 22523 26741
rect 22554 26732 22560 26744
rect 22612 26732 22618 26784
rect 24210 26732 24216 26784
rect 24268 26772 24274 26784
rect 24578 26772 24584 26784
rect 24268 26744 24584 26772
rect 24268 26732 24274 26744
rect 24578 26732 24584 26744
rect 24636 26732 24642 26784
rect 25041 26775 25099 26781
rect 25041 26741 25053 26775
rect 25087 26772 25099 26775
rect 25222 26772 25228 26784
rect 25087 26744 25228 26772
rect 25087 26741 25099 26744
rect 25041 26735 25099 26741
rect 25222 26732 25228 26744
rect 25280 26732 25286 26784
rect 25590 26732 25596 26784
rect 25648 26732 25654 26784
rect 25774 26732 25780 26784
rect 25832 26732 25838 26784
rect 26234 26732 26240 26784
rect 26292 26772 26298 26784
rect 27172 26772 27200 26812
rect 27522 26800 27528 26812
rect 27580 26800 27586 26852
rect 28350 26800 28356 26852
rect 28408 26800 28414 26852
rect 28994 26800 29000 26852
rect 29052 26800 29058 26852
rect 34882 26800 34888 26852
rect 34940 26800 34946 26852
rect 26292 26744 27200 26772
rect 26292 26732 26298 26744
rect 27246 26732 27252 26784
rect 27304 26732 27310 26784
rect 28258 26732 28264 26784
rect 28316 26772 28322 26784
rect 28537 26775 28595 26781
rect 28537 26772 28549 26775
rect 28316 26744 28549 26772
rect 28316 26732 28322 26744
rect 28537 26741 28549 26744
rect 28583 26741 28595 26775
rect 28537 26735 28595 26741
rect 31018 26732 31024 26784
rect 31076 26772 31082 26784
rect 31386 26772 31392 26784
rect 31076 26744 31392 26772
rect 31076 26732 31082 26744
rect 31386 26732 31392 26744
rect 31444 26732 31450 26784
rect 31754 26732 31760 26784
rect 31812 26772 31818 26784
rect 32125 26775 32183 26781
rect 32125 26772 32137 26775
rect 31812 26744 32137 26772
rect 31812 26732 31818 26744
rect 32125 26741 32137 26744
rect 32171 26741 32183 26775
rect 32125 26735 32183 26741
rect 32582 26732 32588 26784
rect 32640 26732 32646 26784
rect 33134 26732 33140 26784
rect 33192 26772 33198 26784
rect 34425 26775 34483 26781
rect 34425 26772 34437 26775
rect 33192 26744 34437 26772
rect 33192 26732 33198 26744
rect 34425 26741 34437 26744
rect 34471 26741 34483 26775
rect 34425 26735 34483 26741
rect 34514 26732 34520 26784
rect 34572 26772 34578 26784
rect 34992 26772 35020 26880
rect 37182 26868 37188 26920
rect 37240 26908 37246 26920
rect 37369 26911 37427 26917
rect 37369 26908 37381 26911
rect 37240 26880 37381 26908
rect 37240 26868 37246 26880
rect 37369 26877 37381 26880
rect 37415 26877 37427 26911
rect 37369 26871 37427 26877
rect 39942 26868 39948 26920
rect 40000 26868 40006 26920
rect 40126 26868 40132 26920
rect 40184 26908 40190 26920
rect 40589 26911 40647 26917
rect 40589 26908 40601 26911
rect 40184 26880 40601 26908
rect 40184 26868 40190 26880
rect 40589 26877 40601 26880
rect 40635 26877 40647 26911
rect 40589 26871 40647 26877
rect 40678 26868 40684 26920
rect 40736 26868 40742 26920
rect 40788 26908 40816 26936
rect 41230 26908 41236 26920
rect 40788 26880 41236 26908
rect 41230 26868 41236 26880
rect 41288 26868 41294 26920
rect 41322 26868 41328 26920
rect 41380 26868 41386 26920
rect 35066 26800 35072 26852
rect 35124 26840 35130 26852
rect 41417 26843 41475 26849
rect 41417 26840 41429 26843
rect 35124 26812 41429 26840
rect 35124 26800 35130 26812
rect 41417 26809 41429 26812
rect 41463 26809 41475 26843
rect 41417 26803 41475 26809
rect 34572 26744 35020 26772
rect 35161 26775 35219 26781
rect 34572 26732 34578 26744
rect 35161 26741 35173 26775
rect 35207 26772 35219 26775
rect 35434 26772 35440 26784
rect 35207 26744 35440 26772
rect 35207 26741 35219 26744
rect 35161 26735 35219 26741
rect 35434 26732 35440 26744
rect 35492 26732 35498 26784
rect 36906 26732 36912 26784
rect 36964 26772 36970 26784
rect 37277 26775 37335 26781
rect 37277 26772 37289 26775
rect 36964 26744 37289 26772
rect 36964 26732 36970 26744
rect 37277 26741 37289 26744
rect 37323 26741 37335 26775
rect 37277 26735 37335 26741
rect 40310 26732 40316 26784
rect 40368 26732 40374 26784
rect 40494 26732 40500 26784
rect 40552 26772 40558 26784
rect 41524 26772 41552 26939
rect 42242 26936 42248 26948
rect 42300 26936 42306 26988
rect 44269 26979 44327 26985
rect 44269 26976 44281 26979
rect 42996 26948 44281 26976
rect 42058 26868 42064 26920
rect 42116 26908 42122 26920
rect 42996 26917 43024 26948
rect 44269 26945 44281 26948
rect 44315 26945 44327 26979
rect 44269 26939 44327 26945
rect 42981 26911 43039 26917
rect 42981 26908 42993 26911
rect 42116 26880 42993 26908
rect 42116 26868 42122 26880
rect 42981 26877 42993 26880
rect 43027 26877 43039 26911
rect 42981 26871 43039 26877
rect 43809 26911 43867 26917
rect 43809 26877 43821 26911
rect 43855 26877 43867 26911
rect 43809 26871 43867 26877
rect 43824 26840 43852 26871
rect 44266 26840 44272 26852
rect 43824 26812 44272 26840
rect 44266 26800 44272 26812
rect 44324 26800 44330 26852
rect 40552 26744 41552 26772
rect 41693 26775 41751 26781
rect 40552 26732 40558 26744
rect 41693 26741 41705 26775
rect 41739 26772 41751 26775
rect 42242 26772 42248 26784
rect 41739 26744 42248 26772
rect 41739 26741 41751 26744
rect 41693 26735 41751 26741
rect 42242 26732 42248 26744
rect 42300 26732 42306 26784
rect 44450 26732 44456 26784
rect 44508 26732 44514 26784
rect 1104 26682 44896 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 44896 26682
rect 1104 26608 44896 26630
rect 10781 26571 10839 26577
rect 10781 26537 10793 26571
rect 10827 26568 10839 26571
rect 10870 26568 10876 26580
rect 10827 26540 10876 26568
rect 10827 26537 10839 26540
rect 10781 26531 10839 26537
rect 10870 26528 10876 26540
rect 10928 26528 10934 26580
rect 10962 26528 10968 26580
rect 11020 26528 11026 26580
rect 11149 26571 11207 26577
rect 11149 26568 11161 26571
rect 11072 26540 11161 26568
rect 9858 26460 9864 26512
rect 9916 26500 9922 26512
rect 10318 26509 10324 26512
rect 10302 26503 10324 26509
rect 10302 26500 10314 26503
rect 9916 26472 10314 26500
rect 9916 26460 9922 26472
rect 10302 26469 10314 26472
rect 10302 26463 10324 26469
rect 10318 26460 10324 26463
rect 10376 26460 10382 26512
rect 10410 26460 10416 26512
rect 10468 26460 10474 26512
rect 11072 26500 11100 26540
rect 11149 26537 11161 26540
rect 11195 26537 11207 26571
rect 11149 26531 11207 26537
rect 11330 26528 11336 26580
rect 11388 26568 11394 26580
rect 12161 26571 12219 26577
rect 12161 26568 12173 26571
rect 11388 26540 12173 26568
rect 11388 26528 11394 26540
rect 12161 26537 12173 26540
rect 12207 26537 12219 26571
rect 12161 26531 12219 26537
rect 12618 26528 12624 26580
rect 12676 26528 12682 26580
rect 14458 26528 14464 26580
rect 14516 26568 14522 26580
rect 14826 26568 14832 26580
rect 14516 26540 14832 26568
rect 14516 26528 14522 26540
rect 14826 26528 14832 26540
rect 14884 26528 14890 26580
rect 15028 26540 15424 26568
rect 15028 26500 15056 26540
rect 10520 26472 11100 26500
rect 11716 26472 15056 26500
rect 15105 26503 15163 26509
rect 10134 26392 10140 26444
rect 10192 26432 10198 26444
rect 10520 26441 10548 26472
rect 11716 26444 11744 26472
rect 15105 26469 15117 26503
rect 15151 26469 15163 26503
rect 15396 26500 15424 26540
rect 15470 26528 15476 26580
rect 15528 26528 15534 26580
rect 15654 26528 15660 26580
rect 15712 26528 15718 26580
rect 17034 26528 17040 26580
rect 17092 26528 17098 26580
rect 17954 26568 17960 26580
rect 17236 26540 17960 26568
rect 16942 26500 16948 26512
rect 15396 26472 16948 26500
rect 15105 26463 15163 26469
rect 10505 26435 10563 26441
rect 10505 26432 10517 26435
rect 10192 26404 10517 26432
rect 10192 26392 10198 26404
rect 10505 26401 10517 26404
rect 10551 26401 10563 26435
rect 10505 26395 10563 26401
rect 11333 26435 11391 26441
rect 11333 26401 11345 26435
rect 11379 26432 11391 26435
rect 11422 26432 11428 26444
rect 11379 26404 11428 26432
rect 11379 26401 11391 26404
rect 11333 26395 11391 26401
rect 11422 26392 11428 26404
rect 11480 26392 11486 26444
rect 11698 26392 11704 26444
rect 11756 26392 11762 26444
rect 12342 26392 12348 26444
rect 12400 26392 12406 26444
rect 13998 26392 14004 26444
rect 14056 26432 14062 26444
rect 14550 26432 14556 26444
rect 14056 26404 14556 26432
rect 14056 26392 14062 26404
rect 14550 26392 14556 26404
rect 14608 26432 14614 26444
rect 14737 26435 14795 26441
rect 14737 26432 14749 26435
rect 14608 26404 14749 26432
rect 14608 26392 14614 26404
rect 14737 26401 14749 26404
rect 14783 26401 14795 26435
rect 14737 26395 14795 26401
rect 7926 26324 7932 26376
rect 7984 26364 7990 26376
rect 8021 26367 8079 26373
rect 8021 26364 8033 26367
rect 7984 26336 8033 26364
rect 7984 26324 7990 26336
rect 8021 26333 8033 26336
rect 8067 26333 8079 26367
rect 8021 26327 8079 26333
rect 8205 26367 8263 26373
rect 8205 26333 8217 26367
rect 8251 26364 8263 26367
rect 10318 26364 10324 26376
rect 8251 26336 10324 26364
rect 8251 26333 8263 26336
rect 8205 26327 8263 26333
rect 10318 26324 10324 26336
rect 10376 26324 10382 26376
rect 11146 26324 11152 26376
rect 11204 26324 11210 26376
rect 11517 26367 11575 26373
rect 11517 26364 11529 26367
rect 11348 26336 11529 26364
rect 6822 26256 6828 26308
rect 6880 26296 6886 26308
rect 7837 26299 7895 26305
rect 7837 26296 7849 26299
rect 6880 26268 7849 26296
rect 6880 26256 6886 26268
rect 7837 26265 7849 26268
rect 7883 26265 7895 26299
rect 7837 26259 7895 26265
rect 10137 26299 10195 26305
rect 10137 26265 10149 26299
rect 10183 26296 10195 26299
rect 11348 26296 11376 26336
rect 11517 26333 11529 26336
rect 11563 26364 11575 26367
rect 11716 26364 11744 26392
rect 11974 26364 11980 26376
rect 11563 26336 11744 26364
rect 11808 26336 11980 26364
rect 11563 26333 11575 26336
rect 11517 26327 11575 26333
rect 10183 26268 11376 26296
rect 11425 26299 11483 26305
rect 10183 26265 10195 26268
rect 10137 26259 10195 26265
rect 11425 26265 11437 26299
rect 11471 26296 11483 26299
rect 11606 26296 11612 26308
rect 11471 26268 11612 26296
rect 11471 26265 11483 26268
rect 11425 26259 11483 26265
rect 11606 26256 11612 26268
rect 11664 26256 11670 26308
rect 11701 26299 11759 26305
rect 11701 26265 11713 26299
rect 11747 26296 11759 26299
rect 11808 26296 11836 26336
rect 11974 26324 11980 26336
rect 12032 26324 12038 26376
rect 12250 26324 12256 26376
rect 12308 26364 12314 26376
rect 12437 26367 12495 26373
rect 12437 26364 12449 26367
rect 12308 26336 12449 26364
rect 12308 26324 12314 26336
rect 12437 26333 12449 26336
rect 12483 26364 12495 26367
rect 13814 26364 13820 26376
rect 12483 26336 13820 26364
rect 12483 26333 12495 26336
rect 12437 26327 12495 26333
rect 13814 26324 13820 26336
rect 13872 26324 13878 26376
rect 14568 26336 14872 26364
rect 11747 26268 11836 26296
rect 11885 26299 11943 26305
rect 11747 26265 11759 26268
rect 11701 26259 11759 26265
rect 11885 26265 11897 26299
rect 11931 26296 11943 26299
rect 12161 26299 12219 26305
rect 12161 26296 12173 26299
rect 11931 26268 12173 26296
rect 11931 26265 11943 26268
rect 11885 26259 11943 26265
rect 12161 26265 12173 26268
rect 12207 26296 12219 26299
rect 14568 26296 14596 26336
rect 12207 26268 14596 26296
rect 12207 26265 12219 26268
rect 12161 26259 12219 26265
rect 14642 26256 14648 26308
rect 14700 26256 14706 26308
rect 14844 26296 14872 26336
rect 14918 26324 14924 26376
rect 14976 26324 14982 26376
rect 15120 26364 15148 26463
rect 16942 26460 16948 26472
rect 17000 26460 17006 26512
rect 15286 26392 15292 26444
rect 15344 26392 15350 26444
rect 17037 26435 17095 26441
rect 17037 26401 17049 26435
rect 17083 26432 17095 26435
rect 17236 26432 17264 26540
rect 17954 26528 17960 26540
rect 18012 26528 18018 26580
rect 18138 26528 18144 26580
rect 18196 26528 18202 26580
rect 18874 26528 18880 26580
rect 18932 26528 18938 26580
rect 19334 26528 19340 26580
rect 19392 26568 19398 26580
rect 20441 26571 20499 26577
rect 20441 26568 20453 26571
rect 19392 26540 20453 26568
rect 19392 26528 19398 26540
rect 20441 26537 20453 26540
rect 20487 26537 20499 26571
rect 20441 26531 20499 26537
rect 20898 26528 20904 26580
rect 20956 26528 20962 26580
rect 22005 26571 22063 26577
rect 22005 26537 22017 26571
rect 22051 26568 22063 26571
rect 22094 26568 22100 26580
rect 22051 26540 22100 26568
rect 22051 26537 22063 26540
rect 22005 26531 22063 26537
rect 22094 26528 22100 26540
rect 22152 26528 22158 26580
rect 22186 26528 22192 26580
rect 22244 26528 22250 26580
rect 23198 26528 23204 26580
rect 23256 26568 23262 26580
rect 23750 26568 23756 26580
rect 23256 26540 23756 26568
rect 23256 26528 23262 26540
rect 23750 26528 23756 26540
rect 23808 26528 23814 26580
rect 25314 26528 25320 26580
rect 25372 26528 25378 26580
rect 25406 26528 25412 26580
rect 25464 26568 25470 26580
rect 26513 26571 26571 26577
rect 26513 26568 26525 26571
rect 25464 26540 26525 26568
rect 25464 26528 25470 26540
rect 26513 26537 26525 26540
rect 26559 26537 26571 26571
rect 26513 26531 26571 26537
rect 26602 26528 26608 26580
rect 26660 26568 26666 26580
rect 29825 26571 29883 26577
rect 29825 26568 29837 26571
rect 26660 26540 29837 26568
rect 26660 26528 26666 26540
rect 29825 26537 29837 26540
rect 29871 26568 29883 26571
rect 30374 26568 30380 26580
rect 29871 26540 30380 26568
rect 29871 26537 29883 26540
rect 29825 26531 29883 26537
rect 30374 26528 30380 26540
rect 30432 26528 30438 26580
rect 31294 26528 31300 26580
rect 31352 26568 31358 26580
rect 31573 26571 31631 26577
rect 31573 26568 31585 26571
rect 31352 26540 31585 26568
rect 31352 26528 31358 26540
rect 31573 26537 31585 26540
rect 31619 26537 31631 26571
rect 31573 26531 31631 26537
rect 32030 26528 32036 26580
rect 32088 26528 32094 26580
rect 32766 26568 32772 26580
rect 32508 26540 32772 26568
rect 17310 26460 17316 26512
rect 17368 26460 17374 26512
rect 17586 26460 17592 26512
rect 17644 26500 17650 26512
rect 18417 26503 18475 26509
rect 18417 26500 18429 26503
rect 17644 26472 18429 26500
rect 17644 26460 17650 26472
rect 18417 26469 18429 26472
rect 18463 26469 18475 26503
rect 21082 26500 21088 26512
rect 18417 26463 18475 26469
rect 18616 26472 21088 26500
rect 17083 26404 17264 26432
rect 17957 26435 18015 26441
rect 17083 26401 17095 26404
rect 17037 26395 17095 26401
rect 17957 26401 17969 26435
rect 18003 26432 18015 26435
rect 18616 26432 18644 26472
rect 21082 26460 21088 26472
rect 21140 26460 21146 26512
rect 23934 26500 23940 26512
rect 21744 26472 23940 26500
rect 18003 26404 18644 26432
rect 18003 26401 18015 26404
rect 17957 26395 18015 26401
rect 18782 26392 18788 26444
rect 18840 26392 18846 26444
rect 19610 26392 19616 26444
rect 19668 26432 19674 26444
rect 21744 26432 21772 26472
rect 23934 26460 23940 26472
rect 23992 26460 23998 26512
rect 24026 26460 24032 26512
rect 24084 26500 24090 26512
rect 26329 26503 26387 26509
rect 24084 26472 26280 26500
rect 24084 26460 24090 26472
rect 19668 26404 21772 26432
rect 19668 26392 19674 26404
rect 21818 26392 21824 26444
rect 21876 26392 21882 26444
rect 22094 26392 22100 26444
rect 22152 26432 22158 26444
rect 25958 26432 25964 26444
rect 22152 26404 25964 26432
rect 22152 26392 22158 26404
rect 25958 26392 25964 26404
rect 26016 26392 26022 26444
rect 26252 26432 26280 26472
rect 26329 26469 26341 26503
rect 26375 26500 26387 26503
rect 26418 26500 26424 26512
rect 26375 26472 26424 26500
rect 26375 26469 26387 26472
rect 26329 26463 26387 26469
rect 26418 26460 26424 26472
rect 26476 26460 26482 26512
rect 29454 26500 29460 26512
rect 27356 26472 29460 26500
rect 27356 26432 27384 26472
rect 29454 26460 29460 26472
rect 29512 26460 29518 26512
rect 32508 26500 32536 26540
rect 32766 26528 32772 26540
rect 32824 26528 32830 26580
rect 33134 26528 33140 26580
rect 33192 26528 33198 26580
rect 33413 26571 33471 26577
rect 33413 26537 33425 26571
rect 33459 26568 33471 26571
rect 35526 26568 35532 26580
rect 33459 26540 35532 26568
rect 33459 26537 33471 26540
rect 33413 26531 33471 26537
rect 35526 26528 35532 26540
rect 35584 26528 35590 26580
rect 37182 26528 37188 26580
rect 37240 26528 37246 26580
rect 37918 26528 37924 26580
rect 37976 26568 37982 26580
rect 40678 26568 40684 26580
rect 37976 26540 40684 26568
rect 37976 26528 37982 26540
rect 40678 26528 40684 26540
rect 40736 26528 40742 26580
rect 42058 26528 42064 26580
rect 42116 26528 42122 26580
rect 43533 26571 43591 26577
rect 43533 26537 43545 26571
rect 43579 26568 43591 26571
rect 44266 26568 44272 26580
rect 43579 26540 44272 26568
rect 43579 26537 43591 26540
rect 43533 26531 43591 26537
rect 44266 26528 44272 26540
rect 44324 26528 44330 26580
rect 31312 26472 32536 26500
rect 26252 26404 27384 26432
rect 27430 26392 27436 26444
rect 27488 26432 27494 26444
rect 29641 26435 29699 26441
rect 29641 26432 29653 26435
rect 27488 26404 29653 26432
rect 27488 26392 27494 26404
rect 29641 26401 29653 26404
rect 29687 26432 29699 26435
rect 29687 26404 31156 26432
rect 29687 26401 29699 26404
rect 29641 26395 29699 26401
rect 15197 26367 15255 26373
rect 15197 26364 15209 26367
rect 15120 26336 15209 26364
rect 15197 26333 15209 26336
rect 15243 26333 15255 26367
rect 15197 26327 15255 26333
rect 15470 26324 15476 26376
rect 15528 26324 15534 26376
rect 16482 26324 16488 26376
rect 16540 26364 16546 26376
rect 16945 26367 17003 26373
rect 16945 26364 16957 26367
rect 16540 26336 16957 26364
rect 16540 26324 16546 26336
rect 16945 26333 16957 26336
rect 16991 26364 17003 26367
rect 18141 26367 18199 26373
rect 16991 26358 18000 26364
rect 18141 26358 18153 26367
rect 16991 26336 18153 26358
rect 16991 26333 17003 26336
rect 16945 26327 17003 26333
rect 17972 26333 18153 26336
rect 18187 26333 18199 26367
rect 17972 26330 18199 26333
rect 18141 26327 18199 26330
rect 18506 26324 18512 26376
rect 18564 26364 18570 26376
rect 18601 26367 18659 26373
rect 18601 26364 18613 26367
rect 18564 26336 18613 26364
rect 18564 26324 18570 26336
rect 18601 26333 18613 26336
rect 18647 26333 18659 26367
rect 18601 26327 18659 26333
rect 20438 26324 20444 26376
rect 20496 26324 20502 26376
rect 20622 26324 20628 26376
rect 20680 26324 20686 26376
rect 20714 26324 20720 26376
rect 20772 26324 20778 26376
rect 21358 26324 21364 26376
rect 21416 26364 21422 26376
rect 22005 26367 22063 26373
rect 22005 26364 22017 26367
rect 21416 26336 22017 26364
rect 21416 26324 21422 26336
rect 22005 26333 22017 26336
rect 22051 26333 22063 26367
rect 24854 26364 24860 26376
rect 22005 26327 22063 26333
rect 23400 26336 24860 26364
rect 17865 26299 17923 26305
rect 17865 26296 17877 26299
rect 14844 26268 17877 26296
rect 17865 26265 17877 26268
rect 17911 26265 17923 26299
rect 17865 26259 17923 26265
rect 18877 26299 18935 26305
rect 18877 26265 18889 26299
rect 18923 26296 18935 26299
rect 19058 26296 19064 26308
rect 18923 26268 19064 26296
rect 18923 26265 18935 26268
rect 18877 26259 18935 26265
rect 19058 26256 19064 26268
rect 19116 26256 19122 26308
rect 19702 26256 19708 26308
rect 19760 26296 19766 26308
rect 21729 26299 21787 26305
rect 21729 26296 21741 26299
rect 19760 26268 21741 26296
rect 19760 26256 19766 26268
rect 21729 26265 21741 26268
rect 21775 26265 21787 26299
rect 21729 26259 21787 26265
rect 10870 26188 10876 26240
rect 10928 26228 10934 26240
rect 12526 26228 12532 26240
rect 10928 26200 12532 26228
rect 10928 26188 10934 26200
rect 12526 26188 12532 26200
rect 12584 26188 12590 26240
rect 12710 26188 12716 26240
rect 12768 26228 12774 26240
rect 15746 26228 15752 26240
rect 12768 26200 15752 26228
rect 12768 26188 12774 26200
rect 15746 26188 15752 26200
rect 15804 26188 15810 26240
rect 18325 26231 18383 26237
rect 18325 26197 18337 26231
rect 18371 26228 18383 26231
rect 18414 26228 18420 26240
rect 18371 26200 18420 26228
rect 18371 26197 18383 26200
rect 18325 26191 18383 26197
rect 18414 26188 18420 26200
rect 18472 26188 18478 26240
rect 18506 26188 18512 26240
rect 18564 26228 18570 26240
rect 23400 26228 23428 26336
rect 24854 26324 24860 26336
rect 24912 26324 24918 26376
rect 25314 26324 25320 26376
rect 25372 26364 25378 26376
rect 25501 26367 25559 26373
rect 25501 26364 25513 26367
rect 25372 26336 25513 26364
rect 25372 26324 25378 26336
rect 25501 26333 25513 26336
rect 25547 26333 25559 26367
rect 25501 26327 25559 26333
rect 25590 26324 25596 26376
rect 25648 26364 25654 26376
rect 25685 26367 25743 26373
rect 25685 26364 25697 26367
rect 25648 26336 25697 26364
rect 25648 26324 25654 26336
rect 25685 26333 25697 26336
rect 25731 26333 25743 26367
rect 25685 26327 25743 26333
rect 26513 26367 26571 26373
rect 26513 26333 26525 26367
rect 26559 26333 26571 26367
rect 26513 26327 26571 26333
rect 26697 26367 26755 26373
rect 26697 26333 26709 26367
rect 26743 26364 26755 26367
rect 26786 26364 26792 26376
rect 26743 26336 26792 26364
rect 26743 26333 26755 26336
rect 26697 26327 26755 26333
rect 23750 26256 23756 26308
rect 23808 26296 23814 26308
rect 26528 26296 26556 26327
rect 26786 26324 26792 26336
rect 26844 26324 26850 26376
rect 29825 26367 29883 26373
rect 29825 26364 29837 26367
rect 28966 26336 29837 26364
rect 23808 26268 26556 26296
rect 23808 26256 23814 26268
rect 18564 26200 23428 26228
rect 18564 26188 18570 26200
rect 23474 26188 23480 26240
rect 23532 26228 23538 26240
rect 28966 26228 28994 26336
rect 29825 26333 29837 26336
rect 29871 26364 29883 26367
rect 30742 26364 30748 26376
rect 29871 26336 30748 26364
rect 29871 26333 29883 26336
rect 29825 26327 29883 26333
rect 30742 26324 30748 26336
rect 30800 26324 30806 26376
rect 31128 26373 31156 26404
rect 31312 26373 31340 26472
rect 32582 26460 32588 26512
rect 32640 26500 32646 26512
rect 37645 26503 37703 26509
rect 32640 26472 37320 26500
rect 32640 26460 32646 26472
rect 31481 26435 31539 26441
rect 31481 26401 31493 26435
rect 31527 26432 31539 26435
rect 31757 26435 31815 26441
rect 31757 26432 31769 26435
rect 31527 26404 31769 26432
rect 31527 26401 31539 26404
rect 31481 26395 31539 26401
rect 31757 26401 31769 26404
rect 31803 26432 31815 26435
rect 31938 26432 31944 26444
rect 31803 26404 31944 26432
rect 31803 26401 31815 26404
rect 31757 26395 31815 26401
rect 31938 26392 31944 26404
rect 31996 26392 32002 26444
rect 33134 26392 33140 26444
rect 33192 26432 33198 26444
rect 33192 26404 33364 26432
rect 33192 26392 33198 26404
rect 31113 26367 31171 26373
rect 31113 26333 31125 26367
rect 31159 26333 31171 26367
rect 31113 26327 31171 26333
rect 31297 26367 31355 26373
rect 31297 26333 31309 26367
rect 31343 26333 31355 26367
rect 31846 26364 31852 26376
rect 31297 26327 31355 26333
rect 31404 26336 31852 26364
rect 29546 26256 29552 26308
rect 29604 26256 29610 26308
rect 31018 26256 31024 26308
rect 31076 26296 31082 26308
rect 31404 26296 31432 26336
rect 31846 26324 31852 26336
rect 31904 26324 31910 26376
rect 32674 26324 32680 26376
rect 32732 26364 32738 26376
rect 33045 26367 33103 26373
rect 33045 26364 33057 26367
rect 32732 26336 33057 26364
rect 32732 26324 32738 26336
rect 33045 26333 33057 26336
rect 33091 26333 33103 26367
rect 33045 26327 33103 26333
rect 33226 26324 33232 26376
rect 33284 26324 33290 26376
rect 33336 26364 33364 26404
rect 33410 26392 33416 26444
rect 33468 26432 33474 26444
rect 36906 26432 36912 26444
rect 33468 26404 36912 26432
rect 33468 26392 33474 26404
rect 36906 26392 36912 26404
rect 36964 26392 36970 26444
rect 37292 26432 37320 26472
rect 37645 26469 37657 26503
rect 37691 26500 37703 26503
rect 39114 26500 39120 26512
rect 37691 26472 39120 26500
rect 37691 26469 37703 26472
rect 37645 26463 37703 26469
rect 39114 26460 39120 26472
rect 39172 26460 39178 26512
rect 44082 26460 44088 26512
rect 44140 26500 44146 26512
rect 44453 26503 44511 26509
rect 44453 26500 44465 26503
rect 44140 26472 44465 26500
rect 44140 26460 44146 26472
rect 44453 26469 44465 26472
rect 44499 26469 44511 26503
rect 44453 26463 44511 26469
rect 39942 26432 39948 26444
rect 37016 26404 37228 26432
rect 37292 26404 39948 26432
rect 37016 26364 37044 26404
rect 33336 26336 37044 26364
rect 37200 26364 37228 26404
rect 39942 26392 39948 26404
rect 40000 26392 40006 26444
rect 40586 26392 40592 26444
rect 40644 26432 40650 26444
rect 40681 26435 40739 26441
rect 40681 26432 40693 26435
rect 40644 26404 40693 26432
rect 40644 26392 40650 26404
rect 40681 26401 40693 26404
rect 40727 26401 40739 26435
rect 40681 26395 40739 26401
rect 37369 26367 37427 26373
rect 37369 26364 37381 26367
rect 37200 26336 37381 26364
rect 37369 26333 37381 26336
rect 37415 26333 37427 26367
rect 37369 26327 37427 26333
rect 37458 26324 37464 26376
rect 37516 26324 37522 26376
rect 40310 26324 40316 26376
rect 40368 26364 40374 26376
rect 40937 26367 40995 26373
rect 40937 26364 40949 26367
rect 40368 26336 40949 26364
rect 40368 26324 40374 26336
rect 40937 26333 40949 26336
rect 40983 26333 40995 26367
rect 40937 26327 40995 26333
rect 41690 26324 41696 26376
rect 41748 26364 41754 26376
rect 42153 26367 42211 26373
rect 42153 26364 42165 26367
rect 41748 26336 42165 26364
rect 41748 26324 41754 26336
rect 42153 26333 42165 26336
rect 42199 26333 42211 26367
rect 42153 26327 42211 26333
rect 42242 26324 42248 26376
rect 42300 26364 42306 26376
rect 42409 26367 42467 26373
rect 42409 26364 42421 26367
rect 42300 26336 42421 26364
rect 42300 26324 42306 26336
rect 42409 26333 42421 26336
rect 42455 26333 42467 26367
rect 42409 26327 42467 26333
rect 43714 26324 43720 26376
rect 43772 26364 43778 26376
rect 44269 26367 44327 26373
rect 44269 26364 44281 26367
rect 43772 26336 44281 26364
rect 43772 26324 43778 26336
rect 44269 26333 44281 26336
rect 44315 26333 44327 26367
rect 44269 26327 44327 26333
rect 31076 26268 31432 26296
rect 31573 26299 31631 26305
rect 31076 26256 31082 26268
rect 31573 26265 31585 26299
rect 31619 26296 31631 26299
rect 31754 26296 31760 26308
rect 31619 26268 31760 26296
rect 31619 26265 31631 26268
rect 31573 26259 31631 26265
rect 31754 26256 31760 26268
rect 31812 26256 31818 26308
rect 32030 26256 32036 26308
rect 32088 26296 32094 26308
rect 32306 26296 32312 26308
rect 32088 26268 32312 26296
rect 32088 26256 32094 26268
rect 32306 26256 32312 26268
rect 32364 26256 32370 26308
rect 37185 26299 37243 26305
rect 37185 26296 37197 26299
rect 32416 26268 37197 26296
rect 23532 26200 28994 26228
rect 23532 26188 23538 26200
rect 29730 26188 29736 26240
rect 29788 26228 29794 26240
rect 30009 26231 30067 26237
rect 30009 26228 30021 26231
rect 29788 26200 30021 26228
rect 29788 26188 29794 26200
rect 30009 26197 30021 26200
rect 30055 26197 30067 26231
rect 30009 26191 30067 26197
rect 30926 26188 30932 26240
rect 30984 26228 30990 26240
rect 32416 26228 32444 26268
rect 37185 26265 37197 26268
rect 37231 26265 37243 26299
rect 40126 26296 40132 26308
rect 37185 26259 37243 26265
rect 37292 26268 40132 26296
rect 30984 26200 32444 26228
rect 30984 26188 30990 26200
rect 34698 26188 34704 26240
rect 34756 26228 34762 26240
rect 35434 26228 35440 26240
rect 34756 26200 35440 26228
rect 34756 26188 34762 26200
rect 35434 26188 35440 26200
rect 35492 26188 35498 26240
rect 36906 26188 36912 26240
rect 36964 26228 36970 26240
rect 37292 26228 37320 26268
rect 40126 26256 40132 26268
rect 40184 26256 40190 26308
rect 36964 26200 37320 26228
rect 36964 26188 36970 26200
rect 1104 26138 44896 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 44896 26138
rect 1104 26064 44896 26086
rect 5442 26024 5448 26036
rect 5000 25996 5448 26024
rect 5000 25888 5028 25996
rect 5442 25984 5448 25996
rect 5500 25984 5506 26036
rect 8205 26027 8263 26033
rect 8205 25993 8217 26027
rect 8251 26024 8263 26027
rect 9401 26027 9459 26033
rect 8251 25996 8984 26024
rect 8251 25993 8263 25996
rect 8205 25987 8263 25993
rect 5077 25959 5135 25965
rect 5077 25925 5089 25959
rect 5123 25956 5135 25959
rect 5350 25956 5356 25968
rect 5123 25928 5356 25956
rect 5123 25925 5135 25928
rect 5077 25919 5135 25925
rect 5350 25916 5356 25928
rect 5408 25916 5414 25968
rect 8956 25965 8984 25996
rect 9401 25993 9413 26027
rect 9447 26024 9459 26027
rect 10870 26024 10876 26036
rect 9447 25996 10876 26024
rect 9447 25993 9459 25996
rect 9401 25987 9459 25993
rect 10870 25984 10876 25996
rect 10928 25984 10934 26036
rect 12434 25984 12440 26036
rect 12492 26024 12498 26036
rect 13078 26024 13084 26036
rect 12492 25996 13084 26024
rect 12492 25984 12498 25996
rect 13078 25984 13084 25996
rect 13136 25984 13142 26036
rect 16482 25984 16488 26036
rect 16540 25984 16546 26036
rect 17218 25984 17224 26036
rect 17276 26024 17282 26036
rect 18506 26024 18512 26036
rect 17276 25996 18512 26024
rect 17276 25984 17282 25996
rect 18506 25984 18512 25996
rect 18564 25984 18570 26036
rect 21818 25984 21824 26036
rect 21876 25984 21882 26036
rect 24949 26027 25007 26033
rect 23216 25996 24532 26024
rect 8941 25959 8999 25965
rect 8941 25925 8953 25959
rect 8987 25925 8999 25959
rect 8941 25919 8999 25925
rect 10502 25916 10508 25968
rect 10560 25956 10566 25968
rect 10560 25928 12434 25956
rect 10560 25916 10566 25928
rect 5166 25888 5172 25900
rect 5000 25860 5172 25888
rect 5166 25848 5172 25860
rect 5224 25888 5230 25900
rect 5261 25891 5319 25897
rect 5261 25888 5273 25891
rect 5224 25860 5273 25888
rect 5224 25848 5230 25860
rect 5261 25857 5273 25860
rect 5307 25857 5319 25891
rect 5261 25851 5319 25857
rect 5442 25848 5448 25900
rect 5500 25848 5506 25900
rect 7098 25848 7104 25900
rect 7156 25888 7162 25900
rect 7742 25888 7748 25900
rect 7156 25860 7748 25888
rect 7156 25848 7162 25860
rect 7742 25848 7748 25860
rect 7800 25848 7806 25900
rect 7834 25848 7840 25900
rect 7892 25888 7898 25900
rect 8021 25891 8079 25897
rect 8021 25888 8033 25891
rect 7892 25860 8033 25888
rect 7892 25848 7898 25860
rect 8021 25857 8033 25860
rect 8067 25857 8079 25891
rect 8021 25851 8079 25857
rect 9214 25848 9220 25900
rect 9272 25848 9278 25900
rect 9858 25848 9864 25900
rect 9916 25888 9922 25900
rect 10137 25891 10195 25897
rect 10137 25888 10149 25891
rect 9916 25860 10149 25888
rect 9916 25848 9922 25860
rect 10137 25857 10149 25860
rect 10183 25857 10195 25891
rect 10137 25851 10195 25857
rect 10226 25848 10232 25900
rect 10284 25888 10290 25900
rect 10321 25891 10379 25897
rect 10321 25888 10333 25891
rect 10284 25860 10333 25888
rect 10284 25848 10290 25860
rect 10321 25857 10333 25860
rect 10367 25857 10379 25891
rect 10321 25851 10379 25857
rect 10594 25848 10600 25900
rect 10652 25848 10658 25900
rect 10870 25848 10876 25900
rect 10928 25848 10934 25900
rect 11974 25848 11980 25900
rect 12032 25848 12038 25900
rect 12250 25848 12256 25900
rect 12308 25848 12314 25900
rect 7650 25780 7656 25832
rect 7708 25820 7714 25832
rect 7852 25820 7880 25848
rect 7708 25792 7880 25820
rect 7708 25780 7714 25792
rect 7926 25780 7932 25832
rect 7984 25780 7990 25832
rect 9030 25780 9036 25832
rect 9088 25780 9094 25832
rect 10686 25780 10692 25832
rect 10744 25820 10750 25832
rect 12069 25823 12127 25829
rect 12069 25820 12081 25823
rect 10744 25792 12081 25820
rect 10744 25780 10750 25792
rect 12069 25789 12081 25792
rect 12115 25789 12127 25823
rect 12406 25820 12434 25928
rect 12526 25916 12532 25968
rect 12584 25956 12590 25968
rect 19334 25956 19340 25968
rect 12584 25928 19340 25956
rect 12584 25916 12590 25928
rect 19334 25916 19340 25928
rect 19392 25916 19398 25968
rect 23216 25965 23244 25996
rect 23201 25959 23259 25965
rect 23201 25925 23213 25959
rect 23247 25925 23259 25959
rect 23201 25919 23259 25925
rect 23750 25916 23756 25968
rect 23808 25916 23814 25968
rect 24504 25965 24532 25996
rect 24949 25993 24961 26027
rect 24995 26024 25007 26027
rect 25038 26024 25044 26036
rect 24995 25996 25044 26024
rect 24995 25993 25007 25996
rect 24949 25987 25007 25993
rect 25038 25984 25044 25996
rect 25096 25984 25102 26036
rect 25406 25984 25412 26036
rect 25464 26024 25470 26036
rect 25590 26024 25596 26036
rect 25464 25996 25596 26024
rect 25464 25984 25470 25996
rect 25590 25984 25596 25996
rect 25648 25984 25654 26036
rect 32030 26024 32036 26036
rect 31864 25996 32036 26024
rect 24489 25959 24547 25965
rect 24489 25925 24501 25959
rect 24535 25925 24547 25959
rect 24489 25919 24547 25925
rect 24854 25916 24860 25968
rect 24912 25956 24918 25968
rect 28445 25959 28503 25965
rect 24912 25928 26924 25956
rect 24912 25916 24918 25928
rect 12894 25848 12900 25900
rect 12952 25848 12958 25900
rect 13078 25848 13084 25900
rect 13136 25888 13142 25900
rect 13630 25888 13636 25900
rect 13136 25860 13636 25888
rect 13136 25848 13142 25860
rect 13630 25848 13636 25860
rect 13688 25848 13694 25900
rect 14734 25848 14740 25900
rect 14792 25848 14798 25900
rect 14826 25848 14832 25900
rect 14884 25888 14890 25900
rect 14921 25891 14979 25897
rect 14921 25888 14933 25891
rect 14884 25860 14933 25888
rect 14884 25848 14890 25860
rect 14921 25857 14933 25860
rect 14967 25888 14979 25891
rect 15746 25888 15752 25900
rect 14967 25860 15752 25888
rect 14967 25857 14979 25860
rect 14921 25851 14979 25857
rect 15746 25848 15752 25860
rect 15804 25848 15810 25900
rect 16022 25848 16028 25900
rect 16080 25888 16086 25900
rect 16117 25891 16175 25897
rect 16117 25888 16129 25891
rect 16080 25860 16129 25888
rect 16080 25848 16086 25860
rect 16117 25857 16129 25860
rect 16163 25857 16175 25891
rect 16117 25851 16175 25857
rect 16301 25891 16359 25897
rect 16301 25857 16313 25891
rect 16347 25857 16359 25891
rect 16301 25851 16359 25857
rect 12986 25820 12992 25832
rect 12406 25792 12992 25820
rect 12069 25783 12127 25789
rect 12986 25780 12992 25792
rect 13044 25780 13050 25832
rect 15764 25820 15792 25848
rect 16316 25820 16344 25851
rect 20714 25848 20720 25900
rect 20772 25888 20778 25900
rect 22189 25891 22247 25897
rect 22189 25888 22201 25891
rect 20772 25860 22201 25888
rect 20772 25848 20778 25860
rect 22189 25857 22201 25860
rect 22235 25857 22247 25891
rect 22189 25851 22247 25857
rect 22646 25848 22652 25900
rect 22704 25888 22710 25900
rect 22833 25891 22891 25897
rect 22833 25888 22845 25891
rect 22704 25860 22845 25888
rect 22704 25848 22710 25860
rect 22833 25857 22845 25860
rect 22879 25857 22891 25891
rect 22833 25851 22891 25857
rect 23017 25891 23075 25897
rect 23017 25857 23029 25891
rect 23063 25888 23075 25891
rect 23290 25888 23296 25900
rect 23063 25860 23296 25888
rect 23063 25857 23075 25860
rect 23017 25851 23075 25857
rect 23290 25848 23296 25860
rect 23348 25848 23354 25900
rect 23474 25848 23480 25900
rect 23532 25848 23538 25900
rect 23569 25891 23627 25897
rect 23569 25857 23581 25891
rect 23615 25857 23627 25891
rect 23569 25851 23627 25857
rect 15764 25792 16344 25820
rect 18874 25780 18880 25832
rect 18932 25820 18938 25832
rect 22094 25820 22100 25832
rect 18932 25792 22100 25820
rect 18932 25780 18938 25792
rect 22094 25780 22100 25792
rect 22152 25780 22158 25832
rect 23584 25820 23612 25851
rect 23658 25848 23664 25900
rect 23716 25888 23722 25900
rect 23845 25891 23903 25897
rect 23845 25888 23857 25891
rect 23716 25860 23857 25888
rect 23716 25848 23722 25860
rect 23845 25857 23857 25860
rect 23891 25857 23903 25891
rect 24121 25891 24179 25897
rect 24121 25888 24133 25891
rect 23845 25851 23903 25857
rect 23952 25860 24133 25888
rect 23499 25792 23612 25820
rect 10318 25712 10324 25764
rect 10376 25752 10382 25764
rect 10870 25752 10876 25764
rect 10376 25724 10876 25752
rect 10376 25712 10382 25724
rect 10870 25712 10876 25724
rect 10928 25712 10934 25764
rect 11057 25755 11115 25761
rect 11057 25721 11069 25755
rect 11103 25752 11115 25755
rect 15102 25752 15108 25764
rect 11103 25724 15108 25752
rect 11103 25721 11115 25724
rect 11057 25715 11115 25721
rect 15102 25712 15108 25724
rect 15160 25712 15166 25764
rect 19518 25712 19524 25764
rect 19576 25752 19582 25764
rect 23293 25755 23351 25761
rect 23293 25752 23305 25755
rect 19576 25724 23305 25752
rect 19576 25712 19582 25724
rect 23293 25721 23305 25724
rect 23339 25721 23351 25755
rect 23293 25715 23351 25721
rect 8021 25687 8079 25693
rect 8021 25653 8033 25687
rect 8067 25684 8079 25687
rect 8202 25684 8208 25696
rect 8067 25656 8208 25684
rect 8067 25653 8079 25656
rect 8021 25647 8079 25653
rect 8202 25644 8208 25656
rect 8260 25644 8266 25696
rect 9217 25687 9275 25693
rect 9217 25653 9229 25687
rect 9263 25684 9275 25687
rect 10042 25684 10048 25696
rect 9263 25656 10048 25684
rect 9263 25653 9275 25656
rect 9217 25647 9275 25653
rect 10042 25644 10048 25656
rect 10100 25644 10106 25696
rect 10134 25644 10140 25696
rect 10192 25684 10198 25696
rect 10597 25687 10655 25693
rect 10597 25684 10609 25687
rect 10192 25656 10609 25684
rect 10192 25644 10198 25656
rect 10597 25653 10609 25656
rect 10643 25653 10655 25687
rect 10597 25647 10655 25653
rect 11882 25644 11888 25696
rect 11940 25684 11946 25696
rect 11977 25687 12035 25693
rect 11977 25684 11989 25687
rect 11940 25656 11989 25684
rect 11940 25644 11946 25656
rect 11977 25653 11989 25656
rect 12023 25653 12035 25687
rect 11977 25647 12035 25653
rect 13081 25687 13139 25693
rect 13081 25653 13093 25687
rect 13127 25684 13139 25687
rect 13170 25684 13176 25696
rect 13127 25656 13176 25684
rect 13127 25653 13139 25656
rect 13081 25647 13139 25653
rect 13170 25644 13176 25656
rect 13228 25644 13234 25696
rect 13262 25644 13268 25696
rect 13320 25644 13326 25696
rect 15013 25687 15071 25693
rect 15013 25653 15025 25687
rect 15059 25684 15071 25687
rect 15194 25684 15200 25696
rect 15059 25656 15200 25684
rect 15059 25653 15071 25656
rect 15013 25647 15071 25653
rect 15194 25644 15200 25656
rect 15252 25644 15258 25696
rect 22189 25687 22247 25693
rect 22189 25653 22201 25687
rect 22235 25684 22247 25687
rect 22370 25684 22376 25696
rect 22235 25656 22376 25684
rect 22235 25653 22247 25656
rect 22189 25647 22247 25653
rect 22370 25644 22376 25656
rect 22428 25684 22434 25696
rect 22830 25684 22836 25696
rect 22428 25656 22836 25684
rect 22428 25644 22434 25656
rect 22830 25644 22836 25656
rect 22888 25644 22894 25696
rect 23198 25644 23204 25696
rect 23256 25684 23262 25696
rect 23499 25684 23527 25792
rect 23952 25752 23980 25860
rect 24121 25857 24133 25860
rect 24167 25888 24179 25891
rect 24167 25860 24716 25888
rect 24167 25857 24179 25860
rect 24121 25851 24179 25857
rect 24029 25823 24087 25829
rect 24029 25789 24041 25823
rect 24075 25820 24087 25823
rect 24075 25792 24256 25820
rect 24075 25789 24087 25792
rect 24029 25783 24087 25789
rect 23676 25724 23980 25752
rect 23676 25693 23704 25724
rect 23256 25656 23527 25684
rect 23661 25687 23719 25693
rect 23256 25644 23262 25656
rect 23661 25653 23673 25687
rect 23707 25653 23719 25687
rect 23661 25647 23719 25653
rect 23750 25644 23756 25696
rect 23808 25684 23814 25696
rect 23845 25687 23903 25693
rect 23845 25684 23857 25687
rect 23808 25656 23857 25684
rect 23808 25644 23814 25656
rect 23845 25653 23857 25656
rect 23891 25653 23903 25687
rect 24228 25684 24256 25792
rect 24394 25780 24400 25832
rect 24452 25820 24458 25832
rect 24581 25823 24639 25829
rect 24581 25820 24593 25823
rect 24452 25792 24593 25820
rect 24452 25780 24458 25792
rect 24581 25789 24593 25792
rect 24627 25789 24639 25823
rect 24688 25820 24716 25860
rect 24762 25848 24768 25900
rect 24820 25848 24826 25900
rect 24946 25848 24952 25900
rect 25004 25888 25010 25900
rect 26234 25888 26240 25900
rect 25004 25860 26240 25888
rect 25004 25848 25010 25860
rect 26234 25848 26240 25860
rect 26292 25888 26298 25900
rect 26421 25891 26479 25897
rect 26421 25888 26433 25891
rect 26292 25860 26433 25888
rect 26292 25848 26298 25860
rect 26421 25857 26433 25860
rect 26467 25857 26479 25891
rect 26421 25851 26479 25857
rect 26602 25848 26608 25900
rect 26660 25848 26666 25900
rect 26786 25848 26792 25900
rect 26844 25848 26850 25900
rect 26896 25888 26924 25928
rect 28445 25925 28457 25959
rect 28491 25956 28503 25959
rect 31864 25956 31892 25996
rect 32030 25984 32036 25996
rect 32088 25984 32094 26036
rect 32766 25984 32772 26036
rect 32824 26024 32830 26036
rect 32824 25996 34744 26024
rect 32824 25984 32830 25996
rect 28491 25928 31892 25956
rect 28491 25925 28503 25928
rect 28445 25919 28503 25925
rect 31938 25916 31944 25968
rect 31996 25956 32002 25968
rect 34716 25956 34744 25996
rect 34790 25984 34796 26036
rect 34848 25984 34854 26036
rect 36630 25984 36636 26036
rect 36688 26024 36694 26036
rect 36906 26024 36912 26036
rect 36688 25996 36912 26024
rect 36688 25984 36694 25996
rect 36906 25984 36912 25996
rect 36964 25984 36970 26036
rect 37090 25984 37096 26036
rect 37148 26024 37154 26036
rect 37458 26024 37464 26036
rect 37148 25996 37464 26024
rect 37148 25984 37154 25996
rect 37458 25984 37464 25996
rect 37516 25984 37522 26036
rect 38933 25959 38991 25965
rect 38933 25956 38945 25959
rect 31996 25928 33824 25956
rect 31996 25916 32002 25928
rect 28629 25891 28687 25897
rect 28629 25888 28641 25891
rect 26896 25860 28641 25888
rect 28629 25857 28641 25860
rect 28675 25857 28687 25891
rect 28629 25851 28687 25857
rect 28721 25891 28779 25897
rect 28721 25857 28733 25891
rect 28767 25888 28779 25891
rect 29178 25888 29184 25900
rect 28767 25860 29184 25888
rect 28767 25857 28779 25860
rect 28721 25851 28779 25857
rect 29178 25848 29184 25860
rect 29236 25848 29242 25900
rect 32858 25848 32864 25900
rect 32916 25848 32922 25900
rect 33796 25897 33824 25928
rect 34256 25928 34560 25956
rect 34716 25928 38945 25956
rect 33781 25891 33839 25897
rect 33781 25857 33793 25891
rect 33827 25857 33839 25891
rect 33781 25851 33839 25857
rect 25590 25820 25596 25832
rect 24688 25792 25596 25820
rect 24581 25783 24639 25789
rect 25590 25780 25596 25792
rect 25648 25780 25654 25832
rect 26050 25780 26056 25832
rect 26108 25820 26114 25832
rect 31478 25820 31484 25832
rect 26108 25792 31484 25820
rect 26108 25780 26114 25792
rect 31478 25780 31484 25792
rect 31536 25780 31542 25832
rect 32030 25780 32036 25832
rect 32088 25820 32094 25832
rect 32953 25823 33011 25829
rect 32953 25820 32965 25823
rect 32088 25792 32965 25820
rect 32088 25780 32094 25792
rect 32953 25789 32965 25792
rect 32999 25789 33011 25823
rect 32953 25783 33011 25789
rect 33134 25780 33140 25832
rect 33192 25820 33198 25832
rect 33873 25823 33931 25829
rect 33873 25820 33885 25823
rect 33192 25792 33885 25820
rect 33192 25780 33198 25792
rect 33873 25789 33885 25792
rect 33919 25789 33931 25823
rect 33873 25783 33931 25789
rect 24305 25755 24363 25761
rect 24305 25721 24317 25755
rect 24351 25752 24363 25755
rect 31938 25752 31944 25764
rect 24351 25724 31944 25752
rect 24351 25721 24363 25724
rect 24305 25715 24363 25721
rect 31938 25712 31944 25724
rect 31996 25712 32002 25764
rect 34256 25752 34284 25928
rect 34422 25848 34428 25900
rect 34480 25848 34486 25900
rect 34532 25888 34560 25928
rect 35345 25891 35403 25897
rect 35345 25888 35357 25891
rect 34532 25860 35357 25888
rect 35345 25857 35357 25860
rect 35391 25857 35403 25891
rect 35345 25851 35403 25857
rect 36078 25848 36084 25900
rect 36136 25888 36142 25900
rect 37277 25891 37335 25897
rect 37277 25888 37289 25891
rect 36136 25860 37289 25888
rect 36136 25848 36142 25860
rect 37277 25857 37289 25860
rect 37323 25857 37335 25891
rect 37277 25851 37335 25857
rect 37458 25848 37464 25900
rect 37516 25848 37522 25900
rect 38381 25891 38439 25897
rect 38381 25888 38393 25891
rect 37660 25860 38393 25888
rect 34517 25823 34575 25829
rect 34517 25789 34529 25823
rect 34563 25789 34575 25823
rect 34517 25783 34575 25789
rect 33796 25724 34284 25752
rect 34532 25752 34560 25783
rect 35158 25780 35164 25832
rect 35216 25820 35222 25832
rect 35437 25823 35495 25829
rect 35437 25820 35449 25823
rect 35216 25792 35449 25820
rect 35216 25780 35222 25792
rect 35437 25789 35449 25792
rect 35483 25789 35495 25823
rect 35437 25783 35495 25789
rect 36446 25752 36452 25764
rect 34532 25724 36452 25752
rect 24394 25684 24400 25696
rect 24228 25656 24400 25684
rect 23845 25647 23903 25653
rect 24394 25644 24400 25656
rect 24452 25644 24458 25696
rect 24486 25644 24492 25696
rect 24544 25644 24550 25696
rect 25038 25644 25044 25696
rect 25096 25684 25102 25696
rect 27614 25684 27620 25696
rect 25096 25656 27620 25684
rect 25096 25644 25102 25656
rect 27614 25644 27620 25656
rect 27672 25644 27678 25696
rect 28258 25644 28264 25696
rect 28316 25684 28322 25696
rect 28445 25687 28503 25693
rect 28445 25684 28457 25687
rect 28316 25656 28457 25684
rect 28316 25644 28322 25656
rect 28445 25653 28457 25656
rect 28491 25684 28503 25687
rect 28534 25684 28540 25696
rect 28491 25656 28540 25684
rect 28491 25653 28503 25656
rect 28445 25647 28503 25653
rect 28534 25644 28540 25656
rect 28592 25644 28598 25696
rect 28905 25687 28963 25693
rect 28905 25653 28917 25687
rect 28951 25684 28963 25687
rect 29546 25684 29552 25696
rect 28951 25656 29552 25684
rect 28951 25653 28963 25656
rect 28905 25647 28963 25653
rect 29546 25644 29552 25656
rect 29604 25644 29610 25696
rect 32306 25644 32312 25696
rect 32364 25684 32370 25696
rect 32861 25687 32919 25693
rect 32861 25684 32873 25687
rect 32364 25656 32873 25684
rect 32364 25644 32370 25656
rect 32861 25653 32873 25656
rect 32907 25653 32919 25687
rect 32861 25647 32919 25653
rect 33229 25687 33287 25693
rect 33229 25653 33241 25687
rect 33275 25684 33287 25687
rect 33410 25684 33416 25696
rect 33275 25656 33416 25684
rect 33275 25653 33287 25656
rect 33229 25647 33287 25653
rect 33410 25644 33416 25656
rect 33468 25644 33474 25696
rect 33594 25644 33600 25696
rect 33652 25684 33658 25696
rect 33796 25693 33824 25724
rect 33781 25687 33839 25693
rect 33781 25684 33793 25687
rect 33652 25656 33793 25684
rect 33652 25644 33658 25656
rect 33781 25653 33793 25656
rect 33827 25653 33839 25687
rect 33781 25647 33839 25653
rect 34146 25644 34152 25696
rect 34204 25644 34210 25696
rect 34425 25687 34483 25693
rect 34425 25653 34437 25687
rect 34471 25684 34483 25687
rect 34514 25684 34520 25696
rect 34471 25656 34520 25684
rect 34471 25653 34483 25656
rect 34425 25647 34483 25653
rect 34514 25644 34520 25656
rect 34572 25644 34578 25696
rect 35360 25693 35388 25724
rect 36446 25712 36452 25724
rect 36504 25712 36510 25764
rect 37274 25712 37280 25764
rect 37332 25752 37338 25764
rect 37660 25761 37688 25860
rect 38381 25857 38393 25860
rect 38427 25857 38439 25891
rect 38381 25851 38439 25857
rect 38562 25848 38568 25900
rect 38620 25888 38626 25900
rect 38657 25891 38715 25897
rect 38657 25888 38669 25891
rect 38620 25860 38669 25888
rect 38620 25848 38626 25860
rect 38657 25857 38669 25860
rect 38703 25857 38715 25891
rect 38657 25851 38715 25857
rect 37918 25780 37924 25832
rect 37976 25820 37982 25832
rect 38473 25823 38531 25829
rect 38473 25820 38485 25823
rect 37976 25792 38485 25820
rect 37976 25780 37982 25792
rect 38473 25789 38485 25792
rect 38519 25789 38531 25823
rect 38473 25783 38531 25789
rect 37645 25755 37703 25761
rect 37645 25752 37657 25755
rect 37332 25724 37657 25752
rect 37332 25712 37338 25724
rect 37645 25721 37657 25724
rect 37691 25721 37703 25755
rect 37645 25715 37703 25721
rect 35345 25687 35403 25693
rect 35345 25653 35357 25687
rect 35391 25653 35403 25687
rect 35345 25647 35403 25653
rect 35434 25644 35440 25696
rect 35492 25684 35498 25696
rect 35713 25687 35771 25693
rect 35713 25684 35725 25687
rect 35492 25656 35725 25684
rect 35492 25644 35498 25656
rect 35713 25653 35725 25656
rect 35759 25653 35771 25687
rect 35713 25647 35771 25653
rect 37458 25644 37464 25696
rect 37516 25684 37522 25696
rect 37737 25687 37795 25693
rect 37737 25684 37749 25687
rect 37516 25656 37749 25684
rect 37516 25644 37522 25656
rect 37737 25653 37749 25656
rect 37783 25653 37795 25687
rect 37737 25647 37795 25653
rect 38378 25644 38384 25696
rect 38436 25644 38442 25696
rect 38764 25684 38792 25928
rect 38933 25925 38945 25928
rect 38979 25925 38991 25959
rect 38933 25919 38991 25925
rect 39114 25916 39120 25968
rect 39172 25916 39178 25968
rect 41690 25956 41696 25968
rect 40512 25928 41696 25956
rect 39393 25891 39451 25897
rect 39393 25857 39405 25891
rect 39439 25888 39451 25891
rect 39850 25888 39856 25900
rect 39439 25860 39856 25888
rect 39439 25857 39451 25860
rect 39393 25851 39451 25857
rect 39850 25848 39856 25860
rect 39908 25848 39914 25900
rect 40512 25897 40540 25928
rect 41690 25916 41696 25928
rect 41748 25916 41754 25968
rect 40497 25891 40555 25897
rect 40497 25857 40509 25891
rect 40543 25857 40555 25891
rect 40497 25851 40555 25857
rect 40586 25848 40592 25900
rect 40644 25888 40650 25900
rect 40753 25891 40811 25897
rect 40753 25888 40765 25891
rect 40644 25860 40765 25888
rect 40644 25848 40650 25860
rect 40753 25857 40765 25860
rect 40799 25857 40811 25891
rect 40753 25851 40811 25857
rect 39209 25823 39267 25829
rect 39209 25789 39221 25823
rect 39255 25789 39267 25823
rect 39209 25783 39267 25789
rect 43073 25823 43131 25829
rect 43073 25789 43085 25823
rect 43119 25820 43131 25823
rect 44174 25820 44180 25832
rect 43119 25792 44180 25820
rect 43119 25789 43131 25792
rect 43073 25783 43131 25789
rect 38841 25755 38899 25761
rect 38841 25721 38853 25755
rect 38887 25752 38899 25755
rect 39224 25752 39252 25783
rect 38887 25724 39252 25752
rect 38887 25721 38899 25724
rect 38841 25715 38899 25721
rect 41506 25712 41512 25764
rect 41564 25752 41570 25764
rect 42429 25755 42487 25761
rect 42429 25752 42441 25755
rect 41564 25724 42441 25752
rect 41564 25712 41570 25724
rect 42429 25721 42441 25724
rect 42475 25721 42487 25755
rect 42429 25715 42487 25721
rect 39117 25687 39175 25693
rect 39117 25684 39129 25687
rect 38764 25656 39129 25684
rect 39117 25653 39129 25656
rect 39163 25653 39175 25687
rect 39117 25647 39175 25653
rect 39577 25687 39635 25693
rect 39577 25653 39589 25687
rect 39623 25684 39635 25687
rect 40678 25684 40684 25696
rect 39623 25656 40684 25684
rect 39623 25653 39635 25656
rect 39577 25647 39635 25653
rect 40678 25644 40684 25656
rect 40736 25644 40742 25696
rect 41877 25687 41935 25693
rect 41877 25653 41889 25687
rect 41923 25684 41935 25687
rect 43088 25684 43116 25783
rect 44174 25780 44180 25792
rect 44232 25780 44238 25832
rect 41923 25656 43116 25684
rect 41923 25653 41935 25656
rect 41877 25647 41935 25653
rect 1104 25594 44896 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 44896 25594
rect 1104 25520 44896 25542
rect 5258 25440 5264 25492
rect 5316 25440 5322 25492
rect 5718 25440 5724 25492
rect 5776 25440 5782 25492
rect 10042 25440 10048 25492
rect 10100 25480 10106 25492
rect 10229 25483 10287 25489
rect 10229 25480 10241 25483
rect 10100 25452 10241 25480
rect 10100 25440 10106 25452
rect 10229 25449 10241 25452
rect 10275 25480 10287 25483
rect 10275 25452 16160 25480
rect 10275 25449 10287 25452
rect 10229 25443 10287 25449
rect 11698 25372 11704 25424
rect 11756 25412 11762 25424
rect 12250 25412 12256 25424
rect 11756 25384 12256 25412
rect 11756 25372 11762 25384
rect 12250 25372 12256 25384
rect 12308 25412 12314 25424
rect 16022 25412 16028 25424
rect 12308 25384 16028 25412
rect 12308 25372 12314 25384
rect 16022 25372 16028 25384
rect 16080 25372 16086 25424
rect 16132 25412 16160 25452
rect 16298 25440 16304 25492
rect 16356 25480 16362 25492
rect 19518 25480 19524 25492
rect 16356 25452 19524 25480
rect 16356 25440 16362 25452
rect 19518 25440 19524 25452
rect 19576 25440 19582 25492
rect 19702 25440 19708 25492
rect 19760 25440 19766 25492
rect 19794 25440 19800 25492
rect 19852 25480 19858 25492
rect 20349 25483 20407 25489
rect 20349 25480 20361 25483
rect 19852 25452 20361 25480
rect 19852 25440 19858 25452
rect 20349 25449 20361 25452
rect 20395 25449 20407 25483
rect 20349 25443 20407 25449
rect 20622 25440 20628 25492
rect 20680 25480 20686 25492
rect 20809 25483 20867 25489
rect 20809 25480 20821 25483
rect 20680 25452 20821 25480
rect 20680 25440 20686 25452
rect 20809 25449 20821 25452
rect 20855 25449 20867 25483
rect 20809 25443 20867 25449
rect 22370 25440 22376 25492
rect 22428 25480 22434 25492
rect 22554 25480 22560 25492
rect 22428 25452 22560 25480
rect 22428 25440 22434 25452
rect 22554 25440 22560 25452
rect 22612 25440 22618 25492
rect 23569 25483 23627 25489
rect 23569 25449 23581 25483
rect 23615 25449 23627 25483
rect 23569 25443 23627 25449
rect 17678 25412 17684 25424
rect 16132 25384 17684 25412
rect 17678 25372 17684 25384
rect 17736 25372 17742 25424
rect 19610 25372 19616 25424
rect 19668 25412 19674 25424
rect 19978 25412 19984 25424
rect 19668 25384 19984 25412
rect 19668 25372 19674 25384
rect 19978 25372 19984 25384
rect 20036 25412 20042 25424
rect 20530 25412 20536 25424
rect 20036 25384 20536 25412
rect 20036 25372 20042 25384
rect 20530 25372 20536 25384
rect 20588 25372 20594 25424
rect 23584 25412 23612 25443
rect 23750 25440 23756 25492
rect 23808 25440 23814 25492
rect 24854 25480 24860 25492
rect 23860 25452 24860 25480
rect 23860 25412 23888 25452
rect 24854 25440 24860 25452
rect 24912 25440 24918 25492
rect 25038 25440 25044 25492
rect 25096 25440 25102 25492
rect 25498 25440 25504 25492
rect 25556 25440 25562 25492
rect 25590 25440 25596 25492
rect 25648 25480 25654 25492
rect 28721 25483 28779 25489
rect 28721 25480 28733 25483
rect 25648 25452 28733 25480
rect 25648 25440 25654 25452
rect 28721 25449 28733 25452
rect 28767 25449 28779 25483
rect 28721 25443 28779 25449
rect 29822 25440 29828 25492
rect 29880 25480 29886 25492
rect 30098 25480 30104 25492
rect 29880 25452 30104 25480
rect 29880 25440 29886 25452
rect 30098 25440 30104 25452
rect 30156 25440 30162 25492
rect 30653 25483 30711 25489
rect 30653 25449 30665 25483
rect 30699 25449 30711 25483
rect 31021 25483 31079 25489
rect 31021 25480 31033 25483
rect 30653 25443 30711 25449
rect 30944 25452 31033 25480
rect 23584 25384 23888 25412
rect 24762 25372 24768 25424
rect 24820 25412 24826 25424
rect 24820 25384 26188 25412
rect 24820 25372 24826 25384
rect 5626 25304 5632 25356
rect 5684 25304 5690 25356
rect 12986 25304 12992 25356
rect 13044 25344 13050 25356
rect 17310 25344 17316 25356
rect 13044 25316 17316 25344
rect 13044 25304 13050 25316
rect 17310 25304 17316 25316
rect 17368 25304 17374 25356
rect 19337 25347 19395 25353
rect 19337 25344 19349 25347
rect 17420 25316 19349 25344
rect 5445 25279 5503 25285
rect 5445 25245 5457 25279
rect 5491 25245 5503 25279
rect 5445 25239 5503 25245
rect 5460 25140 5488 25239
rect 10226 25236 10232 25288
rect 10284 25276 10290 25288
rect 10410 25276 10416 25288
rect 10284 25248 10416 25276
rect 10284 25236 10290 25248
rect 10410 25236 10416 25248
rect 10468 25236 10474 25288
rect 10502 25236 10508 25288
rect 10560 25276 10566 25288
rect 10597 25279 10655 25285
rect 10597 25276 10609 25279
rect 10560 25248 10609 25276
rect 10560 25236 10566 25248
rect 10597 25245 10609 25248
rect 10643 25245 10655 25279
rect 17420 25276 17448 25316
rect 19337 25313 19349 25316
rect 19383 25313 19395 25347
rect 19337 25307 19395 25313
rect 19426 25304 19432 25356
rect 19484 25344 19490 25356
rect 19794 25344 19800 25356
rect 19484 25316 19800 25344
rect 19484 25304 19490 25316
rect 19794 25304 19800 25316
rect 19852 25304 19858 25356
rect 20346 25304 20352 25356
rect 20404 25344 20410 25356
rect 20441 25347 20499 25353
rect 20441 25344 20453 25347
rect 20404 25316 20453 25344
rect 20404 25304 20410 25316
rect 20441 25313 20453 25316
rect 20487 25313 20499 25347
rect 21082 25344 21088 25356
rect 20441 25307 20499 25313
rect 20916 25316 21088 25344
rect 10597 25239 10655 25245
rect 14292 25248 17448 25276
rect 5721 25211 5779 25217
rect 5721 25177 5733 25211
rect 5767 25208 5779 25211
rect 10318 25208 10324 25220
rect 5767 25180 10324 25208
rect 5767 25177 5779 25180
rect 5721 25171 5779 25177
rect 10318 25168 10324 25180
rect 10376 25168 10382 25220
rect 14292 25152 14320 25248
rect 17678 25236 17684 25288
rect 17736 25276 17742 25288
rect 17736 25248 19472 25276
rect 17736 25236 17742 25248
rect 16114 25168 16120 25220
rect 16172 25168 16178 25220
rect 16298 25168 16304 25220
rect 16356 25168 16362 25220
rect 19245 25211 19303 25217
rect 19245 25208 19257 25211
rect 16408 25180 19257 25208
rect 5902 25140 5908 25152
rect 5460 25112 5908 25140
rect 5902 25100 5908 25112
rect 5960 25100 5966 25152
rect 9214 25100 9220 25152
rect 9272 25140 9278 25152
rect 10042 25140 10048 25152
rect 9272 25112 10048 25140
rect 9272 25100 9278 25112
rect 10042 25100 10048 25112
rect 10100 25100 10106 25152
rect 11606 25100 11612 25152
rect 11664 25140 11670 25152
rect 14274 25140 14280 25152
rect 11664 25112 14280 25140
rect 11664 25100 11670 25112
rect 14274 25100 14280 25112
rect 14332 25100 14338 25152
rect 15654 25100 15660 25152
rect 15712 25140 15718 25152
rect 16408 25140 16436 25180
rect 19245 25177 19257 25180
rect 19291 25177 19303 25211
rect 19444 25208 19472 25248
rect 19518 25236 19524 25288
rect 19576 25236 19582 25288
rect 20625 25279 20683 25285
rect 20625 25245 20637 25279
rect 20671 25276 20683 25279
rect 20916 25276 20944 25316
rect 21082 25304 21088 25316
rect 21140 25344 21146 25356
rect 21450 25344 21456 25356
rect 21140 25316 21456 25344
rect 21140 25304 21146 25316
rect 21450 25304 21456 25316
rect 21508 25304 21514 25356
rect 23382 25304 23388 25356
rect 23440 25304 23446 25356
rect 25133 25347 25191 25353
rect 25133 25344 25145 25347
rect 23492 25316 25145 25344
rect 23492 25276 23520 25316
rect 25133 25313 25145 25316
rect 25179 25313 25191 25347
rect 25133 25307 25191 25313
rect 20671 25248 20944 25276
rect 22066 25248 23520 25276
rect 20671 25245 20683 25248
rect 20625 25239 20683 25245
rect 20349 25211 20407 25217
rect 19444 25180 20300 25208
rect 19245 25171 19303 25177
rect 15712 25112 16436 25140
rect 15712 25100 15718 25112
rect 16482 25100 16488 25152
rect 16540 25100 16546 25152
rect 19260 25140 19288 25171
rect 19610 25140 19616 25152
rect 19260 25112 19616 25140
rect 19610 25100 19616 25112
rect 19668 25100 19674 25152
rect 20272 25140 20300 25180
rect 20349 25177 20361 25211
rect 20395 25208 20407 25211
rect 20530 25208 20536 25220
rect 20395 25180 20536 25208
rect 20395 25177 20407 25180
rect 20349 25171 20407 25177
rect 20530 25168 20536 25180
rect 20588 25208 20594 25220
rect 22066 25208 22094 25248
rect 23566 25236 23572 25288
rect 23624 25236 23630 25288
rect 24946 25236 24952 25288
rect 25004 25236 25010 25288
rect 25314 25236 25320 25288
rect 25372 25236 25378 25288
rect 25774 25236 25780 25288
rect 25832 25276 25838 25288
rect 26053 25279 26111 25285
rect 26053 25276 26065 25279
rect 25832 25248 26065 25276
rect 25832 25236 25838 25248
rect 26053 25245 26065 25248
rect 26099 25245 26111 25279
rect 26160 25276 26188 25384
rect 28626 25372 28632 25424
rect 28684 25372 28690 25424
rect 29914 25372 29920 25424
rect 29972 25412 29978 25424
rect 30668 25412 30696 25443
rect 29972 25384 30696 25412
rect 29972 25372 29978 25384
rect 30116 25356 30144 25384
rect 26237 25347 26295 25353
rect 26237 25313 26249 25347
rect 26283 25344 26295 25347
rect 26510 25344 26516 25356
rect 26283 25316 26516 25344
rect 26283 25313 26295 25316
rect 26237 25307 26295 25313
rect 26510 25304 26516 25316
rect 26568 25344 26574 25356
rect 26568 25316 30052 25344
rect 26568 25304 26574 25316
rect 28261 25279 28319 25285
rect 28261 25276 28273 25279
rect 26160 25248 28273 25276
rect 26053 25239 26111 25245
rect 28261 25245 28273 25248
rect 28307 25245 28319 25279
rect 28261 25239 28319 25245
rect 29546 25236 29552 25288
rect 29604 25236 29610 25288
rect 29730 25236 29736 25288
rect 29788 25236 29794 25288
rect 29825 25279 29883 25285
rect 29825 25245 29837 25279
rect 29871 25245 29883 25279
rect 30024 25276 30052 25316
rect 30098 25304 30104 25356
rect 30156 25304 30162 25356
rect 30282 25304 30288 25356
rect 30340 25344 30346 25356
rect 30745 25347 30803 25353
rect 30745 25344 30757 25347
rect 30340 25316 30757 25344
rect 30340 25304 30346 25316
rect 30745 25313 30757 25316
rect 30791 25313 30803 25347
rect 30944 25344 30972 25452
rect 31021 25449 31033 25452
rect 31067 25449 31079 25483
rect 31021 25443 31079 25449
rect 31110 25440 31116 25492
rect 31168 25480 31174 25492
rect 31573 25483 31631 25489
rect 31573 25480 31585 25483
rect 31168 25452 31585 25480
rect 31168 25440 31174 25452
rect 31573 25449 31585 25452
rect 31619 25449 31631 25483
rect 31573 25443 31631 25449
rect 32030 25440 32036 25492
rect 32088 25440 32094 25492
rect 33410 25440 33416 25492
rect 33468 25480 33474 25492
rect 33686 25480 33692 25492
rect 33468 25452 33692 25480
rect 33468 25440 33474 25452
rect 33686 25440 33692 25452
rect 33744 25440 33750 25492
rect 34146 25440 34152 25492
rect 34204 25480 34210 25492
rect 34793 25483 34851 25489
rect 34793 25480 34805 25483
rect 34204 25452 34805 25480
rect 34204 25440 34210 25452
rect 34793 25449 34805 25452
rect 34839 25449 34851 25483
rect 34793 25443 34851 25449
rect 35158 25440 35164 25492
rect 35216 25440 35222 25492
rect 36446 25440 36452 25492
rect 36504 25480 36510 25492
rect 36541 25483 36599 25489
rect 36541 25480 36553 25483
rect 36504 25452 36553 25480
rect 36504 25440 36510 25452
rect 36541 25449 36553 25452
rect 36587 25449 36599 25483
rect 36541 25443 36599 25449
rect 36909 25483 36967 25489
rect 36909 25449 36921 25483
rect 36955 25480 36967 25483
rect 37550 25480 37556 25492
rect 36955 25452 37556 25480
rect 36955 25449 36967 25452
rect 36909 25443 36967 25449
rect 37550 25440 37556 25452
rect 37608 25440 37614 25492
rect 40405 25483 40463 25489
rect 40405 25449 40417 25483
rect 40451 25480 40463 25483
rect 40586 25480 40592 25492
rect 40451 25452 40592 25480
rect 40451 25449 40463 25452
rect 40405 25443 40463 25449
rect 40586 25440 40592 25452
rect 40644 25440 40650 25492
rect 31386 25372 31392 25424
rect 31444 25412 31450 25424
rect 32861 25415 32919 25421
rect 32861 25412 32873 25415
rect 31444 25384 32873 25412
rect 31444 25372 31450 25384
rect 32861 25381 32873 25384
rect 32907 25381 32919 25415
rect 37734 25412 37740 25424
rect 32861 25375 32919 25381
rect 34164 25384 37740 25412
rect 30944 25316 31432 25344
rect 30745 25307 30803 25313
rect 30653 25279 30711 25285
rect 30653 25276 30665 25279
rect 30024 25248 30665 25276
rect 29825 25239 29883 25245
rect 30653 25245 30665 25248
rect 30699 25276 30711 25279
rect 30926 25276 30932 25288
rect 30699 25248 30932 25276
rect 30699 25245 30711 25248
rect 30653 25239 30711 25245
rect 20588 25180 22094 25208
rect 20588 25168 20594 25180
rect 22278 25168 22284 25220
rect 22336 25208 22342 25220
rect 23293 25211 23351 25217
rect 23293 25208 23305 25211
rect 22336 25180 23305 25208
rect 22336 25168 22342 25180
rect 23293 25177 23305 25180
rect 23339 25208 23351 25211
rect 24964 25208 24992 25236
rect 23339 25180 24992 25208
rect 25041 25211 25099 25217
rect 23339 25177 23351 25180
rect 23293 25171 23351 25177
rect 25041 25177 25053 25211
rect 25087 25208 25099 25211
rect 25869 25211 25927 25217
rect 25087 25180 25360 25208
rect 25087 25177 25099 25180
rect 25041 25171 25099 25177
rect 25332 25152 25360 25180
rect 25869 25177 25881 25211
rect 25915 25208 25927 25211
rect 26142 25208 26148 25220
rect 25915 25180 26148 25208
rect 25915 25177 25927 25180
rect 25869 25171 25927 25177
rect 26142 25168 26148 25180
rect 26200 25168 26206 25220
rect 28442 25168 28448 25220
rect 28500 25168 28506 25220
rect 28902 25168 28908 25220
rect 28960 25168 28966 25220
rect 29086 25168 29092 25220
rect 29144 25168 29150 25220
rect 29840 25208 29868 25239
rect 30926 25236 30932 25248
rect 30984 25236 30990 25288
rect 31404 25220 31432 25316
rect 31754 25304 31760 25356
rect 31812 25304 31818 25356
rect 32876 25344 32904 25375
rect 33686 25344 33692 25356
rect 32876 25316 33692 25344
rect 33686 25304 33692 25316
rect 33744 25304 33750 25356
rect 31478 25236 31484 25288
rect 31536 25276 31542 25288
rect 31849 25279 31907 25285
rect 31536 25248 31754 25276
rect 31536 25236 31542 25248
rect 29840 25180 30144 25208
rect 23198 25140 23204 25152
rect 20272 25112 23204 25140
rect 23198 25100 23204 25112
rect 23256 25100 23262 25152
rect 24949 25143 25007 25149
rect 24949 25109 24961 25143
rect 24995 25140 25007 25143
rect 25222 25140 25228 25152
rect 24995 25112 25228 25140
rect 24995 25109 25007 25112
rect 24949 25103 25007 25109
rect 25222 25100 25228 25112
rect 25280 25100 25286 25152
rect 25314 25100 25320 25152
rect 25372 25100 25378 25152
rect 25406 25100 25412 25152
rect 25464 25140 25470 25152
rect 26050 25140 26056 25152
rect 25464 25112 26056 25140
rect 25464 25100 25470 25112
rect 26050 25100 26056 25112
rect 26108 25100 26114 25152
rect 26234 25100 26240 25152
rect 26292 25140 26298 25152
rect 26970 25140 26976 25152
rect 26292 25112 26976 25140
rect 26292 25100 26298 25112
rect 26970 25100 26976 25112
rect 27028 25140 27034 25152
rect 27430 25140 27436 25152
rect 27028 25112 27436 25140
rect 27028 25100 27034 25112
rect 27430 25100 27436 25112
rect 27488 25100 27494 25152
rect 27522 25100 27528 25152
rect 27580 25140 27586 25152
rect 29840 25140 29868 25180
rect 27580 25112 29868 25140
rect 27580 25100 27586 25112
rect 30006 25100 30012 25152
rect 30064 25100 30070 25152
rect 30116 25140 30144 25180
rect 31386 25168 31392 25220
rect 31444 25208 31450 25220
rect 31573 25211 31631 25217
rect 31573 25208 31585 25211
rect 31444 25180 31585 25208
rect 31444 25168 31450 25180
rect 31573 25177 31585 25180
rect 31619 25177 31631 25211
rect 31726 25208 31754 25248
rect 31849 25245 31861 25279
rect 31895 25276 31907 25279
rect 32214 25276 32220 25288
rect 31895 25248 32220 25276
rect 31895 25245 31907 25248
rect 31849 25239 31907 25245
rect 32214 25236 32220 25248
rect 32272 25236 32278 25288
rect 32766 25208 32772 25220
rect 31726 25180 32772 25208
rect 31573 25171 31631 25177
rect 32766 25168 32772 25180
rect 32824 25168 32830 25220
rect 34164 25217 34192 25384
rect 37734 25372 37740 25384
rect 37792 25372 37798 25424
rect 40678 25372 40684 25424
rect 40736 25372 40742 25424
rect 34514 25304 34520 25356
rect 34572 25344 34578 25356
rect 34572 25316 36492 25344
rect 34572 25304 34578 25316
rect 34793 25279 34851 25285
rect 34793 25245 34805 25279
rect 34839 25276 34851 25279
rect 34882 25276 34888 25288
rect 34839 25248 34888 25276
rect 34839 25245 34851 25248
rect 34793 25239 34851 25245
rect 34882 25236 34888 25248
rect 34940 25236 34946 25288
rect 34977 25279 35035 25285
rect 34977 25245 34989 25279
rect 35023 25276 35035 25279
rect 36170 25276 36176 25288
rect 35023 25248 36176 25276
rect 35023 25245 35035 25248
rect 34977 25239 35035 25245
rect 36170 25236 36176 25248
rect 36228 25236 36234 25288
rect 36464 25285 36492 25316
rect 36906 25304 36912 25356
rect 36964 25344 36970 25356
rect 40773 25347 40831 25353
rect 40773 25344 40785 25347
rect 36964 25316 40785 25344
rect 36964 25304 36970 25316
rect 40773 25313 40785 25316
rect 40819 25313 40831 25347
rect 40773 25307 40831 25313
rect 40862 25304 40868 25356
rect 40920 25304 40926 25356
rect 43714 25304 43720 25356
rect 43772 25304 43778 25356
rect 36449 25279 36507 25285
rect 36449 25245 36461 25279
rect 36495 25245 36507 25279
rect 36449 25239 36507 25245
rect 36630 25236 36636 25288
rect 36688 25236 36694 25288
rect 36725 25279 36783 25285
rect 36725 25245 36737 25279
rect 36771 25276 36783 25279
rect 36771 25248 36860 25276
rect 36771 25245 36783 25248
rect 36725 25239 36783 25245
rect 34149 25211 34207 25217
rect 34149 25177 34161 25211
rect 34195 25177 34207 25211
rect 34149 25171 34207 25177
rect 34054 25140 34060 25152
rect 30116 25112 34060 25140
rect 34054 25100 34060 25112
rect 34112 25140 34118 25152
rect 36832 25140 36860 25248
rect 39298 25236 39304 25288
rect 39356 25276 39362 25288
rect 39758 25276 39764 25288
rect 39356 25248 39764 25276
rect 39356 25236 39362 25248
rect 39758 25236 39764 25248
rect 39816 25276 39822 25288
rect 40589 25279 40647 25285
rect 40589 25276 40601 25279
rect 39816 25248 40601 25276
rect 39816 25236 39822 25248
rect 40589 25245 40601 25248
rect 40635 25245 40647 25279
rect 40589 25239 40647 25245
rect 41049 25279 41107 25285
rect 41049 25245 41061 25279
rect 41095 25276 41107 25279
rect 41506 25276 41512 25288
rect 41095 25248 41512 25276
rect 41095 25245 41107 25248
rect 41049 25239 41107 25245
rect 41506 25236 41512 25248
rect 41564 25236 41570 25288
rect 41601 25279 41659 25285
rect 41601 25245 41613 25279
rect 41647 25276 41659 25279
rect 41690 25276 41696 25288
rect 41647 25248 41696 25276
rect 41647 25245 41659 25248
rect 41601 25239 41659 25245
rect 41690 25236 41696 25248
rect 41748 25236 41754 25288
rect 42794 25276 42800 25288
rect 41800 25248 42800 25276
rect 34112 25112 36860 25140
rect 34112 25100 34118 25112
rect 40862 25100 40868 25152
rect 40920 25140 40926 25152
rect 41800 25140 41828 25248
rect 42794 25236 42800 25248
rect 42852 25276 42858 25288
rect 43993 25279 44051 25285
rect 43993 25276 44005 25279
rect 42852 25248 44005 25276
rect 42852 25236 42858 25248
rect 43993 25245 44005 25248
rect 44039 25245 44051 25279
rect 43993 25239 44051 25245
rect 44266 25236 44272 25288
rect 44324 25236 44330 25288
rect 41868 25211 41926 25217
rect 41868 25177 41880 25211
rect 41914 25208 41926 25211
rect 43162 25208 43168 25220
rect 41914 25180 43168 25208
rect 41914 25177 41926 25180
rect 41868 25171 41926 25177
rect 43162 25168 43168 25180
rect 43220 25168 43226 25220
rect 43806 25168 43812 25220
rect 43864 25168 43870 25220
rect 40920 25112 41828 25140
rect 40920 25100 40926 25112
rect 42978 25100 42984 25152
rect 43036 25100 43042 25152
rect 43070 25100 43076 25152
rect 43128 25100 43134 25152
rect 44450 25100 44456 25152
rect 44508 25100 44514 25152
rect 1104 25050 44896 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 44896 25050
rect 1104 24976 44896 24998
rect 5626 24896 5632 24948
rect 5684 24936 5690 24948
rect 5813 24939 5871 24945
rect 5813 24936 5825 24939
rect 5684 24908 5825 24936
rect 5684 24896 5690 24908
rect 5813 24905 5825 24908
rect 5859 24936 5871 24939
rect 5859 24908 13584 24936
rect 5859 24905 5871 24908
rect 5813 24899 5871 24905
rect 13556 24868 13584 24908
rect 13630 24896 13636 24948
rect 13688 24936 13694 24948
rect 15654 24936 15660 24948
rect 13688 24908 15660 24936
rect 13688 24896 13694 24908
rect 15654 24896 15660 24908
rect 15712 24896 15718 24948
rect 16482 24896 16488 24948
rect 16540 24936 16546 24948
rect 16540 24908 19932 24936
rect 16540 24896 16546 24908
rect 19334 24868 19340 24880
rect 11808 24840 12020 24868
rect 13556 24840 19340 24868
rect 5994 24760 6000 24812
rect 6052 24760 6058 24812
rect 6178 24760 6184 24812
rect 6236 24760 6242 24812
rect 6822 24760 6828 24812
rect 6880 24800 6886 24812
rect 8389 24803 8447 24809
rect 8389 24800 8401 24803
rect 6880 24772 8401 24800
rect 6880 24760 6886 24772
rect 8389 24769 8401 24772
rect 8435 24800 8447 24803
rect 10042 24800 10048 24812
rect 8435 24772 10048 24800
rect 8435 24769 8447 24772
rect 8389 24763 8447 24769
rect 10042 24760 10048 24772
rect 10100 24760 10106 24812
rect 10321 24803 10379 24809
rect 10321 24769 10333 24803
rect 10367 24800 10379 24803
rect 11808 24800 11836 24840
rect 10367 24772 11836 24800
rect 11885 24803 11943 24809
rect 10367 24769 10379 24772
rect 10321 24763 10379 24769
rect 11885 24769 11897 24803
rect 11931 24769 11943 24803
rect 11992 24800 12020 24840
rect 19334 24828 19340 24840
rect 19392 24828 19398 24880
rect 19904 24868 19932 24908
rect 20530 24896 20536 24948
rect 20588 24936 20594 24948
rect 20625 24939 20683 24945
rect 20625 24936 20637 24939
rect 20588 24908 20637 24936
rect 20588 24896 20594 24908
rect 20625 24905 20637 24908
rect 20671 24905 20683 24939
rect 20625 24899 20683 24905
rect 23017 24939 23075 24945
rect 23017 24905 23029 24939
rect 23063 24936 23075 24939
rect 24394 24936 24400 24948
rect 23063 24908 24400 24936
rect 23063 24905 23075 24908
rect 23017 24899 23075 24905
rect 24394 24896 24400 24908
rect 24452 24896 24458 24948
rect 24854 24896 24860 24948
rect 24912 24936 24918 24948
rect 26510 24936 26516 24948
rect 24912 24908 26516 24936
rect 24912 24896 24918 24908
rect 26510 24896 26516 24908
rect 26568 24896 26574 24948
rect 29454 24896 29460 24948
rect 29512 24936 29518 24948
rect 30098 24936 30104 24948
rect 29512 24908 30104 24936
rect 29512 24896 29518 24908
rect 30098 24896 30104 24908
rect 30156 24896 30162 24948
rect 31754 24896 31760 24948
rect 31812 24936 31818 24948
rect 32125 24939 32183 24945
rect 32125 24936 32137 24939
rect 31812 24908 32137 24936
rect 31812 24896 31818 24908
rect 32125 24905 32137 24908
rect 32171 24905 32183 24939
rect 32125 24899 32183 24905
rect 32306 24896 32312 24948
rect 32364 24936 32370 24948
rect 32766 24936 32772 24948
rect 32364 24908 32772 24936
rect 32364 24896 32370 24908
rect 32766 24896 32772 24908
rect 32824 24896 32830 24948
rect 34146 24936 34152 24948
rect 33152 24908 34152 24936
rect 24762 24868 24768 24880
rect 19444 24840 19840 24868
rect 19904 24840 24768 24868
rect 12161 24803 12219 24809
rect 11992 24772 12112 24800
rect 11885 24763 11943 24769
rect 8018 24692 8024 24744
rect 8076 24732 8082 24744
rect 8536 24735 8594 24741
rect 8536 24732 8548 24735
rect 8076 24704 8548 24732
rect 8076 24692 8082 24704
rect 8536 24701 8548 24704
rect 8582 24701 8594 24735
rect 8536 24695 8594 24701
rect 8754 24692 8760 24744
rect 8812 24692 8818 24744
rect 10134 24692 10140 24744
rect 10192 24692 10198 24744
rect 11606 24692 11612 24744
rect 11664 24732 11670 24744
rect 11900 24732 11928 24763
rect 11664 24704 11928 24732
rect 11664 24692 11670 24704
rect 11974 24692 11980 24744
rect 12032 24692 12038 24744
rect 12084 24732 12112 24772
rect 12161 24769 12173 24803
rect 12207 24800 12219 24803
rect 13630 24800 13636 24812
rect 12207 24772 13636 24800
rect 12207 24769 12219 24772
rect 12161 24763 12219 24769
rect 13630 24760 13636 24772
rect 13688 24760 13694 24812
rect 13814 24760 13820 24812
rect 13872 24800 13878 24812
rect 14001 24803 14059 24809
rect 14001 24800 14013 24803
rect 13872 24772 14013 24800
rect 13872 24760 13878 24772
rect 14001 24769 14013 24772
rect 14047 24769 14059 24803
rect 14001 24763 14059 24769
rect 14185 24803 14243 24809
rect 14185 24769 14197 24803
rect 14231 24800 14243 24803
rect 14366 24800 14372 24812
rect 14231 24772 14372 24800
rect 14231 24769 14243 24772
rect 14185 24763 14243 24769
rect 14366 24760 14372 24772
rect 14424 24760 14430 24812
rect 15930 24760 15936 24812
rect 15988 24800 15994 24812
rect 16390 24800 16396 24812
rect 15988 24772 16396 24800
rect 15988 24760 15994 24772
rect 16390 24760 16396 24772
rect 16448 24760 16454 24812
rect 17218 24760 17224 24812
rect 17276 24800 17282 24812
rect 17313 24803 17371 24809
rect 17313 24800 17325 24803
rect 17276 24772 17325 24800
rect 17276 24760 17282 24772
rect 17313 24769 17325 24772
rect 17359 24769 17371 24803
rect 17313 24763 17371 24769
rect 17586 24760 17592 24812
rect 17644 24760 17650 24812
rect 17678 24760 17684 24812
rect 17736 24800 17742 24812
rect 17865 24803 17923 24809
rect 17865 24800 17877 24803
rect 17736 24772 17877 24800
rect 17736 24760 17742 24772
rect 17865 24769 17877 24772
rect 17911 24800 17923 24803
rect 18230 24800 18236 24812
rect 17911 24772 18236 24800
rect 17911 24769 17923 24772
rect 17865 24763 17923 24769
rect 18230 24760 18236 24772
rect 18288 24760 18294 24812
rect 18506 24760 18512 24812
rect 18564 24800 18570 24812
rect 19444 24800 19472 24840
rect 18564 24772 19472 24800
rect 18564 24760 18570 24772
rect 19610 24760 19616 24812
rect 19668 24760 19674 24812
rect 19702 24760 19708 24812
rect 19760 24760 19766 24812
rect 19812 24800 19840 24840
rect 24762 24828 24768 24840
rect 24820 24828 24826 24880
rect 26326 24868 26332 24880
rect 25884 24840 26332 24868
rect 20162 24800 20168 24812
rect 19812 24772 20168 24800
rect 20162 24760 20168 24772
rect 20220 24800 20226 24812
rect 20257 24803 20315 24809
rect 20257 24800 20269 24803
rect 20220 24772 20269 24800
rect 20220 24760 20226 24772
rect 20257 24769 20269 24772
rect 20303 24769 20315 24803
rect 20257 24763 20315 24769
rect 20441 24803 20499 24809
rect 20441 24769 20453 24803
rect 20487 24769 20499 24803
rect 20441 24763 20499 24769
rect 16574 24732 16580 24744
rect 12084 24704 16580 24732
rect 16574 24692 16580 24704
rect 16632 24692 16638 24744
rect 16758 24692 16764 24744
rect 16816 24732 16822 24744
rect 17405 24735 17463 24741
rect 17405 24732 17417 24735
rect 16816 24704 17417 24732
rect 16816 24692 16822 24704
rect 17405 24701 17417 24704
rect 17451 24701 17463 24735
rect 17405 24695 17463 24701
rect 17512 24704 17908 24732
rect 10505 24667 10563 24673
rect 10505 24633 10517 24667
rect 10551 24664 10563 24667
rect 13354 24664 13360 24676
rect 10551 24636 13360 24664
rect 10551 24633 10563 24636
rect 10505 24627 10563 24633
rect 13354 24624 13360 24636
rect 13412 24624 13418 24676
rect 13906 24624 13912 24676
rect 13964 24664 13970 24676
rect 17512 24664 17540 24704
rect 13964 24636 17540 24664
rect 13964 24624 13970 24636
rect 17770 24624 17776 24676
rect 17828 24624 17834 24676
rect 17880 24664 17908 24704
rect 17954 24692 17960 24744
rect 18012 24732 18018 24744
rect 18598 24732 18604 24744
rect 18012 24704 18604 24732
rect 18012 24692 18018 24704
rect 18598 24692 18604 24704
rect 18656 24692 18662 24744
rect 20456 24732 20484 24763
rect 20622 24760 20628 24812
rect 20680 24800 20686 24812
rect 20717 24803 20775 24809
rect 20717 24800 20729 24803
rect 20680 24772 20729 24800
rect 20680 24760 20686 24772
rect 20717 24769 20729 24772
rect 20763 24769 20775 24803
rect 20717 24763 20775 24769
rect 20901 24803 20959 24809
rect 20901 24769 20913 24803
rect 20947 24769 20959 24803
rect 20901 24763 20959 24769
rect 19904 24704 20484 24732
rect 20916 24732 20944 24763
rect 22554 24760 22560 24812
rect 22612 24760 22618 24812
rect 22833 24803 22891 24809
rect 22833 24769 22845 24803
rect 22879 24800 22891 24803
rect 22922 24800 22928 24812
rect 22879 24772 22928 24800
rect 22879 24769 22891 24772
rect 22833 24763 22891 24769
rect 22922 24760 22928 24772
rect 22980 24800 22986 24812
rect 25884 24800 25912 24840
rect 26326 24828 26332 24840
rect 26384 24868 26390 24880
rect 27798 24868 27804 24880
rect 26384 24840 27804 24868
rect 26384 24828 26390 24840
rect 27798 24828 27804 24840
rect 27856 24828 27862 24880
rect 28442 24828 28448 24880
rect 28500 24868 28506 24880
rect 28500 24840 32536 24868
rect 28500 24828 28506 24840
rect 32508 24812 32536 24840
rect 26421 24803 26479 24809
rect 26421 24800 26433 24803
rect 22980 24772 25912 24800
rect 25976 24772 26433 24800
rect 22980 24760 22986 24772
rect 21266 24732 21272 24744
rect 20916 24704 21272 24732
rect 17880 24636 18000 24664
rect 8294 24556 8300 24608
rect 8352 24596 8358 24608
rect 8662 24596 8668 24608
rect 8352 24568 8668 24596
rect 8352 24556 8358 24568
rect 8662 24556 8668 24568
rect 8720 24556 8726 24608
rect 9033 24599 9091 24605
rect 9033 24565 9045 24599
rect 9079 24596 9091 24599
rect 9582 24596 9588 24608
rect 9079 24568 9588 24596
rect 9079 24565 9091 24568
rect 9033 24559 9091 24565
rect 9582 24556 9588 24568
rect 9640 24556 9646 24608
rect 9674 24556 9680 24608
rect 9732 24596 9738 24608
rect 9950 24596 9956 24608
rect 9732 24568 9956 24596
rect 9732 24556 9738 24568
rect 9950 24556 9956 24568
rect 10008 24596 10014 24608
rect 10045 24599 10103 24605
rect 10045 24596 10057 24599
rect 10008 24568 10057 24596
rect 10008 24556 10014 24568
rect 10045 24565 10057 24568
rect 10091 24565 10103 24599
rect 10045 24559 10103 24565
rect 10318 24556 10324 24608
rect 10376 24596 10382 24608
rect 11701 24599 11759 24605
rect 11701 24596 11713 24599
rect 10376 24568 11713 24596
rect 10376 24556 10382 24568
rect 11701 24565 11713 24568
rect 11747 24565 11759 24599
rect 11701 24559 11759 24565
rect 11790 24556 11796 24608
rect 11848 24596 11854 24608
rect 11885 24599 11943 24605
rect 11885 24596 11897 24599
rect 11848 24568 11897 24596
rect 11848 24556 11854 24568
rect 11885 24565 11897 24568
rect 11931 24565 11943 24599
rect 11885 24559 11943 24565
rect 14366 24556 14372 24608
rect 14424 24556 14430 24608
rect 16482 24556 16488 24608
rect 16540 24596 16546 24608
rect 17313 24599 17371 24605
rect 17313 24596 17325 24599
rect 16540 24568 17325 24596
rect 16540 24556 16546 24568
rect 17313 24565 17325 24568
rect 17359 24565 17371 24599
rect 17313 24559 17371 24565
rect 17862 24556 17868 24608
rect 17920 24556 17926 24608
rect 17972 24596 18000 24636
rect 18230 24624 18236 24676
rect 18288 24624 18294 24676
rect 18690 24624 18696 24676
rect 18748 24664 18754 24676
rect 19904 24664 19932 24704
rect 21266 24692 21272 24704
rect 21324 24732 21330 24744
rect 22741 24735 22799 24741
rect 22741 24732 22753 24735
rect 21324 24704 22753 24732
rect 21324 24692 21330 24704
rect 22741 24701 22753 24704
rect 22787 24732 22799 24735
rect 25774 24732 25780 24744
rect 22787 24704 25780 24732
rect 22787 24701 22799 24704
rect 22741 24695 22799 24701
rect 25774 24692 25780 24704
rect 25832 24692 25838 24744
rect 18748 24636 19932 24664
rect 19981 24667 20039 24673
rect 18748 24624 18754 24636
rect 19981 24633 19993 24667
rect 20027 24664 20039 24667
rect 25976 24664 26004 24772
rect 26421 24769 26433 24772
rect 26467 24800 26479 24803
rect 31110 24800 31116 24812
rect 26467 24772 31116 24800
rect 26467 24769 26479 24772
rect 26421 24763 26479 24769
rect 31110 24760 31116 24772
rect 31168 24760 31174 24812
rect 31662 24760 31668 24812
rect 31720 24800 31726 24812
rect 32309 24803 32367 24809
rect 32309 24800 32321 24803
rect 31720 24772 32321 24800
rect 31720 24760 31726 24772
rect 32309 24769 32321 24772
rect 32355 24769 32367 24803
rect 32309 24763 32367 24769
rect 32490 24760 32496 24812
rect 32548 24760 32554 24812
rect 32758 24803 32816 24809
rect 32758 24800 32770 24803
rect 32600 24772 32770 24800
rect 26326 24692 26332 24744
rect 26384 24692 26390 24744
rect 26786 24692 26792 24744
rect 26844 24732 26850 24744
rect 31938 24732 31944 24744
rect 26844 24704 31944 24732
rect 26844 24692 26850 24704
rect 31938 24692 31944 24704
rect 31996 24692 32002 24744
rect 20027 24636 26004 24664
rect 20027 24633 20039 24636
rect 19981 24627 20039 24633
rect 26050 24624 26056 24676
rect 26108 24624 26114 24676
rect 26804 24664 26832 24692
rect 26160 24636 26832 24664
rect 19702 24596 19708 24608
rect 17972 24568 19708 24596
rect 19702 24556 19708 24568
rect 19760 24556 19766 24608
rect 19797 24599 19855 24605
rect 19797 24565 19809 24599
rect 19843 24596 19855 24599
rect 20162 24596 20168 24608
rect 19843 24568 20168 24596
rect 19843 24565 19855 24568
rect 19797 24559 19855 24565
rect 20162 24556 20168 24568
rect 20220 24556 20226 24608
rect 21085 24599 21143 24605
rect 21085 24565 21097 24599
rect 21131 24596 21143 24599
rect 21174 24596 21180 24608
rect 21131 24568 21180 24596
rect 21131 24565 21143 24568
rect 21085 24559 21143 24565
rect 21174 24556 21180 24568
rect 21232 24556 21238 24608
rect 22738 24556 22744 24608
rect 22796 24556 22802 24608
rect 22830 24556 22836 24608
rect 22888 24596 22894 24608
rect 26160 24596 26188 24636
rect 26970 24624 26976 24676
rect 27028 24664 27034 24676
rect 27154 24664 27160 24676
rect 27028 24636 27160 24664
rect 27028 24624 27034 24636
rect 27154 24624 27160 24636
rect 27212 24624 27218 24676
rect 27890 24624 27896 24676
rect 27948 24664 27954 24676
rect 30742 24664 30748 24676
rect 27948 24636 30748 24664
rect 27948 24624 27954 24636
rect 30742 24624 30748 24636
rect 30800 24664 30806 24676
rect 31018 24664 31024 24676
rect 30800 24636 31024 24664
rect 30800 24624 30806 24636
rect 31018 24624 31024 24636
rect 31076 24624 31082 24676
rect 32306 24664 32312 24676
rect 31956 24636 32312 24664
rect 22888 24568 26188 24596
rect 26421 24599 26479 24605
rect 22888 24556 22894 24568
rect 26421 24565 26433 24599
rect 26467 24596 26479 24599
rect 26510 24596 26516 24608
rect 26467 24568 26516 24596
rect 26467 24565 26479 24568
rect 26421 24559 26479 24565
rect 26510 24556 26516 24568
rect 26568 24596 26574 24608
rect 27246 24596 27252 24608
rect 26568 24568 27252 24596
rect 26568 24556 26574 24568
rect 27246 24556 27252 24568
rect 27304 24556 27310 24608
rect 28258 24556 28264 24608
rect 28316 24596 28322 24608
rect 31956 24596 31984 24636
rect 32306 24624 32312 24636
rect 32364 24624 32370 24676
rect 28316 24568 31984 24596
rect 28316 24556 28322 24568
rect 32030 24556 32036 24608
rect 32088 24596 32094 24608
rect 32600 24596 32628 24772
rect 32758 24769 32770 24772
rect 32804 24800 32816 24803
rect 32950 24800 32956 24812
rect 32804 24772 32956 24800
rect 32804 24769 32816 24772
rect 32758 24763 32816 24769
rect 32950 24760 32956 24772
rect 33008 24760 33014 24812
rect 33045 24803 33103 24809
rect 33045 24769 33057 24803
rect 33091 24800 33103 24803
rect 33152 24800 33180 24908
rect 34146 24896 34152 24908
rect 34204 24896 34210 24948
rect 35158 24896 35164 24948
rect 35216 24936 35222 24948
rect 41966 24936 41972 24948
rect 35216 24908 41972 24936
rect 35216 24896 35222 24908
rect 41966 24896 41972 24908
rect 42024 24896 42030 24948
rect 43714 24896 43720 24948
rect 43772 24936 43778 24948
rect 43809 24939 43867 24945
rect 43809 24936 43821 24939
rect 43772 24908 43821 24936
rect 43772 24896 43778 24908
rect 43809 24905 43821 24908
rect 43855 24905 43867 24939
rect 43809 24899 43867 24905
rect 33594 24828 33600 24880
rect 33652 24868 33658 24880
rect 33870 24868 33876 24880
rect 33652 24840 33876 24868
rect 33652 24828 33658 24840
rect 33870 24828 33876 24840
rect 33928 24868 33934 24880
rect 35526 24868 35532 24880
rect 33928 24840 34468 24868
rect 33928 24828 33934 24840
rect 33091 24772 33180 24800
rect 33091 24769 33103 24772
rect 33045 24763 33103 24769
rect 33686 24760 33692 24812
rect 33744 24760 33750 24812
rect 34440 24800 34468 24840
rect 35360 24840 35532 24868
rect 35360 24800 35388 24840
rect 35526 24828 35532 24840
rect 35584 24828 35590 24880
rect 41432 24840 42104 24868
rect 34440 24772 35388 24800
rect 35434 24760 35440 24812
rect 35492 24800 35498 24812
rect 38565 24803 38623 24809
rect 38565 24800 38577 24803
rect 35492 24772 38577 24800
rect 35492 24760 35498 24772
rect 38565 24769 38577 24772
rect 38611 24769 38623 24803
rect 38565 24763 38623 24769
rect 38838 24760 38844 24812
rect 38896 24760 38902 24812
rect 32861 24735 32919 24741
rect 32861 24701 32873 24735
rect 32907 24701 32919 24735
rect 33704 24732 33732 24760
rect 35986 24732 35992 24744
rect 33704 24704 35992 24732
rect 32861 24695 32919 24701
rect 32766 24624 32772 24676
rect 32824 24664 32830 24676
rect 32876 24664 32904 24695
rect 35986 24692 35992 24704
rect 36044 24692 36050 24744
rect 38746 24692 38752 24744
rect 38804 24692 38810 24744
rect 41230 24692 41236 24744
rect 41288 24732 41294 24744
rect 41432 24732 41460 24840
rect 41598 24760 41604 24812
rect 41656 24800 41662 24812
rect 42076 24809 42104 24840
rect 41693 24803 41751 24809
rect 41693 24800 41705 24803
rect 41656 24772 41705 24800
rect 41656 24760 41662 24772
rect 41693 24769 41705 24772
rect 41739 24769 41751 24803
rect 41969 24803 42027 24809
rect 41969 24800 41981 24803
rect 41693 24763 41751 24769
rect 41791 24772 41981 24800
rect 41791 24732 41819 24772
rect 41969 24769 41981 24772
rect 42015 24769 42027 24803
rect 41969 24763 42027 24769
rect 42061 24803 42119 24809
rect 42061 24769 42073 24803
rect 42107 24769 42119 24803
rect 42061 24763 42119 24769
rect 42245 24803 42303 24809
rect 42245 24769 42257 24803
rect 42291 24800 42303 24803
rect 42685 24803 42743 24809
rect 42685 24800 42697 24803
rect 42291 24772 42697 24800
rect 42291 24769 42303 24772
rect 42245 24763 42303 24769
rect 42685 24769 42697 24772
rect 42731 24769 42743 24803
rect 42685 24763 42743 24769
rect 42978 24760 42984 24812
rect 43036 24800 43042 24812
rect 44269 24803 44327 24809
rect 44269 24800 44281 24803
rect 43036 24772 44281 24800
rect 43036 24760 43042 24772
rect 44269 24769 44281 24772
rect 44315 24769 44327 24803
rect 44269 24763 44327 24769
rect 41288 24704 41460 24732
rect 41708 24704 41819 24732
rect 41288 24692 41294 24704
rect 32824 24636 32904 24664
rect 32824 24624 32830 24636
rect 33318 24624 33324 24676
rect 33376 24664 33382 24676
rect 33686 24664 33692 24676
rect 33376 24636 33692 24664
rect 33376 24624 33382 24636
rect 33686 24624 33692 24636
rect 33744 24624 33750 24676
rect 36262 24624 36268 24676
rect 36320 24664 36326 24676
rect 36722 24664 36728 24676
rect 36320 24636 36728 24664
rect 36320 24624 36326 24636
rect 36722 24624 36728 24636
rect 36780 24624 36786 24676
rect 41598 24624 41604 24676
rect 41656 24664 41662 24676
rect 41708 24664 41736 24704
rect 41874 24692 41880 24744
rect 41932 24732 41938 24744
rect 42429 24735 42487 24741
rect 42429 24732 42441 24735
rect 41932 24704 42441 24732
rect 41932 24692 41938 24704
rect 42429 24701 42441 24704
rect 42475 24701 42487 24735
rect 42429 24695 42487 24701
rect 41656 24636 41736 24664
rect 41656 24624 41662 24636
rect 32088 24568 32628 24596
rect 32088 24556 32094 24568
rect 32950 24556 32956 24608
rect 33008 24556 33014 24608
rect 33229 24599 33287 24605
rect 33229 24565 33241 24599
rect 33275 24596 33287 24599
rect 33778 24596 33784 24608
rect 33275 24568 33784 24596
rect 33275 24565 33287 24568
rect 33229 24559 33287 24565
rect 33778 24556 33784 24568
rect 33836 24596 33842 24608
rect 35710 24596 35716 24608
rect 33836 24568 35716 24596
rect 33836 24556 33842 24568
rect 35710 24556 35716 24568
rect 35768 24556 35774 24608
rect 38286 24556 38292 24608
rect 38344 24596 38350 24608
rect 38657 24599 38715 24605
rect 38657 24596 38669 24599
rect 38344 24568 38669 24596
rect 38344 24556 38350 24568
rect 38657 24565 38669 24568
rect 38703 24565 38715 24599
rect 38657 24559 38715 24565
rect 39025 24599 39083 24605
rect 39025 24565 39037 24599
rect 39071 24596 39083 24599
rect 39114 24596 39120 24608
rect 39071 24568 39120 24596
rect 39071 24565 39083 24568
rect 39025 24559 39083 24565
rect 39114 24556 39120 24568
rect 39172 24556 39178 24608
rect 41785 24599 41843 24605
rect 41785 24565 41797 24599
rect 41831 24596 41843 24599
rect 43070 24596 43076 24608
rect 41831 24568 43076 24596
rect 41831 24565 41843 24568
rect 41785 24559 41843 24565
rect 43070 24556 43076 24568
rect 43128 24556 43134 24608
rect 44450 24556 44456 24608
rect 44508 24556 44514 24608
rect 1104 24506 44896 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 44896 24506
rect 1104 24432 44896 24454
rect 7837 24395 7895 24401
rect 7837 24361 7849 24395
rect 7883 24392 7895 24395
rect 9674 24392 9680 24404
rect 7883 24364 9680 24392
rect 7883 24361 7895 24364
rect 7837 24355 7895 24361
rect 9674 24352 9680 24364
rect 9732 24352 9738 24404
rect 9766 24352 9772 24404
rect 9824 24392 9830 24404
rect 9950 24392 9956 24404
rect 9824 24364 9956 24392
rect 9824 24352 9830 24364
rect 9950 24352 9956 24364
rect 10008 24352 10014 24404
rect 10781 24395 10839 24401
rect 10781 24361 10793 24395
rect 10827 24392 10839 24395
rect 11698 24392 11704 24404
rect 10827 24364 11704 24392
rect 10827 24361 10839 24364
rect 10781 24355 10839 24361
rect 11698 24352 11704 24364
rect 11756 24352 11762 24404
rect 12802 24352 12808 24404
rect 12860 24352 12866 24404
rect 13354 24352 13360 24404
rect 13412 24352 13418 24404
rect 13814 24352 13820 24404
rect 13872 24392 13878 24404
rect 14182 24392 14188 24404
rect 13872 24364 14188 24392
rect 13872 24352 13878 24364
rect 14182 24352 14188 24364
rect 14240 24352 14246 24404
rect 14366 24352 14372 24404
rect 14424 24392 14430 24404
rect 15105 24395 15163 24401
rect 15105 24392 15117 24395
rect 14424 24364 15117 24392
rect 14424 24352 14430 24364
rect 15105 24361 15117 24364
rect 15151 24361 15163 24395
rect 15105 24355 15163 24361
rect 15381 24395 15439 24401
rect 15381 24361 15393 24395
rect 15427 24392 15439 24395
rect 15470 24392 15476 24404
rect 15427 24364 15476 24392
rect 15427 24361 15439 24364
rect 15381 24355 15439 24361
rect 5442 24284 5448 24336
rect 5500 24324 5506 24336
rect 5500 24296 11008 24324
rect 5500 24284 5506 24296
rect 7282 24216 7288 24268
rect 7340 24256 7346 24268
rect 7745 24259 7803 24265
rect 7745 24256 7757 24259
rect 7340 24228 7757 24256
rect 7340 24216 7346 24228
rect 7745 24225 7757 24228
rect 7791 24225 7803 24259
rect 7745 24219 7803 24225
rect 10042 24216 10048 24268
rect 10100 24216 10106 24268
rect 10410 24256 10416 24268
rect 10152 24228 10416 24256
rect 7466 24148 7472 24200
rect 7524 24188 7530 24200
rect 7653 24191 7711 24197
rect 7653 24188 7665 24191
rect 7524 24160 7665 24188
rect 7524 24148 7530 24160
rect 7653 24157 7665 24160
rect 7699 24157 7711 24191
rect 10152 24188 10180 24228
rect 10410 24216 10416 24228
rect 10468 24216 10474 24268
rect 10686 24216 10692 24268
rect 10744 24216 10750 24268
rect 10870 24256 10876 24268
rect 10796 24228 10876 24256
rect 7653 24151 7711 24157
rect 7852 24160 10180 24188
rect 10229 24191 10287 24197
rect 7742 24080 7748 24132
rect 7800 24120 7806 24132
rect 7852 24120 7880 24160
rect 10229 24157 10241 24191
rect 10275 24188 10287 24191
rect 10318 24188 10324 24200
rect 10275 24160 10324 24188
rect 10275 24157 10287 24160
rect 10229 24151 10287 24157
rect 10318 24148 10324 24160
rect 10376 24148 10382 24200
rect 10796 24197 10824 24228
rect 10870 24216 10876 24228
rect 10928 24216 10934 24268
rect 10774 24191 10832 24197
rect 10428 24160 10640 24188
rect 9766 24120 9772 24132
rect 7800 24092 7880 24120
rect 7944 24092 9772 24120
rect 7800 24080 7806 24092
rect 2774 24012 2780 24064
rect 2832 24052 2838 24064
rect 7944 24052 7972 24092
rect 9766 24080 9772 24092
rect 9824 24080 9830 24132
rect 9953 24123 10011 24129
rect 9953 24089 9965 24123
rect 9999 24120 10011 24123
rect 10428 24120 10456 24160
rect 10612 24132 10640 24160
rect 10774 24157 10786 24191
rect 10820 24157 10832 24191
rect 10980 24188 11008 24296
rect 11606 24284 11612 24336
rect 11664 24324 11670 24336
rect 11790 24324 11796 24336
rect 11664 24296 11796 24324
rect 11664 24284 11670 24296
rect 11790 24284 11796 24296
rect 11848 24324 11854 24336
rect 14918 24324 14924 24336
rect 11848 24296 14924 24324
rect 11848 24284 11854 24296
rect 14918 24284 14924 24296
rect 14976 24284 14982 24336
rect 15120 24324 15148 24355
rect 15470 24352 15476 24364
rect 15528 24352 15534 24404
rect 16298 24352 16304 24404
rect 16356 24352 16362 24404
rect 16482 24352 16488 24404
rect 16540 24352 16546 24404
rect 16942 24352 16948 24404
rect 17000 24352 17006 24404
rect 17218 24352 17224 24404
rect 17276 24352 17282 24404
rect 17865 24395 17923 24401
rect 17865 24361 17877 24395
rect 17911 24392 17923 24395
rect 17911 24364 18092 24392
rect 17911 24361 17923 24364
rect 17865 24355 17923 24361
rect 15120 24296 18000 24324
rect 13541 24259 13599 24265
rect 13541 24225 13553 24259
rect 13587 24256 13599 24259
rect 14090 24256 14096 24268
rect 13587 24228 14096 24256
rect 13587 24225 13599 24228
rect 13541 24219 13599 24225
rect 14090 24216 14096 24228
rect 14148 24216 14154 24268
rect 14182 24216 14188 24268
rect 14240 24256 14246 24268
rect 14826 24256 14832 24268
rect 14240 24228 14832 24256
rect 14240 24216 14246 24228
rect 14826 24216 14832 24228
rect 14884 24216 14890 24268
rect 15028 24228 15240 24256
rect 12710 24188 12716 24200
rect 10980 24160 12716 24188
rect 10774 24151 10832 24157
rect 12710 24148 12716 24160
rect 12768 24148 12774 24200
rect 12894 24148 12900 24200
rect 12952 24148 12958 24200
rect 13633 24191 13691 24197
rect 13633 24157 13645 24191
rect 13679 24188 13691 24191
rect 15028 24188 15056 24228
rect 13679 24160 15056 24188
rect 13679 24157 13691 24160
rect 13633 24151 13691 24157
rect 15102 24148 15108 24200
rect 15160 24148 15166 24200
rect 15212 24197 15240 24228
rect 15930 24216 15936 24268
rect 15988 24256 15994 24268
rect 16117 24259 16175 24265
rect 16117 24256 16129 24259
rect 15988 24228 16129 24256
rect 15988 24216 15994 24228
rect 16117 24225 16129 24228
rect 16163 24225 16175 24259
rect 16390 24256 16396 24268
rect 16117 24219 16175 24225
rect 16224 24228 16396 24256
rect 15197 24191 15255 24197
rect 15197 24157 15209 24191
rect 15243 24188 15255 24191
rect 16224 24188 16252 24228
rect 16390 24216 16396 24228
rect 16448 24216 16454 24268
rect 16850 24216 16856 24268
rect 16908 24216 16914 24268
rect 17218 24256 17224 24268
rect 17052 24228 17224 24256
rect 15243 24160 16252 24188
rect 16301 24191 16359 24197
rect 15243 24157 15255 24160
rect 15197 24151 15255 24157
rect 16301 24157 16313 24191
rect 16347 24157 16359 24191
rect 16301 24151 16359 24157
rect 9999 24092 10456 24120
rect 10505 24123 10563 24129
rect 9999 24089 10011 24092
rect 9953 24083 10011 24089
rect 10505 24089 10517 24123
rect 10551 24089 10563 24123
rect 10505 24083 10563 24089
rect 2832 24024 7972 24052
rect 8021 24055 8079 24061
rect 2832 24012 2838 24024
rect 8021 24021 8033 24055
rect 8067 24052 8079 24055
rect 8110 24052 8116 24064
rect 8067 24024 8116 24052
rect 8067 24021 8079 24024
rect 8021 24015 8079 24021
rect 8110 24012 8116 24024
rect 8168 24012 8174 24064
rect 9858 24012 9864 24064
rect 9916 24052 9922 24064
rect 10318 24052 10324 24064
rect 9916 24024 10324 24052
rect 9916 24012 9922 24024
rect 10318 24012 10324 24024
rect 10376 24012 10382 24064
rect 10413 24055 10471 24061
rect 10413 24021 10425 24055
rect 10459 24052 10471 24055
rect 10520 24052 10548 24083
rect 10594 24080 10600 24132
rect 10652 24080 10658 24132
rect 13357 24123 13415 24129
rect 13357 24089 13369 24123
rect 13403 24089 13415 24123
rect 13357 24083 13415 24089
rect 10459 24024 10548 24052
rect 10459 24021 10471 24024
rect 10413 24015 10471 24021
rect 10962 24012 10968 24064
rect 11020 24012 11026 24064
rect 13081 24055 13139 24061
rect 13081 24021 13093 24055
rect 13127 24052 13139 24055
rect 13372 24052 13400 24083
rect 14274 24080 14280 24132
rect 14332 24120 14338 24132
rect 14369 24123 14427 24129
rect 14369 24120 14381 24123
rect 14332 24092 14381 24120
rect 14332 24080 14338 24092
rect 14369 24089 14381 24092
rect 14415 24089 14427 24123
rect 14369 24083 14427 24089
rect 14550 24080 14556 24132
rect 14608 24080 14614 24132
rect 14737 24123 14795 24129
rect 14737 24089 14749 24123
rect 14783 24120 14795 24123
rect 14921 24123 14979 24129
rect 14921 24120 14933 24123
rect 14783 24092 14933 24120
rect 14783 24089 14795 24092
rect 14737 24083 14795 24089
rect 14921 24089 14933 24092
rect 14967 24120 14979 24123
rect 16025 24123 16083 24129
rect 16025 24120 16037 24123
rect 14967 24092 16037 24120
rect 14967 24089 14979 24092
rect 14921 24083 14979 24089
rect 16025 24089 16037 24092
rect 16071 24089 16083 24123
rect 16025 24083 16083 24089
rect 16206 24080 16212 24132
rect 16264 24120 16270 24132
rect 16316 24120 16344 24151
rect 16574 24148 16580 24200
rect 16632 24188 16638 24200
rect 17052 24197 17080 24228
rect 17218 24216 17224 24228
rect 17276 24216 17282 24268
rect 17678 24216 17684 24268
rect 17736 24256 17742 24268
rect 17773 24259 17831 24265
rect 17773 24256 17785 24259
rect 17736 24228 17785 24256
rect 17736 24216 17742 24228
rect 17773 24225 17785 24228
rect 17819 24225 17831 24259
rect 17773 24219 17831 24225
rect 17037 24191 17095 24197
rect 17037 24188 17049 24191
rect 16632 24160 17049 24188
rect 16632 24148 16638 24160
rect 17037 24157 17049 24160
rect 17083 24157 17095 24191
rect 17037 24151 17095 24157
rect 17494 24148 17500 24200
rect 17552 24188 17558 24200
rect 17862 24188 17868 24200
rect 17552 24160 17868 24188
rect 17552 24148 17558 24160
rect 17862 24148 17868 24160
rect 17920 24148 17926 24200
rect 17972 24197 18000 24296
rect 18064 24268 18092 24364
rect 18230 24352 18236 24404
rect 18288 24352 18294 24404
rect 18782 24352 18788 24404
rect 18840 24392 18846 24404
rect 19794 24392 19800 24404
rect 18840 24364 19800 24392
rect 18840 24352 18846 24364
rect 19794 24352 19800 24364
rect 19852 24352 19858 24404
rect 20070 24352 20076 24404
rect 20128 24392 20134 24404
rect 20254 24392 20260 24404
rect 20128 24364 20260 24392
rect 20128 24352 20134 24364
rect 20254 24352 20260 24364
rect 20312 24352 20318 24404
rect 22830 24352 22836 24404
rect 22888 24352 22894 24404
rect 23753 24395 23811 24401
rect 23753 24361 23765 24395
rect 23799 24392 23811 24395
rect 23842 24392 23848 24404
rect 23799 24364 23848 24392
rect 23799 24361 23811 24364
rect 23753 24355 23811 24361
rect 23842 24352 23848 24364
rect 23900 24352 23906 24404
rect 24118 24352 24124 24404
rect 24176 24392 24182 24404
rect 27890 24392 27896 24404
rect 24176 24364 27896 24392
rect 24176 24352 24182 24364
rect 27890 24352 27896 24364
rect 27948 24352 27954 24404
rect 27985 24395 28043 24401
rect 27985 24361 27997 24395
rect 28031 24361 28043 24395
rect 27985 24355 28043 24361
rect 18141 24327 18199 24333
rect 18141 24293 18153 24327
rect 18187 24324 18199 24327
rect 19058 24324 19064 24336
rect 18187 24296 19064 24324
rect 18187 24293 18199 24296
rect 18141 24287 18199 24293
rect 19058 24284 19064 24296
rect 19116 24284 19122 24336
rect 23017 24327 23075 24333
rect 23017 24293 23029 24327
rect 23063 24293 23075 24327
rect 23017 24287 23075 24293
rect 18046 24216 18052 24268
rect 18104 24256 18110 24268
rect 18322 24256 18328 24268
rect 18104 24228 18328 24256
rect 18104 24216 18110 24228
rect 18322 24216 18328 24228
rect 18380 24216 18386 24268
rect 19794 24216 19800 24268
rect 19852 24256 19858 24268
rect 21450 24256 21456 24268
rect 19852 24228 21456 24256
rect 19852 24216 19858 24228
rect 21450 24216 21456 24228
rect 21508 24216 21514 24268
rect 21542 24216 21548 24268
rect 21600 24256 21606 24268
rect 22278 24256 22284 24268
rect 21600 24228 22284 24256
rect 21600 24216 21606 24228
rect 22278 24216 22284 24228
rect 22336 24256 22342 24268
rect 22649 24259 22707 24265
rect 22649 24256 22661 24259
rect 22336 24228 22661 24256
rect 22336 24216 22342 24228
rect 22649 24225 22661 24228
rect 22695 24225 22707 24259
rect 22649 24219 22707 24225
rect 23032 24200 23060 24287
rect 23106 24284 23112 24336
rect 23164 24324 23170 24336
rect 23293 24327 23351 24333
rect 23293 24324 23305 24327
rect 23164 24296 23305 24324
rect 23164 24284 23170 24296
rect 23293 24293 23305 24296
rect 23339 24293 23351 24327
rect 23860 24324 23888 24352
rect 24762 24324 24768 24336
rect 23860 24296 24768 24324
rect 23293 24287 23351 24293
rect 24762 24284 24768 24296
rect 24820 24284 24826 24336
rect 25590 24284 25596 24336
rect 25648 24324 25654 24336
rect 27522 24324 27528 24336
rect 25648 24296 27528 24324
rect 25648 24284 25654 24296
rect 27522 24284 27528 24296
rect 27580 24284 27586 24336
rect 27614 24284 27620 24336
rect 27672 24324 27678 24336
rect 28000 24324 28028 24355
rect 28258 24352 28264 24404
rect 28316 24352 28322 24404
rect 29270 24352 29276 24404
rect 29328 24392 29334 24404
rect 29733 24395 29791 24401
rect 29733 24392 29745 24395
rect 29328 24364 29745 24392
rect 29328 24352 29334 24364
rect 29733 24361 29745 24364
rect 29779 24392 29791 24395
rect 29822 24392 29828 24404
rect 29779 24364 29828 24392
rect 29779 24361 29791 24364
rect 29733 24355 29791 24361
rect 29822 24352 29828 24364
rect 29880 24352 29886 24404
rect 30742 24352 30748 24404
rect 30800 24392 30806 24404
rect 31021 24395 31079 24401
rect 31021 24392 31033 24395
rect 30800 24364 31033 24392
rect 30800 24352 30806 24364
rect 31021 24361 31033 24364
rect 31067 24361 31079 24395
rect 31573 24395 31631 24401
rect 31573 24392 31585 24395
rect 31021 24355 31079 24361
rect 31305 24364 31585 24392
rect 27672 24296 28028 24324
rect 27672 24284 27678 24296
rect 28074 24284 28080 24336
rect 28132 24324 28138 24336
rect 31305 24324 31333 24364
rect 31573 24361 31585 24364
rect 31619 24361 31631 24395
rect 31573 24355 31631 24361
rect 31754 24352 31760 24404
rect 31812 24352 31818 24404
rect 31938 24352 31944 24404
rect 31996 24392 32002 24404
rect 33318 24392 33324 24404
rect 31996 24364 33324 24392
rect 31996 24352 32002 24364
rect 33318 24352 33324 24364
rect 33376 24352 33382 24404
rect 33870 24352 33876 24404
rect 33928 24392 33934 24404
rect 34057 24395 34115 24401
rect 34057 24392 34069 24395
rect 33928 24364 34069 24392
rect 33928 24352 33934 24364
rect 34057 24361 34069 24364
rect 34103 24392 34115 24395
rect 34330 24392 34336 24404
rect 34103 24364 34336 24392
rect 34103 24361 34115 24364
rect 34057 24355 34115 24361
rect 34330 24352 34336 24364
rect 34388 24352 34394 24404
rect 34422 24352 34428 24404
rect 34480 24392 34486 24404
rect 34701 24395 34759 24401
rect 34701 24392 34713 24395
rect 34480 24364 34713 24392
rect 34480 24352 34486 24364
rect 34701 24361 34713 24364
rect 34747 24361 34759 24395
rect 35253 24395 35311 24401
rect 35253 24392 35265 24395
rect 34701 24355 34759 24361
rect 34808 24364 35265 24392
rect 28132 24296 30880 24324
rect 28132 24284 28138 24296
rect 23198 24216 23204 24268
rect 23256 24256 23262 24268
rect 23566 24256 23572 24268
rect 23256 24228 23572 24256
rect 23256 24216 23262 24228
rect 17957 24191 18015 24197
rect 17957 24157 17969 24191
rect 18003 24157 18015 24191
rect 17957 24151 18015 24157
rect 18340 24160 22784 24188
rect 16264 24092 16344 24120
rect 16264 24080 16270 24092
rect 16666 24080 16672 24132
rect 16724 24120 16730 24132
rect 16761 24123 16819 24129
rect 16761 24120 16773 24123
rect 16724 24092 16773 24120
rect 16724 24080 16730 24092
rect 16761 24089 16773 24092
rect 16807 24120 16819 24123
rect 17681 24123 17739 24129
rect 17681 24120 17693 24123
rect 16807 24092 17693 24120
rect 16807 24089 16819 24092
rect 16761 24083 16819 24089
rect 17681 24089 17693 24092
rect 17727 24089 17739 24123
rect 17681 24083 17739 24089
rect 17770 24080 17776 24132
rect 17828 24120 17834 24132
rect 18340 24120 18368 24160
rect 17828 24092 18368 24120
rect 18417 24123 18475 24129
rect 17828 24080 17834 24092
rect 18417 24089 18429 24123
rect 18463 24120 18475 24123
rect 18506 24120 18512 24132
rect 18463 24092 18512 24120
rect 18463 24089 18475 24092
rect 18417 24083 18475 24089
rect 18506 24080 18512 24092
rect 18564 24080 18570 24132
rect 18601 24123 18659 24129
rect 18601 24089 18613 24123
rect 18647 24120 18659 24123
rect 18874 24120 18880 24132
rect 18647 24092 18880 24120
rect 18647 24089 18659 24092
rect 18601 24083 18659 24089
rect 18874 24080 18880 24092
rect 18932 24080 18938 24132
rect 21174 24080 21180 24132
rect 21232 24120 21238 24132
rect 22557 24123 22615 24129
rect 22557 24120 22569 24123
rect 21232 24092 22569 24120
rect 21232 24080 21238 24092
rect 22557 24089 22569 24092
rect 22603 24120 22615 24123
rect 22646 24120 22652 24132
rect 22603 24092 22652 24120
rect 22603 24089 22615 24092
rect 22557 24083 22615 24089
rect 22646 24080 22652 24092
rect 22704 24080 22710 24132
rect 22756 24120 22784 24160
rect 22830 24148 22836 24200
rect 22888 24148 22894 24200
rect 23014 24148 23020 24200
rect 23072 24148 23078 24200
rect 23492 24197 23520 24228
rect 23566 24216 23572 24228
rect 23624 24216 23630 24268
rect 23661 24259 23719 24265
rect 23661 24225 23673 24259
rect 23707 24256 23719 24259
rect 24670 24256 24676 24268
rect 23707 24228 24676 24256
rect 23707 24225 23719 24228
rect 23661 24219 23719 24225
rect 23477 24191 23535 24197
rect 23477 24157 23489 24191
rect 23523 24157 23535 24191
rect 23477 24151 23535 24157
rect 23676 24120 23704 24219
rect 24670 24216 24676 24228
rect 24728 24216 24734 24268
rect 25222 24216 25228 24268
rect 25280 24256 25286 24268
rect 30098 24256 30104 24268
rect 25280 24228 30104 24256
rect 25280 24216 25286 24228
rect 30098 24216 30104 24228
rect 30156 24216 30162 24268
rect 24854 24148 24860 24200
rect 24912 24188 24918 24200
rect 27614 24188 27620 24200
rect 24912 24160 27620 24188
rect 24912 24148 24918 24160
rect 27614 24148 27620 24160
rect 27672 24148 27678 24200
rect 27982 24148 27988 24200
rect 28040 24148 28046 24200
rect 28077 24191 28135 24197
rect 28077 24157 28089 24191
rect 28123 24157 28135 24191
rect 28077 24151 28135 24157
rect 22756 24092 23704 24120
rect 23753 24123 23811 24129
rect 23753 24089 23765 24123
rect 23799 24120 23811 24123
rect 23842 24120 23848 24132
rect 23799 24092 23848 24120
rect 23799 24089 23811 24092
rect 23753 24083 23811 24089
rect 23842 24080 23848 24092
rect 23900 24080 23906 24132
rect 25130 24080 25136 24132
rect 25188 24120 25194 24132
rect 26050 24120 26056 24132
rect 25188 24092 26056 24120
rect 25188 24080 25194 24092
rect 26050 24080 26056 24092
rect 26108 24080 26114 24132
rect 26418 24120 26424 24132
rect 26160 24092 26424 24120
rect 13127 24024 13400 24052
rect 13127 24021 13139 24024
rect 13081 24015 13139 24021
rect 13814 24012 13820 24064
rect 13872 24012 13878 24064
rect 14090 24012 14096 24064
rect 14148 24052 14154 24064
rect 16942 24052 16948 24064
rect 14148 24024 16948 24052
rect 14148 24012 14154 24024
rect 16942 24012 16948 24024
rect 17000 24012 17006 24064
rect 17218 24012 17224 24064
rect 17276 24052 17282 24064
rect 19426 24052 19432 24064
rect 17276 24024 19432 24052
rect 17276 24012 17282 24024
rect 19426 24012 19432 24024
rect 19484 24012 19490 24064
rect 19702 24012 19708 24064
rect 19760 24052 19766 24064
rect 23382 24052 23388 24064
rect 19760 24024 23388 24052
rect 19760 24012 19766 24024
rect 23382 24012 23388 24024
rect 23440 24012 23446 24064
rect 24118 24012 24124 24064
rect 24176 24052 24182 24064
rect 24394 24052 24400 24064
rect 24176 24024 24400 24052
rect 24176 24012 24182 24024
rect 24394 24012 24400 24024
rect 24452 24012 24458 24064
rect 24486 24012 24492 24064
rect 24544 24052 24550 24064
rect 24762 24052 24768 24064
rect 24544 24024 24768 24052
rect 24544 24012 24550 24024
rect 24762 24012 24768 24024
rect 24820 24012 24826 24064
rect 24946 24012 24952 24064
rect 25004 24052 25010 24064
rect 26160 24052 26188 24092
rect 26418 24080 26424 24092
rect 26476 24080 26482 24132
rect 26878 24080 26884 24132
rect 26936 24120 26942 24132
rect 27154 24120 27160 24132
rect 26936 24092 27160 24120
rect 26936 24080 26942 24092
rect 27154 24080 27160 24092
rect 27212 24120 27218 24132
rect 27801 24123 27859 24129
rect 27801 24120 27813 24123
rect 27212 24092 27813 24120
rect 27212 24080 27218 24092
rect 27801 24089 27813 24092
rect 27847 24089 27859 24123
rect 27801 24083 27859 24089
rect 27890 24080 27896 24132
rect 27948 24120 27954 24132
rect 28092 24120 28120 24151
rect 28350 24148 28356 24200
rect 28408 24148 28414 24200
rect 28534 24148 28540 24200
rect 28592 24148 28598 24200
rect 29546 24148 29552 24200
rect 29604 24148 29610 24200
rect 29733 24191 29791 24197
rect 29733 24157 29745 24191
rect 29779 24157 29791 24191
rect 30852 24188 30880 24296
rect 31220 24296 31333 24324
rect 31481 24327 31539 24333
rect 30926 24216 30932 24268
rect 30984 24256 30990 24268
rect 31220 24265 31248 24296
rect 31481 24293 31493 24327
rect 31527 24324 31539 24327
rect 32122 24324 32128 24336
rect 31527 24296 32128 24324
rect 31527 24293 31539 24296
rect 31481 24287 31539 24293
rect 32122 24284 32128 24296
rect 32180 24284 32186 24336
rect 32214 24284 32220 24336
rect 32272 24324 32278 24336
rect 34808 24324 34836 24364
rect 35253 24361 35265 24364
rect 35299 24392 35311 24395
rect 35618 24392 35624 24404
rect 35299 24364 35624 24392
rect 35299 24361 35311 24364
rect 35253 24355 35311 24361
rect 35618 24352 35624 24364
rect 35676 24352 35682 24404
rect 35713 24395 35771 24401
rect 35713 24361 35725 24395
rect 35759 24392 35771 24395
rect 36265 24395 36323 24401
rect 36265 24392 36277 24395
rect 35759 24364 36277 24392
rect 35759 24361 35771 24364
rect 35713 24355 35771 24361
rect 36265 24361 36277 24364
rect 36311 24361 36323 24395
rect 36265 24355 36323 24361
rect 34974 24324 34980 24336
rect 32272 24296 34836 24324
rect 34900 24296 34980 24324
rect 32272 24284 32278 24296
rect 31205 24259 31263 24265
rect 31205 24256 31217 24259
rect 30984 24228 31217 24256
rect 30984 24216 30990 24228
rect 31205 24225 31217 24228
rect 31251 24225 31263 24259
rect 31662 24256 31668 24268
rect 31205 24219 31263 24225
rect 31305 24228 31668 24256
rect 31305 24198 31333 24228
rect 31662 24216 31668 24228
rect 31720 24216 31726 24268
rect 31846 24216 31852 24268
rect 31904 24216 31910 24268
rect 32490 24216 32496 24268
rect 32548 24256 32554 24268
rect 33870 24256 33876 24268
rect 32548 24228 33876 24256
rect 32548 24216 32554 24228
rect 33870 24216 33876 24228
rect 33928 24216 33934 24268
rect 33962 24216 33968 24268
rect 34020 24256 34026 24268
rect 34900 24265 34928 24296
rect 34974 24284 34980 24296
rect 35032 24284 35038 24336
rect 35161 24327 35219 24333
rect 35161 24293 35173 24327
rect 35207 24324 35219 24327
rect 35207 24296 36400 24324
rect 35207 24293 35219 24296
rect 35161 24287 35219 24293
rect 34149 24259 34207 24265
rect 34149 24256 34161 24259
rect 34020 24228 34161 24256
rect 34020 24216 34026 24228
rect 34149 24225 34161 24228
rect 34195 24225 34207 24259
rect 34149 24219 34207 24225
rect 34885 24259 34943 24265
rect 34885 24225 34897 24259
rect 34931 24225 34943 24259
rect 35710 24256 35716 24268
rect 34885 24219 34943 24225
rect 35268 24228 35716 24256
rect 31305 24197 31340 24198
rect 31297 24191 31355 24197
rect 30852 24160 31248 24188
rect 29733 24151 29791 24157
rect 27948 24092 28120 24120
rect 28721 24123 28779 24129
rect 27948 24080 27954 24092
rect 28721 24089 28733 24123
rect 28767 24120 28779 24123
rect 29086 24120 29092 24132
rect 28767 24092 29092 24120
rect 28767 24089 28779 24092
rect 28721 24083 28779 24089
rect 29086 24080 29092 24092
rect 29144 24080 29150 24132
rect 25004 24024 26188 24052
rect 25004 24012 25010 24024
rect 26326 24012 26332 24064
rect 26384 24052 26390 24064
rect 29748 24052 29776 24151
rect 31021 24123 31079 24129
rect 31021 24120 31033 24123
rect 29932 24092 31033 24120
rect 29932 24061 29960 24092
rect 31021 24089 31033 24092
rect 31067 24089 31079 24123
rect 31220 24120 31248 24160
rect 31297 24157 31309 24191
rect 31343 24157 31355 24191
rect 31297 24151 31355 24157
rect 31941 24191 31999 24197
rect 31941 24157 31953 24191
rect 31987 24188 31999 24191
rect 32306 24188 32312 24200
rect 31987 24160 32312 24188
rect 31987 24157 31999 24160
rect 31941 24151 31999 24157
rect 32306 24148 32312 24160
rect 32364 24148 32370 24200
rect 34333 24191 34391 24197
rect 34333 24157 34345 24191
rect 34379 24188 34391 24191
rect 34379 24160 34928 24188
rect 34379 24157 34391 24160
rect 34333 24151 34391 24157
rect 34057 24123 34115 24129
rect 34057 24120 34069 24123
rect 31220 24092 34069 24120
rect 31021 24083 31079 24089
rect 34057 24089 34069 24092
rect 34103 24120 34115 24123
rect 34701 24123 34759 24129
rect 34701 24120 34713 24123
rect 34103 24092 34713 24120
rect 34103 24089 34115 24092
rect 34057 24083 34115 24089
rect 34701 24089 34713 24092
rect 34747 24089 34759 24123
rect 34701 24083 34759 24089
rect 26384 24024 29776 24052
rect 29917 24055 29975 24061
rect 26384 24012 26390 24024
rect 29917 24021 29929 24055
rect 29963 24021 29975 24055
rect 29917 24015 29975 24021
rect 30098 24012 30104 24064
rect 30156 24052 30162 24064
rect 34146 24052 34152 24064
rect 30156 24024 34152 24052
rect 30156 24012 30162 24024
rect 34146 24012 34152 24024
rect 34204 24012 34210 24064
rect 34517 24055 34575 24061
rect 34517 24021 34529 24055
rect 34563 24052 34575 24055
rect 34606 24052 34612 24064
rect 34563 24024 34612 24052
rect 34563 24021 34575 24024
rect 34517 24015 34575 24021
rect 34606 24012 34612 24024
rect 34664 24012 34670 24064
rect 34900 24052 34928 24160
rect 34974 24148 34980 24200
rect 35032 24148 35038 24200
rect 35268 24197 35296 24228
rect 35710 24216 35716 24228
rect 35768 24216 35774 24268
rect 36372 24265 36400 24296
rect 36357 24259 36415 24265
rect 36357 24225 36369 24259
rect 36403 24225 36415 24259
rect 36357 24219 36415 24225
rect 42978 24216 42984 24268
rect 43036 24216 43042 24268
rect 35253 24191 35311 24197
rect 35253 24157 35265 24191
rect 35299 24157 35311 24191
rect 35253 24151 35311 24157
rect 35434 24148 35440 24200
rect 35492 24148 35498 24200
rect 35526 24148 35532 24200
rect 35584 24148 35590 24200
rect 35618 24148 35624 24200
rect 35676 24188 35682 24200
rect 35805 24191 35863 24197
rect 35805 24188 35817 24191
rect 35676 24160 35817 24188
rect 35676 24148 35682 24160
rect 35805 24157 35817 24160
rect 35851 24157 35863 24191
rect 35805 24151 35863 24157
rect 35989 24191 36047 24197
rect 35989 24157 36001 24191
rect 36035 24188 36047 24191
rect 36078 24188 36084 24200
rect 36035 24160 36084 24188
rect 36035 24157 36047 24160
rect 35989 24151 36047 24157
rect 36078 24148 36084 24160
rect 36136 24148 36142 24200
rect 36262 24148 36268 24200
rect 36320 24148 36326 24200
rect 36814 24148 36820 24200
rect 36872 24188 36878 24200
rect 37734 24188 37740 24200
rect 36872 24160 37740 24188
rect 36872 24148 36878 24160
rect 37734 24148 37740 24160
rect 37792 24148 37798 24200
rect 40310 24148 40316 24200
rect 40368 24188 40374 24200
rect 40589 24191 40647 24197
rect 40589 24188 40601 24191
rect 40368 24160 40601 24188
rect 40368 24148 40374 24160
rect 40589 24157 40601 24160
rect 40635 24188 40647 24191
rect 41782 24188 41788 24200
rect 40635 24160 41788 24188
rect 40635 24157 40647 24160
rect 40589 24151 40647 24157
rect 41782 24148 41788 24160
rect 41840 24148 41846 24200
rect 44269 24191 44327 24197
rect 44269 24188 44281 24191
rect 42996 24160 44281 24188
rect 34992 24120 35020 24148
rect 36998 24120 37004 24132
rect 34992 24092 37004 24120
rect 36998 24080 37004 24092
rect 37056 24080 37062 24132
rect 40856 24123 40914 24129
rect 40856 24089 40868 24123
rect 40902 24120 40914 24123
rect 41046 24120 41052 24132
rect 40902 24092 41052 24120
rect 40902 24089 40914 24092
rect 40856 24083 40914 24089
rect 41046 24080 41052 24092
rect 41104 24080 41110 24132
rect 42996 24064 43024 24160
rect 44269 24157 44281 24160
rect 44315 24157 44327 24191
rect 44269 24151 44327 24157
rect 36173 24055 36231 24061
rect 36173 24052 36185 24055
rect 34900 24024 36185 24052
rect 36173 24021 36185 24024
rect 36219 24052 36231 24055
rect 36538 24052 36544 24064
rect 36219 24024 36544 24052
rect 36219 24021 36231 24024
rect 36173 24015 36231 24021
rect 36538 24012 36544 24024
rect 36596 24012 36602 24064
rect 36633 24055 36691 24061
rect 36633 24021 36645 24055
rect 36679 24052 36691 24055
rect 41874 24052 41880 24064
rect 36679 24024 41880 24052
rect 36679 24021 36691 24024
rect 36633 24015 36691 24021
rect 41874 24012 41880 24024
rect 41932 24012 41938 24064
rect 41969 24055 42027 24061
rect 41969 24021 41981 24055
rect 42015 24052 42027 24055
rect 42978 24052 42984 24064
rect 42015 24024 42984 24052
rect 42015 24021 42027 24024
rect 41969 24015 42027 24021
rect 42978 24012 42984 24024
rect 43036 24012 43042 24064
rect 43622 24012 43628 24064
rect 43680 24012 43686 24064
rect 44450 24012 44456 24064
rect 44508 24012 44514 24064
rect 1104 23962 44896 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 44896 23962
rect 1104 23888 44896 23910
rect 7190 23808 7196 23860
rect 7248 23808 7254 23860
rect 7374 23808 7380 23860
rect 7432 23808 7438 23860
rect 7466 23808 7472 23860
rect 7524 23808 7530 23860
rect 9766 23808 9772 23860
rect 9824 23848 9830 23860
rect 9824 23820 10272 23848
rect 9824 23808 9830 23820
rect 4614 23780 4620 23792
rect 4172 23752 4620 23780
rect 4172 23721 4200 23752
rect 4614 23740 4620 23752
rect 4672 23740 4678 23792
rect 6270 23740 6276 23792
rect 6328 23780 6334 23792
rect 6917 23783 6975 23789
rect 6917 23780 6929 23783
rect 6328 23752 6929 23780
rect 6328 23740 6334 23752
rect 6917 23749 6929 23752
rect 6963 23780 6975 23783
rect 7208 23780 7236 23808
rect 6963 23752 7236 23780
rect 9493 23783 9551 23789
rect 6963 23749 6975 23752
rect 6917 23743 6975 23749
rect 9493 23749 9505 23783
rect 9539 23780 9551 23783
rect 9674 23780 9680 23792
rect 9539 23752 9680 23780
rect 9539 23749 9551 23752
rect 9493 23743 9551 23749
rect 9674 23740 9680 23752
rect 9732 23780 9738 23792
rect 9732 23752 9904 23780
rect 9732 23740 9738 23752
rect 4157 23715 4215 23721
rect 4157 23681 4169 23715
rect 4203 23681 4215 23715
rect 4157 23675 4215 23681
rect 4246 23672 4252 23724
rect 4304 23712 4310 23724
rect 4341 23715 4399 23721
rect 4341 23712 4353 23715
rect 4304 23684 4353 23712
rect 4304 23672 4310 23684
rect 4341 23681 4353 23684
rect 4387 23681 4399 23715
rect 4341 23675 4399 23681
rect 4430 23672 4436 23724
rect 4488 23672 4494 23724
rect 4530 23715 4588 23721
rect 4530 23681 4542 23715
rect 4576 23681 4588 23715
rect 4530 23675 4588 23681
rect 7193 23715 7251 23721
rect 7193 23681 7205 23715
rect 7239 23712 7251 23715
rect 7653 23715 7711 23721
rect 7653 23712 7665 23715
rect 7239 23684 7665 23712
rect 7239 23681 7251 23684
rect 7193 23675 7251 23681
rect 7653 23681 7665 23684
rect 7699 23712 7711 23715
rect 7699 23684 7880 23712
rect 7699 23681 7711 23684
rect 7653 23675 7711 23681
rect 3418 23604 3424 23656
rect 3476 23644 3482 23656
rect 4540 23644 4568 23675
rect 3476 23616 4568 23644
rect 7101 23647 7159 23653
rect 3476 23604 3482 23616
rect 7101 23613 7113 23647
rect 7147 23644 7159 23647
rect 7282 23644 7288 23656
rect 7147 23616 7288 23644
rect 7147 23613 7159 23616
rect 7101 23607 7159 23613
rect 7282 23604 7288 23616
rect 7340 23604 7346 23656
rect 7742 23604 7748 23656
rect 7800 23604 7806 23656
rect 7852 23644 7880 23684
rect 7926 23672 7932 23724
rect 7984 23672 7990 23724
rect 9217 23715 9275 23721
rect 9217 23681 9229 23715
rect 9263 23681 9275 23715
rect 9217 23675 9275 23681
rect 9401 23715 9459 23721
rect 9401 23681 9413 23715
rect 9447 23681 9459 23715
rect 9401 23675 9459 23681
rect 9585 23715 9643 23721
rect 9585 23681 9597 23715
rect 9631 23712 9643 23715
rect 9766 23712 9772 23724
rect 9631 23684 9772 23712
rect 9631 23681 9643 23684
rect 9585 23675 9643 23681
rect 8570 23644 8576 23656
rect 7852 23616 8576 23644
rect 8570 23604 8576 23616
rect 8628 23604 8634 23656
rect 4430 23536 4436 23588
rect 4488 23576 4494 23588
rect 4798 23576 4804 23588
rect 4488 23548 4804 23576
rect 4488 23536 4494 23548
rect 4798 23536 4804 23548
rect 4856 23536 4862 23588
rect 8018 23576 8024 23588
rect 7208 23548 8024 23576
rect 7208 23520 7236 23548
rect 8018 23536 8024 23548
rect 8076 23536 8082 23588
rect 8110 23536 8116 23588
rect 8168 23576 8174 23588
rect 9232 23576 9260 23675
rect 9416 23644 9444 23675
rect 9766 23672 9772 23684
rect 9824 23672 9830 23724
rect 9876 23721 9904 23752
rect 9861 23715 9919 23721
rect 9861 23681 9873 23715
rect 9907 23681 9919 23715
rect 9861 23675 9919 23681
rect 9950 23672 9956 23724
rect 10008 23712 10014 23724
rect 10244 23721 10272 23820
rect 10318 23808 10324 23860
rect 10376 23808 10382 23860
rect 10413 23851 10471 23857
rect 10413 23817 10425 23851
rect 10459 23848 10471 23851
rect 10778 23848 10784 23860
rect 10459 23820 10784 23848
rect 10459 23817 10471 23820
rect 10413 23811 10471 23817
rect 10778 23808 10784 23820
rect 10836 23808 10842 23860
rect 14274 23808 14280 23860
rect 14332 23848 14338 23860
rect 14550 23848 14556 23860
rect 14332 23820 14556 23848
rect 14332 23808 14338 23820
rect 14550 23808 14556 23820
rect 14608 23808 14614 23860
rect 15654 23808 15660 23860
rect 15712 23808 15718 23860
rect 16942 23808 16948 23860
rect 17000 23848 17006 23860
rect 20070 23848 20076 23860
rect 17000 23820 20076 23848
rect 17000 23808 17006 23820
rect 20070 23808 20076 23820
rect 20128 23808 20134 23860
rect 20625 23851 20683 23857
rect 20625 23817 20637 23851
rect 20671 23848 20683 23851
rect 20990 23848 20996 23860
rect 20671 23820 20996 23848
rect 20671 23817 20683 23820
rect 20625 23811 20683 23817
rect 20990 23808 20996 23820
rect 21048 23808 21054 23860
rect 26237 23851 26295 23857
rect 26237 23817 26249 23851
rect 26283 23848 26295 23851
rect 26970 23848 26976 23860
rect 26283 23820 26976 23848
rect 26283 23817 26295 23820
rect 26237 23811 26295 23817
rect 26970 23808 26976 23820
rect 27028 23808 27034 23860
rect 27430 23808 27436 23860
rect 27488 23848 27494 23860
rect 28994 23848 29000 23860
rect 27488 23820 29000 23848
rect 27488 23808 27494 23820
rect 28994 23808 29000 23820
rect 29052 23808 29058 23860
rect 29546 23808 29552 23860
rect 29604 23808 29610 23860
rect 29914 23808 29920 23860
rect 29972 23848 29978 23860
rect 30098 23848 30104 23860
rect 29972 23820 30104 23848
rect 29972 23808 29978 23820
rect 30098 23808 30104 23820
rect 30156 23808 30162 23860
rect 30193 23851 30251 23857
rect 30193 23817 30205 23851
rect 30239 23848 30251 23851
rect 31846 23848 31852 23860
rect 30239 23820 31852 23848
rect 30239 23817 30251 23820
rect 30193 23811 30251 23817
rect 31846 23808 31852 23820
rect 31904 23808 31910 23860
rect 32306 23848 32312 23860
rect 31956 23820 32312 23848
rect 10336 23780 10364 23808
rect 10870 23780 10876 23792
rect 10336 23752 10876 23780
rect 10870 23740 10876 23752
rect 10928 23740 10934 23792
rect 12710 23740 12716 23792
rect 12768 23780 12774 23792
rect 20441 23783 20499 23789
rect 12768 23752 20392 23780
rect 12768 23740 12774 23752
rect 10045 23715 10103 23721
rect 10045 23712 10057 23715
rect 10008 23684 10057 23712
rect 10008 23672 10014 23684
rect 10045 23681 10057 23684
rect 10091 23681 10103 23715
rect 10045 23675 10103 23681
rect 10137 23715 10195 23721
rect 10137 23681 10149 23715
rect 10183 23681 10195 23715
rect 10137 23675 10195 23681
rect 10229 23715 10287 23721
rect 10229 23681 10241 23715
rect 10275 23712 10287 23715
rect 10318 23712 10324 23724
rect 10275 23684 10324 23712
rect 10275 23681 10287 23684
rect 10229 23675 10287 23681
rect 9968 23644 9996 23672
rect 9416 23616 9996 23644
rect 10152 23644 10180 23675
rect 10318 23672 10324 23684
rect 10376 23672 10382 23724
rect 13449 23715 13507 23721
rect 13449 23681 13461 23715
rect 13495 23712 13507 23715
rect 13538 23712 13544 23724
rect 13495 23684 13544 23712
rect 13495 23681 13507 23684
rect 13449 23675 13507 23681
rect 13538 23672 13544 23684
rect 13596 23672 13602 23724
rect 13630 23672 13636 23724
rect 13688 23672 13694 23724
rect 13817 23715 13875 23721
rect 13817 23681 13829 23715
rect 13863 23712 13875 23715
rect 13906 23712 13912 23724
rect 13863 23684 13912 23712
rect 13863 23681 13875 23684
rect 13817 23675 13875 23681
rect 13906 23672 13912 23684
rect 13964 23712 13970 23724
rect 15010 23712 15016 23724
rect 13964 23684 15016 23712
rect 13964 23672 13970 23684
rect 15010 23672 15016 23684
rect 15068 23672 15074 23724
rect 15197 23715 15255 23721
rect 15197 23681 15209 23715
rect 15243 23712 15255 23715
rect 15378 23712 15384 23724
rect 15243 23684 15384 23712
rect 15243 23681 15255 23684
rect 15197 23675 15255 23681
rect 15378 23672 15384 23684
rect 15436 23672 15442 23724
rect 15470 23672 15476 23724
rect 15528 23672 15534 23724
rect 20162 23672 20168 23724
rect 20220 23712 20226 23724
rect 20257 23715 20315 23721
rect 20257 23712 20269 23715
rect 20220 23684 20269 23712
rect 20220 23672 20226 23684
rect 20257 23681 20269 23684
rect 20303 23681 20315 23715
rect 20364 23712 20392 23752
rect 20441 23749 20453 23783
rect 20487 23780 20499 23783
rect 23569 23783 23627 23789
rect 23569 23780 23581 23783
rect 20487 23752 23581 23780
rect 20487 23749 20499 23752
rect 20441 23743 20499 23749
rect 23569 23749 23581 23752
rect 23615 23780 23627 23783
rect 24118 23780 24124 23792
rect 23615 23752 24124 23780
rect 23615 23749 23627 23752
rect 23569 23743 23627 23749
rect 24118 23740 24124 23752
rect 24176 23740 24182 23792
rect 24857 23783 24915 23789
rect 24857 23780 24869 23783
rect 24780 23752 24869 23780
rect 22833 23715 22891 23721
rect 22833 23712 22845 23715
rect 20364 23684 22845 23712
rect 20257 23675 20315 23681
rect 22833 23681 22845 23684
rect 22879 23712 22891 23715
rect 23385 23715 23443 23721
rect 23385 23712 23397 23715
rect 22879 23684 23397 23712
rect 22879 23681 22891 23684
rect 22833 23675 22891 23681
rect 23385 23681 23397 23684
rect 23431 23681 23443 23715
rect 23385 23675 23443 23681
rect 24486 23672 24492 23724
rect 24544 23712 24550 23724
rect 24780 23712 24808 23752
rect 24857 23749 24869 23752
rect 24903 23749 24915 23783
rect 24857 23743 24915 23749
rect 24946 23740 24952 23792
rect 25004 23780 25010 23792
rect 25041 23783 25099 23789
rect 25041 23780 25053 23783
rect 25004 23752 25053 23780
rect 25004 23740 25010 23752
rect 25041 23749 25053 23752
rect 25087 23749 25099 23783
rect 25041 23743 25099 23749
rect 25130 23740 25136 23792
rect 25188 23780 25194 23792
rect 25188 23752 26096 23780
rect 25188 23740 25194 23752
rect 24544 23684 24808 23712
rect 24544 23672 24550 23684
rect 25590 23672 25596 23724
rect 25648 23712 25654 23724
rect 25777 23715 25835 23721
rect 25777 23712 25789 23715
rect 25648 23684 25789 23712
rect 25648 23672 25654 23684
rect 25777 23681 25789 23684
rect 25823 23681 25835 23715
rect 25777 23675 25835 23681
rect 10152 23616 10272 23644
rect 9769 23579 9827 23585
rect 8168 23548 9536 23576
rect 8168 23536 8174 23548
rect 9508 23520 9536 23548
rect 9769 23545 9781 23579
rect 9815 23576 9827 23579
rect 10134 23576 10140 23588
rect 9815 23548 10140 23576
rect 9815 23545 9827 23548
rect 9769 23539 9827 23545
rect 10134 23536 10140 23548
rect 10192 23536 10198 23588
rect 4709 23511 4767 23517
rect 4709 23477 4721 23511
rect 4755 23508 4767 23511
rect 5350 23508 5356 23520
rect 4755 23480 5356 23508
rect 4755 23477 4767 23480
rect 4709 23471 4767 23477
rect 5350 23468 5356 23480
rect 5408 23468 5414 23520
rect 7190 23468 7196 23520
rect 7248 23468 7254 23520
rect 7466 23468 7472 23520
rect 7524 23508 7530 23520
rect 7650 23508 7656 23520
rect 7524 23480 7656 23508
rect 7524 23468 7530 23480
rect 7650 23468 7656 23480
rect 7708 23468 7714 23520
rect 7834 23468 7840 23520
rect 7892 23468 7898 23520
rect 9490 23468 9496 23520
rect 9548 23508 9554 23520
rect 10244 23508 10272 23616
rect 10962 23604 10968 23656
rect 11020 23644 11026 23656
rect 15289 23647 15347 23653
rect 15289 23644 15301 23647
rect 11020 23616 15301 23644
rect 11020 23604 11026 23616
rect 15289 23613 15301 23616
rect 15335 23613 15347 23647
rect 15289 23607 15347 23613
rect 18598 23604 18604 23656
rect 18656 23644 18662 23656
rect 22646 23644 22652 23656
rect 18656 23616 22652 23644
rect 18656 23604 18662 23616
rect 22646 23604 22652 23616
rect 22704 23604 22710 23656
rect 22925 23647 22983 23653
rect 22925 23613 22937 23647
rect 22971 23613 22983 23647
rect 22925 23607 22983 23613
rect 13078 23536 13084 23588
rect 13136 23576 13142 23588
rect 13630 23576 13636 23588
rect 13136 23548 13636 23576
rect 13136 23536 13142 23548
rect 13630 23536 13636 23548
rect 13688 23536 13694 23588
rect 14550 23536 14556 23588
rect 14608 23576 14614 23588
rect 22278 23576 22284 23588
rect 14608 23548 22284 23576
rect 14608 23536 14614 23548
rect 22278 23536 22284 23548
rect 22336 23536 22342 23588
rect 22940 23520 22968 23607
rect 23566 23604 23572 23656
rect 23624 23644 23630 23656
rect 25792 23644 25820 23675
rect 25866 23672 25872 23724
rect 25924 23712 25930 23724
rect 26068 23721 26096 23752
rect 26142 23740 26148 23792
rect 26200 23780 26206 23792
rect 26329 23783 26387 23789
rect 26329 23780 26341 23783
rect 26200 23752 26341 23780
rect 26200 23740 26206 23752
rect 26329 23749 26341 23752
rect 26375 23749 26387 23783
rect 26329 23743 26387 23749
rect 26513 23783 26571 23789
rect 26513 23749 26525 23783
rect 26559 23780 26571 23783
rect 26559 23752 26648 23780
rect 26559 23749 26571 23752
rect 26513 23743 26571 23749
rect 25961 23715 26019 23721
rect 25961 23712 25973 23715
rect 25924 23684 25973 23712
rect 25924 23672 25930 23684
rect 25961 23681 25973 23684
rect 26007 23681 26019 23715
rect 25961 23675 26019 23681
rect 26053 23715 26111 23721
rect 26053 23681 26065 23715
rect 26099 23681 26111 23715
rect 26620 23712 26648 23752
rect 27522 23740 27528 23792
rect 27580 23780 27586 23792
rect 29564 23780 29592 23808
rect 31956 23780 31984 23820
rect 32306 23808 32312 23820
rect 32364 23848 32370 23860
rect 32769 23851 32827 23857
rect 32769 23848 32781 23851
rect 32364 23820 32781 23848
rect 32364 23808 32370 23820
rect 32769 23817 32781 23820
rect 32815 23817 32827 23851
rect 32769 23811 32827 23817
rect 33318 23808 33324 23860
rect 33376 23848 33382 23860
rect 34977 23851 35035 23857
rect 33376 23820 34560 23848
rect 33376 23808 33382 23820
rect 33226 23780 33232 23792
rect 27580 23752 29500 23780
rect 29564 23752 31984 23780
rect 32232 23752 33232 23780
rect 27580 23740 27586 23752
rect 26694 23712 26700 23724
rect 26620 23684 26700 23712
rect 26053 23675 26111 23681
rect 26694 23672 26700 23684
rect 26752 23672 26758 23724
rect 26970 23672 26976 23724
rect 27028 23712 27034 23724
rect 27249 23715 27307 23721
rect 27028 23684 27108 23712
rect 27028 23672 27034 23684
rect 26418 23644 26424 23656
rect 23624 23616 25544 23644
rect 25792 23616 26424 23644
rect 23624 23604 23630 23616
rect 23201 23579 23259 23585
rect 23201 23545 23213 23579
rect 23247 23576 23259 23579
rect 23750 23576 23756 23588
rect 23247 23548 23756 23576
rect 23247 23545 23259 23548
rect 23201 23539 23259 23545
rect 23750 23536 23756 23548
rect 23808 23536 23814 23588
rect 25222 23536 25228 23588
rect 25280 23536 25286 23588
rect 9548 23480 10272 23508
rect 9548 23468 9554 23480
rect 15194 23468 15200 23520
rect 15252 23468 15258 23520
rect 20162 23468 20168 23520
rect 20220 23508 20226 23520
rect 22094 23508 22100 23520
rect 20220 23480 22100 23508
rect 20220 23468 20226 23480
rect 22094 23468 22100 23480
rect 22152 23508 22158 23520
rect 22833 23511 22891 23517
rect 22833 23508 22845 23511
rect 22152 23480 22845 23508
rect 22152 23468 22158 23480
rect 22833 23477 22845 23480
rect 22879 23477 22891 23511
rect 22833 23471 22891 23477
rect 22922 23468 22928 23520
rect 22980 23468 22986 23520
rect 23661 23511 23719 23517
rect 23661 23477 23673 23511
rect 23707 23508 23719 23511
rect 24394 23508 24400 23520
rect 23707 23480 24400 23508
rect 23707 23477 23719 23480
rect 23661 23471 23719 23477
rect 24394 23468 24400 23480
rect 24452 23468 24458 23520
rect 25516 23508 25544 23616
rect 26418 23604 26424 23616
rect 26476 23604 26482 23656
rect 26602 23604 26608 23656
rect 26660 23644 26666 23656
rect 26878 23644 26884 23656
rect 26660 23616 26884 23644
rect 26660 23604 26666 23616
rect 26878 23604 26884 23616
rect 26936 23604 26942 23656
rect 27080 23644 27108 23684
rect 27249 23681 27261 23715
rect 27295 23712 27307 23715
rect 27295 23684 27329 23712
rect 27295 23681 27307 23684
rect 27249 23675 27307 23681
rect 27264 23644 27292 23675
rect 27430 23672 27436 23724
rect 27488 23672 27494 23724
rect 27798 23672 27804 23724
rect 27856 23712 27862 23724
rect 27985 23715 28043 23721
rect 27985 23712 27997 23715
rect 27856 23684 27997 23712
rect 27856 23672 27862 23684
rect 27985 23681 27997 23684
rect 28031 23712 28043 23715
rect 28810 23712 28816 23724
rect 28031 23684 28816 23712
rect 28031 23681 28043 23684
rect 27985 23675 28043 23681
rect 28810 23672 28816 23684
rect 28868 23672 28874 23724
rect 28077 23647 28135 23653
rect 28077 23644 28089 23647
rect 27080 23616 28089 23644
rect 28077 23613 28089 23616
rect 28123 23613 28135 23647
rect 29472 23644 29500 23752
rect 29546 23672 29552 23724
rect 29604 23712 29610 23724
rect 29733 23715 29791 23721
rect 29733 23712 29745 23715
rect 29604 23684 29745 23712
rect 29604 23672 29610 23684
rect 29733 23681 29745 23684
rect 29779 23681 29791 23715
rect 29733 23675 29791 23681
rect 29914 23672 29920 23724
rect 29972 23712 29978 23724
rect 30009 23715 30067 23721
rect 30009 23712 30021 23715
rect 29972 23684 30021 23712
rect 29972 23672 29978 23684
rect 30009 23681 30021 23684
rect 30055 23712 30067 23715
rect 30282 23712 30288 23724
rect 30055 23684 30288 23712
rect 30055 23681 30067 23684
rect 30009 23675 30067 23681
rect 30282 23672 30288 23684
rect 30340 23672 30346 23724
rect 30742 23672 30748 23724
rect 30800 23712 30806 23724
rect 30837 23715 30895 23721
rect 30837 23712 30849 23715
rect 30800 23684 30849 23712
rect 30800 23672 30806 23684
rect 30837 23681 30849 23684
rect 30883 23681 30895 23715
rect 30837 23675 30895 23681
rect 31478 23672 31484 23724
rect 31536 23672 31542 23724
rect 31757 23715 31815 23721
rect 31757 23681 31769 23715
rect 31803 23712 31815 23715
rect 32232 23712 32260 23752
rect 33226 23740 33232 23752
rect 33284 23740 33290 23792
rect 34422 23740 34428 23792
rect 34480 23740 34486 23792
rect 34532 23780 34560 23820
rect 34977 23817 34989 23851
rect 35023 23848 35035 23851
rect 41598 23848 41604 23860
rect 35023 23820 41604 23848
rect 35023 23817 35035 23820
rect 34977 23811 35035 23817
rect 41598 23808 41604 23820
rect 41656 23808 41662 23860
rect 41782 23808 41788 23860
rect 41840 23808 41846 23860
rect 43162 23808 43168 23860
rect 43220 23808 43226 23860
rect 34532 23752 34928 23780
rect 31803 23684 32260 23712
rect 32309 23715 32367 23721
rect 31803 23681 31815 23684
rect 31757 23675 31815 23681
rect 32309 23681 32321 23715
rect 32355 23681 32367 23715
rect 32309 23675 32367 23681
rect 29825 23647 29883 23653
rect 29825 23644 29837 23647
rect 29472 23616 29837 23644
rect 28077 23607 28135 23613
rect 29825 23613 29837 23616
rect 29871 23613 29883 23647
rect 29825 23607 29883 23613
rect 30929 23647 30987 23653
rect 30929 23613 30941 23647
rect 30975 23613 30987 23647
rect 30929 23607 30987 23613
rect 31573 23647 31631 23653
rect 31573 23613 31585 23647
rect 31619 23613 31631 23647
rect 31573 23607 31631 23613
rect 26510 23536 26516 23588
rect 26568 23576 26574 23588
rect 26697 23579 26755 23585
rect 26697 23576 26709 23579
rect 26568 23548 26709 23576
rect 26568 23536 26574 23548
rect 26697 23545 26709 23548
rect 26743 23576 26755 23579
rect 30944 23576 30972 23607
rect 26743 23548 30972 23576
rect 31205 23579 31263 23585
rect 26743 23545 26755 23548
rect 26697 23539 26755 23545
rect 31205 23545 31217 23579
rect 31251 23576 31263 23579
rect 31588 23576 31616 23607
rect 32214 23604 32220 23656
rect 32272 23644 32278 23656
rect 32324 23644 32352 23675
rect 32582 23672 32588 23724
rect 32640 23672 32646 23724
rect 34241 23715 34299 23721
rect 34241 23681 34253 23715
rect 34287 23712 34299 23715
rect 34330 23712 34336 23724
rect 34287 23684 34336 23712
rect 34287 23681 34299 23684
rect 34241 23675 34299 23681
rect 34330 23672 34336 23684
rect 34388 23672 34394 23724
rect 34514 23672 34520 23724
rect 34572 23672 34578 23724
rect 34606 23672 34612 23724
rect 34664 23712 34670 23724
rect 34701 23715 34759 23721
rect 34701 23712 34713 23715
rect 34664 23684 34713 23712
rect 34664 23672 34670 23684
rect 34701 23681 34713 23684
rect 34747 23681 34759 23715
rect 34701 23675 34759 23681
rect 34790 23672 34796 23724
rect 34848 23672 34854 23724
rect 34900 23712 34928 23752
rect 35986 23740 35992 23792
rect 36044 23780 36050 23792
rect 36044 23752 39712 23780
rect 36044 23740 36050 23752
rect 39684 23724 39712 23752
rect 40310 23740 40316 23792
rect 40368 23740 40374 23792
rect 41874 23740 41880 23792
rect 41932 23780 41938 23792
rect 41932 23752 43484 23780
rect 41932 23740 41938 23752
rect 36265 23715 36323 23721
rect 36265 23712 36277 23715
rect 34900 23684 36277 23712
rect 36265 23681 36277 23684
rect 36311 23712 36323 23715
rect 36449 23715 36507 23721
rect 36449 23712 36461 23715
rect 36311 23684 36461 23712
rect 36311 23681 36323 23684
rect 36265 23675 36323 23681
rect 36449 23681 36461 23684
rect 36495 23681 36507 23715
rect 36449 23675 36507 23681
rect 36722 23672 36728 23724
rect 36780 23672 36786 23724
rect 38930 23672 38936 23724
rect 38988 23712 38994 23724
rect 39117 23715 39175 23721
rect 39117 23712 39129 23715
rect 38988 23684 39129 23712
rect 38988 23672 38994 23684
rect 39117 23681 39129 23684
rect 39163 23681 39175 23715
rect 39117 23675 39175 23681
rect 39390 23672 39396 23724
rect 39448 23672 39454 23724
rect 39666 23672 39672 23724
rect 39724 23712 39730 23724
rect 43456 23721 43484 23752
rect 40497 23715 40555 23721
rect 40497 23712 40509 23715
rect 39724 23684 40509 23712
rect 39724 23672 39730 23684
rect 40497 23681 40509 23684
rect 40543 23681 40555 23715
rect 43349 23715 43407 23721
rect 43349 23712 43361 23715
rect 40497 23675 40555 23681
rect 41386 23684 43361 23712
rect 32272 23616 32352 23644
rect 32272 23604 32278 23616
rect 32398 23604 32404 23656
rect 32456 23604 32462 23656
rect 33594 23604 33600 23656
rect 33652 23644 33658 23656
rect 33962 23644 33968 23656
rect 33652 23616 33968 23644
rect 33652 23604 33658 23616
rect 33962 23604 33968 23616
rect 34020 23604 34026 23656
rect 34146 23604 34152 23656
rect 34204 23644 34210 23656
rect 36541 23647 36599 23653
rect 36541 23644 36553 23647
rect 34204 23616 36553 23644
rect 34204 23604 34210 23616
rect 36541 23613 36553 23616
rect 36587 23644 36599 23647
rect 37550 23644 37556 23656
rect 36587 23616 37556 23644
rect 36587 23613 36599 23616
rect 36541 23607 36599 23613
rect 37550 23604 37556 23616
rect 37608 23604 37614 23656
rect 39206 23604 39212 23656
rect 39264 23604 39270 23656
rect 41230 23604 41236 23656
rect 41288 23644 41294 23656
rect 41386 23644 41414 23684
rect 43349 23681 43361 23684
rect 43395 23681 43407 23715
rect 43349 23675 43407 23681
rect 43441 23715 43499 23721
rect 43441 23681 43453 23715
rect 43487 23681 43499 23715
rect 43441 23675 43499 23681
rect 43717 23715 43775 23721
rect 43717 23681 43729 23715
rect 43763 23712 43775 23715
rect 43806 23712 43812 23724
rect 43763 23684 43812 23712
rect 43763 23681 43775 23684
rect 43717 23675 43775 23681
rect 43806 23672 43812 23684
rect 43864 23672 43870 23724
rect 44269 23715 44327 23721
rect 44269 23681 44281 23715
rect 44315 23681 44327 23715
rect 44269 23675 44327 23681
rect 41288 23616 41414 23644
rect 41288 23604 41294 23616
rect 42978 23604 42984 23656
rect 43036 23604 43042 23656
rect 43622 23604 43628 23656
rect 43680 23604 43686 23656
rect 31251 23548 31616 23576
rect 31251 23545 31263 23548
rect 31205 23539 31263 23545
rect 31846 23536 31852 23588
rect 31904 23576 31910 23588
rect 39850 23576 39856 23588
rect 31904 23548 39856 23576
rect 31904 23536 31910 23548
rect 39850 23536 39856 23548
rect 39908 23536 39914 23588
rect 43530 23536 43536 23588
rect 43588 23576 43594 23588
rect 44284 23576 44312 23675
rect 43588 23548 44312 23576
rect 43588 23536 43594 23548
rect 25777 23511 25835 23517
rect 25777 23508 25789 23511
rect 25516 23480 25789 23508
rect 25777 23477 25789 23480
rect 25823 23477 25835 23511
rect 25777 23471 25835 23477
rect 27065 23511 27123 23517
rect 27065 23477 27077 23511
rect 27111 23508 27123 23511
rect 27154 23508 27160 23520
rect 27111 23480 27160 23508
rect 27111 23477 27123 23480
rect 27065 23471 27123 23477
rect 27154 23468 27160 23480
rect 27212 23468 27218 23520
rect 27430 23468 27436 23520
rect 27488 23508 27494 23520
rect 27617 23511 27675 23517
rect 27617 23508 27629 23511
rect 27488 23480 27629 23508
rect 27488 23468 27494 23480
rect 27617 23477 27629 23480
rect 27663 23508 27675 23511
rect 27893 23511 27951 23517
rect 27893 23508 27905 23511
rect 27663 23480 27905 23508
rect 27663 23477 27675 23480
rect 27617 23471 27675 23477
rect 27893 23477 27905 23480
rect 27939 23508 27951 23511
rect 28169 23511 28227 23517
rect 28169 23508 28181 23511
rect 27939 23480 28181 23508
rect 27939 23477 27951 23480
rect 27893 23471 27951 23477
rect 28169 23477 28181 23480
rect 28215 23508 28227 23511
rect 28258 23508 28264 23520
rect 28215 23480 28264 23508
rect 28215 23477 28227 23480
rect 28169 23471 28227 23477
rect 28258 23468 28264 23480
rect 28316 23468 28322 23520
rect 28353 23511 28411 23517
rect 28353 23477 28365 23511
rect 28399 23508 28411 23511
rect 29178 23508 29184 23520
rect 28399 23480 29184 23508
rect 28399 23477 28411 23480
rect 28353 23471 28411 23477
rect 29178 23468 29184 23480
rect 29236 23508 29242 23520
rect 29638 23508 29644 23520
rect 29236 23480 29644 23508
rect 29236 23468 29242 23480
rect 29638 23468 29644 23480
rect 29696 23468 29702 23520
rect 29822 23468 29828 23520
rect 29880 23468 29886 23520
rect 30926 23468 30932 23520
rect 30984 23468 30990 23520
rect 31570 23468 31576 23520
rect 31628 23468 31634 23520
rect 31938 23468 31944 23520
rect 31996 23468 32002 23520
rect 32585 23511 32643 23517
rect 32585 23477 32597 23511
rect 32631 23508 32643 23511
rect 33042 23508 33048 23520
rect 32631 23480 33048 23508
rect 32631 23477 32643 23480
rect 32585 23471 32643 23477
rect 33042 23468 33048 23480
rect 33100 23468 33106 23520
rect 33778 23468 33784 23520
rect 33836 23508 33842 23520
rect 34057 23511 34115 23517
rect 34057 23508 34069 23511
rect 33836 23480 34069 23508
rect 33836 23468 33842 23480
rect 34057 23477 34069 23480
rect 34103 23477 34115 23511
rect 34057 23471 34115 23477
rect 34514 23468 34520 23520
rect 34572 23468 34578 23520
rect 36446 23468 36452 23520
rect 36504 23468 36510 23520
rect 36722 23468 36728 23520
rect 36780 23508 36786 23520
rect 36909 23511 36967 23517
rect 36909 23508 36921 23511
rect 36780 23480 36921 23508
rect 36780 23468 36786 23480
rect 36909 23477 36921 23480
rect 36955 23477 36967 23511
rect 36909 23471 36967 23477
rect 39114 23468 39120 23520
rect 39172 23468 39178 23520
rect 39577 23511 39635 23517
rect 39577 23477 39589 23511
rect 39623 23508 39635 23511
rect 40678 23508 40684 23520
rect 39623 23480 40684 23508
rect 39623 23477 39635 23480
rect 39577 23471 39635 23477
rect 40678 23468 40684 23480
rect 40736 23468 40742 23520
rect 41690 23468 41696 23520
rect 41748 23508 41754 23520
rect 42429 23511 42487 23517
rect 42429 23508 42441 23511
rect 41748 23480 42441 23508
rect 41748 23468 41754 23480
rect 42429 23477 42441 23480
rect 42475 23477 42487 23511
rect 42429 23471 42487 23477
rect 44082 23468 44088 23520
rect 44140 23508 44146 23520
rect 44453 23511 44511 23517
rect 44453 23508 44465 23511
rect 44140 23480 44465 23508
rect 44140 23468 44146 23480
rect 44453 23477 44465 23480
rect 44499 23477 44511 23511
rect 44453 23471 44511 23477
rect 1104 23418 44896 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 44896 23418
rect 1104 23344 44896 23366
rect 3145 23307 3203 23313
rect 3145 23273 3157 23307
rect 3191 23304 3203 23307
rect 5442 23304 5448 23316
rect 3191 23276 5448 23304
rect 3191 23273 3203 23276
rect 3145 23267 3203 23273
rect 5442 23264 5448 23276
rect 5500 23264 5506 23316
rect 5721 23307 5779 23313
rect 5721 23273 5733 23307
rect 5767 23304 5779 23307
rect 6822 23304 6828 23316
rect 5767 23276 6828 23304
rect 5767 23273 5779 23276
rect 5721 23267 5779 23273
rect 6822 23264 6828 23276
rect 6880 23264 6886 23316
rect 10873 23307 10931 23313
rect 6932 23276 10824 23304
rect 3050 23236 3056 23248
rect 2700 23208 3056 23236
rect 2593 23103 2651 23109
rect 2593 23069 2605 23103
rect 2639 23100 2651 23103
rect 2700 23100 2728 23208
rect 3050 23196 3056 23208
rect 3108 23236 3114 23248
rect 3418 23236 3424 23248
rect 3108 23208 3424 23236
rect 3108 23196 3114 23208
rect 3418 23196 3424 23208
rect 3476 23196 3482 23248
rect 4614 23196 4620 23248
rect 4672 23196 4678 23248
rect 5077 23239 5135 23245
rect 5077 23205 5089 23239
rect 5123 23236 5135 23239
rect 5258 23236 5264 23248
rect 5123 23208 5264 23236
rect 5123 23205 5135 23208
rect 5077 23199 5135 23205
rect 5258 23196 5264 23208
rect 5316 23196 5322 23248
rect 5626 23196 5632 23248
rect 5684 23236 5690 23248
rect 6932 23236 6960 23276
rect 5684 23208 6960 23236
rect 5684 23196 5690 23208
rect 7558 23196 7564 23248
rect 7616 23236 7622 23248
rect 7837 23239 7895 23245
rect 7837 23236 7849 23239
rect 7616 23208 7849 23236
rect 7616 23196 7622 23208
rect 7837 23205 7849 23208
rect 7883 23205 7895 23239
rect 7837 23199 7895 23205
rect 8294 23196 8300 23248
rect 8352 23236 8358 23248
rect 9582 23236 9588 23248
rect 8352 23208 9588 23236
rect 8352 23196 8358 23208
rect 9582 23196 9588 23208
rect 9640 23236 9646 23248
rect 9640 23208 10732 23236
rect 9640 23196 9646 23208
rect 3786 23168 3792 23180
rect 2792 23140 3792 23168
rect 2792 23109 2820 23140
rect 3786 23128 3792 23140
rect 3844 23128 3850 23180
rect 4632 23168 4660 23196
rect 4448 23140 5580 23168
rect 2639 23072 2728 23100
rect 2777 23103 2835 23109
rect 2639 23069 2651 23072
rect 2593 23063 2651 23069
rect 2777 23069 2789 23103
rect 2823 23069 2835 23103
rect 2777 23063 2835 23069
rect 3013 23103 3071 23109
rect 3013 23069 3025 23103
rect 3059 23100 3071 23103
rect 4338 23100 4344 23112
rect 3059 23072 4344 23100
rect 3059 23069 3071 23072
rect 3013 23063 3071 23069
rect 4338 23060 4344 23072
rect 4396 23060 4402 23112
rect 4448 23109 4476 23140
rect 4433 23103 4491 23109
rect 4433 23069 4445 23103
rect 4479 23069 4491 23103
rect 4433 23063 4491 23069
rect 4617 23103 4675 23109
rect 4617 23069 4629 23103
rect 4663 23069 4675 23103
rect 4617 23063 4675 23069
rect 2130 22992 2136 23044
rect 2188 23032 2194 23044
rect 2869 23035 2927 23041
rect 2188 23004 2774 23032
rect 2188 22992 2194 23004
rect 2746 22964 2774 23004
rect 2869 23001 2881 23035
rect 2915 23001 2927 23035
rect 4632 23032 4660 23063
rect 4706 23060 4712 23112
rect 4764 23100 4770 23112
rect 4893 23103 4951 23109
rect 4893 23100 4905 23103
rect 4764 23072 4905 23100
rect 4764 23060 4770 23072
rect 4893 23069 4905 23072
rect 4939 23069 4951 23103
rect 4893 23063 4951 23069
rect 5169 23103 5227 23109
rect 5169 23069 5181 23103
rect 5215 23100 5227 23103
rect 5258 23100 5264 23112
rect 5215 23072 5264 23100
rect 5215 23069 5227 23072
rect 5169 23063 5227 23069
rect 5258 23060 5264 23072
rect 5316 23060 5322 23112
rect 5552 23109 5580 23140
rect 9214 23128 9220 23180
rect 9272 23168 9278 23180
rect 9272 23140 10640 23168
rect 9272 23128 9278 23140
rect 5537 23103 5595 23109
rect 5537 23069 5549 23103
rect 5583 23100 5595 23103
rect 6638 23100 6644 23112
rect 5583 23072 6644 23100
rect 5583 23069 5595 23072
rect 5537 23063 5595 23069
rect 6638 23060 6644 23072
rect 6696 23100 6702 23112
rect 7285 23103 7343 23109
rect 7285 23100 7297 23103
rect 6696 23072 7297 23100
rect 6696 23060 6702 23072
rect 7285 23069 7297 23072
rect 7331 23069 7343 23103
rect 7561 23103 7619 23109
rect 7561 23100 7573 23103
rect 7285 23063 7343 23069
rect 7392 23072 7573 23100
rect 4798 23032 4804 23044
rect 4632 23004 4804 23032
rect 2869 22995 2927 23001
rect 2884 22964 2912 22995
rect 4798 22992 4804 23004
rect 4856 23032 4862 23044
rect 5353 23035 5411 23041
rect 5353 23032 5365 23035
rect 4856 23004 5365 23032
rect 4856 22992 4862 23004
rect 5353 23001 5365 23004
rect 5399 23001 5411 23035
rect 5353 22995 5411 23001
rect 4062 22964 4068 22976
rect 2746 22936 4068 22964
rect 4062 22924 4068 22936
rect 4120 22924 4126 22976
rect 5368 22964 5396 22995
rect 5442 22992 5448 23044
rect 5500 22992 5506 23044
rect 6730 23032 6736 23044
rect 5552 23004 6736 23032
rect 5552 22964 5580 23004
rect 6730 22992 6736 23004
rect 6788 23032 6794 23044
rect 7392 23032 7420 23072
rect 7561 23069 7573 23072
rect 7607 23069 7619 23103
rect 7561 23063 7619 23069
rect 7705 23103 7763 23109
rect 7705 23069 7717 23103
rect 7751 23100 7763 23103
rect 8294 23100 8300 23112
rect 7751 23072 8300 23100
rect 7751 23069 7763 23072
rect 7705 23063 7763 23069
rect 8294 23060 8300 23072
rect 8352 23060 8358 23112
rect 9493 23103 9551 23109
rect 9493 23069 9505 23103
rect 9539 23069 9551 23103
rect 9493 23063 9551 23069
rect 9677 23103 9735 23109
rect 9677 23069 9689 23103
rect 9723 23100 9735 23103
rect 9858 23100 9864 23112
rect 9723 23072 9864 23100
rect 9723 23069 9735 23072
rect 9677 23063 9735 23069
rect 6788 23004 7420 23032
rect 7469 23035 7527 23041
rect 6788 22992 6794 23004
rect 7469 23001 7481 23035
rect 7515 23032 7527 23035
rect 9398 23032 9404 23044
rect 7515 23004 9404 23032
rect 7515 23001 7527 23004
rect 7469 22995 7527 23001
rect 9398 22992 9404 23004
rect 9456 22992 9462 23044
rect 9508 23032 9536 23063
rect 9858 23060 9864 23072
rect 9916 23060 9922 23112
rect 10045 23103 10103 23109
rect 10045 23069 10057 23103
rect 10091 23100 10103 23103
rect 10226 23100 10232 23112
rect 10091 23072 10232 23100
rect 10091 23069 10103 23072
rect 10045 23063 10103 23069
rect 10226 23060 10232 23072
rect 10284 23060 10290 23112
rect 10321 23103 10379 23109
rect 10321 23069 10333 23103
rect 10367 23100 10379 23103
rect 10410 23100 10416 23112
rect 10367 23072 10416 23100
rect 10367 23069 10379 23072
rect 10321 23063 10379 23069
rect 10410 23060 10416 23072
rect 10468 23060 10474 23112
rect 10612 23109 10640 23140
rect 10704 23109 10732 23208
rect 10597 23103 10655 23109
rect 10597 23069 10609 23103
rect 10643 23069 10655 23103
rect 10597 23063 10655 23069
rect 10694 23103 10752 23109
rect 10694 23069 10706 23103
rect 10740 23069 10752 23103
rect 10694 23063 10752 23069
rect 9766 23032 9772 23044
rect 9508 23004 9772 23032
rect 9766 22992 9772 23004
rect 9824 22992 9830 23044
rect 10505 23035 10563 23041
rect 9876 23004 10180 23032
rect 5368 22936 5580 22964
rect 9416 22964 9444 22992
rect 9876 22964 9904 23004
rect 9416 22936 9904 22964
rect 9953 22967 10011 22973
rect 9953 22933 9965 22967
rect 9999 22964 10011 22967
rect 10042 22964 10048 22976
rect 9999 22936 10048 22964
rect 9999 22933 10011 22936
rect 9953 22927 10011 22933
rect 10042 22924 10048 22936
rect 10100 22924 10106 22976
rect 10152 22964 10180 23004
rect 10505 23001 10517 23035
rect 10551 23001 10563 23035
rect 10796 23032 10824 23276
rect 10873 23273 10885 23307
rect 10919 23304 10931 23307
rect 11238 23304 11244 23316
rect 10919 23276 11244 23304
rect 10919 23273 10931 23276
rect 10873 23267 10931 23273
rect 11238 23264 11244 23276
rect 11296 23264 11302 23316
rect 12710 23264 12716 23316
rect 12768 23304 12774 23316
rect 12805 23307 12863 23313
rect 12805 23304 12817 23307
rect 12768 23276 12817 23304
rect 12768 23264 12774 23276
rect 12805 23273 12817 23276
rect 12851 23273 12863 23307
rect 12805 23267 12863 23273
rect 12894 23264 12900 23316
rect 12952 23304 12958 23316
rect 12952 23276 14412 23304
rect 12952 23264 12958 23276
rect 11698 23196 11704 23248
rect 11756 23236 11762 23248
rect 11756 23208 14320 23236
rect 11756 23196 11762 23208
rect 12268 23140 14228 23168
rect 12268 23112 12296 23140
rect 11238 23060 11244 23112
rect 11296 23100 11302 23112
rect 12066 23100 12072 23112
rect 11296 23072 12072 23100
rect 11296 23060 11302 23072
rect 12066 23060 12072 23072
rect 12124 23060 12130 23112
rect 12250 23060 12256 23112
rect 12308 23060 12314 23112
rect 12618 23060 12624 23112
rect 12676 23060 12682 23112
rect 14093 23103 14151 23109
rect 14093 23069 14105 23103
rect 14139 23069 14151 23103
rect 14093 23063 14151 23069
rect 12437 23035 12495 23041
rect 12437 23032 12449 23035
rect 10796 23004 12449 23032
rect 10505 22995 10563 23001
rect 12437 23001 12449 23004
rect 12483 23001 12495 23035
rect 12437 22995 12495 23001
rect 12529 23035 12587 23041
rect 12529 23001 12541 23035
rect 12575 23032 12587 23035
rect 13078 23032 13084 23044
rect 12575 23004 13084 23032
rect 12575 23001 12587 23004
rect 12529 22995 12587 23001
rect 10520 22964 10548 22995
rect 13078 22992 13084 23004
rect 13136 23032 13142 23044
rect 14108 23032 14136 23063
rect 13136 23004 14136 23032
rect 14200 23032 14228 23140
rect 14292 23109 14320 23208
rect 14384 23168 14412 23276
rect 14642 23264 14648 23316
rect 14700 23264 14706 23316
rect 15013 23307 15071 23313
rect 15013 23273 15025 23307
rect 15059 23304 15071 23307
rect 15102 23304 15108 23316
rect 15059 23276 15108 23304
rect 15059 23273 15071 23276
rect 15013 23267 15071 23273
rect 15028 23236 15056 23267
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 15194 23264 15200 23316
rect 15252 23264 15258 23316
rect 18601 23307 18659 23313
rect 18601 23273 18613 23307
rect 18647 23304 18659 23307
rect 18874 23304 18880 23316
rect 18647 23276 18880 23304
rect 18647 23273 18659 23276
rect 18601 23267 18659 23273
rect 18874 23264 18880 23276
rect 18932 23304 18938 23316
rect 18932 23276 22324 23304
rect 18932 23264 18938 23276
rect 18785 23239 18843 23245
rect 15028 23208 18552 23236
rect 18524 23168 18552 23208
rect 18785 23205 18797 23239
rect 18831 23236 18843 23239
rect 22186 23236 22192 23248
rect 18831 23208 22192 23236
rect 18831 23205 18843 23208
rect 18785 23199 18843 23205
rect 22186 23196 22192 23208
rect 22244 23196 22250 23248
rect 22296 23236 22324 23276
rect 22646 23264 22652 23316
rect 22704 23304 22710 23316
rect 23569 23307 23627 23313
rect 23569 23304 23581 23307
rect 22704 23276 23581 23304
rect 22704 23264 22710 23276
rect 23569 23273 23581 23276
rect 23615 23273 23627 23307
rect 23569 23267 23627 23273
rect 23750 23264 23756 23316
rect 23808 23304 23814 23316
rect 23937 23307 23995 23313
rect 23937 23304 23949 23307
rect 23808 23276 23949 23304
rect 23808 23264 23814 23276
rect 23937 23273 23949 23276
rect 23983 23304 23995 23307
rect 25130 23304 25136 23316
rect 23983 23276 25136 23304
rect 23983 23273 23995 23276
rect 23937 23267 23995 23273
rect 25130 23264 25136 23276
rect 25188 23264 25194 23316
rect 26510 23304 26516 23316
rect 25332 23276 26516 23304
rect 25222 23236 25228 23248
rect 22296 23208 25228 23236
rect 25222 23196 25228 23208
rect 25280 23196 25286 23248
rect 19334 23168 19340 23180
rect 14384 23140 17954 23168
rect 18524 23140 19340 23168
rect 14277 23103 14335 23109
rect 14277 23069 14289 23103
rect 14323 23069 14335 23103
rect 14277 23063 14335 23069
rect 14466 23103 14524 23109
rect 14466 23069 14478 23103
rect 14512 23069 14524 23103
rect 14466 23063 14524 23069
rect 14369 23035 14427 23041
rect 14369 23032 14381 23035
rect 14200 23004 14381 23032
rect 13136 22992 13142 23004
rect 14369 23001 14381 23004
rect 14415 23001 14427 23035
rect 14369 22995 14427 23001
rect 10152 22936 10548 22964
rect 11974 22924 11980 22976
rect 12032 22964 12038 22976
rect 12618 22964 12624 22976
rect 12032 22936 12624 22964
rect 12032 22924 12038 22936
rect 12618 22924 12624 22936
rect 12676 22964 12682 22976
rect 12986 22964 12992 22976
rect 12676 22936 12992 22964
rect 12676 22924 12682 22936
rect 12986 22924 12992 22936
rect 13044 22964 13050 22976
rect 14481 22964 14509 23063
rect 14826 23060 14832 23112
rect 14884 23060 14890 23112
rect 15013 23103 15071 23109
rect 15013 23069 15025 23103
rect 15059 23100 15071 23103
rect 15194 23100 15200 23112
rect 15059 23072 15200 23100
rect 15059 23069 15071 23072
rect 15013 23063 15071 23069
rect 15194 23060 15200 23072
rect 15252 23100 15258 23112
rect 16206 23100 16212 23112
rect 15252 23072 16212 23100
rect 15252 23060 15258 23072
rect 16206 23060 16212 23072
rect 16264 23060 16270 23112
rect 17926 23100 17954 23140
rect 19334 23128 19340 23140
rect 19392 23128 19398 23180
rect 20346 23128 20352 23180
rect 20404 23168 20410 23180
rect 20441 23171 20499 23177
rect 20441 23168 20453 23171
rect 20404 23140 20453 23168
rect 20404 23128 20410 23140
rect 20441 23137 20453 23140
rect 20487 23137 20499 23171
rect 20441 23131 20499 23137
rect 20548 23140 20852 23168
rect 18417 23103 18475 23109
rect 18417 23100 18429 23103
rect 17926 23072 18429 23100
rect 18417 23069 18429 23072
rect 18463 23069 18475 23103
rect 18417 23063 18475 23069
rect 18432 23032 18460 23063
rect 18506 23060 18512 23112
rect 18564 23060 18570 23112
rect 20073 23103 20131 23109
rect 20073 23069 20085 23103
rect 20119 23100 20131 23103
rect 20548 23100 20576 23140
rect 20119 23072 20576 23100
rect 20119 23069 20131 23072
rect 20073 23063 20131 23069
rect 20088 23032 20116 23063
rect 20622 23060 20628 23112
rect 20680 23100 20686 23112
rect 20717 23103 20775 23109
rect 20717 23100 20729 23103
rect 20680 23072 20729 23100
rect 20680 23060 20686 23072
rect 20717 23069 20729 23072
rect 20763 23069 20775 23103
rect 20717 23063 20775 23069
rect 18432 23004 20116 23032
rect 20257 23035 20315 23041
rect 20257 23001 20269 23035
rect 20303 23001 20315 23035
rect 20257 22995 20315 23001
rect 13044 22936 14509 22964
rect 13044 22924 13050 22936
rect 19242 22924 19248 22976
rect 19300 22964 19306 22976
rect 20272 22964 20300 22995
rect 20530 22992 20536 23044
rect 20588 22992 20594 23044
rect 20824 23032 20852 23140
rect 23382 23128 23388 23180
rect 23440 23168 23446 23180
rect 24854 23168 24860 23180
rect 23440 23140 24860 23168
rect 23440 23128 23446 23140
rect 24854 23128 24860 23140
rect 24912 23128 24918 23180
rect 24946 23128 24952 23180
rect 25004 23168 25010 23180
rect 25332 23168 25360 23276
rect 26510 23264 26516 23276
rect 26568 23264 26574 23316
rect 26878 23264 26884 23316
rect 26936 23304 26942 23316
rect 27062 23304 27068 23316
rect 26936 23276 27068 23304
rect 26936 23264 26942 23276
rect 27062 23264 27068 23276
rect 27120 23304 27126 23316
rect 27522 23304 27528 23316
rect 27120 23276 27528 23304
rect 27120 23264 27126 23276
rect 27522 23264 27528 23276
rect 27580 23264 27586 23316
rect 27890 23264 27896 23316
rect 27948 23304 27954 23316
rect 29733 23307 29791 23313
rect 29733 23304 29745 23307
rect 27948 23276 29745 23304
rect 27948 23264 27954 23276
rect 29733 23273 29745 23276
rect 29779 23273 29791 23307
rect 29733 23267 29791 23273
rect 31018 23264 31024 23316
rect 31076 23304 31082 23316
rect 32858 23304 32864 23316
rect 31076 23276 32864 23304
rect 31076 23264 31082 23276
rect 32858 23264 32864 23276
rect 32916 23264 32922 23316
rect 33594 23264 33600 23316
rect 33652 23304 33658 23316
rect 33689 23307 33747 23313
rect 33689 23304 33701 23307
rect 33652 23276 33701 23304
rect 33652 23264 33658 23276
rect 33689 23273 33701 23276
rect 33735 23273 33747 23307
rect 33689 23267 33747 23273
rect 34149 23307 34207 23313
rect 34149 23273 34161 23307
rect 34195 23304 34207 23307
rect 34514 23304 34520 23316
rect 34195 23276 34520 23304
rect 34195 23273 34207 23276
rect 34149 23267 34207 23273
rect 34514 23264 34520 23276
rect 34572 23264 34578 23316
rect 34606 23264 34612 23316
rect 34664 23304 34670 23316
rect 34701 23307 34759 23313
rect 34701 23304 34713 23307
rect 34664 23276 34713 23304
rect 34664 23264 34670 23276
rect 34701 23273 34713 23276
rect 34747 23273 34759 23307
rect 34701 23267 34759 23273
rect 37090 23264 37096 23316
rect 37148 23264 37154 23316
rect 37274 23264 37280 23316
rect 37332 23304 37338 23316
rect 37369 23307 37427 23313
rect 37369 23304 37381 23307
rect 37332 23276 37381 23304
rect 37332 23264 37338 23276
rect 37369 23273 37381 23276
rect 37415 23273 37427 23307
rect 37369 23267 37427 23273
rect 37458 23264 37464 23316
rect 37516 23304 37522 23316
rect 38010 23304 38016 23316
rect 37516 23276 38016 23304
rect 37516 23264 37522 23276
rect 38010 23264 38016 23276
rect 38068 23264 38074 23316
rect 38102 23264 38108 23316
rect 38160 23304 38166 23316
rect 38197 23307 38255 23313
rect 38197 23304 38209 23307
rect 38160 23276 38209 23304
rect 38160 23264 38166 23276
rect 38197 23273 38209 23276
rect 38243 23273 38255 23307
rect 38197 23267 38255 23273
rect 38657 23307 38715 23313
rect 38657 23273 38669 23307
rect 38703 23304 38715 23307
rect 39206 23304 39212 23316
rect 38703 23276 39212 23304
rect 38703 23273 38715 23276
rect 38657 23267 38715 23273
rect 39206 23264 39212 23276
rect 39264 23264 39270 23316
rect 39758 23264 39764 23316
rect 39816 23304 39822 23316
rect 39853 23307 39911 23313
rect 39853 23304 39865 23307
rect 39816 23276 39865 23304
rect 39816 23264 39822 23276
rect 39853 23273 39865 23276
rect 39899 23273 39911 23307
rect 39853 23267 39911 23273
rect 39942 23264 39948 23316
rect 40000 23304 40006 23316
rect 40000 23276 41368 23304
rect 40000 23264 40006 23276
rect 25958 23196 25964 23248
rect 26016 23236 26022 23248
rect 26602 23236 26608 23248
rect 26016 23208 26608 23236
rect 26016 23196 26022 23208
rect 26602 23196 26608 23208
rect 26660 23196 26666 23248
rect 26786 23196 26792 23248
rect 26844 23236 26850 23248
rect 27341 23239 27399 23245
rect 27341 23236 27353 23239
rect 26844 23208 27353 23236
rect 26844 23196 26850 23208
rect 27341 23205 27353 23208
rect 27387 23205 27399 23239
rect 27341 23199 27399 23205
rect 28994 23196 29000 23248
rect 29052 23236 29058 23248
rect 29052 23208 29408 23236
rect 29052 23196 29058 23208
rect 29086 23168 29092 23180
rect 25004 23140 25360 23168
rect 26252 23140 29092 23168
rect 25004 23128 25010 23140
rect 20990 23060 20996 23112
rect 21048 23100 21054 23112
rect 23474 23100 23480 23112
rect 21048 23072 23480 23100
rect 21048 23060 21054 23072
rect 23474 23060 23480 23072
rect 23532 23100 23538 23112
rect 23569 23103 23627 23109
rect 23569 23100 23581 23103
rect 23532 23072 23581 23100
rect 23532 23060 23538 23072
rect 23569 23069 23581 23072
rect 23615 23069 23627 23103
rect 23569 23063 23627 23069
rect 23658 23060 23664 23112
rect 23716 23100 23722 23112
rect 26252 23100 26280 23140
rect 29086 23128 29092 23140
rect 29144 23168 29150 23180
rect 29270 23168 29276 23180
rect 29144 23140 29276 23168
rect 29144 23128 29150 23140
rect 29270 23128 29276 23140
rect 29328 23128 29334 23180
rect 29380 23168 29408 23208
rect 29546 23196 29552 23248
rect 29604 23196 29610 23248
rect 29638 23196 29644 23248
rect 29696 23236 29702 23248
rect 29822 23236 29828 23248
rect 29696 23208 29828 23236
rect 29696 23196 29702 23208
rect 29822 23196 29828 23208
rect 29880 23196 29886 23248
rect 31202 23196 31208 23248
rect 31260 23236 31266 23248
rect 32582 23236 32588 23248
rect 31260 23208 32588 23236
rect 31260 23196 31266 23208
rect 32582 23196 32588 23208
rect 32640 23236 32646 23248
rect 34882 23236 34888 23248
rect 32640 23208 34888 23236
rect 32640 23196 32646 23208
rect 34882 23196 34888 23208
rect 34940 23196 34946 23248
rect 35161 23239 35219 23245
rect 35161 23205 35173 23239
rect 35207 23236 35219 23239
rect 39390 23236 39396 23248
rect 35207 23208 39396 23236
rect 35207 23205 35219 23208
rect 35161 23199 35219 23205
rect 39390 23196 39396 23208
rect 39448 23196 39454 23248
rect 40221 23239 40279 23245
rect 40221 23205 40233 23239
rect 40267 23236 40279 23239
rect 40589 23239 40647 23245
rect 40589 23236 40601 23239
rect 40267 23208 40601 23236
rect 40267 23205 40279 23208
rect 40221 23199 40279 23205
rect 40589 23205 40601 23208
rect 40635 23205 40647 23239
rect 40589 23199 40647 23205
rect 41046 23196 41052 23248
rect 41104 23196 41110 23248
rect 41340 23245 41368 23276
rect 41325 23239 41383 23245
rect 41325 23205 41337 23239
rect 41371 23205 41383 23239
rect 41325 23199 41383 23205
rect 29917 23171 29975 23177
rect 29917 23168 29929 23171
rect 29380 23140 29929 23168
rect 29917 23137 29929 23140
rect 29963 23168 29975 23171
rect 29963 23140 31248 23168
rect 29963 23137 29975 23140
rect 29917 23131 29975 23137
rect 31220 23112 31248 23140
rect 32766 23128 32772 23180
rect 32824 23168 32830 23180
rect 33781 23171 33839 23177
rect 33781 23168 33793 23171
rect 32824 23140 33793 23168
rect 32824 23128 32830 23140
rect 33781 23137 33793 23140
rect 33827 23137 33839 23171
rect 33781 23131 33839 23137
rect 34146 23128 34152 23180
rect 34204 23168 34210 23180
rect 34793 23171 34851 23177
rect 34793 23168 34805 23171
rect 34204 23140 34805 23168
rect 34204 23128 34210 23140
rect 34793 23137 34805 23140
rect 34839 23168 34851 23171
rect 35434 23168 35440 23180
rect 34839 23140 35440 23168
rect 34839 23137 34851 23140
rect 34793 23131 34851 23137
rect 35434 23128 35440 23140
rect 35492 23128 35498 23180
rect 37550 23168 37556 23180
rect 37384 23140 37556 23168
rect 23716 23072 26280 23100
rect 26421 23103 26479 23109
rect 23716 23060 23722 23072
rect 26421 23069 26433 23103
rect 26467 23100 26479 23103
rect 26878 23100 26884 23112
rect 26467 23072 26884 23100
rect 26467 23069 26479 23072
rect 26421 23063 26479 23069
rect 26878 23060 26884 23072
rect 26936 23060 26942 23112
rect 27154 23060 27160 23112
rect 27212 23100 27218 23112
rect 29733 23103 29791 23109
rect 29733 23100 29745 23103
rect 27212 23072 29745 23100
rect 27212 23060 27218 23072
rect 29733 23069 29745 23072
rect 29779 23069 29791 23103
rect 29733 23063 29791 23069
rect 31202 23060 31208 23112
rect 31260 23060 31266 23112
rect 32585 23103 32643 23109
rect 32585 23069 32597 23103
rect 32631 23100 32643 23103
rect 33226 23100 33232 23112
rect 32631 23072 33232 23100
rect 32631 23069 32643 23072
rect 32585 23063 32643 23069
rect 33226 23060 33232 23072
rect 33284 23060 33290 23112
rect 33502 23060 33508 23112
rect 33560 23100 33566 23112
rect 33689 23103 33747 23109
rect 33689 23100 33701 23103
rect 33560 23072 33701 23100
rect 33560 23060 33566 23072
rect 33689 23069 33701 23072
rect 33735 23069 33747 23103
rect 33689 23063 33747 23069
rect 33962 23060 33968 23112
rect 34020 23060 34026 23112
rect 34882 23060 34888 23112
rect 34940 23100 34946 23112
rect 34977 23103 35035 23109
rect 34977 23100 34989 23103
rect 34940 23072 34989 23100
rect 34940 23060 34946 23072
rect 34977 23069 34989 23072
rect 35023 23100 35035 23103
rect 35618 23100 35624 23112
rect 35023 23072 35624 23100
rect 35023 23069 35035 23072
rect 34977 23063 35035 23069
rect 35618 23060 35624 23072
rect 35676 23060 35682 23112
rect 36170 23060 36176 23112
rect 36228 23100 36234 23112
rect 36906 23100 36912 23112
rect 36228 23072 36912 23100
rect 36228 23060 36234 23072
rect 36906 23060 36912 23072
rect 36964 23100 36970 23112
rect 37001 23103 37059 23109
rect 37001 23100 37013 23103
rect 36964 23072 37013 23100
rect 36964 23060 36970 23072
rect 37001 23069 37013 23072
rect 37047 23069 37059 23103
rect 37001 23063 37059 23069
rect 37182 23060 37188 23112
rect 37240 23060 37246 23112
rect 37384 23109 37412 23140
rect 37550 23128 37556 23140
rect 37608 23128 37614 23180
rect 39945 23171 40003 23177
rect 39945 23168 39957 23171
rect 38672 23140 39957 23168
rect 37369 23103 37427 23109
rect 37369 23069 37381 23103
rect 37415 23069 37427 23103
rect 37369 23063 37427 23069
rect 37458 23060 37464 23112
rect 37516 23060 37522 23112
rect 38381 23103 38439 23109
rect 38381 23100 38393 23103
rect 37568 23072 38393 23100
rect 26050 23032 26056 23044
rect 20824 23004 26056 23032
rect 26050 22992 26056 23004
rect 26108 22992 26114 23044
rect 26142 22992 26148 23044
rect 26200 23032 26206 23044
rect 26237 23035 26295 23041
rect 26237 23032 26249 23035
rect 26200 23004 26249 23032
rect 26200 22992 26206 23004
rect 26237 23001 26249 23004
rect 26283 23001 26295 23035
rect 26237 22995 26295 23001
rect 26510 22992 26516 23044
rect 26568 23032 26574 23044
rect 27525 23035 27583 23041
rect 27525 23032 27537 23035
rect 26568 23004 27537 23032
rect 26568 22992 26574 23004
rect 27525 23001 27537 23004
rect 27571 23001 27583 23035
rect 27525 22995 27583 23001
rect 27709 23035 27767 23041
rect 27709 23001 27721 23035
rect 27755 23032 27767 23035
rect 27798 23032 27804 23044
rect 27755 23004 27804 23032
rect 27755 23001 27767 23004
rect 27709 22995 27767 23001
rect 27798 22992 27804 23004
rect 27856 22992 27862 23044
rect 28074 22992 28080 23044
rect 28132 23032 28138 23044
rect 28132 23004 28488 23032
rect 28132 22992 28138 23004
rect 20806 22964 20812 22976
rect 19300 22936 20812 22964
rect 19300 22924 19306 22936
rect 20806 22924 20812 22936
rect 20864 22924 20870 22976
rect 20901 22967 20959 22973
rect 20901 22933 20913 22967
rect 20947 22964 20959 22967
rect 23474 22964 23480 22976
rect 20947 22936 23480 22964
rect 20947 22933 20959 22936
rect 20901 22927 20959 22933
rect 23474 22924 23480 22936
rect 23532 22924 23538 22976
rect 23658 22924 23664 22976
rect 23716 22964 23722 22976
rect 23842 22964 23848 22976
rect 23716 22936 23848 22964
rect 23716 22924 23722 22936
rect 23842 22924 23848 22936
rect 23900 22964 23906 22976
rect 26878 22964 26884 22976
rect 23900 22936 26884 22964
rect 23900 22924 23906 22936
rect 26878 22924 26884 22936
rect 26936 22924 26942 22976
rect 28460 22964 28488 23004
rect 28994 22992 29000 23044
rect 29052 23032 29058 23044
rect 30009 23035 30067 23041
rect 30009 23032 30021 23035
rect 29052 23004 30021 23032
rect 29052 22992 29058 23004
rect 30009 23001 30021 23004
rect 30055 23032 30067 23035
rect 31018 23032 31024 23044
rect 30055 23004 31024 23032
rect 30055 23001 30067 23004
rect 30009 22995 30067 23001
rect 31018 22992 31024 23004
rect 31076 22992 31082 23044
rect 31386 22992 31392 23044
rect 31444 23032 31450 23044
rect 32769 23035 32827 23041
rect 32769 23032 32781 23035
rect 31444 23004 32781 23032
rect 31444 22992 31450 23004
rect 32769 23001 32781 23004
rect 32815 23001 32827 23035
rect 32769 22995 32827 23001
rect 32950 22992 32956 23044
rect 33008 22992 33014 23044
rect 33778 22992 33784 23044
rect 33836 23032 33842 23044
rect 34701 23035 34759 23041
rect 34701 23032 34713 23035
rect 33836 23004 34713 23032
rect 33836 22992 33842 23004
rect 34701 23001 34713 23004
rect 34747 23001 34759 23035
rect 34701 22995 34759 23001
rect 35434 22992 35440 23044
rect 35492 23032 35498 23044
rect 37568 23032 37596 23072
rect 38381 23069 38393 23072
rect 38427 23069 38439 23103
rect 38381 23063 38439 23069
rect 38473 23103 38531 23109
rect 38473 23069 38485 23103
rect 38519 23100 38531 23103
rect 38562 23100 38568 23112
rect 38519 23072 38568 23100
rect 38519 23069 38531 23072
rect 38473 23063 38531 23069
rect 38562 23060 38568 23072
rect 38620 23060 38626 23112
rect 35492 23004 37596 23032
rect 38197 23035 38255 23041
rect 35492 22992 35498 23004
rect 38197 23001 38209 23035
rect 38243 23001 38255 23035
rect 38672 23032 38700 23140
rect 39945 23137 39957 23140
rect 39991 23137 40003 23171
rect 39945 23131 40003 23137
rect 40678 23128 40684 23180
rect 40736 23128 40742 23180
rect 40770 23128 40776 23180
rect 40828 23168 40834 23180
rect 40828 23140 41092 23168
rect 40828 23128 40834 23140
rect 39850 23060 39856 23112
rect 39908 23060 39914 23112
rect 40497 23103 40555 23109
rect 40497 23069 40509 23103
rect 40543 23100 40555 23103
rect 40862 23100 40868 23112
rect 40543 23072 40868 23100
rect 40543 23069 40555 23072
rect 40497 23063 40555 23069
rect 40862 23060 40868 23072
rect 40920 23060 40926 23112
rect 40957 23103 41015 23109
rect 40957 23069 40969 23103
rect 41003 23069 41015 23103
rect 41064 23100 41092 23140
rect 41138 23128 41144 23180
rect 41196 23168 41202 23180
rect 41417 23171 41475 23177
rect 41417 23168 41429 23171
rect 41196 23140 41429 23168
rect 41196 23128 41202 23140
rect 41417 23137 41429 23140
rect 41463 23137 41475 23171
rect 41417 23131 41475 23137
rect 41506 23128 41512 23180
rect 41564 23128 41570 23180
rect 41064 23072 41184 23100
rect 40957 23063 41015 23069
rect 38197 22995 38255 23001
rect 38626 23004 38700 23032
rect 31846 22964 31852 22976
rect 28460 22936 31852 22964
rect 31846 22924 31852 22936
rect 31904 22924 31910 22976
rect 32122 22924 32128 22976
rect 32180 22964 32186 22976
rect 34606 22964 34612 22976
rect 32180 22936 34612 22964
rect 32180 22924 32186 22936
rect 34606 22924 34612 22936
rect 34664 22924 34670 22976
rect 35618 22924 35624 22976
rect 35676 22964 35682 22976
rect 36817 22967 36875 22973
rect 36817 22964 36829 22967
rect 35676 22936 36829 22964
rect 35676 22924 35682 22936
rect 36817 22933 36829 22936
rect 36863 22933 36875 22967
rect 36817 22927 36875 22933
rect 37737 22967 37795 22973
rect 37737 22933 37749 22967
rect 37783 22964 37795 22967
rect 38212 22964 38240 22995
rect 37783 22936 38240 22964
rect 37783 22933 37795 22936
rect 37737 22927 37795 22933
rect 38470 22924 38476 22976
rect 38528 22964 38534 22976
rect 38626 22964 38654 23004
rect 38528 22936 38654 22964
rect 40313 22967 40371 22973
rect 38528 22924 38534 22936
rect 40313 22933 40325 22967
rect 40359 22964 40371 22967
rect 40402 22964 40408 22976
rect 40359 22936 40408 22964
rect 40359 22933 40371 22936
rect 40313 22927 40371 22933
rect 40402 22924 40408 22936
rect 40460 22924 40466 22976
rect 40972 22964 41000 23063
rect 41156 23032 41184 23072
rect 41230 23060 41236 23112
rect 41288 23060 41294 23112
rect 41340 23100 41451 23102
rect 41524 23100 41552 23128
rect 41340 23074 41552 23100
rect 41340 23032 41368 23074
rect 41423 23072 41552 23074
rect 41690 23060 41696 23112
rect 41748 23060 41754 23112
rect 42426 23060 42432 23112
rect 42484 23060 42490 23112
rect 41156 23004 41368 23032
rect 41785 22967 41843 22973
rect 41785 22964 41797 22967
rect 40972 22936 41797 22964
rect 41785 22933 41797 22936
rect 41831 22933 41843 22967
rect 41785 22927 41843 22933
rect 1104 22874 44896 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 44896 22874
rect 1104 22800 44896 22822
rect 5258 22760 5264 22772
rect 4724 22732 5264 22760
rect 4724 22633 4752 22732
rect 5258 22720 5264 22732
rect 5316 22760 5322 22772
rect 8941 22763 8999 22769
rect 5316 22732 5764 22760
rect 5316 22720 5322 22732
rect 4985 22695 5043 22701
rect 4985 22661 4997 22695
rect 5031 22692 5043 22695
rect 5031 22664 5488 22692
rect 5031 22661 5043 22664
rect 4985 22655 5043 22661
rect 5460 22636 5488 22664
rect 5626 22652 5632 22704
rect 5684 22652 5690 22704
rect 5736 22701 5764 22732
rect 8941 22729 8953 22763
rect 8987 22760 8999 22763
rect 9030 22760 9036 22772
rect 8987 22732 9036 22760
rect 8987 22729 8999 22732
rect 8941 22723 8999 22729
rect 9030 22720 9036 22732
rect 9088 22720 9094 22772
rect 9122 22720 9128 22772
rect 9180 22760 9186 22772
rect 9180 22732 12434 22760
rect 9180 22720 9186 22732
rect 5721 22695 5779 22701
rect 5721 22661 5733 22695
rect 5767 22692 5779 22695
rect 8110 22692 8116 22704
rect 5767 22664 8116 22692
rect 5767 22661 5779 22664
rect 5721 22655 5779 22661
rect 8110 22652 8116 22664
rect 8168 22652 8174 22704
rect 9398 22692 9404 22704
rect 9048 22664 9404 22692
rect 9048 22636 9076 22664
rect 9398 22652 9404 22664
rect 9456 22652 9462 22704
rect 9493 22695 9551 22701
rect 9493 22661 9505 22695
rect 9539 22692 9551 22695
rect 10321 22695 10379 22701
rect 9539 22664 10180 22692
rect 9539 22661 9551 22664
rect 9493 22655 9551 22661
rect 10152 22636 10180 22664
rect 10321 22661 10333 22695
rect 10367 22692 10379 22695
rect 11882 22692 11888 22704
rect 10367 22664 11888 22692
rect 10367 22661 10379 22664
rect 10321 22655 10379 22661
rect 11882 22652 11888 22664
rect 11940 22652 11946 22704
rect 12406 22692 12434 22732
rect 13354 22720 13360 22772
rect 13412 22720 13418 22772
rect 14461 22763 14519 22769
rect 14461 22729 14473 22763
rect 14507 22760 14519 22763
rect 14826 22760 14832 22772
rect 14507 22732 14832 22760
rect 14507 22729 14519 22732
rect 14461 22723 14519 22729
rect 14826 22720 14832 22732
rect 14884 22720 14890 22772
rect 15010 22720 15016 22772
rect 15068 22760 15074 22772
rect 21085 22763 21143 22769
rect 15068 22732 19748 22760
rect 15068 22720 15074 22732
rect 14001 22695 14059 22701
rect 14001 22692 14013 22695
rect 12406 22664 14013 22692
rect 14001 22661 14013 22664
rect 14047 22661 14059 22695
rect 16301 22695 16359 22701
rect 16301 22692 16313 22695
rect 14001 22655 14059 22661
rect 14200 22664 16313 22692
rect 4709 22627 4767 22633
rect 4709 22593 4721 22627
rect 4755 22624 4767 22627
rect 4798 22624 4804 22636
rect 4755 22596 4804 22624
rect 4755 22593 4767 22596
rect 4709 22587 4767 22593
rect 4798 22584 4804 22596
rect 4856 22584 4862 22636
rect 5166 22633 5172 22636
rect 4893 22627 4951 22633
rect 4893 22593 4905 22627
rect 4939 22593 4951 22627
rect 4893 22587 4951 22593
rect 5123 22627 5172 22633
rect 5123 22593 5135 22627
rect 5169 22593 5172 22627
rect 5123 22587 5172 22593
rect 3786 22516 3792 22568
rect 3844 22556 3850 22568
rect 4908 22556 4936 22587
rect 5166 22584 5172 22587
rect 5224 22584 5230 22636
rect 5442 22584 5448 22636
rect 5500 22584 5506 22636
rect 5810 22584 5816 22636
rect 5868 22584 5874 22636
rect 8386 22584 8392 22636
rect 8444 22624 8450 22636
rect 8481 22627 8539 22633
rect 8481 22624 8493 22627
rect 8444 22596 8493 22624
rect 8444 22584 8450 22596
rect 8481 22593 8493 22596
rect 8527 22593 8539 22627
rect 8481 22587 8539 22593
rect 8757 22627 8815 22633
rect 8757 22593 8769 22627
rect 8803 22624 8815 22627
rect 8803 22596 8984 22624
rect 8803 22593 8815 22596
rect 8757 22587 8815 22593
rect 5460 22556 5488 22584
rect 8202 22556 8208 22568
rect 3844 22528 5028 22556
rect 5460 22528 8208 22556
rect 3844 22516 3850 22528
rect 5000 22488 5028 22528
rect 8202 22516 8208 22528
rect 8260 22516 8266 22568
rect 8665 22559 8723 22565
rect 8665 22525 8677 22559
rect 8711 22556 8723 22559
rect 8846 22556 8852 22568
rect 8711 22528 8852 22556
rect 8711 22525 8723 22528
rect 8665 22519 8723 22525
rect 8846 22516 8852 22528
rect 8904 22516 8910 22568
rect 8956 22556 8984 22596
rect 9030 22584 9036 22636
rect 9088 22584 9094 22636
rect 9214 22584 9220 22636
rect 9272 22584 9278 22636
rect 9582 22624 9588 22636
rect 9640 22633 9646 22636
rect 9548 22596 9588 22624
rect 9582 22584 9588 22596
rect 9640 22587 9648 22633
rect 9640 22584 9646 22587
rect 9766 22584 9772 22636
rect 9824 22624 9830 22636
rect 9950 22624 9956 22636
rect 9824 22596 9956 22624
rect 9824 22584 9830 22596
rect 9950 22584 9956 22596
rect 10008 22584 10014 22636
rect 10042 22584 10048 22636
rect 10100 22584 10106 22636
rect 10134 22584 10140 22636
rect 10192 22624 10198 22636
rect 10229 22627 10287 22633
rect 10229 22624 10241 22627
rect 10192 22596 10241 22624
rect 10192 22584 10198 22596
rect 10229 22593 10241 22596
rect 10275 22593 10287 22627
rect 10418 22627 10476 22633
rect 10418 22624 10430 22627
rect 10229 22587 10287 22593
rect 10336 22596 10430 22624
rect 9122 22556 9128 22568
rect 8956 22528 9128 22556
rect 9122 22516 9128 22528
rect 9180 22516 9186 22568
rect 9232 22556 9260 22584
rect 10336 22568 10364 22596
rect 10418 22593 10430 22596
rect 10464 22593 10476 22627
rect 10418 22587 10476 22593
rect 10686 22584 10692 22636
rect 10744 22624 10750 22636
rect 11793 22627 11851 22633
rect 11793 22624 11805 22627
rect 10744 22596 11805 22624
rect 10744 22584 10750 22596
rect 11793 22593 11805 22596
rect 11839 22593 11851 22627
rect 11793 22587 11851 22593
rect 11977 22627 12035 22633
rect 11977 22593 11989 22627
rect 12023 22593 12035 22627
rect 11977 22587 12035 22593
rect 12253 22627 12311 22633
rect 12253 22593 12265 22627
rect 12299 22624 12311 22627
rect 12434 22624 12440 22636
rect 12299 22596 12440 22624
rect 12299 22593 12311 22596
rect 12253 22587 12311 22593
rect 9398 22556 9404 22568
rect 9232 22528 9404 22556
rect 9398 22516 9404 22528
rect 9456 22516 9462 22568
rect 10318 22516 10324 22568
rect 10376 22516 10382 22568
rect 11698 22516 11704 22568
rect 11756 22556 11762 22568
rect 11992 22556 12020 22587
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 12713 22627 12771 22633
rect 12713 22593 12725 22627
rect 12759 22624 12771 22627
rect 12802 22624 12808 22636
rect 12759 22596 12808 22624
rect 12759 22593 12771 22596
rect 12713 22587 12771 22593
rect 12802 22584 12808 22596
rect 12860 22584 12866 22636
rect 14200 22624 14228 22664
rect 16301 22661 16313 22664
rect 16347 22692 16359 22695
rect 19334 22692 19340 22704
rect 16347 22664 19340 22692
rect 16347 22661 16359 22664
rect 16301 22655 16359 22661
rect 19334 22652 19340 22664
rect 19392 22652 19398 22704
rect 13096 22596 14228 22624
rect 14277 22627 14335 22633
rect 11756 22528 12020 22556
rect 11756 22516 11762 22528
rect 12158 22516 12164 22568
rect 12216 22556 12222 22568
rect 13096 22565 13124 22596
rect 14277 22593 14289 22627
rect 14323 22624 14335 22627
rect 14366 22624 14372 22636
rect 14323 22596 14372 22624
rect 14323 22593 14335 22596
rect 14277 22587 14335 22593
rect 14366 22584 14372 22596
rect 14424 22584 14430 22636
rect 14550 22584 14556 22636
rect 14608 22624 14614 22636
rect 16485 22627 16543 22633
rect 16485 22624 16497 22627
rect 14608 22596 16497 22624
rect 14608 22584 14614 22596
rect 16485 22593 16497 22596
rect 16531 22624 16543 22627
rect 18506 22624 18512 22636
rect 16531 22596 18512 22624
rect 16531 22593 16543 22596
rect 16485 22587 16543 22593
rect 18506 22584 18512 22596
rect 18564 22584 18570 22636
rect 13081 22559 13139 22565
rect 13081 22556 13093 22559
rect 12216 22528 13093 22556
rect 12216 22516 12222 22528
rect 13081 22525 13093 22528
rect 13127 22525 13139 22559
rect 13081 22519 13139 22525
rect 13814 22516 13820 22568
rect 13872 22556 13878 22568
rect 13872 22528 14136 22556
rect 13872 22516 13878 22528
rect 5626 22488 5632 22500
rect 5000 22460 5632 22488
rect 5626 22448 5632 22460
rect 5684 22448 5690 22500
rect 5994 22448 6000 22500
rect 6052 22488 6058 22500
rect 12989 22491 13047 22497
rect 12989 22488 13001 22491
rect 6052 22460 13001 22488
rect 6052 22448 6058 22460
rect 12989 22457 13001 22460
rect 13035 22488 13047 22491
rect 13538 22488 13544 22500
rect 13035 22460 13544 22488
rect 13035 22457 13047 22460
rect 12989 22451 13047 22457
rect 13538 22448 13544 22460
rect 13596 22448 13602 22500
rect 5074 22380 5080 22432
rect 5132 22420 5138 22432
rect 5261 22423 5319 22429
rect 5261 22420 5273 22423
rect 5132 22392 5273 22420
rect 5132 22380 5138 22392
rect 5261 22389 5273 22392
rect 5307 22389 5319 22423
rect 5261 22383 5319 22389
rect 8662 22380 8668 22432
rect 8720 22380 8726 22432
rect 9769 22423 9827 22429
rect 9769 22389 9781 22423
rect 9815 22420 9827 22423
rect 10502 22420 10508 22432
rect 9815 22392 10508 22420
rect 9815 22389 9827 22392
rect 9769 22383 9827 22389
rect 10502 22380 10508 22392
rect 10560 22380 10566 22432
rect 10597 22423 10655 22429
rect 10597 22389 10609 22423
rect 10643 22420 10655 22423
rect 10778 22420 10784 22432
rect 10643 22392 10784 22420
rect 10643 22389 10655 22392
rect 10597 22383 10655 22389
rect 10778 22380 10784 22392
rect 10836 22380 10842 22432
rect 12437 22423 12495 22429
rect 12437 22389 12449 22423
rect 12483 22420 12495 22423
rect 12710 22420 12716 22432
rect 12483 22392 12716 22420
rect 12483 22389 12495 22392
rect 12437 22383 12495 22389
rect 12710 22380 12716 22392
rect 12768 22380 12774 22432
rect 12878 22423 12936 22429
rect 12878 22389 12890 22423
rect 12924 22420 12936 22423
rect 13170 22420 13176 22432
rect 12924 22392 13176 22420
rect 12924 22389 12936 22392
rect 12878 22383 12936 22389
rect 13170 22380 13176 22392
rect 13228 22380 13234 22432
rect 14108 22429 14136 22528
rect 14182 22516 14188 22568
rect 14240 22516 14246 22568
rect 14366 22448 14372 22500
rect 14424 22488 14430 22500
rect 16942 22488 16948 22500
rect 14424 22460 16948 22488
rect 14424 22448 14430 22460
rect 16942 22448 16948 22460
rect 17000 22448 17006 22500
rect 19720 22488 19748 22732
rect 21085 22729 21097 22763
rect 21131 22760 21143 22763
rect 23658 22760 23664 22772
rect 21131 22732 21956 22760
rect 21131 22729 21143 22732
rect 21085 22723 21143 22729
rect 20346 22652 20352 22704
rect 20404 22692 20410 22704
rect 21177 22695 21235 22701
rect 21177 22692 21189 22695
rect 20404 22664 21189 22692
rect 20404 22652 20410 22664
rect 21177 22661 21189 22664
rect 21223 22661 21235 22695
rect 21542 22692 21548 22704
rect 21177 22655 21235 22661
rect 21376 22664 21548 22692
rect 19794 22584 19800 22636
rect 19852 22624 19858 22636
rect 20625 22627 20683 22633
rect 20625 22624 20637 22627
rect 19852 22596 20637 22624
rect 19852 22584 19858 22596
rect 20625 22593 20637 22596
rect 20671 22593 20683 22627
rect 20625 22587 20683 22593
rect 20806 22584 20812 22636
rect 20864 22584 20870 22636
rect 21376 22633 21404 22664
rect 21542 22652 21548 22664
rect 21600 22652 21606 22704
rect 21928 22701 21956 22732
rect 22020 22732 23664 22760
rect 21913 22695 21971 22701
rect 21913 22661 21925 22695
rect 21959 22661 21971 22695
rect 21913 22655 21971 22661
rect 20901 22627 20959 22633
rect 20901 22593 20913 22627
rect 20947 22624 20959 22627
rect 21361 22627 21419 22633
rect 20947 22596 21036 22624
rect 20947 22593 20959 22596
rect 20901 22587 20959 22593
rect 21008 22568 21036 22596
rect 21361 22593 21373 22627
rect 21407 22593 21419 22627
rect 21361 22587 21419 22593
rect 21450 22584 21456 22636
rect 21508 22624 21514 22636
rect 22020 22624 22048 22732
rect 23658 22720 23664 22732
rect 23716 22720 23722 22772
rect 26697 22763 26755 22769
rect 26697 22729 26709 22763
rect 26743 22729 26755 22763
rect 26697 22723 26755 22729
rect 29457 22763 29515 22769
rect 29457 22729 29469 22763
rect 29503 22760 29515 22763
rect 29503 22732 31754 22760
rect 29503 22729 29515 22732
rect 29457 22723 29515 22729
rect 22094 22652 22100 22704
rect 22152 22692 22158 22704
rect 24486 22692 24492 22704
rect 22152 22664 24492 22692
rect 22152 22652 22158 22664
rect 24486 22652 24492 22664
rect 24544 22652 24550 22704
rect 26712 22692 26740 22723
rect 27338 22692 27344 22704
rect 26712 22664 27344 22692
rect 27338 22652 27344 22664
rect 27396 22652 27402 22704
rect 28997 22695 29055 22701
rect 28997 22661 29009 22695
rect 29043 22692 29055 22695
rect 29086 22692 29092 22704
rect 29043 22664 29092 22692
rect 29043 22661 29055 22664
rect 28997 22655 29055 22661
rect 29086 22652 29092 22664
rect 29144 22652 29150 22704
rect 29362 22652 29368 22704
rect 29420 22692 29426 22704
rect 29546 22692 29552 22704
rect 29420 22664 29552 22692
rect 29420 22652 29426 22664
rect 29546 22652 29552 22664
rect 29604 22652 29610 22704
rect 29822 22652 29828 22704
rect 29880 22692 29886 22704
rect 31478 22692 31484 22704
rect 29880 22664 31484 22692
rect 29880 22652 29886 22664
rect 31478 22652 31484 22664
rect 31536 22652 31542 22704
rect 31726 22692 31754 22732
rect 31846 22720 31852 22772
rect 31904 22760 31910 22772
rect 32950 22760 32956 22772
rect 31904 22732 32956 22760
rect 31904 22720 31910 22732
rect 32950 22720 32956 22732
rect 33008 22720 33014 22772
rect 33410 22720 33416 22772
rect 33468 22760 33474 22772
rect 33962 22760 33968 22772
rect 33468 22732 33968 22760
rect 33468 22720 33474 22732
rect 33962 22720 33968 22732
rect 34020 22720 34026 22772
rect 36538 22720 36544 22772
rect 36596 22760 36602 22772
rect 38470 22760 38476 22772
rect 36596 22732 38476 22760
rect 36596 22720 36602 22732
rect 38470 22720 38476 22732
rect 38528 22720 38534 22772
rect 41693 22763 41751 22769
rect 41693 22729 41705 22763
rect 41739 22760 41751 22763
rect 42426 22760 42432 22772
rect 41739 22732 42432 22760
rect 41739 22729 41751 22732
rect 41693 22723 41751 22729
rect 42426 22720 42432 22732
rect 42484 22720 42490 22772
rect 33318 22692 33324 22704
rect 31726 22664 33324 22692
rect 33318 22652 33324 22664
rect 33376 22652 33382 22704
rect 36354 22652 36360 22704
rect 36412 22692 36418 22704
rect 38102 22692 38108 22704
rect 36412 22664 38108 22692
rect 36412 22652 36418 22664
rect 38102 22652 38108 22664
rect 38160 22652 38166 22704
rect 40862 22652 40868 22704
rect 40920 22692 40926 22704
rect 41782 22692 41788 22704
rect 40920 22664 41788 22692
rect 40920 22652 40926 22664
rect 41782 22652 41788 22664
rect 41840 22652 41846 22704
rect 21508 22596 22048 22624
rect 21508 22584 21514 22596
rect 22186 22584 22192 22636
rect 22244 22624 22250 22636
rect 22830 22624 22836 22636
rect 22244 22596 22836 22624
rect 22244 22584 22250 22596
rect 22830 22584 22836 22596
rect 22888 22584 22894 22636
rect 24305 22627 24363 22633
rect 24305 22593 24317 22627
rect 24351 22624 24363 22627
rect 24394 22624 24400 22636
rect 24351 22596 24400 22624
rect 24351 22593 24363 22596
rect 24305 22587 24363 22593
rect 24394 22584 24400 22596
rect 24452 22584 24458 22636
rect 25222 22584 25228 22636
rect 25280 22624 25286 22636
rect 26142 22624 26148 22636
rect 25280 22596 26148 22624
rect 25280 22584 25286 22596
rect 26142 22584 26148 22596
rect 26200 22584 26206 22636
rect 26234 22584 26240 22636
rect 26292 22584 26298 22636
rect 26510 22584 26516 22636
rect 26568 22584 26574 22636
rect 26878 22584 26884 22636
rect 26936 22624 26942 22636
rect 26936 22596 29224 22624
rect 26936 22584 26942 22596
rect 20990 22516 20996 22568
rect 21048 22516 21054 22568
rect 22005 22559 22063 22565
rect 22005 22525 22017 22559
rect 22051 22525 22063 22559
rect 22005 22519 22063 22525
rect 21637 22491 21695 22497
rect 19720 22460 21496 22488
rect 14093 22423 14151 22429
rect 14093 22389 14105 22423
rect 14139 22389 14151 22423
rect 14093 22383 14151 22389
rect 16209 22423 16267 22429
rect 16209 22389 16221 22423
rect 16255 22420 16267 22423
rect 16298 22420 16304 22432
rect 16255 22392 16304 22420
rect 16255 22389 16267 22392
rect 16209 22383 16267 22389
rect 16298 22380 16304 22392
rect 16356 22420 16362 22432
rect 20530 22420 20536 22432
rect 16356 22392 20536 22420
rect 16356 22380 16362 22392
rect 20530 22380 20536 22392
rect 20588 22380 20594 22432
rect 20806 22380 20812 22432
rect 20864 22380 20870 22432
rect 21468 22429 21496 22460
rect 21637 22457 21649 22491
rect 21683 22488 21695 22491
rect 22020 22488 22048 22519
rect 24854 22516 24860 22568
rect 24912 22556 24918 22568
rect 26050 22556 26056 22568
rect 24912 22528 26056 22556
rect 24912 22516 24918 22528
rect 26050 22516 26056 22528
rect 26108 22516 26114 22568
rect 26326 22556 26332 22568
rect 26160 22528 26332 22556
rect 21683 22460 22048 22488
rect 21683 22457 21695 22460
rect 21637 22451 21695 22457
rect 21453 22423 21511 22429
rect 21453 22389 21465 22423
rect 21499 22420 21511 22423
rect 21818 22420 21824 22432
rect 21499 22392 21824 22420
rect 21499 22389 21511 22392
rect 21453 22383 21511 22389
rect 21818 22380 21824 22392
rect 21876 22380 21882 22432
rect 22189 22423 22247 22429
rect 22189 22389 22201 22423
rect 22235 22420 22247 22423
rect 22278 22420 22284 22432
rect 22235 22392 22284 22420
rect 22235 22389 22247 22392
rect 22189 22383 22247 22389
rect 22278 22380 22284 22392
rect 22336 22380 22342 22432
rect 22370 22380 22376 22432
rect 22428 22380 22434 22432
rect 23934 22380 23940 22432
rect 23992 22420 23998 22432
rect 24673 22423 24731 22429
rect 24673 22420 24685 22423
rect 23992 22392 24685 22420
rect 23992 22380 23998 22392
rect 24673 22389 24685 22392
rect 24719 22420 24731 22423
rect 25590 22420 25596 22432
rect 24719 22392 25596 22420
rect 24719 22389 24731 22392
rect 24673 22383 24731 22389
rect 25590 22380 25596 22392
rect 25648 22380 25654 22432
rect 26160 22420 26188 22528
rect 26326 22516 26332 22528
rect 26384 22516 26390 22568
rect 27338 22516 27344 22568
rect 27396 22556 27402 22568
rect 28994 22556 29000 22568
rect 27396 22528 29000 22556
rect 27396 22516 27402 22528
rect 28994 22516 29000 22528
rect 29052 22516 29058 22568
rect 29089 22559 29147 22565
rect 29089 22525 29101 22559
rect 29135 22525 29147 22559
rect 29196 22556 29224 22596
rect 29270 22584 29276 22636
rect 29328 22584 29334 22636
rect 31018 22584 31024 22636
rect 31076 22584 31082 22636
rect 31202 22584 31208 22636
rect 31260 22584 31266 22636
rect 31294 22584 31300 22636
rect 31352 22624 31358 22636
rect 31757 22627 31815 22633
rect 31757 22624 31769 22627
rect 31352 22596 31769 22624
rect 31352 22584 31358 22596
rect 31757 22593 31769 22596
rect 31803 22593 31815 22627
rect 31757 22587 31815 22593
rect 31941 22627 31999 22633
rect 31941 22593 31953 22627
rect 31987 22624 31999 22627
rect 35618 22624 35624 22636
rect 31987 22596 35624 22624
rect 31987 22593 31999 22596
rect 31941 22587 31999 22593
rect 35618 22584 35624 22596
rect 35676 22584 35682 22636
rect 38010 22584 38016 22636
rect 38068 22624 38074 22636
rect 38378 22624 38384 22636
rect 38068 22596 38384 22624
rect 38068 22584 38074 22596
rect 38378 22584 38384 22596
rect 38436 22584 38442 22636
rect 40310 22584 40316 22636
rect 40368 22584 40374 22636
rect 40402 22584 40408 22636
rect 40460 22624 40466 22636
rect 40569 22627 40627 22633
rect 40569 22624 40581 22627
rect 40460 22596 40581 22624
rect 40460 22584 40466 22596
rect 40569 22593 40581 22596
rect 40615 22593 40627 22627
rect 40569 22587 40627 22593
rect 42426 22584 42432 22636
rect 42484 22624 42490 22636
rect 44269 22627 44327 22633
rect 44269 22624 44281 22627
rect 42484 22596 44281 22624
rect 42484 22584 42490 22596
rect 44269 22593 44281 22596
rect 44315 22593 44327 22627
rect 44269 22587 44327 22593
rect 30926 22556 30932 22568
rect 29196 22528 30932 22556
rect 29089 22519 29147 22525
rect 26326 22420 26332 22432
rect 26160 22392 26332 22420
rect 26326 22380 26332 22392
rect 26384 22380 26390 22432
rect 26513 22423 26571 22429
rect 26513 22389 26525 22423
rect 26559 22420 26571 22423
rect 27430 22420 27436 22432
rect 26559 22392 27436 22420
rect 26559 22389 26571 22392
rect 26513 22383 26571 22389
rect 27430 22380 27436 22392
rect 27488 22380 27494 22432
rect 28994 22380 29000 22432
rect 29052 22420 29058 22432
rect 29104 22420 29132 22519
rect 30926 22516 30932 22528
rect 30984 22516 30990 22568
rect 29270 22448 29276 22500
rect 29328 22488 29334 22500
rect 29730 22488 29736 22500
rect 29328 22460 29736 22488
rect 29328 22448 29334 22460
rect 29730 22448 29736 22460
rect 29788 22448 29794 22500
rect 31036 22488 31064 22584
rect 32950 22516 32956 22568
rect 33008 22556 33014 22568
rect 37918 22556 37924 22568
rect 33008 22528 37924 22556
rect 33008 22516 33014 22528
rect 37918 22516 37924 22528
rect 37976 22516 37982 22568
rect 31036 22460 31800 22488
rect 29052 22392 29132 22420
rect 29052 22380 29058 22392
rect 29178 22380 29184 22432
rect 29236 22380 29242 22432
rect 30926 22380 30932 22432
rect 30984 22420 30990 22432
rect 31021 22423 31079 22429
rect 31021 22420 31033 22423
rect 30984 22392 31033 22420
rect 30984 22380 30990 22392
rect 31021 22389 31033 22392
rect 31067 22420 31079 22423
rect 31294 22420 31300 22432
rect 31067 22392 31300 22420
rect 31067 22389 31079 22392
rect 31021 22383 31079 22389
rect 31294 22380 31300 22392
rect 31352 22380 31358 22432
rect 31386 22380 31392 22432
rect 31444 22380 31450 22432
rect 31478 22380 31484 22432
rect 31536 22420 31542 22432
rect 31772 22429 31800 22460
rect 33410 22448 33416 22500
rect 33468 22488 33474 22500
rect 35526 22488 35532 22500
rect 33468 22460 35532 22488
rect 33468 22448 33474 22460
rect 35526 22448 35532 22460
rect 35584 22448 35590 22500
rect 44450 22448 44456 22500
rect 44508 22448 44514 22500
rect 31573 22423 31631 22429
rect 31573 22420 31585 22423
rect 31536 22392 31585 22420
rect 31536 22380 31542 22392
rect 31573 22389 31585 22392
rect 31619 22389 31631 22423
rect 31573 22383 31631 22389
rect 31757 22423 31815 22429
rect 31757 22389 31769 22423
rect 31803 22389 31815 22423
rect 31757 22383 31815 22389
rect 32030 22380 32036 22432
rect 32088 22420 32094 22432
rect 36814 22420 36820 22432
rect 32088 22392 36820 22420
rect 32088 22380 32094 22392
rect 36814 22380 36820 22392
rect 36872 22420 36878 22432
rect 39758 22420 39764 22432
rect 36872 22392 39764 22420
rect 36872 22380 36878 22392
rect 39758 22380 39764 22392
rect 39816 22380 39822 22432
rect 1104 22330 44896 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 44896 22330
rect 1104 22256 44896 22278
rect 5353 22219 5411 22225
rect 5353 22185 5365 22219
rect 5399 22216 5411 22219
rect 5718 22216 5724 22228
rect 5399 22188 5724 22216
rect 5399 22185 5411 22188
rect 5353 22179 5411 22185
rect 5718 22176 5724 22188
rect 5776 22176 5782 22228
rect 7285 22219 7343 22225
rect 7285 22185 7297 22219
rect 7331 22216 7343 22219
rect 7374 22216 7380 22228
rect 7331 22188 7380 22216
rect 7331 22185 7343 22188
rect 7285 22179 7343 22185
rect 7374 22176 7380 22188
rect 7432 22176 7438 22228
rect 7742 22216 7748 22228
rect 7484 22188 7748 22216
rect 5810 22108 5816 22160
rect 5868 22148 5874 22160
rect 7484 22148 7512 22188
rect 7742 22176 7748 22188
rect 7800 22216 7806 22228
rect 10686 22216 10692 22228
rect 7800 22188 10692 22216
rect 7800 22176 7806 22188
rect 10686 22176 10692 22188
rect 10744 22176 10750 22228
rect 13538 22176 13544 22228
rect 13596 22216 13602 22228
rect 14550 22216 14556 22228
rect 13596 22188 14556 22216
rect 13596 22176 13602 22188
rect 14550 22176 14556 22188
rect 14608 22176 14614 22228
rect 14918 22176 14924 22228
rect 14976 22176 14982 22228
rect 15197 22219 15255 22225
rect 15197 22185 15209 22219
rect 15243 22216 15255 22219
rect 15562 22216 15568 22228
rect 15243 22188 15568 22216
rect 15243 22185 15255 22188
rect 15197 22179 15255 22185
rect 15562 22176 15568 22188
rect 15620 22176 15626 22228
rect 15838 22176 15844 22228
rect 15896 22216 15902 22228
rect 16298 22216 16304 22228
rect 15896 22188 16304 22216
rect 15896 22176 15902 22188
rect 16298 22176 16304 22188
rect 16356 22216 16362 22228
rect 16356 22188 16804 22216
rect 16356 22176 16362 22188
rect 5868 22120 7512 22148
rect 5868 22108 5874 22120
rect 10134 22108 10140 22160
rect 10192 22148 10198 22160
rect 10410 22148 10416 22160
rect 10192 22120 10416 22148
rect 10192 22108 10198 22120
rect 10410 22108 10416 22120
rect 10468 22108 10474 22160
rect 12158 22108 12164 22160
rect 12216 22108 12222 22160
rect 12805 22151 12863 22157
rect 12805 22148 12817 22151
rect 12783 22120 12817 22148
rect 12805 22117 12817 22120
rect 12851 22117 12863 22151
rect 12805 22111 12863 22117
rect 6454 22040 6460 22092
rect 6512 22080 6518 22092
rect 7193 22083 7251 22089
rect 7193 22080 7205 22083
rect 6512 22052 7205 22080
rect 6512 22040 6518 22052
rect 7193 22049 7205 22052
rect 7239 22080 7251 22083
rect 7239 22052 7788 22080
rect 7239 22049 7251 22052
rect 7193 22043 7251 22049
rect 5074 21972 5080 22024
rect 5132 21972 5138 22024
rect 5258 21972 5264 22024
rect 5316 21972 5322 22024
rect 5353 22015 5411 22021
rect 5353 21981 5365 22015
rect 5399 22012 5411 22015
rect 5902 22012 5908 22024
rect 5399 21984 5908 22012
rect 5399 21981 5411 21984
rect 5353 21975 5411 21981
rect 5902 21972 5908 21984
rect 5960 22012 5966 22024
rect 6472 22012 6500 22040
rect 7760 22021 7788 22052
rect 7926 22040 7932 22092
rect 7984 22040 7990 22092
rect 11054 22040 11060 22092
rect 11112 22080 11118 22092
rect 11330 22080 11336 22092
rect 11112 22052 11336 22080
rect 11112 22040 11118 22052
rect 11330 22040 11336 22052
rect 11388 22040 11394 22092
rect 12820 22080 12848 22111
rect 13906 22108 13912 22160
rect 13964 22108 13970 22160
rect 13998 22108 14004 22160
rect 14056 22148 14062 22160
rect 14274 22148 14280 22160
rect 14056 22120 14280 22148
rect 14056 22108 14062 22120
rect 14274 22108 14280 22120
rect 14332 22108 14338 22160
rect 13924 22080 13952 22108
rect 11624 22052 12480 22080
rect 12820 22052 13952 22080
rect 5960 21984 6500 22012
rect 7101 22015 7159 22021
rect 5960 21972 5966 21984
rect 7101 21981 7113 22015
rect 7147 21981 7159 22015
rect 7101 21975 7159 21981
rect 7745 22015 7803 22021
rect 7745 21981 7757 22015
rect 7791 21981 7803 22015
rect 7745 21975 7803 21981
rect 6641 21947 6699 21953
rect 6641 21913 6653 21947
rect 6687 21913 6699 21947
rect 6641 21907 6699 21913
rect 6825 21947 6883 21953
rect 6825 21913 6837 21947
rect 6871 21944 6883 21947
rect 6914 21944 6920 21956
rect 6871 21916 6920 21944
rect 6871 21913 6883 21916
rect 6825 21907 6883 21913
rect 5534 21836 5540 21888
rect 5592 21836 5598 21888
rect 6656 21876 6684 21907
rect 6914 21904 6920 21916
rect 6972 21904 6978 21956
rect 7006 21904 7012 21956
rect 7064 21904 7070 21956
rect 7116 21876 7144 21975
rect 10042 21972 10048 22024
rect 10100 22012 10106 22024
rect 10410 22012 10416 22024
rect 10100 21984 10416 22012
rect 10100 21972 10106 21984
rect 10410 21972 10416 21984
rect 10468 22012 10474 22024
rect 11624 22021 11652 22052
rect 12452 22024 12480 22052
rect 15838 22040 15844 22092
rect 15896 22080 15902 22092
rect 16482 22080 16488 22092
rect 15896 22052 16488 22080
rect 15896 22040 15902 22052
rect 16482 22040 16488 22052
rect 16540 22040 16546 22092
rect 11609 22015 11667 22021
rect 11609 22012 11621 22015
rect 10468 21984 11621 22012
rect 10468 21972 10474 21984
rect 11609 21981 11621 21984
rect 11655 21981 11667 22015
rect 11609 21975 11667 21981
rect 11974 21972 11980 22024
rect 12032 21972 12038 22024
rect 12066 21972 12072 22024
rect 12124 22012 12130 22024
rect 12253 22015 12311 22021
rect 12253 22012 12265 22015
rect 12124 21984 12265 22012
rect 12124 21972 12130 21984
rect 12253 21981 12265 21984
rect 12299 21981 12311 22015
rect 12253 21975 12311 21981
rect 12434 21972 12440 22024
rect 12492 21972 12498 22024
rect 12621 22015 12679 22021
rect 12621 21981 12633 22015
rect 12667 21981 12679 22015
rect 12621 21975 12679 21981
rect 7374 21904 7380 21956
rect 7432 21944 7438 21956
rect 7561 21947 7619 21953
rect 7561 21944 7573 21947
rect 7432 21916 7573 21944
rect 7432 21904 7438 21916
rect 7561 21913 7573 21916
rect 7607 21913 7619 21947
rect 7561 21907 7619 21913
rect 8202 21904 8208 21956
rect 8260 21944 8266 21956
rect 9674 21944 9680 21956
rect 8260 21916 9680 21944
rect 8260 21904 8266 21916
rect 9674 21904 9680 21916
rect 9732 21944 9738 21956
rect 10870 21944 10876 21956
rect 9732 21916 10876 21944
rect 9732 21904 9738 21916
rect 10870 21904 10876 21916
rect 10928 21904 10934 21956
rect 11330 21904 11336 21956
rect 11388 21944 11394 21956
rect 11698 21944 11704 21956
rect 11388 21916 11704 21944
rect 11388 21904 11394 21916
rect 11698 21904 11704 21916
rect 11756 21944 11762 21956
rect 11793 21947 11851 21953
rect 11793 21944 11805 21947
rect 11756 21916 11805 21944
rect 11756 21904 11762 21916
rect 11793 21913 11805 21916
rect 11839 21913 11851 21947
rect 11793 21907 11851 21913
rect 11882 21904 11888 21956
rect 11940 21904 11946 21956
rect 12526 21904 12532 21956
rect 12584 21904 12590 21956
rect 7282 21876 7288 21888
rect 6656 21848 7288 21876
rect 7282 21836 7288 21848
rect 7340 21836 7346 21888
rect 7469 21879 7527 21885
rect 7469 21845 7481 21879
rect 7515 21876 7527 21879
rect 8478 21876 8484 21888
rect 7515 21848 8484 21876
rect 7515 21845 7527 21848
rect 7469 21839 7527 21845
rect 8478 21836 8484 21848
rect 8536 21836 8542 21888
rect 11900 21876 11928 21904
rect 12636 21876 12664 21975
rect 14918 21972 14924 22024
rect 14976 21972 14982 22024
rect 15010 21972 15016 22024
rect 15068 21972 15074 22024
rect 15746 21972 15752 22024
rect 15804 22012 15810 22024
rect 16776 22021 16804 22188
rect 17126 22176 17132 22228
rect 17184 22216 17190 22228
rect 17773 22219 17831 22225
rect 17773 22216 17785 22219
rect 17184 22188 17785 22216
rect 17184 22176 17190 22188
rect 17773 22185 17785 22188
rect 17819 22185 17831 22219
rect 17773 22179 17831 22185
rect 19337 22219 19395 22225
rect 19337 22185 19349 22219
rect 19383 22216 19395 22219
rect 20806 22216 20812 22228
rect 19383 22188 20812 22216
rect 19383 22185 19395 22188
rect 19337 22179 19395 22185
rect 16942 22108 16948 22160
rect 17000 22148 17006 22160
rect 19352 22148 19380 22179
rect 20806 22176 20812 22188
rect 20864 22176 20870 22228
rect 21174 22176 21180 22228
rect 21232 22216 21238 22228
rect 21542 22216 21548 22228
rect 21232 22188 21548 22216
rect 21232 22176 21238 22188
rect 21542 22176 21548 22188
rect 21600 22176 21606 22228
rect 25130 22176 25136 22228
rect 25188 22176 25194 22228
rect 25222 22176 25228 22228
rect 25280 22216 25286 22228
rect 25685 22219 25743 22225
rect 25685 22216 25697 22219
rect 25280 22188 25697 22216
rect 25280 22176 25286 22188
rect 25685 22185 25697 22188
rect 25731 22185 25743 22219
rect 25685 22179 25743 22185
rect 17000 22120 19380 22148
rect 17000 22108 17006 22120
rect 19610 22108 19616 22160
rect 19668 22148 19674 22160
rect 20438 22148 20444 22160
rect 19668 22120 20444 22148
rect 19668 22108 19674 22120
rect 20438 22108 20444 22120
rect 20496 22108 20502 22160
rect 24670 22148 24676 22160
rect 24228 22120 24676 22148
rect 18046 22040 18052 22092
rect 18104 22080 18110 22092
rect 18693 22083 18751 22089
rect 18693 22080 18705 22083
rect 18104 22052 18705 22080
rect 18104 22040 18110 22052
rect 18693 22049 18705 22052
rect 18739 22049 18751 22083
rect 18693 22043 18751 22049
rect 19429 22083 19487 22089
rect 19429 22049 19441 22083
rect 19475 22080 19487 22083
rect 21266 22080 21272 22092
rect 19475 22052 21272 22080
rect 19475 22049 19487 22052
rect 19429 22043 19487 22049
rect 21266 22040 21272 22052
rect 21324 22080 21330 22092
rect 21634 22080 21640 22092
rect 21324 22052 21640 22080
rect 21324 22040 21330 22052
rect 21634 22040 21640 22052
rect 21692 22040 21698 22092
rect 24228 22024 24256 22120
rect 24670 22108 24676 22120
rect 24728 22108 24734 22160
rect 25700 22148 25728 22179
rect 26050 22176 26056 22228
rect 26108 22216 26114 22228
rect 26108 22188 26740 22216
rect 26108 22176 26114 22188
rect 26326 22148 26332 22160
rect 25700 22120 26332 22148
rect 26326 22108 26332 22120
rect 26384 22108 26390 22160
rect 26418 22108 26424 22160
rect 26476 22148 26482 22160
rect 26602 22148 26608 22160
rect 26476 22120 26608 22148
rect 26476 22108 26482 22120
rect 26602 22108 26608 22120
rect 26660 22108 26666 22160
rect 26712 22148 26740 22188
rect 26786 22176 26792 22228
rect 26844 22176 26850 22228
rect 27246 22176 27252 22228
rect 27304 22216 27310 22228
rect 27798 22216 27804 22228
rect 27304 22188 27804 22216
rect 27304 22176 27310 22188
rect 27798 22176 27804 22188
rect 27856 22176 27862 22228
rect 27982 22176 27988 22228
rect 28040 22216 28046 22228
rect 28166 22216 28172 22228
rect 28040 22188 28172 22216
rect 28040 22176 28046 22188
rect 28166 22176 28172 22188
rect 28224 22216 28230 22228
rect 28353 22219 28411 22225
rect 28353 22216 28365 22219
rect 28224 22188 28365 22216
rect 28224 22176 28230 22188
rect 28353 22185 28365 22188
rect 28399 22185 28411 22219
rect 28353 22179 28411 22185
rect 28442 22176 28448 22228
rect 28500 22216 28506 22228
rect 32677 22219 32735 22225
rect 32677 22216 32689 22219
rect 28500 22188 32689 22216
rect 28500 22176 28506 22188
rect 32677 22185 32689 22188
rect 32723 22185 32735 22219
rect 32677 22179 32735 22185
rect 33042 22176 33048 22228
rect 33100 22216 33106 22228
rect 33137 22219 33195 22225
rect 33137 22216 33149 22219
rect 33100 22188 33149 22216
rect 33100 22176 33106 22188
rect 33137 22185 33149 22188
rect 33183 22185 33195 22219
rect 33137 22179 33195 22185
rect 33226 22176 33232 22228
rect 33284 22176 33290 22228
rect 33502 22176 33508 22228
rect 33560 22216 33566 22228
rect 33560 22188 34284 22216
rect 33560 22176 33566 22188
rect 27816 22148 27844 22176
rect 26712 22120 27476 22148
rect 27816 22120 28304 22148
rect 24578 22040 24584 22092
rect 24636 22080 24642 22092
rect 24765 22083 24823 22089
rect 24765 22080 24777 22083
rect 24636 22052 24777 22080
rect 24636 22040 24642 22052
rect 24765 22049 24777 22052
rect 24811 22049 24823 22083
rect 25593 22083 25651 22089
rect 24765 22043 24823 22049
rect 24964 22052 25544 22080
rect 15933 22015 15991 22021
rect 15933 22012 15945 22015
rect 15804 21984 15945 22012
rect 15804 21972 15810 21984
rect 15933 21981 15945 21984
rect 15979 21981 15991 22015
rect 15933 21975 15991 21981
rect 16761 22015 16819 22021
rect 16761 21981 16773 22015
rect 16807 21981 16819 22015
rect 16761 21975 16819 21981
rect 16850 21972 16856 22024
rect 16908 22012 16914 22024
rect 17773 22015 17831 22021
rect 17773 22012 17785 22015
rect 16908 21984 17785 22012
rect 16908 21972 16914 21984
rect 17773 21981 17785 21984
rect 17819 21981 17831 22015
rect 17773 21975 17831 21981
rect 17865 22015 17923 22021
rect 17865 21981 17877 22015
rect 17911 22012 17923 22015
rect 18230 22012 18236 22024
rect 17911 21984 18236 22012
rect 17911 21981 17923 21984
rect 17865 21975 17923 21981
rect 18230 21972 18236 21984
rect 18288 22012 18294 22024
rect 19150 22012 19156 22024
rect 18288 21984 19156 22012
rect 18288 21972 18294 21984
rect 19150 21972 19156 21984
rect 19208 21972 19214 22024
rect 19242 21972 19248 22024
rect 19300 21972 19306 22024
rect 19518 21972 19524 22024
rect 19576 22012 19582 22024
rect 21174 22012 21180 22024
rect 19576 21984 21180 22012
rect 19576 21972 19582 21984
rect 21174 21972 21180 21984
rect 21232 21972 21238 22024
rect 24210 21972 24216 22024
rect 24268 21972 24274 22024
rect 24964 22012 24992 22052
rect 24320 21984 24992 22012
rect 25041 22015 25099 22021
rect 14550 21904 14556 21956
rect 14608 21944 14614 21956
rect 14737 21947 14795 21953
rect 14737 21944 14749 21947
rect 14608 21916 14749 21944
rect 14608 21904 14614 21916
rect 14737 21913 14749 21916
rect 14783 21913 14795 21947
rect 14737 21907 14795 21913
rect 14826 21904 14832 21956
rect 14884 21944 14890 21956
rect 15657 21947 15715 21953
rect 15657 21944 15669 21947
rect 14884 21916 15669 21944
rect 14884 21904 14890 21916
rect 15657 21913 15669 21916
rect 15703 21913 15715 21947
rect 15657 21907 15715 21913
rect 16482 21904 16488 21956
rect 16540 21944 16546 21956
rect 16577 21947 16635 21953
rect 16577 21944 16589 21947
rect 16540 21916 16589 21944
rect 16540 21904 16546 21916
rect 16577 21913 16589 21916
rect 16623 21913 16635 21947
rect 16577 21907 16635 21913
rect 16942 21904 16948 21956
rect 17000 21904 17006 21956
rect 18064 21916 18276 21944
rect 12710 21876 12716 21888
rect 11900 21848 12716 21876
rect 12710 21836 12716 21848
rect 12768 21836 12774 21888
rect 12802 21836 12808 21888
rect 12860 21876 12866 21888
rect 13538 21876 13544 21888
rect 12860 21848 13544 21876
rect 12860 21836 12866 21848
rect 13538 21836 13544 21848
rect 13596 21836 13602 21888
rect 16117 21879 16175 21885
rect 16117 21845 16129 21879
rect 16163 21876 16175 21879
rect 18064 21876 18092 21916
rect 16163 21848 18092 21876
rect 16163 21845 16175 21848
rect 16117 21839 16175 21845
rect 18138 21836 18144 21888
rect 18196 21836 18202 21888
rect 18248 21876 18276 21916
rect 18322 21904 18328 21956
rect 18380 21904 18386 21956
rect 18506 21904 18512 21956
rect 18564 21904 18570 21956
rect 18874 21904 18880 21956
rect 18932 21944 18938 21956
rect 19260 21944 19288 21972
rect 24320 21944 24348 21984
rect 25041 21981 25053 22015
rect 25087 21981 25099 22015
rect 25041 21975 25099 21981
rect 18932 21916 19288 21944
rect 19628 21916 24348 21944
rect 18932 21904 18938 21916
rect 19628 21876 19656 21916
rect 24394 21904 24400 21956
rect 24452 21904 24458 21956
rect 24581 21947 24639 21953
rect 24581 21913 24593 21947
rect 24627 21913 24639 21947
rect 24581 21907 24639 21913
rect 18248 21848 19656 21876
rect 19705 21879 19763 21885
rect 19705 21845 19717 21879
rect 19751 21876 19763 21879
rect 20622 21876 20628 21888
rect 19751 21848 20628 21876
rect 19751 21845 19763 21848
rect 19705 21839 19763 21845
rect 20622 21836 20628 21848
rect 20680 21836 20686 21888
rect 21818 21836 21824 21888
rect 21876 21876 21882 21888
rect 24486 21876 24492 21888
rect 21876 21848 24492 21876
rect 21876 21836 21882 21848
rect 24486 21836 24492 21848
rect 24544 21836 24550 21888
rect 24596 21876 24624 21907
rect 24854 21904 24860 21956
rect 24912 21904 24918 21956
rect 25056 21944 25084 21975
rect 25130 21972 25136 22024
rect 25188 21972 25194 22024
rect 25222 21944 25228 21956
rect 25056 21916 25228 21944
rect 25222 21904 25228 21916
rect 25280 21904 25286 21956
rect 25409 21947 25467 21953
rect 25409 21944 25421 21947
rect 25332 21916 25421 21944
rect 25038 21876 25044 21888
rect 24596 21848 25044 21876
rect 25038 21836 25044 21848
rect 25096 21836 25102 21888
rect 25332 21885 25360 21916
rect 25409 21913 25421 21916
rect 25455 21913 25467 21947
rect 25409 21907 25467 21913
rect 25317 21879 25375 21885
rect 25317 21845 25329 21879
rect 25363 21845 25375 21879
rect 25516 21876 25544 22052
rect 25593 22049 25605 22083
rect 25639 22080 25651 22083
rect 25958 22080 25964 22092
rect 25639 22052 25964 22080
rect 25639 22049 25651 22052
rect 25593 22043 25651 22049
rect 25958 22040 25964 22052
rect 26016 22040 26022 22092
rect 26142 22040 26148 22092
rect 26200 22040 26206 22092
rect 27154 22080 27160 22092
rect 26344 22052 27160 22080
rect 25685 22015 25743 22021
rect 25685 21981 25697 22015
rect 25731 22012 25743 22015
rect 26160 22012 26188 22040
rect 26344 22021 26372 22052
rect 27154 22040 27160 22052
rect 27212 22040 27218 22092
rect 25731 21984 26188 22012
rect 26329 22015 26387 22021
rect 25731 21981 25743 21984
rect 25685 21975 25743 21981
rect 26329 21981 26341 22015
rect 26375 21981 26387 22015
rect 26605 22015 26663 22021
rect 26605 22012 26617 22015
rect 26329 21975 26387 21981
rect 26436 21984 26617 22012
rect 25958 21904 25964 21956
rect 26016 21944 26022 21956
rect 26053 21947 26111 21953
rect 26053 21944 26065 21947
rect 26016 21916 26065 21944
rect 26016 21904 26022 21916
rect 26053 21913 26065 21916
rect 26099 21913 26111 21947
rect 26053 21907 26111 21913
rect 25682 21876 25688 21888
rect 25516 21848 25688 21876
rect 25317 21839 25375 21845
rect 25682 21836 25688 21848
rect 25740 21836 25746 21888
rect 25869 21879 25927 21885
rect 25869 21845 25881 21879
rect 25915 21876 25927 21879
rect 26436 21876 26464 21984
rect 26605 21981 26617 21984
rect 26651 21981 26663 22015
rect 26605 21975 26663 21981
rect 26786 21972 26792 22024
rect 26844 21972 26850 22024
rect 27448 22012 27476 22120
rect 27982 22040 27988 22092
rect 28040 22040 28046 22092
rect 28276 22080 28304 22120
rect 30558 22108 30564 22160
rect 30616 22148 30622 22160
rect 31110 22148 31116 22160
rect 30616 22120 31116 22148
rect 30616 22108 30622 22120
rect 31110 22108 31116 22120
rect 31168 22108 31174 22160
rect 31202 22108 31208 22160
rect 31260 22148 31266 22160
rect 31478 22148 31484 22160
rect 31260 22120 31484 22148
rect 31260 22108 31266 22120
rect 31478 22108 31484 22120
rect 31536 22108 31542 22160
rect 34146 22148 34152 22160
rect 33060 22120 34152 22148
rect 28276 22052 28994 22080
rect 28966 22024 28994 22052
rect 31018 22040 31024 22092
rect 31076 22080 31082 22092
rect 33060 22080 33088 22120
rect 34146 22108 34152 22120
rect 34204 22108 34210 22160
rect 34256 22080 34284 22188
rect 34514 22176 34520 22228
rect 34572 22216 34578 22228
rect 34701 22219 34759 22225
rect 34701 22216 34713 22219
rect 34572 22188 34713 22216
rect 34572 22176 34578 22188
rect 34701 22185 34713 22188
rect 34747 22185 34759 22219
rect 34701 22179 34759 22185
rect 35158 22176 35164 22228
rect 35216 22216 35222 22228
rect 35434 22216 35440 22228
rect 35216 22188 35440 22216
rect 35216 22176 35222 22188
rect 35434 22176 35440 22188
rect 35492 22176 35498 22228
rect 35805 22219 35863 22225
rect 35805 22185 35817 22219
rect 35851 22216 35863 22219
rect 36354 22216 36360 22228
rect 35851 22188 36360 22216
rect 35851 22185 35863 22188
rect 35805 22179 35863 22185
rect 36354 22176 36360 22188
rect 36412 22176 36418 22228
rect 41230 22216 41236 22228
rect 40236 22188 41236 22216
rect 35250 22108 35256 22160
rect 35308 22148 35314 22160
rect 36078 22148 36084 22160
rect 35308 22120 36084 22148
rect 35308 22108 35314 22120
rect 36078 22108 36084 22120
rect 36136 22108 36142 22160
rect 31076 22052 33088 22080
rect 33244 22052 33456 22080
rect 34256 22052 35020 22080
rect 31076 22040 31082 22052
rect 27448 21984 28028 22012
rect 27801 21947 27859 21953
rect 27801 21944 27813 21947
rect 26528 21916 27813 21944
rect 26528 21885 26556 21916
rect 27801 21913 27813 21916
rect 27847 21913 27859 21947
rect 28000 21944 28028 21984
rect 28074 21972 28080 22024
rect 28132 22012 28138 22024
rect 28353 22015 28411 22021
rect 28353 22012 28365 22015
rect 28132 21984 28365 22012
rect 28132 21972 28138 21984
rect 28353 21981 28365 21984
rect 28399 21981 28411 22015
rect 28353 21975 28411 21981
rect 28445 22015 28503 22021
rect 28445 21981 28457 22015
rect 28491 21981 28503 22015
rect 28966 21984 29000 22024
rect 28445 21975 28503 21981
rect 28460 21944 28488 21975
rect 28994 21972 29000 21984
rect 29052 21972 29058 22024
rect 33244 22021 33272 22052
rect 33428 22022 33456 22052
rect 32861 22015 32919 22021
rect 32861 22012 32873 22015
rect 31726 21984 32873 22012
rect 31726 21944 31754 21984
rect 32861 21981 32873 21984
rect 32907 21981 32919 22015
rect 32861 21975 32919 21981
rect 32953 22015 33011 22021
rect 32953 21981 32965 22015
rect 32999 21981 33011 22015
rect 32953 21975 33011 21981
rect 33229 22015 33287 22021
rect 33229 21981 33241 22015
rect 33275 21981 33287 22015
rect 33229 21975 33287 21981
rect 33321 22015 33379 22021
rect 33321 21981 33333 22015
rect 33367 21981 33379 22015
rect 33428 22012 33640 22022
rect 33686 22012 33692 22024
rect 33428 21994 33692 22012
rect 33612 21984 33692 21994
rect 33321 21975 33379 21981
rect 28000 21916 28488 21944
rect 28644 21916 31754 21944
rect 27801 21907 27859 21913
rect 25915 21848 26464 21876
rect 26513 21879 26571 21885
rect 25915 21845 25927 21848
rect 25869 21839 25927 21845
rect 26513 21845 26525 21879
rect 26559 21845 26571 21879
rect 26513 21839 26571 21845
rect 26970 21836 26976 21888
rect 27028 21836 27034 21888
rect 28261 21879 28319 21885
rect 28261 21845 28273 21879
rect 28307 21876 28319 21879
rect 28644 21876 28672 21916
rect 32490 21904 32496 21956
rect 32548 21944 32554 21956
rect 32677 21947 32735 21953
rect 32677 21944 32689 21947
rect 32548 21916 32689 21944
rect 32548 21904 32554 21916
rect 32677 21913 32689 21916
rect 32723 21913 32735 21947
rect 32677 21907 32735 21913
rect 28307 21848 28672 21876
rect 28721 21879 28779 21885
rect 28307 21845 28319 21848
rect 28261 21839 28319 21845
rect 28721 21845 28733 21879
rect 28767 21876 28779 21879
rect 32030 21876 32036 21888
rect 28767 21848 32036 21876
rect 28767 21845 28779 21848
rect 28721 21839 28779 21845
rect 32030 21836 32036 21848
rect 32088 21836 32094 21888
rect 32968 21876 32996 21975
rect 33042 21904 33048 21956
rect 33100 21944 33106 21956
rect 33336 21944 33364 21975
rect 33686 21972 33692 21984
rect 33744 21972 33750 22024
rect 34992 22021 35020 22052
rect 35526 22040 35532 22092
rect 35584 22080 35590 22092
rect 35621 22083 35679 22089
rect 35621 22080 35633 22083
rect 35584 22052 35633 22080
rect 35584 22040 35590 22052
rect 35621 22049 35633 22052
rect 35667 22080 35679 22083
rect 38378 22080 38384 22092
rect 35667 22052 38384 22080
rect 35667 22049 35679 22052
rect 35621 22043 35679 22049
rect 38378 22040 38384 22052
rect 38436 22040 38442 22092
rect 34885 22015 34943 22021
rect 34885 21981 34897 22015
rect 34931 21981 34943 22015
rect 34885 21975 34943 21981
rect 34977 22015 35035 22021
rect 34977 21981 34989 22015
rect 35023 21981 35035 22015
rect 34977 21975 35035 21981
rect 33100 21916 33364 21944
rect 33100 21904 33106 21916
rect 34054 21904 34060 21956
rect 34112 21944 34118 21956
rect 34514 21944 34520 21956
rect 34112 21916 34520 21944
rect 34112 21904 34118 21916
rect 34514 21904 34520 21916
rect 34572 21904 34578 21956
rect 34698 21904 34704 21956
rect 34756 21904 34762 21956
rect 33597 21879 33655 21885
rect 33597 21876 33609 21879
rect 32968 21848 33609 21876
rect 33597 21845 33609 21848
rect 33643 21876 33655 21879
rect 34900 21876 34928 21975
rect 35434 21972 35440 22024
rect 35492 22012 35498 22024
rect 35805 22015 35863 22021
rect 35805 22012 35817 22015
rect 35492 21984 35817 22012
rect 35492 21972 35498 21984
rect 35805 21981 35817 21984
rect 35851 21981 35863 22015
rect 35805 21975 35863 21981
rect 40034 21972 40040 22024
rect 40092 22012 40098 22024
rect 40236 22012 40264 22188
rect 41230 22176 41236 22188
rect 41288 22176 41294 22228
rect 40310 22108 40316 22160
rect 40368 22108 40374 22160
rect 40328 22080 40356 22108
rect 41509 22083 41567 22089
rect 41509 22080 41521 22083
rect 40328 22052 41521 22080
rect 41509 22049 41521 22052
rect 41555 22049 41567 22083
rect 41509 22043 41567 22049
rect 40313 22015 40371 22021
rect 40313 22012 40325 22015
rect 40092 21984 40325 22012
rect 40092 21972 40098 21984
rect 40313 21981 40325 21984
rect 40359 21981 40371 22015
rect 40313 21975 40371 21981
rect 40402 21972 40408 22024
rect 40460 21972 40466 22024
rect 40497 22015 40555 22021
rect 40497 21981 40509 22015
rect 40543 21981 40555 22015
rect 40497 21975 40555 21981
rect 40589 22015 40647 22021
rect 40589 21981 40601 22015
rect 40635 22012 40647 22015
rect 40678 22012 40684 22024
rect 40635 21984 40684 22012
rect 40635 21981 40647 21984
rect 40589 21975 40647 21981
rect 35526 21904 35532 21956
rect 35584 21904 35590 21956
rect 38654 21944 38660 21956
rect 35912 21916 38660 21944
rect 33643 21848 34928 21876
rect 35161 21879 35219 21885
rect 33643 21845 33655 21848
rect 33597 21839 33655 21845
rect 35161 21845 35173 21879
rect 35207 21876 35219 21879
rect 35912 21876 35940 21916
rect 38654 21904 38660 21916
rect 38712 21904 38718 21956
rect 38930 21904 38936 21956
rect 38988 21944 38994 21956
rect 40512 21944 40540 21975
rect 40678 21972 40684 21984
rect 40736 21972 40742 22024
rect 40773 22015 40831 22021
rect 40773 21981 40785 22015
rect 40819 22012 40831 22015
rect 42981 22015 43039 22021
rect 42981 22012 42993 22015
rect 40819 21984 42993 22012
rect 40819 21981 40831 21984
rect 40773 21975 40831 21981
rect 42981 21981 42993 21984
rect 43027 21981 43039 22015
rect 42981 21975 43039 21981
rect 43530 21972 43536 22024
rect 43588 21972 43594 22024
rect 44269 22015 44327 22021
rect 44269 21981 44281 22015
rect 44315 21981 44327 22015
rect 44269 21975 44327 21981
rect 38988 21916 40540 21944
rect 41776 21947 41834 21953
rect 38988 21904 38994 21916
rect 41776 21913 41788 21947
rect 41822 21944 41834 21947
rect 43346 21944 43352 21956
rect 41822 21916 43352 21944
rect 41822 21913 41834 21916
rect 41776 21907 41834 21913
rect 43346 21904 43352 21916
rect 43404 21904 43410 21956
rect 35207 21848 35940 21876
rect 35207 21845 35219 21848
rect 35161 21839 35219 21845
rect 35986 21836 35992 21888
rect 36044 21836 36050 21888
rect 36446 21836 36452 21888
rect 36504 21876 36510 21888
rect 39942 21876 39948 21888
rect 36504 21848 39948 21876
rect 36504 21836 36510 21848
rect 39942 21836 39948 21848
rect 40000 21836 40006 21888
rect 40126 21836 40132 21888
rect 40184 21836 40190 21888
rect 42889 21879 42947 21885
rect 42889 21845 42901 21879
rect 42935 21876 42947 21879
rect 43070 21876 43076 21888
rect 42935 21848 43076 21876
rect 42935 21845 42947 21848
rect 42889 21839 42947 21845
rect 43070 21836 43076 21848
rect 43128 21876 43134 21888
rect 44284 21876 44312 21975
rect 43128 21848 44312 21876
rect 43128 21836 43134 21848
rect 44450 21836 44456 21888
rect 44508 21836 44514 21888
rect 1104 21786 44896 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 44896 21786
rect 1104 21712 44896 21734
rect 6181 21675 6239 21681
rect 6181 21641 6193 21675
rect 6227 21672 6239 21675
rect 6914 21672 6920 21684
rect 6227 21644 6920 21672
rect 6227 21641 6239 21644
rect 6181 21635 6239 21641
rect 6914 21632 6920 21644
rect 6972 21672 6978 21684
rect 7374 21672 7380 21684
rect 6972 21644 7380 21672
rect 6972 21632 6978 21644
rect 7374 21632 7380 21644
rect 7432 21672 7438 21684
rect 7834 21672 7840 21684
rect 7432 21644 7840 21672
rect 7432 21632 7438 21644
rect 7834 21632 7840 21644
rect 7892 21632 7898 21684
rect 8478 21632 8484 21684
rect 8536 21672 8542 21684
rect 9030 21672 9036 21684
rect 8536 21644 9036 21672
rect 8536 21632 8542 21644
rect 9030 21632 9036 21644
rect 9088 21632 9094 21684
rect 9858 21632 9864 21684
rect 9916 21632 9922 21684
rect 11054 21672 11060 21684
rect 9968 21644 11060 21672
rect 2869 21607 2927 21613
rect 2869 21573 2881 21607
rect 2915 21604 2927 21607
rect 3970 21604 3976 21616
rect 2915 21576 3976 21604
rect 2915 21573 2927 21576
rect 2869 21567 2927 21573
rect 3970 21564 3976 21576
rect 4028 21564 4034 21616
rect 9968 21604 9996 21644
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 12802 21672 12808 21684
rect 11532 21644 12020 21672
rect 8220 21576 9996 21604
rect 2682 21496 2688 21548
rect 2740 21496 2746 21548
rect 2961 21539 3019 21545
rect 2961 21505 2973 21539
rect 3007 21505 3019 21539
rect 2961 21499 3019 21505
rect 3053 21539 3111 21545
rect 3053 21505 3065 21539
rect 3099 21536 3111 21539
rect 3099 21508 4936 21536
rect 3099 21505 3111 21508
rect 3053 21499 3111 21505
rect 2498 21428 2504 21480
rect 2556 21468 2562 21480
rect 2976 21468 3004 21499
rect 4908 21480 4936 21508
rect 5626 21496 5632 21548
rect 5684 21496 5690 21548
rect 5810 21496 5816 21548
rect 5868 21496 5874 21548
rect 5902 21496 5908 21548
rect 5960 21496 5966 21548
rect 5997 21539 6055 21545
rect 5997 21505 6009 21539
rect 6043 21505 6055 21539
rect 5997 21499 6055 21505
rect 2556 21440 3004 21468
rect 2556 21428 2562 21440
rect 4890 21428 4896 21480
rect 4948 21468 4954 21480
rect 6012 21468 6040 21499
rect 6362 21496 6368 21548
rect 6420 21536 6426 21548
rect 8220 21536 8248 21576
rect 10042 21564 10048 21616
rect 10100 21604 10106 21616
rect 10229 21607 10287 21613
rect 10229 21604 10241 21607
rect 10100 21576 10241 21604
rect 10100 21564 10106 21576
rect 10229 21573 10241 21576
rect 10275 21604 10287 21607
rect 11532 21604 11560 21644
rect 10275 21576 11560 21604
rect 10275 21573 10287 21576
rect 10229 21567 10287 21573
rect 11606 21564 11612 21616
rect 11664 21604 11670 21616
rect 11882 21604 11888 21616
rect 11664 21576 11888 21604
rect 11664 21564 11670 21576
rect 11882 21564 11888 21576
rect 11940 21564 11946 21616
rect 11992 21604 12020 21644
rect 12452 21644 12808 21672
rect 12452 21604 12480 21644
rect 12802 21632 12808 21644
rect 12860 21632 12866 21684
rect 12897 21675 12955 21681
rect 12897 21641 12909 21675
rect 12943 21672 12955 21675
rect 14366 21672 14372 21684
rect 12943 21644 14372 21672
rect 12943 21641 12955 21644
rect 12897 21635 12955 21641
rect 14366 21632 14372 21644
rect 14424 21632 14430 21684
rect 20806 21632 20812 21684
rect 20864 21632 20870 21684
rect 31018 21672 31024 21684
rect 20916 21644 31024 21672
rect 11992 21576 12480 21604
rect 12621 21607 12679 21613
rect 12621 21573 12633 21607
rect 12667 21604 12679 21607
rect 13722 21604 13728 21616
rect 12667 21576 13728 21604
rect 12667 21573 12679 21576
rect 12621 21567 12679 21573
rect 13722 21564 13728 21576
rect 13780 21564 13786 21616
rect 14550 21564 14556 21616
rect 14608 21604 14614 21616
rect 14608 21576 18092 21604
rect 14608 21564 14614 21576
rect 6420 21508 8248 21536
rect 6420 21496 6426 21508
rect 8754 21496 8760 21548
rect 8812 21536 8818 21548
rect 9677 21539 9735 21545
rect 9677 21536 9689 21539
rect 8812 21508 9689 21536
rect 8812 21496 8818 21508
rect 9677 21505 9689 21508
rect 9723 21505 9735 21539
rect 9677 21499 9735 21505
rect 9950 21496 9956 21548
rect 10008 21496 10014 21548
rect 10137 21539 10195 21545
rect 10137 21505 10149 21539
rect 10183 21505 10195 21539
rect 10137 21499 10195 21505
rect 10321 21539 10379 21545
rect 10321 21505 10333 21539
rect 10367 21536 10379 21539
rect 10686 21536 10692 21548
rect 10367 21508 10692 21536
rect 10367 21505 10379 21508
rect 10321 21499 10379 21505
rect 4948 21440 6040 21468
rect 4948 21428 4954 21440
rect 9490 21428 9496 21480
rect 9548 21468 9554 21480
rect 10152 21468 10180 21499
rect 10686 21496 10692 21508
rect 10744 21496 10750 21548
rect 12158 21496 12164 21548
rect 12216 21536 12222 21548
rect 12345 21539 12403 21545
rect 12345 21536 12357 21539
rect 12216 21508 12357 21536
rect 12216 21496 12222 21508
rect 12345 21505 12357 21508
rect 12391 21505 12403 21539
rect 12345 21499 12403 21505
rect 12434 21496 12440 21548
rect 12492 21536 12498 21548
rect 12529 21539 12587 21545
rect 12529 21536 12541 21539
rect 12492 21508 12541 21536
rect 12492 21496 12498 21508
rect 12529 21505 12541 21508
rect 12575 21505 12587 21539
rect 12529 21499 12587 21505
rect 12710 21496 12716 21548
rect 12768 21496 12774 21548
rect 13262 21496 13268 21548
rect 13320 21536 13326 21548
rect 17678 21536 17684 21548
rect 13320 21508 17684 21536
rect 13320 21496 13326 21508
rect 17678 21496 17684 21508
rect 17736 21496 17742 21548
rect 18064 21536 18092 21576
rect 18138 21564 18144 21616
rect 18196 21604 18202 21616
rect 20916 21604 20944 21644
rect 31018 21632 31024 21644
rect 31076 21632 31082 21684
rect 32030 21632 32036 21684
rect 32088 21672 32094 21684
rect 32306 21672 32312 21684
rect 32088 21644 32312 21672
rect 32088 21632 32094 21644
rect 32306 21632 32312 21644
rect 32364 21632 32370 21684
rect 33042 21672 33048 21684
rect 32508 21644 33048 21672
rect 18196 21576 20944 21604
rect 18196 21564 18202 21576
rect 23934 21564 23940 21616
rect 23992 21564 23998 21616
rect 24489 21607 24547 21613
rect 24489 21573 24501 21607
rect 24535 21604 24547 21607
rect 24578 21604 24584 21616
rect 24535 21576 24584 21604
rect 24535 21573 24547 21576
rect 24489 21567 24547 21573
rect 24578 21564 24584 21576
rect 24636 21564 24642 21616
rect 25148 21576 30512 21604
rect 20441 21539 20499 21545
rect 20441 21536 20453 21539
rect 18064 21508 20453 21536
rect 20441 21505 20453 21508
rect 20487 21505 20499 21539
rect 20441 21499 20499 21505
rect 10962 21468 10968 21480
rect 9548 21440 10968 21468
rect 9548 21428 9554 21440
rect 10962 21428 10968 21440
rect 11020 21468 11026 21480
rect 14826 21468 14832 21480
rect 11020 21440 14832 21468
rect 11020 21428 11026 21440
rect 14826 21428 14832 21440
rect 14884 21428 14890 21480
rect 14918 21428 14924 21480
rect 14976 21468 14982 21480
rect 17494 21468 17500 21480
rect 14976 21440 17500 21468
rect 14976 21428 14982 21440
rect 17494 21428 17500 21440
rect 17552 21428 17558 21480
rect 20456 21468 20484 21499
rect 20622 21496 20628 21548
rect 20680 21536 20686 21548
rect 21177 21539 21235 21545
rect 21177 21536 21189 21539
rect 20680 21508 21189 21536
rect 20680 21496 20686 21508
rect 21177 21505 21189 21508
rect 21223 21505 21235 21539
rect 21177 21499 21235 21505
rect 21266 21496 21272 21548
rect 21324 21536 21330 21548
rect 21361 21539 21419 21545
rect 21361 21536 21373 21539
rect 21324 21508 21373 21536
rect 21324 21496 21330 21508
rect 21361 21505 21373 21508
rect 21407 21505 21419 21539
rect 23842 21536 23848 21548
rect 21361 21499 21419 21505
rect 21468 21508 23848 21536
rect 20714 21468 20720 21480
rect 20456 21440 20720 21468
rect 20714 21428 20720 21440
rect 20772 21468 20778 21480
rect 21468 21468 21496 21508
rect 23842 21496 23848 21508
rect 23900 21536 23906 21548
rect 24213 21539 24271 21545
rect 24213 21536 24225 21539
rect 23900 21508 24225 21536
rect 23900 21496 23906 21508
rect 24213 21505 24225 21508
rect 24259 21505 24271 21539
rect 24213 21499 24271 21505
rect 24394 21496 24400 21548
rect 24452 21536 24458 21548
rect 24670 21536 24676 21548
rect 24452 21508 24532 21536
rect 24452 21496 24458 21508
rect 20772 21440 21496 21468
rect 20772 21428 20778 21440
rect 23106 21428 23112 21480
rect 23164 21468 23170 21480
rect 24029 21471 24087 21477
rect 24029 21468 24041 21471
rect 23164 21440 24041 21468
rect 23164 21428 23170 21440
rect 24029 21437 24041 21440
rect 24075 21437 24087 21471
rect 24029 21431 24087 21437
rect 3237 21403 3295 21409
rect 3237 21369 3249 21403
rect 3283 21400 3295 21403
rect 9674 21400 9680 21412
rect 3283 21372 9680 21400
rect 3283 21369 3295 21372
rect 3237 21363 3295 21369
rect 9674 21360 9680 21372
rect 9732 21360 9738 21412
rect 11974 21360 11980 21412
rect 12032 21400 12038 21412
rect 15470 21400 15476 21412
rect 12032 21372 15476 21400
rect 12032 21360 12038 21372
rect 15470 21360 15476 21372
rect 15528 21360 15534 21412
rect 17218 21360 17224 21412
rect 17276 21400 17282 21412
rect 23842 21400 23848 21412
rect 17276 21372 23848 21400
rect 17276 21360 17282 21372
rect 23842 21360 23848 21372
rect 23900 21360 23906 21412
rect 24394 21360 24400 21412
rect 24452 21360 24458 21412
rect 24504 21400 24532 21508
rect 24596 21508 24676 21536
rect 24596 21480 24624 21508
rect 24670 21496 24676 21508
rect 24728 21496 24734 21548
rect 24765 21539 24823 21545
rect 24765 21505 24777 21539
rect 24811 21505 24823 21539
rect 24765 21499 24823 21505
rect 24578 21428 24584 21480
rect 24636 21428 24642 21480
rect 24780 21412 24808 21499
rect 24854 21496 24860 21548
rect 24912 21526 24918 21548
rect 25148 21536 25176 21576
rect 24964 21526 25176 21536
rect 24912 21508 25176 21526
rect 24912 21498 24992 21508
rect 24912 21496 24918 21498
rect 26970 21496 26976 21548
rect 27028 21536 27034 21548
rect 30484 21545 30512 21576
rect 29813 21539 29871 21545
rect 29813 21536 29825 21539
rect 27028 21508 29825 21536
rect 27028 21496 27034 21508
rect 29813 21505 29825 21508
rect 29859 21505 29871 21539
rect 29813 21499 29871 21505
rect 30469 21539 30527 21545
rect 30469 21505 30481 21539
rect 30515 21536 30527 21539
rect 30558 21536 30564 21548
rect 30515 21508 30564 21536
rect 30515 21505 30527 21508
rect 30469 21499 30527 21505
rect 30558 21496 30564 21508
rect 30616 21496 30622 21548
rect 30742 21496 30748 21548
rect 30800 21496 30806 21548
rect 30834 21496 30840 21548
rect 30892 21536 30898 21548
rect 30892 21508 31064 21536
rect 30892 21496 30898 21508
rect 25958 21428 25964 21480
rect 26016 21468 26022 21480
rect 27798 21468 27804 21480
rect 26016 21440 27804 21468
rect 26016 21428 26022 21440
rect 27798 21428 27804 21440
rect 27856 21428 27862 21480
rect 29917 21471 29975 21477
rect 29917 21437 29929 21471
rect 29963 21468 29975 21471
rect 30653 21471 30711 21477
rect 29963 21440 30420 21468
rect 29963 21437 29975 21440
rect 29917 21431 29975 21437
rect 24504 21372 24624 21400
rect 5626 21292 5632 21344
rect 5684 21332 5690 21344
rect 6362 21332 6368 21344
rect 5684 21304 6368 21332
rect 5684 21292 5690 21304
rect 6362 21292 6368 21304
rect 6420 21292 6426 21344
rect 8570 21292 8576 21344
rect 8628 21332 8634 21344
rect 8846 21332 8852 21344
rect 8628 21304 8852 21332
rect 8628 21292 8634 21304
rect 8846 21292 8852 21304
rect 8904 21332 8910 21344
rect 10226 21332 10232 21344
rect 8904 21304 10232 21332
rect 8904 21292 8910 21304
rect 10226 21292 10232 21304
rect 10284 21292 10290 21344
rect 10505 21335 10563 21341
rect 10505 21301 10517 21335
rect 10551 21332 10563 21335
rect 11422 21332 11428 21344
rect 10551 21304 11428 21332
rect 10551 21301 10563 21304
rect 10505 21295 10563 21301
rect 11422 21292 11428 21304
rect 11480 21332 11486 21344
rect 14918 21332 14924 21344
rect 11480 21304 14924 21332
rect 11480 21292 11486 21304
rect 14918 21292 14924 21304
rect 14976 21292 14982 21344
rect 15010 21292 15016 21344
rect 15068 21332 15074 21344
rect 19518 21332 19524 21344
rect 15068 21304 19524 21332
rect 15068 21292 15074 21304
rect 19518 21292 19524 21304
rect 19576 21292 19582 21344
rect 19610 21292 19616 21344
rect 19668 21332 19674 21344
rect 20070 21332 20076 21344
rect 19668 21304 20076 21332
rect 19668 21292 19674 21304
rect 20070 21292 20076 21304
rect 20128 21292 20134 21344
rect 20806 21292 20812 21344
rect 20864 21332 20870 21344
rect 20990 21332 20996 21344
rect 20864 21304 20996 21332
rect 20864 21292 20870 21304
rect 20990 21292 20996 21304
rect 21048 21292 21054 21344
rect 21542 21292 21548 21344
rect 21600 21292 21606 21344
rect 23474 21292 23480 21344
rect 23532 21332 23538 21344
rect 23937 21335 23995 21341
rect 23937 21332 23949 21335
rect 23532 21304 23949 21332
rect 23532 21292 23538 21304
rect 23937 21301 23949 21304
rect 23983 21332 23995 21335
rect 24026 21332 24032 21344
rect 23983 21304 24032 21332
rect 23983 21301 23995 21304
rect 23937 21295 23995 21301
rect 24026 21292 24032 21304
rect 24084 21292 24090 21344
rect 24210 21292 24216 21344
rect 24268 21332 24274 21344
rect 24489 21335 24547 21341
rect 24489 21332 24501 21335
rect 24268 21304 24501 21332
rect 24268 21292 24274 21304
rect 24489 21301 24501 21304
rect 24535 21301 24547 21335
rect 24596 21332 24624 21372
rect 24762 21360 24768 21412
rect 24820 21360 24826 21412
rect 24854 21360 24860 21412
rect 24912 21400 24918 21412
rect 24949 21403 25007 21409
rect 24949 21400 24961 21403
rect 24912 21372 24961 21400
rect 24912 21360 24918 21372
rect 24949 21369 24961 21372
rect 24995 21369 25007 21403
rect 24949 21363 25007 21369
rect 27062 21360 27068 21412
rect 27120 21400 27126 21412
rect 29730 21400 29736 21412
rect 27120 21372 29736 21400
rect 27120 21360 27126 21372
rect 29730 21360 29736 21372
rect 29788 21360 29794 21412
rect 27338 21332 27344 21344
rect 24596 21304 27344 21332
rect 24489 21295 24547 21301
rect 27338 21292 27344 21304
rect 27396 21292 27402 21344
rect 30006 21292 30012 21344
rect 30064 21292 30070 21344
rect 30190 21292 30196 21344
rect 30248 21292 30254 21344
rect 30285 21335 30343 21341
rect 30285 21301 30297 21335
rect 30331 21332 30343 21335
rect 30392 21332 30420 21440
rect 30653 21437 30665 21471
rect 30699 21468 30711 21471
rect 30926 21468 30932 21480
rect 30699 21440 30932 21468
rect 30699 21437 30711 21440
rect 30653 21431 30711 21437
rect 30926 21428 30932 21440
rect 30984 21428 30990 21480
rect 31036 21468 31064 21508
rect 31202 21496 31208 21548
rect 31260 21496 31266 21548
rect 31481 21539 31539 21545
rect 31481 21505 31493 21539
rect 31527 21536 31539 21539
rect 31570 21536 31576 21548
rect 31527 21508 31576 21536
rect 31527 21505 31539 21508
rect 31481 21499 31539 21505
rect 31570 21496 31576 21508
rect 31628 21496 31634 21548
rect 32306 21496 32312 21548
rect 32364 21536 32370 21548
rect 32508 21545 32536 21644
rect 33042 21632 33048 21644
rect 33100 21632 33106 21684
rect 33226 21632 33232 21684
rect 33284 21632 33290 21684
rect 34701 21675 34759 21681
rect 33520 21644 34468 21672
rect 33520 21604 33548 21644
rect 32968 21576 33548 21604
rect 32493 21539 32551 21545
rect 32493 21536 32505 21539
rect 32364 21508 32505 21536
rect 32364 21496 32370 21508
rect 32493 21505 32505 21508
rect 32539 21505 32551 21539
rect 32493 21499 32551 21505
rect 31297 21471 31355 21477
rect 31297 21468 31309 21471
rect 31036 21440 31309 21468
rect 31297 21437 31309 21440
rect 31343 21437 31355 21471
rect 31297 21431 31355 21437
rect 32398 21428 32404 21480
rect 32456 21468 32462 21480
rect 32968 21468 32996 21576
rect 33502 21496 33508 21548
rect 33560 21496 33566 21548
rect 33689 21539 33747 21545
rect 33689 21505 33701 21539
rect 33735 21536 33747 21539
rect 34333 21539 34391 21545
rect 34333 21536 34345 21539
rect 33735 21508 34345 21536
rect 33735 21505 33747 21508
rect 33689 21499 33747 21505
rect 34333 21505 34345 21508
rect 34379 21505 34391 21539
rect 34440 21536 34468 21644
rect 34701 21641 34713 21675
rect 34747 21672 34759 21675
rect 35342 21672 35348 21684
rect 34747 21644 35348 21672
rect 34747 21641 34759 21644
rect 34701 21635 34759 21641
rect 35342 21632 35348 21644
rect 35400 21632 35406 21684
rect 37200 21644 37964 21672
rect 35066 21564 35072 21616
rect 35124 21604 35130 21616
rect 37200 21604 37228 21644
rect 35124 21576 37228 21604
rect 35124 21564 35130 21576
rect 37274 21564 37280 21616
rect 37332 21564 37338 21616
rect 37366 21564 37372 21616
rect 37424 21604 37430 21616
rect 37936 21613 37964 21644
rect 38930 21632 38936 21684
rect 38988 21632 38994 21684
rect 41693 21675 41751 21681
rect 41693 21641 41705 21675
rect 41739 21672 41751 21675
rect 43530 21672 43536 21684
rect 41739 21644 43536 21672
rect 41739 21641 41751 21644
rect 41693 21635 41751 21641
rect 43530 21632 43536 21644
rect 43588 21632 43594 21684
rect 37921 21607 37979 21613
rect 37424 21576 37872 21604
rect 37424 21564 37430 21576
rect 34517 21539 34575 21545
rect 34517 21536 34529 21539
rect 34440 21508 34529 21536
rect 34333 21499 34391 21505
rect 34517 21505 34529 21508
rect 34563 21536 34575 21539
rect 35250 21536 35256 21548
rect 34563 21508 35256 21536
rect 34563 21505 34575 21508
rect 34517 21499 34575 21505
rect 32456 21440 32996 21468
rect 32456 21428 32462 21440
rect 33042 21428 33048 21480
rect 33100 21468 33106 21480
rect 33704 21468 33732 21499
rect 35250 21496 35256 21508
rect 35308 21496 35314 21548
rect 37458 21496 37464 21548
rect 37516 21536 37522 21548
rect 37553 21539 37611 21545
rect 37553 21536 37565 21539
rect 37516 21508 37565 21536
rect 37516 21496 37522 21508
rect 37553 21505 37565 21508
rect 37599 21505 37611 21539
rect 37844 21536 37872 21576
rect 37921 21573 37933 21607
rect 37967 21573 37979 21607
rect 37921 21567 37979 21573
rect 38102 21564 38108 21616
rect 38160 21604 38166 21616
rect 38473 21607 38531 21613
rect 38473 21604 38485 21607
rect 38160 21576 38485 21604
rect 38160 21564 38166 21576
rect 38473 21573 38485 21576
rect 38519 21573 38531 21607
rect 38473 21567 38531 21573
rect 40126 21564 40132 21616
rect 40184 21604 40190 21616
rect 40558 21607 40616 21613
rect 40558 21604 40570 21607
rect 40184 21576 40570 21604
rect 40184 21564 40190 21576
rect 40558 21573 40570 21576
rect 40604 21573 40616 21607
rect 40558 21567 40616 21573
rect 38197 21539 38255 21545
rect 37844 21508 38148 21536
rect 37553 21499 37611 21505
rect 33100 21440 33732 21468
rect 33100 21428 33106 21440
rect 35158 21428 35164 21480
rect 35216 21468 35222 21480
rect 35526 21468 35532 21480
rect 35216 21440 35532 21468
rect 35216 21428 35222 21440
rect 35526 21428 35532 21440
rect 35584 21428 35590 21480
rect 37369 21471 37427 21477
rect 37369 21437 37381 21471
rect 37415 21468 37427 21471
rect 37734 21468 37740 21480
rect 37415 21440 37740 21468
rect 37415 21437 37427 21440
rect 37369 21431 37427 21437
rect 37734 21428 37740 21440
rect 37792 21428 37798 21480
rect 38010 21428 38016 21480
rect 38068 21428 38074 21480
rect 38120 21468 38148 21508
rect 38197 21505 38209 21539
rect 38243 21536 38255 21539
rect 38286 21536 38292 21548
rect 38243 21508 38292 21536
rect 38243 21505 38255 21508
rect 38197 21499 38255 21505
rect 38286 21496 38292 21508
rect 38344 21496 38350 21548
rect 38746 21496 38752 21548
rect 38804 21496 38810 21548
rect 38838 21496 38844 21548
rect 38896 21536 38902 21548
rect 39025 21539 39083 21545
rect 39025 21536 39037 21539
rect 38896 21508 39037 21536
rect 38896 21496 38902 21508
rect 39025 21505 39037 21508
rect 39071 21505 39083 21539
rect 40402 21536 40408 21548
rect 39025 21499 39083 21505
rect 39224 21508 40408 21536
rect 38565 21471 38623 21477
rect 38565 21468 38577 21471
rect 38120 21440 38577 21468
rect 38565 21437 38577 21440
rect 38611 21437 38623 21471
rect 38565 21431 38623 21437
rect 39114 21428 39120 21480
rect 39172 21428 39178 21480
rect 31665 21403 31723 21409
rect 30576 21372 31333 21400
rect 30331 21304 30420 21332
rect 30331 21301 30343 21304
rect 30285 21295 30343 21301
rect 30466 21292 30472 21344
rect 30524 21332 30530 21344
rect 30576 21332 30604 21372
rect 30524 21304 30604 21332
rect 30524 21292 30530 21304
rect 31018 21292 31024 21344
rect 31076 21332 31082 21344
rect 31205 21335 31263 21341
rect 31205 21332 31217 21335
rect 31076 21304 31217 21332
rect 31076 21292 31082 21304
rect 31205 21301 31217 21304
rect 31251 21301 31263 21335
rect 31305 21332 31333 21372
rect 31665 21369 31677 21403
rect 31711 21400 31723 21403
rect 39224 21400 39252 21508
rect 40402 21496 40408 21508
rect 40460 21496 40466 21548
rect 42794 21496 42800 21548
rect 42852 21496 42858 21548
rect 43070 21496 43076 21548
rect 43128 21496 43134 21548
rect 44174 21496 44180 21548
rect 44232 21536 44238 21548
rect 44269 21539 44327 21545
rect 44269 21536 44281 21539
rect 44232 21508 44281 21536
rect 44232 21496 44238 21508
rect 44269 21505 44281 21508
rect 44315 21505 44327 21539
rect 44269 21499 44327 21505
rect 40310 21428 40316 21480
rect 40368 21428 40374 21480
rect 31711 21372 39252 21400
rect 31711 21369 31723 21372
rect 31665 21363 31723 21369
rect 41322 21360 41328 21412
rect 41380 21400 41386 21412
rect 42613 21403 42671 21409
rect 42613 21400 42625 21403
rect 41380 21372 42625 21400
rect 41380 21360 41386 21372
rect 42613 21369 42625 21372
rect 42659 21400 42671 21403
rect 43898 21400 43904 21412
rect 42659 21372 43904 21400
rect 42659 21369 42671 21372
rect 42613 21363 42671 21369
rect 43898 21360 43904 21372
rect 43956 21360 43962 21412
rect 32125 21335 32183 21341
rect 32125 21332 32137 21335
rect 31305 21304 32137 21332
rect 31205 21295 31263 21301
rect 32125 21301 32137 21304
rect 32171 21301 32183 21335
rect 32125 21295 32183 21301
rect 32306 21292 32312 21344
rect 32364 21332 32370 21344
rect 33042 21332 33048 21344
rect 32364 21304 33048 21332
rect 32364 21292 32370 21304
rect 33042 21292 33048 21304
rect 33100 21292 33106 21344
rect 33321 21335 33379 21341
rect 33321 21301 33333 21335
rect 33367 21332 33379 21335
rect 33686 21332 33692 21344
rect 33367 21304 33692 21332
rect 33367 21301 33379 21304
rect 33321 21295 33379 21301
rect 33686 21292 33692 21304
rect 33744 21332 33750 21344
rect 37366 21332 37372 21344
rect 33744 21304 37372 21332
rect 33744 21292 33750 21304
rect 37366 21292 37372 21304
rect 37424 21292 37430 21344
rect 37550 21292 37556 21344
rect 37608 21292 37614 21344
rect 37737 21335 37795 21341
rect 37737 21301 37749 21335
rect 37783 21332 37795 21335
rect 38102 21332 38108 21344
rect 37783 21304 38108 21332
rect 37783 21301 37795 21304
rect 37737 21295 37795 21301
rect 38102 21292 38108 21304
rect 38160 21292 38166 21344
rect 38197 21335 38255 21341
rect 38197 21301 38209 21335
rect 38243 21332 38255 21335
rect 38286 21332 38292 21344
rect 38243 21304 38292 21332
rect 38243 21301 38255 21304
rect 38197 21295 38255 21301
rect 38286 21292 38292 21304
rect 38344 21292 38350 21344
rect 38378 21292 38384 21344
rect 38436 21332 38442 21344
rect 38473 21335 38531 21341
rect 38473 21332 38485 21335
rect 38436 21304 38485 21332
rect 38436 21292 38442 21304
rect 38473 21301 38485 21304
rect 38519 21301 38531 21335
rect 38473 21295 38531 21301
rect 39022 21292 39028 21344
rect 39080 21292 39086 21344
rect 39390 21292 39396 21344
rect 39448 21292 39454 21344
rect 43625 21335 43683 21341
rect 43625 21301 43637 21335
rect 43671 21332 43683 21335
rect 43806 21332 43812 21344
rect 43671 21304 43812 21332
rect 43671 21301 43683 21304
rect 43625 21295 43683 21301
rect 43806 21292 43812 21304
rect 43864 21292 43870 21344
rect 44450 21292 44456 21344
rect 44508 21292 44514 21344
rect 1104 21242 44896 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 44896 21242
rect 1104 21168 44896 21190
rect 3970 21088 3976 21140
rect 4028 21128 4034 21140
rect 4614 21128 4620 21140
rect 4028 21100 4620 21128
rect 4028 21088 4034 21100
rect 4614 21088 4620 21100
rect 4672 21128 4678 21140
rect 5810 21128 5816 21140
rect 4672 21100 5816 21128
rect 4672 21088 4678 21100
rect 5810 21088 5816 21100
rect 5868 21088 5874 21140
rect 7190 21128 7196 21140
rect 7116 21100 7196 21128
rect 4341 21063 4399 21069
rect 4341 21029 4353 21063
rect 4387 21060 4399 21063
rect 7116 21060 7144 21100
rect 7190 21088 7196 21100
rect 7248 21128 7254 21140
rect 7377 21131 7435 21137
rect 7248 21100 7328 21128
rect 7248 21088 7254 21100
rect 4387 21032 7144 21060
rect 4387 21029 4399 21032
rect 4341 21023 4399 21029
rect 3050 20992 3056 21004
rect 2424 20964 3056 20992
rect 2130 20884 2136 20936
rect 2188 20884 2194 20936
rect 2424 20933 2452 20964
rect 3050 20952 3056 20964
rect 3108 20952 3114 21004
rect 7300 21001 7328 21100
rect 7377 21097 7389 21131
rect 7423 21128 7435 21131
rect 7834 21128 7840 21140
rect 7423 21100 7840 21128
rect 7423 21097 7435 21100
rect 7377 21091 7435 21097
rect 7834 21088 7840 21100
rect 7892 21088 7898 21140
rect 8757 21131 8815 21137
rect 8757 21097 8769 21131
rect 8803 21128 8815 21131
rect 8846 21128 8852 21140
rect 8803 21100 8852 21128
rect 8803 21097 8815 21100
rect 8757 21091 8815 21097
rect 8846 21088 8852 21100
rect 8904 21088 8910 21140
rect 9766 21088 9772 21140
rect 9824 21088 9830 21140
rect 11425 21131 11483 21137
rect 11425 21097 11437 21131
rect 11471 21128 11483 21131
rect 11514 21128 11520 21140
rect 11471 21100 11520 21128
rect 11471 21097 11483 21100
rect 11425 21091 11483 21097
rect 11514 21088 11520 21100
rect 11572 21088 11578 21140
rect 13078 21088 13084 21140
rect 13136 21088 13142 21140
rect 13262 21088 13268 21140
rect 13320 21128 13326 21140
rect 13320 21100 13400 21128
rect 13320 21088 13326 21100
rect 9490 21060 9496 21072
rect 8501 21032 9496 21060
rect 7285 20995 7343 21001
rect 7285 20961 7297 20995
rect 7331 20961 7343 20995
rect 7285 20955 7343 20961
rect 2409 20927 2467 20933
rect 2409 20893 2421 20927
rect 2455 20893 2467 20927
rect 2409 20887 2467 20893
rect 2501 20927 2559 20933
rect 2501 20893 2513 20927
rect 2547 20924 2559 20927
rect 2590 20924 2596 20936
rect 2547 20896 2596 20924
rect 2547 20893 2559 20896
rect 2501 20887 2559 20893
rect 2590 20884 2596 20896
rect 2648 20884 2654 20936
rect 3234 20884 3240 20936
rect 3292 20924 3298 20936
rect 3789 20927 3847 20933
rect 3789 20924 3801 20927
rect 3292 20896 3801 20924
rect 3292 20884 3298 20896
rect 3789 20893 3801 20896
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 3878 20884 3884 20936
rect 3936 20924 3942 20936
rect 3936 20896 4108 20924
rect 3936 20884 3942 20896
rect 2317 20859 2375 20865
rect 2317 20825 2329 20859
rect 2363 20856 2375 20859
rect 3970 20856 3976 20868
rect 2363 20828 3976 20856
rect 2363 20825 2375 20828
rect 2317 20819 2375 20825
rect 3970 20816 3976 20828
rect 4028 20816 4034 20868
rect 4080 20865 4108 20896
rect 4154 20884 4160 20936
rect 4212 20933 4218 20936
rect 4212 20927 4267 20933
rect 4212 20893 4221 20927
rect 4255 20924 4267 20927
rect 4890 20924 4896 20936
rect 4255 20896 4896 20924
rect 4255 20893 4267 20896
rect 4212 20887 4267 20893
rect 4212 20884 4218 20887
rect 4890 20884 4896 20896
rect 4948 20924 4954 20936
rect 5258 20924 5264 20936
rect 4948 20896 5264 20924
rect 4948 20884 4954 20896
rect 5258 20884 5264 20896
rect 5316 20884 5322 20936
rect 5626 20884 5632 20936
rect 5684 20924 5690 20936
rect 6454 20924 6460 20936
rect 5684 20896 6460 20924
rect 5684 20884 5690 20896
rect 6454 20884 6460 20896
rect 6512 20924 6518 20936
rect 7377 20927 7435 20933
rect 7377 20924 7389 20927
rect 6512 20896 7389 20924
rect 6512 20884 6518 20896
rect 7377 20893 7389 20896
rect 7423 20893 7435 20927
rect 7377 20887 7435 20893
rect 8202 20884 8208 20936
rect 8260 20884 8266 20936
rect 8389 20927 8447 20933
rect 8389 20893 8401 20927
rect 8435 20924 8447 20927
rect 8501 20924 8529 21032
rect 9490 21020 9496 21032
rect 9548 21020 9554 21072
rect 9600 21032 9996 21060
rect 9122 20952 9128 21004
rect 9180 20992 9186 21004
rect 9600 20992 9628 21032
rect 9968 21001 9996 21032
rect 10870 21020 10876 21072
rect 10928 21020 10934 21072
rect 12066 21060 12072 21072
rect 11900 21032 12072 21060
rect 9180 20964 9628 20992
rect 9953 20995 10011 21001
rect 9180 20952 9186 20964
rect 9953 20961 9965 20995
rect 9999 20961 10011 20995
rect 9953 20955 10011 20961
rect 10229 20995 10287 21001
rect 10229 20961 10241 20995
rect 10275 20992 10287 20995
rect 10318 20992 10324 21004
rect 10275 20964 10324 20992
rect 10275 20961 10287 20964
rect 10229 20955 10287 20961
rect 10318 20952 10324 20964
rect 10376 20952 10382 21004
rect 10888 20992 10916 21020
rect 10888 20964 11192 20992
rect 8435 20896 8529 20924
rect 8573 20927 8631 20933
rect 8435 20893 8447 20896
rect 8389 20887 8447 20893
rect 8573 20893 8585 20927
rect 8619 20924 8631 20927
rect 9217 20927 9275 20933
rect 9217 20924 9229 20927
rect 8619 20896 9229 20924
rect 8619 20893 8631 20896
rect 8573 20887 8631 20893
rect 9217 20893 9229 20896
rect 9263 20893 9275 20927
rect 9217 20887 9275 20893
rect 4065 20859 4123 20865
rect 4065 20825 4077 20859
rect 4111 20825 4123 20859
rect 4065 20819 4123 20825
rect 7101 20859 7159 20865
rect 7101 20825 7113 20859
rect 7147 20856 7159 20859
rect 7282 20856 7288 20868
rect 7147 20828 7288 20856
rect 7147 20825 7159 20828
rect 7101 20819 7159 20825
rect 2685 20791 2743 20797
rect 2685 20757 2697 20791
rect 2731 20788 2743 20791
rect 7116 20788 7144 20819
rect 7282 20816 7288 20828
rect 7340 20816 7346 20868
rect 8481 20859 8539 20865
rect 8481 20825 8493 20859
rect 8527 20856 8539 20859
rect 8846 20856 8852 20868
rect 8527 20828 8852 20856
rect 8527 20825 8539 20828
rect 8481 20819 8539 20825
rect 8846 20816 8852 20828
rect 8904 20816 8910 20868
rect 2731 20760 7144 20788
rect 7561 20791 7619 20797
rect 2731 20757 2743 20760
rect 2685 20751 2743 20757
rect 7561 20757 7573 20791
rect 7607 20788 7619 20791
rect 8202 20788 8208 20800
rect 7607 20760 8208 20788
rect 7607 20757 7619 20760
rect 7561 20751 7619 20757
rect 8202 20748 8208 20760
rect 8260 20748 8266 20800
rect 8938 20748 8944 20800
rect 8996 20788 9002 20800
rect 9232 20788 9260 20887
rect 9490 20884 9496 20936
rect 9548 20884 9554 20936
rect 9674 20933 9680 20936
rect 9637 20927 9680 20933
rect 9637 20893 9649 20927
rect 9637 20887 9680 20893
rect 9674 20884 9680 20887
rect 9732 20884 9738 20936
rect 9766 20884 9772 20936
rect 9824 20924 9830 20936
rect 10873 20927 10931 20933
rect 10873 20924 10885 20927
rect 9824 20896 10885 20924
rect 9824 20884 9830 20896
rect 10873 20893 10885 20896
rect 10919 20893 10931 20927
rect 10873 20887 10931 20893
rect 10962 20884 10968 20936
rect 11020 20924 11026 20936
rect 11164 20933 11192 20964
rect 11057 20927 11115 20933
rect 11057 20924 11069 20927
rect 11020 20896 11069 20924
rect 11020 20884 11026 20896
rect 11057 20893 11069 20896
rect 11103 20893 11115 20927
rect 11057 20887 11115 20893
rect 11149 20927 11207 20933
rect 11149 20893 11161 20927
rect 11195 20893 11207 20927
rect 11149 20887 11207 20893
rect 11293 20927 11351 20933
rect 11293 20893 11305 20927
rect 11339 20893 11351 20927
rect 11293 20887 11351 20893
rect 11793 20927 11851 20933
rect 11793 20893 11805 20927
rect 11839 20924 11851 20927
rect 11900 20924 11928 21032
rect 12066 21020 12072 21032
rect 12124 21020 12130 21072
rect 12250 21020 12256 21072
rect 12308 21020 12314 21072
rect 12345 21063 12403 21069
rect 12345 21029 12357 21063
rect 12391 21060 12403 21063
rect 12391 21032 12480 21060
rect 12391 21029 12403 21032
rect 12345 21023 12403 21029
rect 12268 20992 12296 21020
rect 12452 21004 12480 21032
rect 12802 21020 12808 21072
rect 12860 21020 12866 21072
rect 13372 21060 13400 21100
rect 13446 21088 13452 21140
rect 13504 21128 13510 21140
rect 13633 21131 13691 21137
rect 13633 21128 13645 21131
rect 13504 21100 13645 21128
rect 13504 21088 13510 21100
rect 13633 21097 13645 21100
rect 13679 21097 13691 21131
rect 13633 21091 13691 21097
rect 14642 21088 14648 21140
rect 14700 21128 14706 21140
rect 14737 21131 14795 21137
rect 14737 21128 14749 21131
rect 14700 21100 14749 21128
rect 14700 21088 14706 21100
rect 14737 21097 14749 21100
rect 14783 21128 14795 21131
rect 17126 21128 17132 21140
rect 14783 21100 17132 21128
rect 14783 21097 14795 21100
rect 14737 21091 14795 21097
rect 17126 21088 17132 21100
rect 17184 21128 17190 21140
rect 17405 21131 17463 21137
rect 17405 21128 17417 21131
rect 17184 21100 17417 21128
rect 17184 21088 17190 21100
rect 17405 21097 17417 21100
rect 17451 21097 17463 21131
rect 17405 21091 17463 21097
rect 18138 21088 18144 21140
rect 18196 21088 18202 21140
rect 19242 21088 19248 21140
rect 19300 21088 19306 21140
rect 19702 21088 19708 21140
rect 19760 21088 19766 21140
rect 20806 21088 20812 21140
rect 20864 21128 20870 21140
rect 20901 21131 20959 21137
rect 20901 21128 20913 21131
rect 20864 21100 20913 21128
rect 20864 21088 20870 21100
rect 20901 21097 20913 21100
rect 20947 21097 20959 21131
rect 21453 21131 21511 21137
rect 21453 21128 21465 21131
rect 20901 21091 20959 21097
rect 21008 21100 21465 21128
rect 14090 21060 14096 21072
rect 13372 21032 14096 21060
rect 14090 21020 14096 21032
rect 14148 21020 14154 21072
rect 15010 21020 15016 21072
rect 15068 21060 15074 21072
rect 15381 21063 15439 21069
rect 15381 21060 15393 21063
rect 15068 21032 15393 21060
rect 15068 21020 15074 21032
rect 15381 21029 15393 21032
rect 15427 21029 15439 21063
rect 15381 21023 15439 21029
rect 15470 21020 15476 21072
rect 15528 21060 15534 21072
rect 20824 21060 20852 21088
rect 15528 21032 20852 21060
rect 15528 21020 15534 21032
rect 11992 20964 12296 20992
rect 11992 20933 12020 20964
rect 12434 20952 12440 21004
rect 12492 20952 12498 21004
rect 12820 20992 12848 21020
rect 12544 20964 12848 20992
rect 12250 20933 12256 20936
rect 11839 20896 11928 20924
rect 11977 20927 12035 20933
rect 11839 20893 11851 20896
rect 11793 20887 11851 20893
rect 11977 20893 11989 20927
rect 12023 20893 12035 20927
rect 11977 20887 12035 20893
rect 12213 20927 12256 20933
rect 12213 20893 12225 20927
rect 12213 20887 12256 20893
rect 9398 20816 9404 20868
rect 9456 20856 9462 20868
rect 10410 20856 10416 20868
rect 9456 20828 10416 20856
rect 9456 20816 9462 20828
rect 10410 20816 10416 20828
rect 10468 20816 10474 20868
rect 10686 20816 10692 20868
rect 10744 20856 10750 20868
rect 11308 20856 11336 20887
rect 12250 20884 12256 20887
rect 12308 20884 12314 20936
rect 12544 20933 12572 20964
rect 13998 20952 14004 21004
rect 14056 20992 14062 21004
rect 14056 20964 14596 20992
rect 14056 20952 14062 20964
rect 12529 20927 12587 20933
rect 12529 20893 12541 20927
rect 12575 20893 12587 20927
rect 12529 20887 12587 20893
rect 12802 20884 12808 20936
rect 12860 20884 12866 20936
rect 12949 20927 13007 20933
rect 12949 20893 12961 20927
rect 12995 20902 13007 20927
rect 13354 20924 13360 20936
rect 13096 20902 13360 20924
rect 12995 20896 13360 20902
rect 12995 20893 13124 20896
rect 12949 20887 13124 20893
rect 12964 20874 13124 20887
rect 13354 20884 13360 20896
rect 13412 20884 13418 20936
rect 13538 20884 13544 20936
rect 13596 20884 13602 20936
rect 13814 20884 13820 20936
rect 13872 20924 13878 20936
rect 14093 20927 14151 20933
rect 14093 20924 14105 20927
rect 13872 20896 14105 20924
rect 13872 20884 13878 20896
rect 14093 20893 14105 20896
rect 14139 20893 14151 20927
rect 14093 20887 14151 20893
rect 14277 20927 14335 20933
rect 14277 20893 14289 20927
rect 14323 20924 14335 20927
rect 14458 20924 14464 20936
rect 14323 20896 14464 20924
rect 14323 20893 14335 20896
rect 14277 20887 14335 20893
rect 14458 20884 14464 20896
rect 14516 20884 14522 20936
rect 14568 20933 14596 20964
rect 18414 20952 18420 21004
rect 18472 20992 18478 21004
rect 19337 20995 19395 21001
rect 19337 20992 19349 20995
rect 18472 20964 19349 20992
rect 18472 20952 18478 20964
rect 19337 20961 19349 20964
rect 19383 20961 19395 20995
rect 19337 20955 19395 20961
rect 20898 20952 20904 21004
rect 20956 20992 20962 21004
rect 21008 21001 21036 21100
rect 21453 21097 21465 21100
rect 21499 21097 21511 21131
rect 21453 21091 21511 21097
rect 21821 21131 21879 21137
rect 21821 21097 21833 21131
rect 21867 21128 21879 21131
rect 24578 21128 24584 21140
rect 21867 21100 24584 21128
rect 21867 21097 21879 21100
rect 21821 21091 21879 21097
rect 24578 21088 24584 21100
rect 24636 21088 24642 21140
rect 24765 21131 24823 21137
rect 24765 21097 24777 21131
rect 24811 21128 24823 21131
rect 24854 21128 24860 21140
rect 24811 21100 24860 21128
rect 24811 21097 24823 21100
rect 24765 21091 24823 21097
rect 24854 21088 24860 21100
rect 24912 21088 24918 21140
rect 26970 21088 26976 21140
rect 27028 21088 27034 21140
rect 30558 21088 30564 21140
rect 30616 21128 30622 21140
rect 34054 21128 34060 21140
rect 30616 21100 34060 21128
rect 30616 21088 30622 21100
rect 34054 21088 34060 21100
rect 34112 21088 34118 21140
rect 34882 21088 34888 21140
rect 34940 21128 34946 21140
rect 34977 21131 35035 21137
rect 34977 21128 34989 21131
rect 34940 21100 34989 21128
rect 34940 21088 34946 21100
rect 34977 21097 34989 21100
rect 35023 21128 35035 21131
rect 35526 21128 35532 21140
rect 35023 21100 35532 21128
rect 35023 21097 35035 21100
rect 34977 21091 35035 21097
rect 35526 21088 35532 21100
rect 35584 21088 35590 21140
rect 35986 21088 35992 21140
rect 36044 21088 36050 21140
rect 36262 21088 36268 21140
rect 36320 21128 36326 21140
rect 36449 21131 36507 21137
rect 36449 21128 36461 21131
rect 36320 21100 36461 21128
rect 36320 21088 36326 21100
rect 36449 21097 36461 21100
rect 36495 21097 36507 21131
rect 36449 21091 36507 21097
rect 38378 21088 38384 21140
rect 38436 21088 38442 21140
rect 38565 21131 38623 21137
rect 38565 21097 38577 21131
rect 38611 21128 38623 21131
rect 38838 21128 38844 21140
rect 38611 21100 38844 21128
rect 38611 21097 38623 21100
rect 38565 21091 38623 21097
rect 38838 21088 38844 21100
rect 38896 21088 38902 21140
rect 39390 21088 39396 21140
rect 39448 21128 39454 21140
rect 39448 21100 43668 21128
rect 39448 21088 39454 21100
rect 21542 21020 21548 21072
rect 21600 21060 21606 21072
rect 33410 21060 33416 21072
rect 21600 21032 33416 21060
rect 21600 21020 21606 21032
rect 33410 21020 33416 21032
rect 33468 21020 33474 21072
rect 33962 21020 33968 21072
rect 34020 21060 34026 21072
rect 36354 21060 36360 21072
rect 34020 21032 36360 21060
rect 34020 21020 34026 21032
rect 36354 21020 36360 21032
rect 36412 21060 36418 21072
rect 37090 21060 37096 21072
rect 36412 21032 37096 21060
rect 36412 21020 36418 21032
rect 37090 21020 37096 21032
rect 37148 21020 37154 21072
rect 42521 21063 42579 21069
rect 42521 21029 42533 21063
rect 42567 21029 42579 21063
rect 42521 21023 42579 21029
rect 20993 20995 21051 21001
rect 20993 20992 21005 20995
rect 20956 20964 21005 20992
rect 20956 20952 20962 20964
rect 20993 20961 21005 20964
rect 21039 20961 21051 20995
rect 20993 20955 21051 20961
rect 21100 20964 21680 20992
rect 14553 20927 14611 20933
rect 14553 20893 14565 20927
rect 14599 20924 14611 20927
rect 14734 20924 14740 20936
rect 14599 20896 14740 20924
rect 14599 20893 14611 20896
rect 14553 20887 14611 20893
rect 14734 20884 14740 20896
rect 14792 20884 14798 20936
rect 14829 20927 14887 20933
rect 14829 20893 14841 20927
rect 14875 20893 14887 20927
rect 14829 20887 14887 20893
rect 15197 20927 15255 20933
rect 15197 20893 15209 20927
rect 15243 20924 15255 20927
rect 15286 20924 15292 20936
rect 15243 20896 15292 20924
rect 15243 20893 15255 20896
rect 15197 20887 15255 20893
rect 11882 20856 11888 20868
rect 10744 20828 11888 20856
rect 10744 20816 10750 20828
rect 11882 20816 11888 20828
rect 11940 20816 11946 20868
rect 12069 20859 12127 20865
rect 12069 20856 12081 20859
rect 11992 20828 12081 20856
rect 10704 20788 10732 20816
rect 11992 20800 12020 20828
rect 12069 20825 12081 20828
rect 12115 20825 12127 20859
rect 12069 20819 12127 20825
rect 12434 20816 12440 20868
rect 12492 20856 12498 20868
rect 12713 20859 12771 20865
rect 12713 20856 12725 20859
rect 12492 20828 12725 20856
rect 12492 20816 12498 20828
rect 12713 20825 12725 20828
rect 12759 20825 12771 20859
rect 12713 20819 12771 20825
rect 13170 20816 13176 20868
rect 13228 20856 13234 20868
rect 13265 20859 13323 20865
rect 13265 20856 13277 20859
rect 13228 20828 13277 20856
rect 13228 20816 13234 20828
rect 13265 20825 13277 20828
rect 13311 20825 13323 20859
rect 13265 20819 13323 20825
rect 13446 20816 13452 20868
rect 13504 20816 13510 20868
rect 13556 20856 13584 20884
rect 14844 20856 14872 20887
rect 15286 20884 15292 20896
rect 15344 20884 15350 20936
rect 17218 20884 17224 20936
rect 17276 20924 17282 20936
rect 17405 20927 17463 20933
rect 17405 20924 17417 20927
rect 17276 20896 17417 20924
rect 17276 20884 17282 20896
rect 17405 20893 17417 20896
rect 17451 20893 17463 20927
rect 17405 20887 17463 20893
rect 17586 20884 17592 20936
rect 17644 20884 17650 20936
rect 17678 20884 17684 20936
rect 17736 20884 17742 20936
rect 18233 20927 18291 20933
rect 18233 20893 18245 20927
rect 18279 20893 18291 20927
rect 18233 20887 18291 20893
rect 13556 20828 14872 20856
rect 15013 20859 15071 20865
rect 14108 20800 14136 20828
rect 15013 20825 15025 20859
rect 15059 20825 15071 20859
rect 15013 20819 15071 20825
rect 8996 20760 10732 20788
rect 8996 20748 9002 20760
rect 10962 20748 10968 20800
rect 11020 20788 11026 20800
rect 11422 20788 11428 20800
rect 11020 20760 11428 20788
rect 11020 20748 11026 20760
rect 11422 20748 11428 20760
rect 11480 20748 11486 20800
rect 11974 20748 11980 20800
rect 12032 20748 12038 20800
rect 12618 20748 12624 20800
rect 12676 20788 12682 20800
rect 13538 20788 13544 20800
rect 12676 20760 13544 20788
rect 12676 20748 12682 20760
rect 13538 20748 13544 20760
rect 13596 20748 13602 20800
rect 14090 20748 14096 20800
rect 14148 20748 14154 20800
rect 14826 20748 14832 20800
rect 14884 20788 14890 20800
rect 15028 20788 15056 20819
rect 15102 20816 15108 20868
rect 15160 20816 15166 20868
rect 18049 20859 18107 20865
rect 18049 20825 18061 20859
rect 18095 20825 18107 20859
rect 18248 20856 18276 20887
rect 18322 20884 18328 20936
rect 18380 20884 18386 20936
rect 19426 20884 19432 20936
rect 19484 20924 19490 20936
rect 19521 20927 19579 20933
rect 19521 20924 19533 20927
rect 19484 20896 19533 20924
rect 19484 20884 19490 20896
rect 19521 20893 19533 20896
rect 19567 20924 19579 20927
rect 21100 20924 21128 20964
rect 19567 20896 21128 20924
rect 19567 20893 19579 20896
rect 19521 20887 19579 20893
rect 21174 20884 21180 20936
rect 21232 20884 21238 20936
rect 21453 20927 21511 20933
rect 21453 20893 21465 20927
rect 21499 20893 21511 20927
rect 21453 20887 21511 20893
rect 18690 20856 18696 20868
rect 18248 20828 18696 20856
rect 18049 20819 18107 20825
rect 14884 20760 15056 20788
rect 17865 20791 17923 20797
rect 14884 20748 14890 20760
rect 17865 20757 17877 20791
rect 17911 20788 17923 20791
rect 18064 20788 18092 20819
rect 18340 20800 18368 20828
rect 18690 20816 18696 20828
rect 18748 20816 18754 20868
rect 19245 20859 19303 20865
rect 19245 20825 19257 20859
rect 19291 20825 19303 20859
rect 20622 20856 20628 20868
rect 19245 20819 19303 20825
rect 19536 20828 20628 20856
rect 17911 20760 18092 20788
rect 17911 20757 17923 20760
rect 17865 20751 17923 20757
rect 18322 20748 18328 20800
rect 18380 20748 18386 20800
rect 18509 20791 18567 20797
rect 18509 20757 18521 20791
rect 18555 20788 18567 20791
rect 19260 20788 19288 20819
rect 19536 20800 19564 20828
rect 20622 20816 20628 20828
rect 20680 20856 20686 20868
rect 20901 20859 20959 20865
rect 20901 20856 20913 20859
rect 20680 20828 20913 20856
rect 20680 20816 20686 20828
rect 20901 20825 20913 20828
rect 20947 20856 20959 20859
rect 21468 20856 21496 20887
rect 21542 20884 21548 20936
rect 21600 20884 21606 20936
rect 20947 20828 21496 20856
rect 21652 20856 21680 20964
rect 21726 20952 21732 21004
rect 21784 20992 21790 21004
rect 23106 20992 23112 21004
rect 21784 20964 23112 20992
rect 21784 20952 21790 20964
rect 23106 20952 23112 20964
rect 23164 20952 23170 21004
rect 24578 20952 24584 21004
rect 24636 20952 24642 21004
rect 24688 20964 24992 20992
rect 23290 20884 23296 20936
rect 23348 20884 23354 20936
rect 24394 20884 24400 20936
rect 24452 20924 24458 20936
rect 24489 20927 24547 20933
rect 24489 20924 24501 20927
rect 24452 20896 24501 20924
rect 24452 20884 24458 20896
rect 24489 20893 24501 20896
rect 24535 20893 24547 20927
rect 24489 20887 24547 20893
rect 23477 20859 23535 20865
rect 21652 20828 22094 20856
rect 20947 20825 20959 20828
rect 20901 20819 20959 20825
rect 18555 20760 19288 20788
rect 18555 20757 18567 20760
rect 18509 20751 18567 20757
rect 19518 20748 19524 20800
rect 19576 20748 19582 20800
rect 19886 20748 19892 20800
rect 19944 20788 19950 20800
rect 20806 20788 20812 20800
rect 19944 20760 20812 20788
rect 19944 20748 19950 20760
rect 20806 20748 20812 20760
rect 20864 20748 20870 20800
rect 21358 20748 21364 20800
rect 21416 20788 21422 20800
rect 21818 20788 21824 20800
rect 21416 20760 21824 20788
rect 21416 20748 21422 20760
rect 21818 20748 21824 20760
rect 21876 20748 21882 20800
rect 22066 20788 22094 20828
rect 23477 20825 23489 20859
rect 23523 20856 23535 20859
rect 23658 20856 23664 20868
rect 23523 20828 23664 20856
rect 23523 20825 23535 20828
rect 23477 20819 23535 20825
rect 23658 20816 23664 20828
rect 23716 20856 23722 20868
rect 24688 20856 24716 20964
rect 24765 20927 24823 20933
rect 24765 20893 24777 20927
rect 24811 20924 24823 20927
rect 24854 20924 24860 20936
rect 24811 20896 24860 20924
rect 24811 20893 24823 20896
rect 24765 20887 24823 20893
rect 23716 20828 24716 20856
rect 23716 20816 23722 20828
rect 24780 20788 24808 20887
rect 24854 20884 24860 20896
rect 24912 20884 24918 20936
rect 24964 20924 24992 20964
rect 25314 20952 25320 21004
rect 25372 20992 25378 21004
rect 25372 20964 26832 20992
rect 25372 20952 25378 20964
rect 24964 20896 26280 20924
rect 25314 20816 25320 20868
rect 25372 20856 25378 20868
rect 25774 20856 25780 20868
rect 25372 20828 25780 20856
rect 25372 20816 25378 20828
rect 25774 20816 25780 20828
rect 25832 20816 25838 20868
rect 22066 20760 24808 20788
rect 24949 20791 25007 20797
rect 24949 20757 24961 20791
rect 24995 20788 25007 20791
rect 25130 20788 25136 20800
rect 24995 20760 25136 20788
rect 24995 20757 25007 20760
rect 24949 20751 25007 20757
rect 25130 20748 25136 20760
rect 25188 20748 25194 20800
rect 26252 20788 26280 20896
rect 26326 20884 26332 20936
rect 26384 20884 26390 20936
rect 26804 20933 26832 20964
rect 30190 20952 30196 21004
rect 30248 20992 30254 21004
rect 33686 20992 33692 21004
rect 30248 20964 33692 20992
rect 30248 20952 30254 20964
rect 33686 20952 33692 20964
rect 33744 20952 33750 21004
rect 35161 20995 35219 21001
rect 35161 20961 35173 20995
rect 35207 20992 35219 20995
rect 35342 20992 35348 21004
rect 35207 20964 35348 20992
rect 35207 20961 35219 20964
rect 35161 20955 35219 20961
rect 35342 20952 35348 20964
rect 35400 20952 35406 21004
rect 40310 20952 40316 21004
rect 40368 20992 40374 21004
rect 41141 20995 41199 21001
rect 41141 20992 41153 20995
rect 40368 20964 41153 20992
rect 40368 20952 40374 20964
rect 41141 20961 41153 20964
rect 41187 20961 41199 20995
rect 41141 20955 41199 20961
rect 26789 20927 26847 20933
rect 26789 20893 26801 20927
rect 26835 20893 26847 20927
rect 26789 20887 26847 20893
rect 26973 20927 27031 20933
rect 26973 20893 26985 20927
rect 27019 20924 27031 20927
rect 27062 20924 27068 20936
rect 27019 20896 27068 20924
rect 27019 20893 27031 20896
rect 26973 20887 27031 20893
rect 27062 20884 27068 20896
rect 27120 20884 27126 20936
rect 27798 20884 27804 20936
rect 27856 20924 27862 20936
rect 30834 20924 30840 20936
rect 27856 20896 30840 20924
rect 27856 20884 27862 20896
rect 30834 20884 30840 20896
rect 30892 20884 30898 20936
rect 34606 20884 34612 20936
rect 34664 20924 34670 20936
rect 35253 20927 35311 20933
rect 35253 20924 35265 20927
rect 34664 20896 35265 20924
rect 34664 20884 34670 20896
rect 35253 20893 35265 20896
rect 35299 20893 35311 20927
rect 35253 20887 35311 20893
rect 36170 20884 36176 20936
rect 36228 20884 36234 20936
rect 36262 20884 36268 20936
rect 36320 20884 36326 20936
rect 38194 20884 38200 20936
rect 38252 20884 38258 20936
rect 38286 20884 38292 20936
rect 38344 20884 38350 20936
rect 42536 20924 42564 21023
rect 43346 21020 43352 21072
rect 43404 21020 43410 21072
rect 43254 20924 43260 20936
rect 42536 20896 43260 20924
rect 43254 20884 43260 20896
rect 43312 20884 43318 20936
rect 43640 20933 43668 21100
rect 43806 21088 43812 21140
rect 43864 21088 43870 21140
rect 43533 20927 43591 20933
rect 43533 20893 43545 20927
rect 43579 20893 43591 20927
rect 43533 20887 43591 20893
rect 43625 20927 43683 20933
rect 43625 20893 43637 20927
rect 43671 20893 43683 20927
rect 43625 20887 43683 20893
rect 26510 20816 26516 20868
rect 26568 20816 26574 20868
rect 26697 20859 26755 20865
rect 26697 20825 26709 20859
rect 26743 20856 26755 20859
rect 26743 20828 29684 20856
rect 26743 20825 26755 20828
rect 26697 20819 26755 20825
rect 27062 20788 27068 20800
rect 26252 20760 27068 20788
rect 27062 20748 27068 20760
rect 27120 20748 27126 20800
rect 27157 20791 27215 20797
rect 27157 20757 27169 20791
rect 27203 20788 27215 20791
rect 27614 20788 27620 20800
rect 27203 20760 27620 20788
rect 27203 20757 27215 20760
rect 27157 20751 27215 20757
rect 27614 20748 27620 20760
rect 27672 20748 27678 20800
rect 29656 20788 29684 20828
rect 29730 20816 29736 20868
rect 29788 20856 29794 20868
rect 34882 20856 34888 20868
rect 29788 20828 34888 20856
rect 29788 20816 29794 20828
rect 34882 20816 34888 20828
rect 34940 20816 34946 20868
rect 34977 20859 35035 20865
rect 34977 20825 34989 20859
rect 35023 20856 35035 20859
rect 35342 20856 35348 20868
rect 35023 20828 35348 20856
rect 35023 20825 35035 20828
rect 34977 20819 35035 20825
rect 35342 20816 35348 20828
rect 35400 20816 35406 20868
rect 35989 20859 36047 20865
rect 35989 20825 36001 20859
rect 36035 20825 36047 20859
rect 35989 20819 36047 20825
rect 41408 20859 41466 20865
rect 41408 20825 41420 20859
rect 41454 20856 41466 20859
rect 41598 20856 41604 20868
rect 41454 20828 41604 20856
rect 41454 20825 41466 20828
rect 41408 20819 41466 20825
rect 31018 20788 31024 20800
rect 29656 20760 31024 20788
rect 31018 20748 31024 20760
rect 31076 20748 31082 20800
rect 35437 20791 35495 20797
rect 35437 20757 35449 20791
rect 35483 20788 35495 20791
rect 36004 20788 36032 20819
rect 41598 20816 41604 20828
rect 41656 20816 41662 20868
rect 41782 20816 41788 20868
rect 41840 20856 41846 20868
rect 43548 20856 43576 20887
rect 43898 20884 43904 20936
rect 43956 20884 43962 20936
rect 44266 20884 44272 20936
rect 44324 20884 44330 20936
rect 41840 20828 43576 20856
rect 41840 20816 41846 20828
rect 35483 20760 36032 20788
rect 35483 20757 35495 20760
rect 35437 20751 35495 20757
rect 42610 20748 42616 20800
rect 42668 20748 42674 20800
rect 44082 20748 44088 20800
rect 44140 20788 44146 20800
rect 44453 20791 44511 20797
rect 44453 20788 44465 20791
rect 44140 20760 44465 20788
rect 44140 20748 44146 20760
rect 44453 20757 44465 20760
rect 44499 20757 44511 20791
rect 44453 20751 44511 20757
rect 1104 20698 44896 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 44896 20698
rect 1104 20624 44896 20646
rect 6086 20544 6092 20596
rect 6144 20544 6150 20596
rect 8570 20544 8576 20596
rect 8628 20584 8634 20596
rect 8628 20556 10272 20584
rect 8628 20544 8634 20556
rect 2682 20476 2688 20528
rect 2740 20516 2746 20528
rect 8478 20516 8484 20528
rect 2740 20488 8484 20516
rect 2740 20476 2746 20488
rect 8478 20476 8484 20488
rect 8536 20516 8542 20528
rect 9030 20516 9036 20528
rect 8536 20488 9036 20516
rect 8536 20476 8542 20488
rect 9030 20476 9036 20488
rect 9088 20476 9094 20528
rect 9493 20519 9551 20525
rect 9493 20485 9505 20519
rect 9539 20516 9551 20519
rect 9858 20516 9864 20528
rect 9539 20488 9864 20516
rect 9539 20485 9551 20488
rect 9493 20479 9551 20485
rect 9858 20476 9864 20488
rect 9916 20516 9922 20528
rect 10137 20519 10195 20525
rect 10137 20516 10149 20519
rect 9916 20488 10149 20516
rect 9916 20476 9922 20488
rect 10137 20485 10149 20488
rect 10183 20485 10195 20519
rect 10244 20516 10272 20556
rect 11330 20544 11336 20596
rect 11388 20584 11394 20596
rect 12434 20584 12440 20596
rect 11388 20556 12440 20584
rect 11388 20544 11394 20556
rect 12434 20544 12440 20556
rect 12492 20544 12498 20596
rect 12914 20587 12972 20593
rect 12914 20553 12926 20587
rect 12960 20584 12972 20587
rect 13262 20584 13268 20596
rect 12960 20556 13268 20584
rect 12960 20553 12972 20556
rect 12914 20547 12972 20553
rect 13262 20544 13268 20556
rect 13320 20544 13326 20596
rect 13354 20544 13360 20596
rect 13412 20584 13418 20596
rect 14550 20584 14556 20596
rect 13412 20556 14556 20584
rect 13412 20544 13418 20556
rect 14550 20544 14556 20556
rect 14608 20544 14614 20596
rect 16022 20544 16028 20596
rect 16080 20584 16086 20596
rect 19518 20584 19524 20596
rect 16080 20556 19524 20584
rect 16080 20544 16086 20556
rect 19518 20544 19524 20556
rect 19576 20544 19582 20596
rect 19981 20587 20039 20593
rect 19981 20553 19993 20587
rect 20027 20553 20039 20587
rect 19981 20547 20039 20553
rect 10244 20488 10548 20516
rect 10137 20479 10195 20485
rect 3326 20408 3332 20460
rect 3384 20448 3390 20460
rect 3697 20451 3755 20457
rect 3697 20448 3709 20451
rect 3384 20420 3709 20448
rect 3384 20408 3390 20420
rect 3697 20417 3709 20420
rect 3743 20448 3755 20451
rect 4154 20448 4160 20460
rect 3743 20420 4160 20448
rect 3743 20417 3755 20420
rect 3697 20411 3755 20417
rect 4154 20408 4160 20420
rect 4212 20408 4218 20460
rect 5718 20408 5724 20460
rect 5776 20408 5782 20460
rect 5902 20408 5908 20460
rect 5960 20448 5966 20460
rect 7558 20448 7564 20460
rect 5960 20420 7564 20448
rect 5960 20408 5966 20420
rect 7558 20408 7564 20420
rect 7616 20408 7622 20460
rect 9309 20451 9367 20457
rect 9309 20417 9321 20451
rect 9355 20448 9367 20451
rect 9355 20420 9536 20448
rect 9355 20417 9367 20420
rect 9309 20411 9367 20417
rect 3418 20340 3424 20392
rect 3476 20340 3482 20392
rect 5994 20340 6000 20392
rect 6052 20380 6058 20392
rect 8110 20380 8116 20392
rect 6052 20352 8116 20380
rect 6052 20340 6058 20352
rect 8110 20340 8116 20352
rect 8168 20340 8174 20392
rect 9508 20312 9536 20420
rect 9582 20408 9588 20460
rect 9640 20408 9646 20460
rect 9677 20451 9735 20457
rect 9677 20417 9689 20451
rect 9723 20417 9735 20451
rect 9677 20411 9735 20417
rect 9692 20380 9720 20411
rect 9766 20408 9772 20460
rect 9824 20448 9830 20460
rect 9953 20451 10011 20457
rect 9953 20448 9965 20451
rect 9824 20420 9965 20448
rect 9824 20408 9830 20420
rect 9953 20417 9965 20420
rect 9999 20448 10011 20451
rect 10042 20448 10048 20460
rect 9999 20420 10048 20448
rect 9999 20417 10011 20420
rect 9953 20411 10011 20417
rect 10042 20408 10048 20420
rect 10100 20408 10106 20460
rect 10226 20408 10232 20460
rect 10284 20408 10290 20460
rect 10318 20408 10324 20460
rect 10376 20457 10382 20460
rect 10376 20448 10384 20457
rect 10376 20420 10421 20448
rect 10376 20411 10384 20420
rect 10376 20408 10382 20411
rect 10336 20380 10364 20408
rect 9692 20352 10364 20380
rect 10520 20380 10548 20488
rect 10962 20476 10968 20528
rect 11020 20516 11026 20528
rect 12529 20519 12587 20525
rect 12529 20516 12541 20519
rect 11020 20488 12541 20516
rect 11020 20476 11026 20488
rect 12529 20485 12541 20488
rect 12575 20485 12587 20519
rect 12529 20479 12587 20485
rect 12621 20519 12679 20525
rect 12621 20485 12633 20519
rect 12667 20516 12679 20519
rect 13170 20516 13176 20528
rect 12667 20488 13176 20516
rect 12667 20485 12679 20488
rect 12621 20479 12679 20485
rect 13170 20476 13176 20488
rect 13228 20476 13234 20528
rect 15381 20519 15439 20525
rect 15381 20516 15393 20519
rect 13464 20488 15393 20516
rect 11882 20408 11888 20460
rect 11940 20448 11946 20460
rect 12345 20451 12403 20457
rect 12345 20448 12357 20451
rect 11940 20420 12357 20448
rect 11940 20408 11946 20420
rect 12345 20417 12357 20420
rect 12391 20417 12403 20451
rect 12345 20411 12403 20417
rect 12718 20451 12776 20457
rect 12718 20417 12730 20451
rect 12764 20417 12776 20451
rect 12718 20411 12776 20417
rect 10520 20352 10640 20380
rect 9950 20312 9956 20324
rect 9508 20284 9956 20312
rect 9950 20272 9956 20284
rect 10008 20312 10014 20324
rect 10226 20312 10232 20324
rect 10008 20284 10232 20312
rect 10008 20272 10014 20284
rect 10226 20272 10232 20284
rect 10284 20272 10290 20324
rect 10502 20272 10508 20324
rect 10560 20272 10566 20324
rect 10612 20312 10640 20352
rect 10686 20340 10692 20392
rect 10744 20380 10750 20392
rect 12728 20380 12756 20411
rect 13078 20408 13084 20460
rect 13136 20448 13142 20460
rect 13464 20448 13492 20488
rect 15381 20485 15393 20488
rect 15427 20516 15439 20519
rect 15562 20516 15568 20528
rect 15427 20488 15568 20516
rect 15427 20485 15439 20488
rect 15381 20479 15439 20485
rect 15562 20476 15568 20488
rect 15620 20476 15626 20528
rect 18141 20519 18199 20525
rect 15672 20488 16252 20516
rect 15672 20460 15700 20488
rect 13136 20420 13492 20448
rect 13541 20451 13599 20457
rect 13136 20408 13142 20420
rect 13541 20417 13553 20451
rect 13587 20448 13599 20451
rect 13722 20448 13728 20460
rect 13587 20420 13728 20448
rect 13587 20417 13599 20420
rect 13541 20411 13599 20417
rect 13722 20408 13728 20420
rect 13780 20408 13786 20460
rect 13906 20408 13912 20460
rect 13964 20448 13970 20460
rect 14461 20451 14519 20457
rect 14461 20448 14473 20451
rect 13964 20420 14473 20448
rect 13964 20408 13970 20420
rect 14461 20417 14473 20420
rect 14507 20417 14519 20451
rect 14461 20411 14519 20417
rect 14734 20408 14740 20460
rect 14792 20408 14798 20460
rect 15654 20408 15660 20460
rect 15712 20408 15718 20460
rect 15838 20408 15844 20460
rect 15896 20448 15902 20460
rect 16224 20457 16252 20488
rect 18141 20485 18153 20519
rect 18187 20516 18199 20519
rect 18230 20516 18236 20528
rect 18187 20488 18236 20516
rect 18187 20485 18199 20488
rect 18141 20479 18199 20485
rect 18230 20476 18236 20488
rect 18288 20476 18294 20528
rect 19334 20476 19340 20528
rect 19392 20516 19398 20528
rect 19996 20516 20024 20547
rect 20530 20544 20536 20596
rect 20588 20584 20594 20596
rect 23106 20584 23112 20596
rect 20588 20556 23112 20584
rect 20588 20544 20594 20556
rect 23106 20544 23112 20556
rect 23164 20544 23170 20596
rect 23293 20587 23351 20593
rect 23293 20553 23305 20587
rect 23339 20584 23351 20587
rect 23658 20584 23664 20596
rect 23339 20556 23664 20584
rect 23339 20553 23351 20556
rect 23293 20547 23351 20553
rect 23658 20544 23664 20556
rect 23716 20544 23722 20596
rect 24210 20544 24216 20596
rect 24268 20544 24274 20596
rect 24854 20544 24860 20596
rect 24912 20584 24918 20596
rect 26510 20584 26516 20596
rect 24912 20556 26516 20584
rect 24912 20544 24918 20556
rect 26510 20544 26516 20556
rect 26568 20544 26574 20596
rect 26602 20544 26608 20596
rect 26660 20584 26666 20596
rect 27433 20587 27491 20593
rect 26660 20556 27292 20584
rect 26660 20544 26666 20556
rect 26973 20519 27031 20525
rect 26973 20516 26985 20519
rect 19392 20488 19840 20516
rect 19996 20488 26985 20516
rect 19392 20476 19398 20488
rect 16117 20451 16175 20457
rect 16117 20448 16129 20451
rect 15896 20420 16129 20448
rect 15896 20408 15902 20420
rect 16117 20417 16129 20420
rect 16163 20417 16175 20451
rect 16117 20411 16175 20417
rect 16209 20451 16267 20457
rect 16209 20417 16221 20451
rect 16255 20417 16267 20451
rect 16209 20411 16267 20417
rect 18414 20408 18420 20460
rect 18472 20408 18478 20460
rect 19521 20451 19579 20457
rect 19521 20417 19533 20451
rect 19567 20448 19579 20451
rect 19702 20448 19708 20460
rect 19567 20420 19708 20448
rect 19567 20417 19579 20420
rect 19521 20411 19579 20417
rect 19702 20408 19708 20420
rect 19760 20408 19766 20460
rect 19812 20457 19840 20488
rect 26973 20485 26985 20488
rect 27019 20485 27031 20519
rect 26973 20479 27031 20485
rect 19797 20451 19855 20457
rect 19797 20417 19809 20451
rect 19843 20448 19855 20451
rect 19886 20448 19892 20460
rect 19843 20420 19892 20448
rect 19843 20417 19855 20420
rect 19797 20411 19855 20417
rect 19886 20408 19892 20420
rect 19944 20408 19950 20460
rect 19978 20408 19984 20460
rect 20036 20408 20042 20460
rect 20898 20408 20904 20460
rect 20956 20448 20962 20460
rect 20993 20451 21051 20457
rect 20993 20448 21005 20451
rect 20956 20420 21005 20448
rect 20956 20408 20962 20420
rect 20993 20417 21005 20420
rect 21039 20417 21051 20451
rect 20993 20411 21051 20417
rect 21174 20408 21180 20460
rect 21232 20448 21238 20460
rect 21542 20448 21548 20460
rect 21232 20420 21548 20448
rect 21232 20408 21238 20420
rect 21542 20408 21548 20420
rect 21600 20408 21606 20460
rect 22094 20408 22100 20460
rect 22152 20448 22158 20460
rect 22646 20448 22652 20460
rect 22152 20420 22652 20448
rect 22152 20408 22158 20420
rect 22646 20408 22652 20420
rect 22704 20448 22710 20460
rect 22925 20451 22983 20457
rect 22925 20448 22937 20451
rect 22704 20420 22937 20448
rect 22704 20408 22710 20420
rect 22925 20417 22937 20420
rect 22971 20417 22983 20451
rect 22925 20411 22983 20417
rect 23109 20451 23167 20457
rect 23109 20417 23121 20451
rect 23155 20448 23167 20451
rect 23382 20448 23388 20460
rect 23155 20420 23388 20448
rect 23155 20417 23167 20420
rect 23109 20411 23167 20417
rect 23382 20408 23388 20420
rect 23440 20408 23446 20460
rect 23750 20408 23756 20460
rect 23808 20408 23814 20460
rect 24026 20408 24032 20460
rect 24084 20408 24090 20460
rect 25590 20408 25596 20460
rect 25648 20448 25654 20460
rect 25777 20451 25835 20457
rect 25777 20448 25789 20451
rect 25648 20420 25789 20448
rect 25648 20408 25654 20420
rect 25777 20417 25789 20420
rect 25823 20448 25835 20451
rect 25823 20420 26004 20448
rect 25823 20417 25835 20420
rect 25777 20411 25835 20417
rect 10744 20352 12756 20380
rect 13265 20383 13323 20389
rect 10744 20340 10750 20352
rect 13265 20349 13277 20383
rect 13311 20349 13323 20383
rect 13265 20343 13323 20349
rect 13280 20312 13308 20343
rect 13630 20340 13636 20392
rect 13688 20380 13694 20392
rect 14553 20383 14611 20389
rect 14553 20380 14565 20383
rect 13688 20352 14565 20380
rect 13688 20340 13694 20352
rect 14553 20349 14565 20352
rect 14599 20349 14611 20383
rect 14553 20343 14611 20349
rect 15470 20340 15476 20392
rect 15528 20380 15534 20392
rect 15528 20352 17264 20380
rect 15528 20340 15534 20352
rect 15841 20315 15899 20321
rect 10612 20284 13308 20312
rect 13372 20284 15424 20312
rect 5905 20247 5963 20253
rect 5905 20213 5917 20247
rect 5951 20244 5963 20247
rect 5994 20244 6000 20256
rect 5951 20216 6000 20244
rect 5951 20213 5963 20216
rect 5905 20207 5963 20213
rect 5994 20204 6000 20216
rect 6052 20204 6058 20256
rect 6546 20204 6552 20256
rect 6604 20244 6610 20256
rect 9766 20244 9772 20256
rect 6604 20216 9772 20244
rect 6604 20204 6610 20216
rect 9766 20204 9772 20216
rect 9824 20204 9830 20256
rect 9861 20247 9919 20253
rect 9861 20213 9873 20247
rect 9907 20244 9919 20247
rect 10778 20244 10784 20256
rect 9907 20216 10784 20244
rect 9907 20213 9919 20216
rect 9861 20207 9919 20213
rect 10778 20204 10784 20216
rect 10836 20244 10842 20256
rect 13372 20244 13400 20284
rect 10836 20216 13400 20244
rect 10836 20204 10842 20216
rect 14642 20204 14648 20256
rect 14700 20204 14706 20256
rect 14918 20204 14924 20256
rect 14976 20204 14982 20256
rect 15396 20253 15424 20284
rect 15841 20281 15853 20315
rect 15887 20312 15899 20315
rect 16485 20315 16543 20321
rect 15887 20284 16436 20312
rect 15887 20281 15899 20284
rect 15841 20275 15899 20281
rect 15381 20247 15439 20253
rect 15381 20213 15393 20247
rect 15427 20213 15439 20247
rect 15381 20207 15439 20213
rect 16298 20204 16304 20256
rect 16356 20204 16362 20256
rect 16408 20244 16436 20284
rect 16485 20281 16497 20315
rect 16531 20312 16543 20315
rect 16850 20312 16856 20324
rect 16531 20284 16856 20312
rect 16531 20281 16543 20284
rect 16485 20275 16543 20281
rect 16850 20272 16856 20284
rect 16908 20272 16914 20324
rect 17236 20312 17264 20352
rect 17494 20340 17500 20392
rect 17552 20380 17558 20392
rect 18233 20383 18291 20389
rect 18233 20380 18245 20383
rect 17552 20352 18245 20380
rect 17552 20340 17558 20352
rect 18233 20349 18245 20352
rect 18279 20349 18291 20383
rect 18233 20343 18291 20349
rect 18690 20340 18696 20392
rect 18748 20380 18754 20392
rect 18966 20380 18972 20392
rect 18748 20352 18972 20380
rect 18748 20340 18754 20352
rect 18966 20340 18972 20352
rect 19024 20340 19030 20392
rect 19613 20383 19671 20389
rect 19613 20349 19625 20383
rect 19659 20380 19671 20383
rect 19996 20380 20024 20408
rect 20346 20380 20352 20392
rect 19659 20352 20352 20380
rect 19659 20349 19671 20352
rect 19613 20343 19671 20349
rect 20346 20340 20352 20352
rect 20404 20340 20410 20392
rect 21358 20340 21364 20392
rect 21416 20380 21422 20392
rect 22002 20380 22008 20392
rect 21416 20352 22008 20380
rect 21416 20340 21422 20352
rect 22002 20340 22008 20352
rect 22060 20340 22066 20392
rect 23014 20340 23020 20392
rect 23072 20380 23078 20392
rect 23937 20383 23995 20389
rect 23937 20380 23949 20383
rect 23072 20352 23949 20380
rect 23072 20340 23078 20352
rect 23937 20349 23949 20352
rect 23983 20380 23995 20383
rect 24118 20380 24124 20392
rect 23983 20352 24124 20380
rect 23983 20349 23995 20352
rect 23937 20343 23995 20349
rect 24118 20340 24124 20352
rect 24176 20340 24182 20392
rect 25130 20340 25136 20392
rect 25188 20380 25194 20392
rect 25869 20383 25927 20389
rect 25869 20380 25881 20383
rect 25188 20352 25881 20380
rect 25188 20340 25194 20352
rect 25869 20349 25881 20352
rect 25915 20349 25927 20383
rect 25976 20380 26004 20420
rect 26050 20408 26056 20460
rect 26108 20408 26114 20460
rect 26326 20408 26332 20460
rect 26384 20408 26390 20460
rect 26605 20451 26663 20457
rect 26605 20417 26617 20451
rect 26651 20448 26663 20451
rect 26786 20448 26792 20460
rect 26651 20420 26792 20448
rect 26651 20417 26663 20420
rect 26605 20411 26663 20417
rect 26786 20408 26792 20420
rect 26844 20448 26850 20460
rect 27264 20457 27292 20556
rect 27433 20553 27445 20587
rect 27479 20584 27491 20587
rect 27479 20556 27568 20584
rect 27479 20553 27491 20556
rect 27433 20547 27491 20553
rect 27540 20525 27568 20556
rect 27982 20544 27988 20596
rect 28040 20544 28046 20596
rect 29086 20544 29092 20596
rect 29144 20584 29150 20596
rect 29365 20587 29423 20593
rect 29365 20584 29377 20587
rect 29144 20556 29377 20584
rect 29144 20544 29150 20556
rect 29365 20553 29377 20556
rect 29411 20553 29423 20587
rect 29365 20547 29423 20553
rect 29457 20587 29515 20593
rect 29457 20553 29469 20587
rect 29503 20584 29515 20587
rect 29503 20556 29960 20584
rect 29503 20553 29515 20556
rect 29457 20547 29515 20553
rect 27525 20519 27583 20525
rect 27525 20485 27537 20519
rect 27571 20485 27583 20519
rect 28718 20516 28724 20528
rect 27525 20479 27583 20485
rect 27632 20488 28724 20516
rect 27249 20451 27307 20457
rect 26844 20420 27200 20448
rect 26844 20408 26850 20420
rect 26142 20380 26148 20392
rect 25976 20352 26148 20380
rect 25869 20343 25927 20349
rect 26142 20340 26148 20352
rect 26200 20340 26206 20392
rect 26418 20340 26424 20392
rect 26476 20340 26482 20392
rect 27065 20383 27123 20389
rect 27065 20380 27077 20383
rect 26712 20352 27077 20380
rect 18601 20315 18659 20321
rect 17236 20284 18460 20312
rect 17770 20244 17776 20256
rect 16408 20216 17776 20244
rect 17770 20204 17776 20216
rect 17828 20204 17834 20256
rect 18432 20253 18460 20284
rect 18601 20281 18613 20315
rect 18647 20312 18659 20315
rect 19978 20312 19984 20324
rect 18647 20284 19984 20312
rect 18647 20281 18659 20284
rect 18601 20275 18659 20281
rect 19978 20272 19984 20284
rect 20036 20272 20042 20324
rect 21450 20312 21456 20324
rect 20916 20284 21456 20312
rect 18417 20247 18475 20253
rect 18417 20213 18429 20247
rect 18463 20244 18475 20247
rect 18506 20244 18512 20256
rect 18463 20216 18512 20244
rect 18463 20213 18475 20216
rect 18417 20207 18475 20213
rect 18506 20204 18512 20216
rect 18564 20204 18570 20256
rect 19610 20204 19616 20256
rect 19668 20244 19674 20256
rect 19797 20247 19855 20253
rect 19797 20244 19809 20247
rect 19668 20216 19809 20244
rect 19668 20204 19674 20216
rect 19797 20213 19809 20216
rect 19843 20244 19855 20247
rect 20916 20244 20944 20284
rect 21450 20272 21456 20284
rect 21508 20272 21514 20324
rect 22066 20284 23060 20312
rect 19843 20216 20944 20244
rect 19843 20213 19855 20216
rect 19797 20207 19855 20213
rect 20990 20204 20996 20256
rect 21048 20204 21054 20256
rect 21361 20247 21419 20253
rect 21361 20213 21373 20247
rect 21407 20244 21419 20247
rect 22066 20244 22094 20284
rect 21407 20216 22094 20244
rect 21407 20213 21419 20216
rect 21361 20207 21419 20213
rect 22646 20204 22652 20256
rect 22704 20244 22710 20256
rect 22741 20247 22799 20253
rect 22741 20244 22753 20247
rect 22704 20216 22753 20244
rect 22704 20204 22710 20216
rect 22741 20213 22753 20216
rect 22787 20213 22799 20247
rect 23032 20244 23060 20284
rect 23106 20272 23112 20324
rect 23164 20312 23170 20324
rect 24854 20312 24860 20324
rect 23164 20284 24860 20312
rect 23164 20272 23170 20284
rect 23658 20244 23664 20256
rect 23032 20216 23664 20244
rect 22741 20207 22799 20213
rect 23658 20204 23664 20216
rect 23716 20204 23722 20256
rect 23768 20253 23796 20284
rect 24854 20272 24860 20284
rect 24912 20272 24918 20324
rect 25038 20272 25044 20324
rect 25096 20312 25102 20324
rect 26237 20315 26295 20321
rect 25096 20284 26096 20312
rect 25096 20272 25102 20284
rect 26068 20256 26096 20284
rect 26237 20281 26249 20315
rect 26283 20312 26295 20315
rect 26712 20312 26740 20352
rect 27065 20349 27077 20352
rect 27111 20349 27123 20383
rect 27172 20380 27200 20420
rect 27249 20417 27261 20451
rect 27295 20417 27307 20451
rect 27632 20448 27660 20488
rect 28718 20476 28724 20488
rect 28776 20476 28782 20528
rect 29730 20516 29736 20528
rect 29012 20488 29736 20516
rect 29012 20460 29040 20488
rect 29730 20476 29736 20488
rect 29788 20516 29794 20528
rect 29932 20525 29960 20556
rect 33594 20544 33600 20596
rect 33652 20584 33658 20596
rect 33870 20584 33876 20596
rect 33652 20556 33876 20584
rect 33652 20544 33658 20556
rect 33870 20544 33876 20556
rect 33928 20544 33934 20596
rect 36170 20544 36176 20596
rect 36228 20584 36234 20596
rect 36541 20587 36599 20593
rect 36541 20584 36553 20587
rect 36228 20556 36553 20584
rect 36228 20544 36234 20556
rect 36541 20553 36553 20556
rect 36587 20553 36599 20587
rect 38286 20584 38292 20596
rect 36541 20547 36599 20553
rect 36648 20556 38292 20584
rect 29825 20519 29883 20525
rect 29825 20516 29837 20519
rect 29788 20488 29837 20516
rect 29788 20476 29794 20488
rect 29825 20485 29837 20488
rect 29871 20485 29883 20519
rect 29825 20479 29883 20485
rect 29917 20519 29975 20525
rect 29917 20485 29929 20519
rect 29963 20485 29975 20519
rect 29917 20479 29975 20485
rect 27249 20411 27307 20417
rect 27356 20420 27660 20448
rect 27801 20451 27859 20457
rect 27356 20380 27384 20420
rect 27801 20417 27813 20451
rect 27847 20417 27859 20451
rect 27801 20411 27859 20417
rect 27172 20352 27384 20380
rect 27617 20383 27675 20389
rect 27065 20343 27123 20349
rect 27617 20349 27629 20383
rect 27663 20349 27675 20383
rect 27816 20380 27844 20411
rect 28074 20408 28080 20460
rect 28132 20408 28138 20460
rect 28258 20408 28264 20460
rect 28316 20408 28322 20460
rect 28994 20408 29000 20460
rect 29052 20408 29058 20460
rect 29270 20408 29276 20460
rect 29328 20448 29334 20460
rect 29641 20451 29699 20457
rect 29641 20448 29653 20451
rect 29328 20420 29653 20448
rect 29328 20408 29334 20420
rect 29641 20417 29653 20420
rect 29687 20417 29699 20451
rect 29641 20411 29699 20417
rect 27816 20352 28488 20380
rect 27617 20343 27675 20349
rect 26283 20284 26740 20312
rect 26789 20315 26847 20321
rect 26283 20281 26295 20284
rect 26237 20275 26295 20281
rect 26789 20281 26801 20315
rect 26835 20312 26847 20315
rect 27632 20312 27660 20343
rect 28460 20321 28488 20352
rect 29086 20340 29092 20392
rect 29144 20340 29150 20392
rect 26835 20284 27660 20312
rect 28445 20315 28503 20321
rect 26835 20281 26847 20284
rect 26789 20275 26847 20281
rect 28445 20281 28457 20315
rect 28491 20312 28503 20315
rect 29730 20312 29736 20324
rect 28491 20284 29736 20312
rect 28491 20281 28503 20284
rect 28445 20275 28503 20281
rect 29730 20272 29736 20284
rect 29788 20272 29794 20324
rect 29932 20312 29960 20479
rect 30190 20476 30196 20528
rect 30248 20516 30254 20528
rect 32398 20516 32404 20528
rect 30248 20488 32404 20516
rect 30248 20476 30254 20488
rect 32398 20476 32404 20488
rect 32456 20476 32462 20528
rect 32674 20476 32680 20528
rect 32732 20516 32738 20528
rect 36648 20516 36676 20556
rect 38286 20544 38292 20556
rect 38344 20544 38350 20596
rect 38841 20587 38899 20593
rect 38841 20553 38853 20587
rect 38887 20584 38899 20587
rect 39114 20584 39120 20596
rect 38887 20556 39120 20584
rect 38887 20553 38899 20556
rect 38841 20547 38899 20553
rect 39114 20544 39120 20556
rect 39172 20544 39178 20596
rect 41598 20544 41604 20596
rect 41656 20544 41662 20596
rect 36814 20516 36820 20528
rect 32732 20488 36676 20516
rect 36747 20488 36820 20516
rect 32732 20476 32738 20488
rect 30101 20451 30159 20457
rect 30101 20417 30113 20451
rect 30147 20417 30159 20451
rect 30101 20411 30159 20417
rect 30006 20312 30012 20324
rect 29932 20284 30012 20312
rect 30006 20272 30012 20284
rect 30064 20272 30070 20324
rect 23753 20247 23811 20253
rect 23753 20213 23765 20247
rect 23799 20213 23811 20247
rect 23753 20207 23811 20213
rect 23842 20204 23848 20256
rect 23900 20244 23906 20256
rect 25777 20247 25835 20253
rect 25777 20244 25789 20247
rect 23900 20216 25789 20244
rect 23900 20204 23906 20216
rect 25777 20213 25789 20216
rect 25823 20244 25835 20247
rect 25958 20244 25964 20256
rect 25823 20216 25964 20244
rect 25823 20213 25835 20216
rect 25777 20207 25835 20213
rect 25958 20204 25964 20216
rect 26016 20204 26022 20256
rect 26050 20204 26056 20256
rect 26108 20244 26114 20256
rect 26329 20247 26387 20253
rect 26329 20244 26341 20247
rect 26108 20216 26341 20244
rect 26108 20204 26114 20216
rect 26329 20213 26341 20216
rect 26375 20213 26387 20247
rect 26329 20207 26387 20213
rect 26970 20204 26976 20256
rect 27028 20204 27034 20256
rect 27614 20204 27620 20256
rect 27672 20204 27678 20256
rect 28994 20204 29000 20256
rect 29052 20244 29058 20256
rect 29270 20244 29276 20256
rect 29052 20216 29276 20244
rect 29052 20204 29058 20216
rect 29270 20204 29276 20216
rect 29328 20204 29334 20256
rect 29362 20204 29368 20256
rect 29420 20244 29426 20256
rect 30116 20244 30144 20411
rect 34422 20408 34428 20460
rect 34480 20448 34486 20460
rect 36747 20457 36775 20488
rect 36814 20476 36820 20488
rect 36872 20476 36878 20528
rect 38381 20519 38439 20525
rect 38381 20485 38393 20519
rect 38427 20516 38439 20519
rect 38470 20516 38476 20528
rect 38427 20488 38476 20516
rect 38427 20485 38439 20488
rect 38381 20479 38439 20485
rect 38470 20476 38476 20488
rect 38528 20476 38534 20528
rect 40770 20476 40776 20528
rect 40828 20516 40834 20528
rect 40828 20488 42196 20516
rect 40828 20476 40834 20488
rect 34701 20451 34759 20457
rect 34701 20448 34713 20451
rect 34480 20420 34713 20448
rect 34480 20408 34486 20420
rect 34701 20417 34713 20420
rect 34747 20417 34759 20451
rect 34701 20411 34759 20417
rect 36725 20451 36783 20457
rect 36725 20417 36737 20451
rect 36771 20417 36783 20451
rect 37001 20451 37059 20457
rect 37001 20448 37013 20451
rect 36725 20411 36783 20417
rect 36832 20420 37013 20448
rect 34606 20340 34612 20392
rect 34664 20380 34670 20392
rect 34793 20383 34851 20389
rect 34793 20380 34805 20383
rect 34664 20352 34805 20380
rect 34664 20340 34670 20352
rect 34793 20349 34805 20352
rect 34839 20349 34851 20383
rect 34793 20343 34851 20349
rect 36170 20340 36176 20392
rect 36228 20380 36234 20392
rect 36832 20380 36860 20420
rect 37001 20417 37013 20420
rect 37047 20417 37059 20451
rect 37001 20411 37059 20417
rect 37090 20408 37096 20460
rect 37148 20448 37154 20460
rect 38657 20451 38715 20457
rect 38657 20448 38669 20451
rect 37148 20420 38669 20448
rect 37148 20408 37154 20420
rect 38657 20417 38669 20420
rect 38703 20417 38715 20451
rect 38657 20411 38715 20417
rect 41782 20408 41788 20460
rect 41840 20408 41846 20460
rect 41877 20451 41935 20457
rect 41877 20417 41889 20451
rect 41923 20448 41935 20451
rect 41966 20448 41972 20460
rect 41923 20420 41972 20448
rect 41923 20417 41935 20420
rect 41877 20411 41935 20417
rect 41966 20408 41972 20420
rect 42024 20408 42030 20460
rect 42168 20457 42196 20488
rect 42153 20451 42211 20457
rect 42153 20417 42165 20451
rect 42199 20417 42211 20451
rect 42153 20411 42211 20417
rect 36228 20352 36860 20380
rect 36228 20340 36234 20352
rect 36906 20340 36912 20392
rect 36964 20380 36970 20392
rect 37182 20380 37188 20392
rect 36964 20352 37188 20380
rect 36964 20340 36970 20352
rect 37182 20340 37188 20352
rect 37240 20340 37246 20392
rect 37918 20340 37924 20392
rect 37976 20380 37982 20392
rect 38473 20383 38531 20389
rect 38473 20380 38485 20383
rect 37976 20352 38485 20380
rect 37976 20340 37982 20352
rect 38473 20349 38485 20352
rect 38519 20349 38531 20383
rect 38473 20343 38531 20349
rect 42061 20383 42119 20389
rect 42061 20349 42073 20383
rect 42107 20380 42119 20383
rect 42610 20380 42616 20392
rect 42107 20352 42616 20380
rect 42107 20349 42119 20352
rect 42061 20343 42119 20349
rect 31846 20272 31852 20324
rect 31904 20312 31910 20324
rect 38488 20312 38516 20343
rect 42610 20340 42616 20352
rect 42668 20340 42674 20392
rect 38654 20312 38660 20324
rect 31904 20284 38424 20312
rect 38488 20284 38660 20312
rect 31904 20272 31910 20284
rect 29420 20216 30144 20244
rect 29420 20204 29426 20216
rect 30282 20204 30288 20256
rect 30340 20204 30346 20256
rect 30834 20204 30840 20256
rect 30892 20244 30898 20256
rect 31662 20244 31668 20256
rect 30892 20216 31668 20244
rect 30892 20204 30898 20216
rect 31662 20204 31668 20216
rect 31720 20204 31726 20256
rect 33870 20204 33876 20256
rect 33928 20244 33934 20256
rect 34701 20247 34759 20253
rect 34701 20244 34713 20247
rect 33928 20216 34713 20244
rect 33928 20204 33934 20216
rect 34701 20213 34713 20216
rect 34747 20213 34759 20247
rect 34701 20207 34759 20213
rect 34790 20204 34796 20256
rect 34848 20244 34854 20256
rect 35069 20247 35127 20253
rect 35069 20244 35081 20247
rect 34848 20216 35081 20244
rect 34848 20204 34854 20216
rect 35069 20213 35081 20216
rect 35115 20213 35127 20247
rect 35069 20207 35127 20213
rect 36354 20204 36360 20256
rect 36412 20244 36418 20256
rect 38396 20253 38424 20284
rect 38654 20272 38660 20284
rect 38712 20272 38718 20324
rect 36725 20247 36783 20253
rect 36725 20244 36737 20247
rect 36412 20216 36737 20244
rect 36412 20204 36418 20216
rect 36725 20213 36737 20216
rect 36771 20213 36783 20247
rect 36725 20207 36783 20213
rect 38381 20247 38439 20253
rect 38381 20213 38393 20247
rect 38427 20213 38439 20247
rect 38381 20207 38439 20213
rect 1104 20154 44896 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 44896 20154
rect 1104 20080 44896 20102
rect 5353 20043 5411 20049
rect 5353 20009 5365 20043
rect 5399 20040 5411 20043
rect 5902 20040 5908 20052
rect 5399 20012 5908 20040
rect 5399 20009 5411 20012
rect 5353 20003 5411 20009
rect 5902 20000 5908 20012
rect 5960 20000 5966 20052
rect 9214 20000 9220 20052
rect 9272 20040 9278 20052
rect 9398 20040 9404 20052
rect 9272 20012 9404 20040
rect 9272 20000 9278 20012
rect 9398 20000 9404 20012
rect 9456 20040 9462 20052
rect 9493 20043 9551 20049
rect 9493 20040 9505 20043
rect 9456 20012 9505 20040
rect 9456 20000 9462 20012
rect 9493 20009 9505 20012
rect 9539 20009 9551 20043
rect 9493 20003 9551 20009
rect 10226 20000 10232 20052
rect 10284 20040 10290 20052
rect 12710 20040 12716 20052
rect 10284 20012 12716 20040
rect 10284 20000 10290 20012
rect 12710 20000 12716 20012
rect 12768 20000 12774 20052
rect 13354 20040 13360 20052
rect 13004 20012 13360 20040
rect 3513 19975 3571 19981
rect 3513 19941 3525 19975
rect 3559 19972 3571 19975
rect 5718 19972 5724 19984
rect 3559 19944 5724 19972
rect 3559 19941 3571 19944
rect 3513 19935 3571 19941
rect 5718 19932 5724 19944
rect 5776 19932 5782 19984
rect 7392 19944 9536 19972
rect 3878 19904 3884 19916
rect 2976 19876 3884 19904
rect 2976 19845 3004 19876
rect 3878 19864 3884 19876
rect 3936 19864 3942 19916
rect 6549 19907 6607 19913
rect 6549 19873 6561 19907
rect 6595 19904 6607 19907
rect 6638 19904 6644 19916
rect 6595 19876 6644 19904
rect 6595 19873 6607 19876
rect 6549 19867 6607 19873
rect 6638 19864 6644 19876
rect 6696 19864 6702 19916
rect 6730 19864 6736 19916
rect 6788 19864 6794 19916
rect 2961 19839 3019 19845
rect 2961 19805 2973 19839
rect 3007 19805 3019 19839
rect 2961 19799 3019 19805
rect 3326 19796 3332 19848
rect 3384 19796 3390 19848
rect 4798 19796 4804 19848
rect 4856 19796 4862 19848
rect 5258 19845 5264 19848
rect 5221 19839 5264 19845
rect 5221 19805 5233 19839
rect 5221 19799 5264 19805
rect 5258 19796 5264 19799
rect 5316 19796 5322 19848
rect 6362 19796 6368 19848
rect 6420 19836 6426 19848
rect 6457 19839 6515 19845
rect 6457 19836 6469 19839
rect 6420 19808 6469 19836
rect 6420 19796 6426 19808
rect 6457 19805 6469 19808
rect 6503 19805 6515 19839
rect 6457 19799 6515 19805
rect 6825 19839 6883 19845
rect 6825 19805 6837 19839
rect 6871 19836 6883 19839
rect 7392 19836 7420 19944
rect 7466 19864 7472 19916
rect 7524 19864 7530 19916
rect 8294 19864 8300 19916
rect 8352 19904 8358 19916
rect 8846 19904 8852 19916
rect 8352 19876 8852 19904
rect 8352 19864 8358 19876
rect 8846 19864 8852 19876
rect 8904 19904 8910 19916
rect 8904 19876 9352 19904
rect 8904 19864 8910 19876
rect 8205 19839 8263 19845
rect 8205 19836 8217 19839
rect 6871 19808 7420 19836
rect 7484 19808 8217 19836
rect 6871 19805 6883 19808
rect 6825 19799 6883 19805
rect 3145 19771 3203 19777
rect 3145 19737 3157 19771
rect 3191 19737 3203 19771
rect 3145 19731 3203 19737
rect 2406 19660 2412 19712
rect 2464 19700 2470 19712
rect 3160 19700 3188 19731
rect 3234 19728 3240 19780
rect 3292 19728 3298 19780
rect 4062 19728 4068 19780
rect 4120 19768 4126 19780
rect 4614 19768 4620 19780
rect 4120 19740 4620 19768
rect 4120 19728 4126 19740
rect 4614 19728 4620 19740
rect 4672 19768 4678 19780
rect 4985 19771 5043 19777
rect 4985 19768 4997 19771
rect 4672 19740 4997 19768
rect 4672 19728 4678 19740
rect 4985 19737 4997 19740
rect 5031 19737 5043 19771
rect 4985 19731 5043 19737
rect 5077 19771 5135 19777
rect 5077 19737 5089 19771
rect 5123 19768 5135 19771
rect 5350 19768 5356 19780
rect 5123 19740 5356 19768
rect 5123 19737 5135 19740
rect 5077 19731 5135 19737
rect 5350 19728 5356 19740
rect 5408 19728 5414 19780
rect 6546 19728 6552 19780
rect 6604 19768 6610 19780
rect 6840 19768 6868 19799
rect 7484 19780 7512 19808
rect 8205 19805 8217 19808
rect 8251 19805 8263 19839
rect 8205 19799 8263 19805
rect 8478 19796 8484 19848
rect 8536 19836 8542 19848
rect 8573 19839 8631 19845
rect 8573 19836 8585 19839
rect 8536 19808 8585 19836
rect 8536 19796 8542 19808
rect 8573 19805 8585 19808
rect 8619 19805 8631 19839
rect 8573 19799 8631 19805
rect 8757 19839 8815 19845
rect 8757 19805 8769 19839
rect 8803 19805 8815 19839
rect 8757 19799 8815 19805
rect 6604 19740 6868 19768
rect 6604 19728 6610 19740
rect 7466 19728 7472 19780
rect 7524 19728 7530 19780
rect 8772 19768 8800 19799
rect 8938 19796 8944 19848
rect 8996 19796 9002 19848
rect 9030 19796 9036 19848
rect 9088 19836 9094 19848
rect 9324 19845 9352 19876
rect 9508 19848 9536 19944
rect 10870 19932 10876 19984
rect 10928 19972 10934 19984
rect 13004 19972 13032 20012
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 13449 20043 13507 20049
rect 13449 20009 13461 20043
rect 13495 20040 13507 20043
rect 13630 20040 13636 20052
rect 13495 20012 13636 20040
rect 13495 20009 13507 20012
rect 13449 20003 13507 20009
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 14553 20043 14611 20049
rect 14553 20009 14565 20043
rect 14599 20040 14611 20043
rect 14734 20040 14740 20052
rect 14599 20012 14740 20040
rect 14599 20009 14611 20012
rect 14553 20003 14611 20009
rect 14734 20000 14740 20012
rect 14792 20000 14798 20052
rect 15378 20000 15384 20052
rect 15436 20040 15442 20052
rect 15657 20043 15715 20049
rect 15657 20040 15669 20043
rect 15436 20012 15669 20040
rect 15436 20000 15442 20012
rect 15657 20009 15669 20012
rect 15703 20009 15715 20043
rect 15657 20003 15715 20009
rect 16022 20000 16028 20052
rect 16080 20000 16086 20052
rect 16482 20000 16488 20052
rect 16540 20040 16546 20052
rect 18325 20043 18383 20049
rect 18325 20040 18337 20043
rect 16540 20012 18337 20040
rect 16540 20000 16546 20012
rect 18325 20009 18337 20012
rect 18371 20040 18383 20043
rect 18966 20040 18972 20052
rect 18371 20012 18972 20040
rect 18371 20009 18383 20012
rect 18325 20003 18383 20009
rect 18966 20000 18972 20012
rect 19024 20000 19030 20052
rect 23569 20043 23627 20049
rect 23569 20009 23581 20043
rect 23615 20040 23627 20043
rect 23842 20040 23848 20052
rect 23615 20012 23848 20040
rect 23615 20009 23627 20012
rect 23569 20003 23627 20009
rect 23842 20000 23848 20012
rect 23900 20040 23906 20052
rect 24302 20040 24308 20052
rect 23900 20012 24308 20040
rect 23900 20000 23906 20012
rect 24302 20000 24308 20012
rect 24360 20000 24366 20052
rect 25498 20000 25504 20052
rect 25556 20000 25562 20052
rect 25590 20000 25596 20052
rect 25648 20040 25654 20052
rect 25866 20040 25872 20052
rect 25648 20012 25872 20040
rect 25648 20000 25654 20012
rect 25866 20000 25872 20012
rect 25924 20000 25930 20052
rect 25961 20043 26019 20049
rect 25961 20009 25973 20043
rect 26007 20040 26019 20043
rect 26326 20040 26332 20052
rect 26007 20012 26332 20040
rect 26007 20009 26019 20012
rect 25961 20003 26019 20009
rect 26326 20000 26332 20012
rect 26384 20000 26390 20052
rect 26510 20000 26516 20052
rect 26568 20000 26574 20052
rect 28810 20000 28816 20052
rect 28868 20040 28874 20052
rect 30009 20043 30067 20049
rect 28868 20012 29960 20040
rect 28868 20000 28874 20012
rect 10928 19944 13032 19972
rect 10928 19932 10934 19944
rect 13078 19932 13084 19984
rect 13136 19972 13142 19984
rect 13722 19972 13728 19984
rect 13136 19944 13728 19972
rect 13136 19932 13142 19944
rect 13722 19932 13728 19944
rect 13780 19932 13786 19984
rect 13814 19932 13820 19984
rect 13872 19972 13878 19984
rect 14369 19975 14427 19981
rect 14369 19972 14381 19975
rect 13872 19944 14381 19972
rect 13872 19932 13878 19944
rect 14369 19941 14381 19944
rect 14415 19941 14427 19975
rect 14369 19935 14427 19941
rect 18506 19932 18512 19984
rect 18564 19972 18570 19984
rect 24765 19975 24823 19981
rect 18564 19944 24440 19972
rect 18564 19932 18570 19944
rect 9766 19864 9772 19916
rect 9824 19904 9830 19916
rect 11514 19904 11520 19916
rect 9824 19876 11520 19904
rect 9824 19864 9830 19876
rect 11514 19864 11520 19876
rect 11572 19864 11578 19916
rect 14458 19904 14464 19916
rect 12912 19876 14464 19904
rect 9125 19839 9183 19845
rect 9125 19836 9137 19839
rect 9088 19808 9137 19836
rect 9088 19796 9094 19808
rect 9125 19805 9137 19808
rect 9171 19805 9183 19839
rect 9125 19799 9183 19805
rect 9314 19839 9372 19845
rect 9314 19805 9326 19839
rect 9360 19805 9372 19839
rect 9314 19799 9372 19805
rect 9490 19796 9496 19848
rect 9548 19836 9554 19848
rect 10410 19836 10416 19848
rect 9548 19808 10416 19836
rect 9548 19796 9554 19808
rect 10410 19796 10416 19808
rect 10468 19836 10474 19848
rect 10962 19836 10968 19848
rect 10468 19808 10968 19836
rect 10468 19796 10474 19808
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 12158 19796 12164 19848
rect 12216 19836 12222 19848
rect 12912 19845 12940 19876
rect 14458 19864 14464 19876
rect 14516 19864 14522 19916
rect 14550 19864 14556 19916
rect 14608 19904 14614 19916
rect 15102 19904 15108 19916
rect 14608 19876 15108 19904
rect 14608 19864 14614 19876
rect 15102 19864 15108 19876
rect 15160 19864 15166 19916
rect 15562 19864 15568 19916
rect 15620 19904 15626 19916
rect 19610 19904 19616 19916
rect 15620 19876 18460 19904
rect 15620 19864 15626 19876
rect 12897 19839 12955 19845
rect 12897 19836 12909 19839
rect 12216 19808 12909 19836
rect 12216 19796 12222 19808
rect 12897 19805 12909 19808
rect 12943 19805 12955 19839
rect 12897 19799 12955 19805
rect 13078 19796 13084 19848
rect 13136 19796 13142 19848
rect 13317 19839 13375 19845
rect 13317 19805 13329 19839
rect 13363 19836 13375 19839
rect 15194 19836 15200 19848
rect 13363 19808 15200 19836
rect 13363 19805 13375 19808
rect 13317 19799 13375 19805
rect 15194 19796 15200 19808
rect 15252 19796 15258 19848
rect 15930 19796 15936 19848
rect 15988 19796 15994 19848
rect 16025 19839 16083 19845
rect 16025 19805 16037 19839
rect 16071 19836 16083 19839
rect 16482 19836 16488 19848
rect 16071 19808 16488 19836
rect 16071 19805 16083 19808
rect 16025 19799 16083 19805
rect 16482 19796 16488 19808
rect 16540 19796 16546 19848
rect 18046 19796 18052 19848
rect 18104 19796 18110 19848
rect 18230 19796 18236 19848
rect 18288 19796 18294 19848
rect 18325 19839 18383 19845
rect 18325 19805 18337 19839
rect 18371 19805 18383 19839
rect 18325 19799 18383 19805
rect 9217 19771 9275 19777
rect 9217 19768 9229 19771
rect 8220 19740 9229 19768
rect 4080 19700 4108 19728
rect 8220 19712 8248 19740
rect 9217 19737 9229 19740
rect 9263 19768 9275 19771
rect 9398 19768 9404 19780
rect 9263 19740 9404 19768
rect 9263 19737 9275 19740
rect 9217 19731 9275 19737
rect 9398 19728 9404 19740
rect 9456 19728 9462 19780
rect 13173 19771 13231 19777
rect 13173 19737 13185 19771
rect 13219 19768 13231 19771
rect 13814 19768 13820 19780
rect 13219 19740 13820 19768
rect 13219 19737 13231 19740
rect 13173 19731 13231 19737
rect 13814 19728 13820 19740
rect 13872 19728 13878 19780
rect 14093 19771 14151 19777
rect 14093 19737 14105 19771
rect 14139 19768 14151 19771
rect 15010 19768 15016 19780
rect 14139 19740 15016 19768
rect 14139 19737 14151 19740
rect 14093 19731 14151 19737
rect 15010 19728 15016 19740
rect 15068 19728 15074 19780
rect 15838 19728 15844 19780
rect 15896 19768 15902 19780
rect 16390 19768 16396 19780
rect 15896 19740 16396 19768
rect 15896 19728 15902 19740
rect 16390 19728 16396 19740
rect 16448 19728 16454 19780
rect 2464 19672 4108 19700
rect 2464 19660 2470 19672
rect 8202 19660 8208 19712
rect 8260 19660 8266 19712
rect 8294 19660 8300 19712
rect 8352 19660 8358 19712
rect 8386 19660 8392 19712
rect 8444 19700 8450 19712
rect 15654 19700 15660 19712
rect 8444 19672 15660 19700
rect 8444 19660 8450 19672
rect 15654 19660 15660 19672
rect 15712 19660 15718 19712
rect 17862 19660 17868 19712
rect 17920 19700 17926 19712
rect 18340 19700 18368 19799
rect 18432 19768 18460 19876
rect 19306 19876 19616 19904
rect 18506 19796 18512 19848
rect 18564 19836 18570 19848
rect 19306 19836 19334 19876
rect 19610 19864 19616 19876
rect 19668 19864 19674 19916
rect 19794 19864 19800 19916
rect 19852 19904 19858 19916
rect 20070 19904 20076 19916
rect 19852 19876 20076 19904
rect 19852 19864 19858 19876
rect 20070 19864 20076 19876
rect 20128 19864 20134 19916
rect 23385 19907 23443 19913
rect 23385 19873 23397 19907
rect 23431 19904 23443 19907
rect 24118 19904 24124 19916
rect 23431 19876 24124 19904
rect 23431 19873 23443 19876
rect 23385 19867 23443 19873
rect 24118 19864 24124 19876
rect 24176 19864 24182 19916
rect 18564 19808 19334 19836
rect 23201 19839 23259 19845
rect 18564 19796 18570 19808
rect 23201 19805 23213 19839
rect 23247 19836 23259 19839
rect 23474 19836 23480 19848
rect 23247 19808 23480 19836
rect 23247 19805 23259 19808
rect 23201 19799 23259 19805
rect 23474 19796 23480 19808
rect 23532 19796 23538 19848
rect 23566 19796 23572 19848
rect 23624 19796 23630 19848
rect 23750 19796 23756 19848
rect 23808 19796 23814 19848
rect 24412 19845 24440 19944
rect 24765 19941 24777 19975
rect 24811 19972 24823 19975
rect 25406 19972 25412 19984
rect 24811 19944 25412 19972
rect 24811 19941 24823 19944
rect 24765 19935 24823 19941
rect 25406 19932 25412 19944
rect 25464 19932 25470 19984
rect 29549 19975 29607 19981
rect 29549 19972 29561 19975
rect 25608 19944 29561 19972
rect 24578 19864 24584 19916
rect 24636 19904 24642 19916
rect 25608 19904 25636 19944
rect 29549 19941 29561 19944
rect 29595 19941 29607 19975
rect 29549 19935 29607 19941
rect 24636 19876 25636 19904
rect 24636 19864 24642 19876
rect 25682 19864 25688 19916
rect 25740 19864 25746 19916
rect 26418 19864 26424 19916
rect 26476 19904 26482 19916
rect 26605 19907 26663 19913
rect 26605 19904 26617 19907
rect 26476 19876 26617 19904
rect 26476 19864 26482 19876
rect 26605 19873 26617 19876
rect 26651 19873 26663 19907
rect 27246 19904 27252 19916
rect 26605 19867 26663 19873
rect 26712 19876 27252 19904
rect 24397 19839 24455 19845
rect 24397 19805 24409 19839
rect 24443 19805 24455 19839
rect 24397 19799 24455 19805
rect 25501 19839 25559 19845
rect 25501 19805 25513 19839
rect 25547 19836 25559 19839
rect 25590 19836 25596 19848
rect 25547 19808 25596 19836
rect 25547 19805 25559 19808
rect 25501 19799 25559 19805
rect 25590 19796 25596 19808
rect 25648 19796 25654 19848
rect 25774 19796 25780 19848
rect 25832 19796 25838 19848
rect 26513 19839 26571 19845
rect 26513 19805 26525 19839
rect 26559 19836 26571 19839
rect 26712 19836 26740 19876
rect 27246 19864 27252 19876
rect 27304 19904 27310 19916
rect 29362 19904 29368 19916
rect 27304 19876 29368 19904
rect 27304 19864 27310 19876
rect 29362 19864 29368 19876
rect 29420 19864 29426 19916
rect 29822 19864 29828 19916
rect 29880 19864 29886 19916
rect 29932 19904 29960 20012
rect 30009 20009 30021 20043
rect 30055 20009 30067 20043
rect 30009 20003 30067 20009
rect 30024 19972 30052 20003
rect 30558 20000 30564 20052
rect 30616 20040 30622 20052
rect 31297 20043 31355 20049
rect 31297 20040 31309 20043
rect 30616 20012 31309 20040
rect 30616 20000 30622 20012
rect 31297 20009 31309 20012
rect 31343 20009 31355 20043
rect 31297 20003 31355 20009
rect 31386 20000 31392 20052
rect 31444 20040 31450 20052
rect 32309 20043 32367 20049
rect 32309 20040 32321 20043
rect 31444 20012 32321 20040
rect 31444 20000 31450 20012
rect 32309 20009 32321 20012
rect 32355 20009 32367 20043
rect 32309 20003 32367 20009
rect 33594 20000 33600 20052
rect 33652 20000 33658 20052
rect 33870 20000 33876 20052
rect 33928 20040 33934 20052
rect 33965 20043 34023 20049
rect 33965 20040 33977 20043
rect 33928 20012 33977 20040
rect 33928 20000 33934 20012
rect 33965 20009 33977 20012
rect 34011 20040 34023 20043
rect 35434 20040 35440 20052
rect 34011 20012 35440 20040
rect 34011 20009 34023 20012
rect 33965 20003 34023 20009
rect 35434 20000 35440 20012
rect 35492 20000 35498 20052
rect 35526 20000 35532 20052
rect 35584 20000 35590 20052
rect 36998 20000 37004 20052
rect 37056 20040 37062 20052
rect 37093 20043 37151 20049
rect 37093 20040 37105 20043
rect 37056 20012 37105 20040
rect 37056 20000 37062 20012
rect 37093 20009 37105 20012
rect 37139 20040 37151 20043
rect 37182 20040 37188 20052
rect 37139 20012 37188 20040
rect 37139 20009 37151 20012
rect 37093 20003 37151 20009
rect 37182 20000 37188 20012
rect 37240 20000 37246 20052
rect 30282 19972 30288 19984
rect 30024 19944 30288 19972
rect 30282 19932 30288 19944
rect 30340 19972 30346 19984
rect 30340 19944 37136 19972
rect 30340 19932 30346 19944
rect 31570 19904 31576 19916
rect 29932 19876 31576 19904
rect 26559 19808 26740 19836
rect 26559 19805 26571 19808
rect 26513 19799 26571 19805
rect 26786 19796 26792 19848
rect 26844 19796 26850 19848
rect 28902 19796 28908 19848
rect 28960 19836 28966 19848
rect 31312 19845 31340 19876
rect 31570 19864 31576 19876
rect 31628 19864 31634 19916
rect 32214 19864 32220 19916
rect 32272 19904 32278 19916
rect 32401 19907 32459 19913
rect 32401 19904 32413 19907
rect 32272 19876 32413 19904
rect 32272 19864 32278 19876
rect 32401 19873 32413 19876
rect 32447 19873 32459 19907
rect 32674 19904 32680 19916
rect 32401 19867 32459 19873
rect 32508 19876 32680 19904
rect 29733 19839 29791 19845
rect 29733 19836 29745 19839
rect 28960 19808 29745 19836
rect 28960 19796 28966 19808
rect 29733 19805 29745 19808
rect 29779 19805 29791 19839
rect 29733 19799 29791 19805
rect 31297 19839 31355 19845
rect 31297 19805 31309 19839
rect 31343 19805 31355 19839
rect 31297 19799 31355 19805
rect 31389 19839 31447 19845
rect 31389 19805 31401 19839
rect 31435 19805 31447 19839
rect 32309 19839 32367 19845
rect 32309 19836 32321 19839
rect 31389 19799 31447 19805
rect 31680 19808 32321 19836
rect 22094 19768 22100 19780
rect 18432 19740 22100 19768
rect 22094 19728 22100 19740
rect 22152 19728 22158 19780
rect 22186 19728 22192 19780
rect 22244 19768 22250 19780
rect 22833 19771 22891 19777
rect 22833 19768 22845 19771
rect 22244 19740 22845 19768
rect 22244 19728 22250 19740
rect 22833 19737 22845 19740
rect 22879 19737 22891 19771
rect 22833 19731 22891 19737
rect 23017 19771 23075 19777
rect 23017 19737 23029 19771
rect 23063 19768 23075 19771
rect 23106 19768 23112 19780
rect 23063 19740 23112 19768
rect 23063 19737 23075 19740
rect 23017 19731 23075 19737
rect 17920 19672 18368 19700
rect 18509 19703 18567 19709
rect 17920 19660 17926 19672
rect 18509 19669 18521 19703
rect 18555 19700 18567 19703
rect 19150 19700 19156 19712
rect 18555 19672 19156 19700
rect 18555 19669 18567 19672
rect 18509 19663 18567 19669
rect 19150 19660 19156 19672
rect 19208 19660 19214 19712
rect 20990 19660 20996 19712
rect 21048 19700 21054 19712
rect 22002 19700 22008 19712
rect 21048 19672 22008 19700
rect 21048 19660 21054 19672
rect 22002 19660 22008 19672
rect 22060 19700 22066 19712
rect 23032 19700 23060 19731
rect 23106 19728 23112 19740
rect 23164 19728 23170 19780
rect 23293 19771 23351 19777
rect 23293 19737 23305 19771
rect 23339 19768 23351 19771
rect 23382 19768 23388 19780
rect 23339 19740 23388 19768
rect 23339 19737 23351 19740
rect 23293 19731 23351 19737
rect 23382 19728 23388 19740
rect 23440 19728 23446 19780
rect 23768 19709 23796 19796
rect 24578 19728 24584 19780
rect 24636 19728 24642 19780
rect 28994 19728 29000 19780
rect 29052 19728 29058 19780
rect 29086 19728 29092 19780
rect 29144 19768 29150 19780
rect 29181 19771 29239 19777
rect 29181 19768 29193 19771
rect 29144 19740 29193 19768
rect 29144 19728 29150 19740
rect 29181 19737 29193 19740
rect 29227 19737 29239 19771
rect 29181 19731 29239 19737
rect 30006 19728 30012 19780
rect 30064 19728 30070 19780
rect 30466 19728 30472 19780
rect 30524 19768 30530 19780
rect 31404 19768 31432 19799
rect 30524 19740 31432 19768
rect 30524 19728 30530 19740
rect 22060 19672 23060 19700
rect 23753 19703 23811 19709
rect 22060 19660 22066 19672
rect 23753 19669 23765 19703
rect 23799 19669 23811 19703
rect 23753 19663 23811 19669
rect 26326 19660 26332 19712
rect 26384 19660 26390 19712
rect 26510 19660 26516 19712
rect 26568 19700 26574 19712
rect 30190 19700 30196 19712
rect 26568 19672 30196 19700
rect 26568 19660 26574 19672
rect 30190 19660 30196 19672
rect 30248 19660 30254 19712
rect 31680 19709 31708 19808
rect 32309 19805 32321 19808
rect 32355 19836 32367 19839
rect 32508 19836 32536 19876
rect 32674 19864 32680 19876
rect 32732 19864 32738 19916
rect 34054 19864 34060 19916
rect 34112 19864 34118 19916
rect 34514 19904 34520 19916
rect 34164 19876 34520 19904
rect 32355 19808 32536 19836
rect 32585 19839 32643 19845
rect 32355 19805 32367 19808
rect 32309 19799 32367 19805
rect 32585 19805 32597 19839
rect 32631 19836 32643 19839
rect 33134 19836 33140 19848
rect 32631 19808 33140 19836
rect 32631 19805 32643 19808
rect 32585 19799 32643 19805
rect 33134 19796 33140 19808
rect 33192 19836 33198 19848
rect 33410 19836 33416 19848
rect 33192 19808 33416 19836
rect 33192 19796 33198 19808
rect 33410 19796 33416 19808
rect 33468 19796 33474 19848
rect 33502 19796 33508 19848
rect 33560 19796 33566 19848
rect 33597 19839 33655 19845
rect 33597 19805 33609 19839
rect 33643 19836 33655 19839
rect 34164 19836 34192 19876
rect 34514 19864 34520 19876
rect 34572 19864 34578 19916
rect 34606 19864 34612 19916
rect 34664 19904 34670 19916
rect 35529 19907 35587 19913
rect 35529 19904 35541 19907
rect 34664 19876 35541 19904
rect 34664 19864 34670 19876
rect 35529 19873 35541 19876
rect 35575 19873 35587 19907
rect 35529 19867 35587 19873
rect 33643 19808 34192 19836
rect 34241 19839 34299 19845
rect 33643 19805 33655 19808
rect 33597 19799 33655 19805
rect 34241 19805 34253 19839
rect 34287 19836 34299 19839
rect 34422 19836 34428 19848
rect 34287 19808 34428 19836
rect 34287 19805 34299 19808
rect 34241 19799 34299 19805
rect 34422 19796 34428 19808
rect 34480 19796 34486 19848
rect 35434 19796 35440 19848
rect 35492 19796 35498 19848
rect 37108 19845 37136 19944
rect 37185 19907 37243 19913
rect 37185 19873 37197 19907
rect 37231 19904 37243 19907
rect 38746 19904 38752 19916
rect 37231 19876 38752 19904
rect 37231 19873 37243 19876
rect 37185 19867 37243 19873
rect 37093 19839 37151 19845
rect 37093 19805 37105 19839
rect 37139 19805 37151 19839
rect 37093 19799 37151 19805
rect 32214 19728 32220 19780
rect 32272 19768 32278 19780
rect 32272 19740 32904 19768
rect 32272 19728 32278 19740
rect 31665 19703 31723 19709
rect 31665 19669 31677 19703
rect 31711 19669 31723 19703
rect 31665 19663 31723 19669
rect 32766 19660 32772 19712
rect 32824 19660 32830 19712
rect 32876 19700 32904 19740
rect 32950 19728 32956 19780
rect 33008 19768 33014 19780
rect 33321 19771 33379 19777
rect 33321 19768 33333 19771
rect 33008 19740 33333 19768
rect 33008 19728 33014 19740
rect 33321 19737 33333 19740
rect 33367 19737 33379 19771
rect 33321 19731 33379 19737
rect 33962 19728 33968 19780
rect 34020 19728 34026 19780
rect 34440 19768 34468 19796
rect 35526 19768 35532 19780
rect 34440 19740 35532 19768
rect 35526 19728 35532 19740
rect 35584 19728 35590 19780
rect 33042 19700 33048 19712
rect 32876 19672 33048 19700
rect 33042 19660 33048 19672
rect 33100 19660 33106 19712
rect 33781 19703 33839 19709
rect 33781 19669 33793 19703
rect 33827 19700 33839 19703
rect 34054 19700 34060 19712
rect 33827 19672 34060 19700
rect 33827 19669 33839 19672
rect 33781 19663 33839 19669
rect 34054 19660 34060 19672
rect 34112 19660 34118 19712
rect 34238 19660 34244 19712
rect 34296 19700 34302 19712
rect 34425 19703 34483 19709
rect 34425 19700 34437 19703
rect 34296 19672 34437 19700
rect 34296 19660 34302 19672
rect 34425 19669 34437 19672
rect 34471 19669 34483 19703
rect 34425 19663 34483 19669
rect 35805 19703 35863 19709
rect 35805 19669 35817 19703
rect 35851 19700 35863 19703
rect 37200 19700 37228 19867
rect 38746 19864 38752 19876
rect 38804 19864 38810 19916
rect 44174 19904 44180 19916
rect 41386 19876 44180 19904
rect 39666 19796 39672 19848
rect 39724 19796 39730 19848
rect 40770 19796 40776 19848
rect 40828 19836 40834 19848
rect 41386 19836 41414 19876
rect 44174 19864 44180 19876
rect 44232 19864 44238 19916
rect 40828 19808 41414 19836
rect 40828 19796 40834 19808
rect 43254 19796 43260 19848
rect 43312 19836 43318 19848
rect 44269 19839 44327 19845
rect 44269 19836 44281 19839
rect 43312 19808 44281 19836
rect 43312 19796 43318 19808
rect 44269 19805 44281 19808
rect 44315 19805 44327 19839
rect 44269 19799 44327 19805
rect 35851 19672 37228 19700
rect 35851 19669 35863 19672
rect 35805 19663 35863 19669
rect 37458 19660 37464 19712
rect 37516 19660 37522 19712
rect 38381 19703 38439 19709
rect 38381 19669 38393 19703
rect 38427 19700 38439 19703
rect 38562 19700 38568 19712
rect 38427 19672 38568 19700
rect 38427 19669 38439 19672
rect 38381 19663 38439 19669
rect 38562 19660 38568 19672
rect 38620 19660 38626 19712
rect 40221 19703 40279 19709
rect 40221 19669 40233 19703
rect 40267 19700 40279 19703
rect 40402 19700 40408 19712
rect 40267 19672 40408 19700
rect 40267 19669 40279 19672
rect 40221 19663 40279 19669
rect 40402 19660 40408 19672
rect 40460 19660 40466 19712
rect 44450 19660 44456 19712
rect 44508 19660 44514 19712
rect 1104 19610 44896 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 44896 19610
rect 1104 19536 44896 19558
rect 2682 19456 2688 19508
rect 2740 19496 2746 19508
rect 6917 19499 6975 19505
rect 2740 19468 2820 19496
rect 2740 19456 2746 19468
rect 2406 19388 2412 19440
rect 2464 19388 2470 19440
rect 2501 19431 2559 19437
rect 2501 19397 2513 19431
rect 2547 19428 2559 19431
rect 2792 19428 2820 19468
rect 6917 19465 6929 19499
rect 6963 19496 6975 19499
rect 8386 19496 8392 19508
rect 6963 19468 8392 19496
rect 6963 19465 6975 19468
rect 6917 19459 6975 19465
rect 8386 19456 8392 19468
rect 8444 19456 8450 19508
rect 8757 19499 8815 19505
rect 8757 19465 8769 19499
rect 8803 19496 8815 19499
rect 8938 19496 8944 19508
rect 8803 19468 8944 19496
rect 8803 19465 8815 19468
rect 8757 19459 8815 19465
rect 8938 19456 8944 19468
rect 8996 19456 9002 19508
rect 9766 19456 9772 19508
rect 9824 19496 9830 19508
rect 10686 19496 10692 19508
rect 9824 19468 10692 19496
rect 9824 19456 9830 19468
rect 10686 19456 10692 19468
rect 10744 19456 10750 19508
rect 12158 19456 12164 19508
rect 12216 19496 12222 19508
rect 12434 19496 12440 19508
rect 12216 19468 12440 19496
rect 12216 19456 12222 19468
rect 12434 19456 12440 19468
rect 12492 19496 12498 19508
rect 12621 19499 12679 19505
rect 12621 19496 12633 19499
rect 12492 19468 12633 19496
rect 12492 19456 12498 19468
rect 12621 19465 12633 19468
rect 12667 19465 12679 19499
rect 12621 19459 12679 19465
rect 12802 19456 12808 19508
rect 12860 19496 12866 19508
rect 18414 19496 18420 19508
rect 12860 19468 18420 19496
rect 12860 19456 12866 19468
rect 2961 19431 3019 19437
rect 2961 19428 2973 19431
rect 2547 19400 2973 19428
rect 2547 19397 2559 19400
rect 2501 19391 2559 19397
rect 2961 19397 2973 19400
rect 3007 19397 3019 19431
rect 2961 19391 3019 19397
rect 6178 19388 6184 19440
rect 6236 19428 6242 19440
rect 6641 19431 6699 19437
rect 6641 19428 6653 19431
rect 6236 19400 6653 19428
rect 6236 19388 6242 19400
rect 6641 19397 6653 19400
rect 6687 19397 6699 19431
rect 6641 19391 6699 19397
rect 8018 19388 8024 19440
rect 8076 19428 8082 19440
rect 12529 19431 12587 19437
rect 12529 19428 12541 19431
rect 8076 19400 12541 19428
rect 8076 19388 8082 19400
rect 12529 19397 12541 19400
rect 12575 19397 12587 19431
rect 13265 19431 13323 19437
rect 13265 19428 13277 19431
rect 12529 19391 12587 19397
rect 12636 19400 13277 19428
rect 2225 19363 2283 19369
rect 2225 19360 2237 19363
rect 2203 19332 2237 19360
rect 2225 19329 2237 19332
rect 2271 19329 2283 19363
rect 2225 19323 2283 19329
rect 2240 19292 2268 19323
rect 2590 19320 2596 19372
rect 2648 19369 2654 19372
rect 2648 19360 2656 19369
rect 2648 19332 2693 19360
rect 2648 19323 2656 19332
rect 2648 19320 2654 19323
rect 2774 19320 2780 19372
rect 2832 19369 2838 19372
rect 2832 19363 2852 19369
rect 2840 19329 2852 19363
rect 2832 19323 2852 19329
rect 2832 19320 2838 19323
rect 3142 19320 3148 19372
rect 3200 19360 3206 19372
rect 3329 19363 3387 19369
rect 3329 19360 3341 19363
rect 3200 19332 3341 19360
rect 3200 19320 3206 19332
rect 3329 19329 3341 19332
rect 3375 19329 3387 19363
rect 3329 19323 3387 19329
rect 6365 19363 6423 19369
rect 6365 19329 6377 19363
rect 6411 19360 6423 19363
rect 6454 19360 6460 19372
rect 6411 19332 6460 19360
rect 6411 19329 6423 19332
rect 6365 19323 6423 19329
rect 6454 19320 6460 19332
rect 6512 19320 6518 19372
rect 6546 19320 6552 19372
rect 6604 19320 6610 19372
rect 6730 19320 6736 19372
rect 6788 19320 6794 19372
rect 8570 19320 8576 19372
rect 8628 19320 8634 19372
rect 10134 19320 10140 19372
rect 10192 19360 10198 19372
rect 10229 19363 10287 19369
rect 10229 19360 10241 19363
rect 10192 19332 10241 19360
rect 10192 19320 10198 19332
rect 10229 19329 10241 19332
rect 10275 19329 10287 19363
rect 10229 19323 10287 19329
rect 10410 19320 10416 19372
rect 10468 19320 10474 19372
rect 10686 19369 10692 19372
rect 10505 19363 10563 19369
rect 10505 19329 10517 19363
rect 10551 19329 10563 19363
rect 10505 19323 10563 19329
rect 10649 19363 10692 19369
rect 10649 19329 10661 19363
rect 10649 19323 10692 19329
rect 2498 19292 2504 19304
rect 2240 19264 2504 19292
rect 2498 19252 2504 19264
rect 2556 19252 2562 19304
rect 8478 19252 8484 19304
rect 8536 19292 8542 19304
rect 9306 19292 9312 19304
rect 8536 19264 9312 19292
rect 8536 19252 8542 19264
rect 9306 19252 9312 19264
rect 9364 19292 9370 19304
rect 9674 19292 9680 19304
rect 9364 19264 9680 19292
rect 9364 19252 9370 19264
rect 9674 19252 9680 19264
rect 9732 19292 9738 19304
rect 10520 19292 10548 19323
rect 10686 19320 10692 19323
rect 10744 19320 10750 19372
rect 10870 19360 10876 19372
rect 10796 19332 10876 19360
rect 9732 19264 10548 19292
rect 9732 19252 9738 19264
rect 3602 19184 3608 19236
rect 3660 19224 3666 19236
rect 5994 19224 6000 19236
rect 3660 19196 6000 19224
rect 3660 19184 3666 19196
rect 5994 19184 6000 19196
rect 6052 19184 6058 19236
rect 6086 19184 6092 19236
rect 6144 19224 6150 19236
rect 6638 19224 6644 19236
rect 6144 19196 6644 19224
rect 6144 19184 6150 19196
rect 6638 19184 6644 19196
rect 6696 19184 6702 19236
rect 10796 19233 10824 19332
rect 10870 19320 10876 19332
rect 10928 19320 10934 19372
rect 12066 19320 12072 19372
rect 12124 19360 12130 19372
rect 12124 19332 12480 19360
rect 12124 19320 12130 19332
rect 12452 19292 12480 19332
rect 12636 19292 12664 19400
rect 13265 19397 13277 19400
rect 13311 19397 13323 19431
rect 13265 19391 13323 19397
rect 13650 19431 13708 19437
rect 13650 19397 13662 19431
rect 13696 19428 13708 19431
rect 14366 19428 14372 19440
rect 13696 19400 14372 19428
rect 13696 19397 13708 19400
rect 13650 19391 13708 19397
rect 14366 19388 14372 19400
rect 14424 19388 14430 19440
rect 14642 19388 14648 19440
rect 14700 19428 14706 19440
rect 15672 19437 15700 19468
rect 18414 19456 18420 19468
rect 18472 19456 18478 19508
rect 19061 19499 19119 19505
rect 19061 19465 19073 19499
rect 19107 19465 19119 19499
rect 19061 19459 19119 19465
rect 19153 19499 19211 19505
rect 19153 19465 19165 19499
rect 19199 19496 19211 19499
rect 19242 19496 19248 19508
rect 19199 19468 19248 19496
rect 19199 19465 19211 19468
rect 19153 19459 19211 19465
rect 15013 19431 15071 19437
rect 15013 19428 15025 19431
rect 14700 19400 15025 19428
rect 14700 19388 14706 19400
rect 15013 19397 15025 19400
rect 15059 19397 15071 19431
rect 15013 19391 15071 19397
rect 15306 19431 15364 19437
rect 15306 19397 15318 19431
rect 15352 19428 15364 19431
rect 15657 19431 15715 19437
rect 15352 19400 15608 19428
rect 15352 19397 15364 19400
rect 15306 19391 15364 19397
rect 12710 19320 12716 19372
rect 12768 19360 12774 19372
rect 13538 19369 13544 19372
rect 13081 19363 13139 19369
rect 12768 19332 13032 19360
rect 12768 19320 12774 19332
rect 12452 19264 12664 19292
rect 10781 19227 10839 19233
rect 10781 19193 10793 19227
rect 10827 19193 10839 19227
rect 10781 19187 10839 19193
rect 12158 19184 12164 19236
rect 12216 19224 12222 19236
rect 12618 19224 12624 19236
rect 12216 19196 12624 19224
rect 12216 19184 12222 19196
rect 12618 19184 12624 19196
rect 12676 19184 12682 19236
rect 13004 19224 13032 19332
rect 13081 19329 13093 19363
rect 13127 19360 13139 19363
rect 13357 19363 13415 19369
rect 13127 19332 13308 19360
rect 13127 19329 13139 19332
rect 13081 19323 13139 19329
rect 13280 19304 13308 19332
rect 13357 19329 13369 19363
rect 13403 19329 13415 19363
rect 13357 19323 13415 19329
rect 13501 19363 13544 19369
rect 13501 19329 13513 19363
rect 13501 19323 13544 19329
rect 13262 19252 13268 19304
rect 13320 19252 13326 19304
rect 13372 19292 13400 19323
rect 13538 19320 13544 19323
rect 13596 19320 13602 19372
rect 13814 19320 13820 19372
rect 13872 19360 13878 19372
rect 14737 19363 14795 19369
rect 14737 19360 14749 19363
rect 13872 19332 14749 19360
rect 13872 19320 13878 19332
rect 14737 19329 14749 19332
rect 14783 19360 14795 19363
rect 14826 19360 14832 19372
rect 14783 19332 14832 19360
rect 14783 19329 14795 19332
rect 14737 19323 14795 19329
rect 14826 19320 14832 19332
rect 14884 19320 14890 19372
rect 15194 19369 15200 19372
rect 14921 19363 14979 19369
rect 14921 19329 14933 19363
rect 14967 19329 14979 19363
rect 14921 19323 14979 19329
rect 15157 19363 15200 19369
rect 15157 19329 15169 19363
rect 15157 19323 15200 19329
rect 14550 19292 14556 19304
rect 13372 19264 14556 19292
rect 13372 19224 13400 19264
rect 14550 19252 14556 19264
rect 14608 19252 14614 19304
rect 13004 19196 13400 19224
rect 13722 19184 13728 19236
rect 13780 19224 13786 19236
rect 14936 19224 14964 19323
rect 15172 19292 15200 19323
rect 15252 19320 15258 19372
rect 15470 19320 15476 19372
rect 15528 19320 15534 19372
rect 15286 19292 15292 19304
rect 15172 19264 15292 19292
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 15580 19292 15608 19400
rect 15657 19397 15669 19431
rect 15703 19397 15715 19431
rect 16666 19428 16672 19440
rect 15657 19391 15715 19397
rect 15764 19400 16672 19428
rect 15764 19292 15792 19400
rect 16666 19388 16672 19400
rect 16724 19428 16730 19440
rect 18601 19431 18659 19437
rect 18601 19428 18613 19431
rect 16724 19400 18613 19428
rect 16724 19388 16730 19400
rect 18601 19397 18613 19400
rect 18647 19397 18659 19431
rect 19076 19428 19104 19459
rect 19242 19456 19248 19468
rect 19300 19456 19306 19508
rect 20162 19456 20168 19508
rect 20220 19456 20226 19508
rect 20714 19456 20720 19508
rect 20772 19496 20778 19508
rect 20772 19468 22324 19496
rect 20772 19456 20778 19468
rect 21542 19428 21548 19440
rect 18601 19391 18659 19397
rect 18708 19400 19012 19428
rect 19076 19400 21548 19428
rect 15841 19363 15899 19369
rect 15841 19329 15853 19363
rect 15887 19360 15899 19363
rect 15930 19360 15936 19372
rect 15887 19332 15936 19360
rect 15887 19329 15899 19332
rect 15841 19323 15899 19329
rect 15930 19320 15936 19332
rect 15988 19360 15994 19372
rect 18708 19360 18736 19400
rect 15988 19332 18736 19360
rect 15988 19320 15994 19332
rect 18782 19320 18788 19372
rect 18840 19320 18846 19372
rect 18874 19320 18880 19372
rect 18932 19320 18938 19372
rect 18984 19360 19012 19400
rect 19337 19363 19395 19369
rect 19337 19360 19349 19363
rect 18984 19332 19349 19360
rect 19337 19329 19349 19332
rect 19383 19329 19395 19363
rect 19337 19323 19395 19329
rect 19429 19363 19487 19369
rect 19429 19329 19441 19363
rect 19475 19360 19487 19363
rect 19518 19360 19524 19372
rect 19475 19332 19524 19360
rect 19475 19329 19487 19332
rect 19429 19323 19487 19329
rect 19518 19320 19524 19332
rect 19576 19320 19582 19372
rect 19610 19320 19616 19372
rect 19668 19320 19674 19372
rect 19904 19369 19932 19400
rect 21542 19388 21548 19400
rect 21600 19388 21606 19440
rect 22296 19437 22324 19468
rect 23658 19456 23664 19508
rect 23716 19496 23722 19508
rect 24578 19496 24584 19508
rect 23716 19468 24584 19496
rect 23716 19456 23722 19468
rect 24578 19456 24584 19468
rect 24636 19456 24642 19508
rect 29914 19456 29920 19508
rect 29972 19496 29978 19508
rect 32122 19496 32128 19508
rect 29972 19468 32128 19496
rect 29972 19456 29978 19468
rect 32122 19456 32128 19468
rect 32180 19456 32186 19508
rect 32398 19456 32404 19508
rect 32456 19496 32462 19508
rect 32493 19499 32551 19505
rect 32493 19496 32505 19499
rect 32456 19468 32505 19496
rect 32456 19456 32462 19468
rect 32493 19465 32505 19468
rect 32539 19465 32551 19499
rect 32493 19459 32551 19465
rect 34517 19499 34575 19505
rect 34517 19465 34529 19499
rect 34563 19496 34575 19499
rect 34698 19496 34704 19508
rect 34563 19468 34704 19496
rect 34563 19465 34575 19468
rect 34517 19459 34575 19465
rect 34698 19456 34704 19468
rect 34756 19456 34762 19508
rect 39945 19499 40003 19505
rect 39945 19465 39957 19499
rect 39991 19496 40003 19499
rect 40770 19496 40776 19508
rect 39991 19468 40776 19496
rect 39991 19465 40003 19468
rect 39945 19459 40003 19465
rect 40770 19456 40776 19468
rect 40828 19456 40834 19508
rect 44082 19456 44088 19508
rect 44140 19496 44146 19508
rect 44453 19499 44511 19505
rect 44453 19496 44465 19499
rect 44140 19468 44465 19496
rect 44140 19456 44146 19468
rect 44453 19465 44465 19468
rect 44499 19465 44511 19499
rect 44453 19459 44511 19465
rect 22281 19431 22339 19437
rect 21652 19400 22140 19428
rect 19705 19363 19763 19369
rect 19705 19329 19717 19363
rect 19751 19334 19763 19363
rect 19889 19363 19947 19369
rect 19751 19329 19840 19334
rect 19705 19323 19840 19329
rect 19889 19329 19901 19363
rect 19935 19329 19947 19363
rect 19889 19323 19947 19329
rect 19720 19306 19840 19323
rect 19978 19320 19984 19372
rect 20036 19320 20042 19372
rect 20714 19320 20720 19372
rect 20772 19360 20778 19372
rect 20901 19363 20959 19369
rect 20901 19360 20913 19363
rect 20772 19332 20913 19360
rect 20772 19320 20778 19332
rect 20901 19329 20913 19332
rect 20947 19329 20959 19363
rect 21085 19363 21143 19369
rect 21085 19360 21097 19363
rect 20901 19323 20959 19329
rect 21008 19332 21097 19360
rect 19812 19292 19840 19306
rect 20162 19292 20168 19304
rect 15580 19264 15792 19292
rect 16500 19264 19656 19292
rect 19812 19264 20168 19292
rect 15930 19224 15936 19236
rect 13780 19196 15936 19224
rect 13780 19184 13786 19196
rect 15930 19184 15936 19196
rect 15988 19184 15994 19236
rect 4614 19116 4620 19168
rect 4672 19156 4678 19168
rect 8294 19156 8300 19168
rect 4672 19128 8300 19156
rect 4672 19116 4678 19128
rect 8294 19116 8300 19128
rect 8352 19116 8358 19168
rect 11698 19116 11704 19168
rect 11756 19156 11762 19168
rect 16500 19156 16528 19264
rect 16850 19184 16856 19236
rect 16908 19224 16914 19236
rect 17402 19224 17408 19236
rect 16908 19196 17408 19224
rect 16908 19184 16914 19196
rect 17402 19184 17408 19196
rect 17460 19184 17466 19236
rect 18138 19184 18144 19236
rect 18196 19224 18202 19236
rect 19518 19224 19524 19236
rect 18196 19196 19524 19224
rect 18196 19184 18202 19196
rect 19518 19184 19524 19196
rect 19576 19184 19582 19236
rect 11756 19128 16528 19156
rect 11756 19116 11762 19128
rect 16574 19116 16580 19168
rect 16632 19156 16638 19168
rect 18506 19156 18512 19168
rect 16632 19128 18512 19156
rect 16632 19116 16638 19128
rect 18506 19116 18512 19128
rect 18564 19116 18570 19168
rect 18598 19116 18604 19168
rect 18656 19116 18662 19168
rect 19242 19116 19248 19168
rect 19300 19156 19306 19168
rect 19337 19159 19395 19165
rect 19337 19156 19349 19159
rect 19300 19128 19349 19156
rect 19300 19116 19306 19128
rect 19337 19125 19349 19128
rect 19383 19125 19395 19159
rect 19628 19156 19656 19264
rect 20162 19252 20168 19264
rect 20220 19252 20226 19304
rect 20622 19252 20628 19304
rect 20680 19292 20686 19304
rect 21008 19292 21036 19332
rect 21085 19329 21097 19332
rect 21131 19360 21143 19363
rect 21652 19360 21680 19400
rect 21131 19332 21680 19360
rect 21131 19329 21143 19332
rect 21085 19323 21143 19329
rect 22002 19320 22008 19372
rect 22060 19320 22066 19372
rect 22112 19369 22140 19400
rect 22281 19397 22293 19431
rect 22327 19397 22339 19431
rect 22281 19391 22339 19397
rect 23106 19388 23112 19440
rect 23164 19428 23170 19440
rect 23382 19428 23388 19440
rect 23164 19400 23388 19428
rect 23164 19388 23170 19400
rect 23382 19388 23388 19400
rect 23440 19428 23446 19440
rect 33502 19428 33508 19440
rect 23440 19400 33508 19428
rect 23440 19388 23446 19400
rect 33502 19388 33508 19400
rect 33560 19388 33566 19440
rect 34054 19388 34060 19440
rect 34112 19388 34118 19440
rect 34146 19388 34152 19440
rect 34204 19428 34210 19440
rect 41046 19428 41052 19440
rect 34204 19400 34376 19428
rect 34204 19388 34210 19400
rect 22097 19363 22155 19369
rect 22097 19329 22109 19363
rect 22143 19360 22155 19363
rect 22186 19360 22192 19372
rect 22143 19332 22192 19360
rect 22143 19329 22155 19332
rect 22097 19323 22155 19329
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 25958 19320 25964 19372
rect 26016 19360 26022 19372
rect 26970 19360 26976 19372
rect 26016 19332 26976 19360
rect 26016 19320 26022 19332
rect 26970 19320 26976 19332
rect 27028 19360 27034 19372
rect 27798 19360 27804 19372
rect 27028 19332 27804 19360
rect 27028 19320 27034 19332
rect 27798 19320 27804 19332
rect 27856 19360 27862 19372
rect 27982 19360 27988 19372
rect 27856 19332 27988 19360
rect 27856 19320 27862 19332
rect 27982 19320 27988 19332
rect 28040 19320 28046 19372
rect 31294 19320 31300 19372
rect 31352 19360 31358 19372
rect 31389 19363 31447 19369
rect 31389 19360 31401 19363
rect 31352 19332 31401 19360
rect 31352 19320 31358 19332
rect 31389 19329 31401 19332
rect 31435 19360 31447 19363
rect 32125 19363 32183 19369
rect 32125 19360 32137 19363
rect 31435 19332 32137 19360
rect 31435 19329 31447 19332
rect 31389 19323 31447 19329
rect 32125 19329 32137 19332
rect 32171 19329 32183 19363
rect 32125 19323 32183 19329
rect 34238 19320 34244 19372
rect 34296 19320 34302 19372
rect 34348 19369 34376 19400
rect 38580 19400 41052 19428
rect 38580 19372 38608 19400
rect 41046 19388 41052 19400
rect 41104 19428 41110 19440
rect 41104 19400 42472 19428
rect 41104 19388 41110 19400
rect 42444 19372 42472 19400
rect 34333 19363 34391 19369
rect 34333 19329 34345 19363
rect 34379 19329 34391 19363
rect 34333 19323 34391 19329
rect 38562 19320 38568 19372
rect 38620 19320 38626 19372
rect 38654 19320 38660 19372
rect 38712 19360 38718 19372
rect 38821 19363 38879 19369
rect 38821 19360 38833 19363
rect 38712 19332 38833 19360
rect 38712 19320 38718 19332
rect 38821 19329 38833 19332
rect 38867 19329 38879 19363
rect 38821 19323 38879 19329
rect 40221 19363 40279 19369
rect 40221 19329 40233 19363
rect 40267 19360 40279 19363
rect 40310 19360 40316 19372
rect 40267 19332 40316 19360
rect 40267 19329 40279 19332
rect 40221 19323 40279 19329
rect 40310 19320 40316 19332
rect 40368 19320 40374 19372
rect 40402 19320 40408 19372
rect 40460 19320 40466 19372
rect 42426 19320 42432 19372
rect 42484 19320 42490 19372
rect 42702 19369 42708 19372
rect 42696 19323 42708 19369
rect 42702 19320 42708 19323
rect 42760 19320 42766 19372
rect 44269 19363 44327 19369
rect 44269 19360 44281 19363
rect 43824 19332 44281 19360
rect 22922 19292 22928 19304
rect 20680 19264 21036 19292
rect 21376 19264 22928 19292
rect 20680 19252 20686 19264
rect 21376 19224 21404 19264
rect 22922 19252 22928 19264
rect 22980 19292 22986 19304
rect 24026 19292 24032 19304
rect 22980 19264 24032 19292
rect 22980 19252 22986 19264
rect 24026 19252 24032 19264
rect 24084 19292 24090 19304
rect 26234 19292 26240 19304
rect 24084 19264 26240 19292
rect 24084 19252 24090 19264
rect 26234 19252 26240 19264
rect 26292 19252 26298 19304
rect 27890 19252 27896 19304
rect 27948 19292 27954 19304
rect 28074 19292 28080 19304
rect 27948 19264 28080 19292
rect 27948 19252 27954 19264
rect 28074 19252 28080 19264
rect 28132 19252 28138 19304
rect 28994 19252 29000 19304
rect 29052 19292 29058 19304
rect 31481 19295 31539 19301
rect 31481 19292 31493 19295
rect 29052 19264 31493 19292
rect 29052 19252 29058 19264
rect 31481 19261 31493 19264
rect 31527 19292 31539 19295
rect 31527 19264 32168 19292
rect 31527 19261 31539 19264
rect 31481 19255 31539 19261
rect 19904 19196 21404 19224
rect 19904 19156 19932 19196
rect 21450 19184 21456 19236
rect 21508 19224 21514 19236
rect 21508 19196 22232 19224
rect 21508 19184 21514 19196
rect 19628 19128 19932 19156
rect 19981 19159 20039 19165
rect 19337 19119 19395 19125
rect 19981 19125 19993 19159
rect 20027 19156 20039 19159
rect 21266 19156 21272 19168
rect 20027 19128 21272 19156
rect 20027 19125 20039 19128
rect 19981 19119 20039 19125
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 21726 19116 21732 19168
rect 21784 19156 21790 19168
rect 21821 19159 21879 19165
rect 21821 19156 21833 19159
rect 21784 19128 21833 19156
rect 21784 19116 21790 19128
rect 21821 19125 21833 19128
rect 21867 19156 21879 19159
rect 21910 19156 21916 19168
rect 21867 19128 21916 19156
rect 21867 19125 21879 19128
rect 21821 19119 21879 19125
rect 21910 19116 21916 19128
rect 21968 19116 21974 19168
rect 22094 19116 22100 19168
rect 22152 19116 22158 19168
rect 22204 19156 22232 19196
rect 22278 19184 22284 19236
rect 22336 19224 22342 19236
rect 31662 19224 31668 19236
rect 22336 19196 31668 19224
rect 22336 19184 22342 19196
rect 31662 19184 31668 19196
rect 31720 19184 31726 19236
rect 31757 19227 31815 19233
rect 31757 19193 31769 19227
rect 31803 19224 31815 19227
rect 31846 19224 31852 19236
rect 31803 19196 31852 19224
rect 31803 19193 31815 19196
rect 31757 19187 31815 19193
rect 31846 19184 31852 19196
rect 31904 19184 31910 19236
rect 32140 19224 32168 19264
rect 32214 19252 32220 19304
rect 32272 19252 32278 19304
rect 36538 19252 36544 19304
rect 36596 19292 36602 19304
rect 38286 19292 38292 19304
rect 36596 19264 38292 19292
rect 36596 19252 36602 19264
rect 38286 19252 38292 19264
rect 38344 19252 38350 19304
rect 43824 19236 43852 19332
rect 44269 19329 44281 19332
rect 44315 19329 44327 19363
rect 44269 19323 44327 19329
rect 38470 19224 38476 19236
rect 32140 19196 38476 19224
rect 38470 19184 38476 19196
rect 38528 19224 38534 19236
rect 38528 19196 38608 19224
rect 38528 19184 38534 19196
rect 25130 19156 25136 19168
rect 22204 19128 25136 19156
rect 25130 19116 25136 19128
rect 25188 19156 25194 19168
rect 25682 19156 25688 19168
rect 25188 19128 25688 19156
rect 25188 19116 25194 19128
rect 25682 19116 25688 19128
rect 25740 19116 25746 19168
rect 27062 19116 27068 19168
rect 27120 19156 27126 19168
rect 31386 19156 31392 19168
rect 27120 19128 31392 19156
rect 27120 19116 27126 19128
rect 31386 19116 31392 19128
rect 31444 19116 31450 19168
rect 31478 19116 31484 19168
rect 31536 19116 31542 19168
rect 32122 19116 32128 19168
rect 32180 19116 32186 19168
rect 33502 19116 33508 19168
rect 33560 19156 33566 19168
rect 34057 19159 34115 19165
rect 34057 19156 34069 19159
rect 33560 19128 34069 19156
rect 33560 19116 33566 19128
rect 34057 19125 34069 19128
rect 34103 19125 34115 19159
rect 38580 19156 38608 19196
rect 43806 19184 43812 19236
rect 43864 19184 43870 19236
rect 38838 19156 38844 19168
rect 38580 19128 38844 19156
rect 34057 19119 34115 19125
rect 38838 19116 38844 19128
rect 38896 19116 38902 19168
rect 40034 19116 40040 19168
rect 40092 19116 40098 19168
rect 1104 19066 44896 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 44896 19066
rect 1104 18992 44896 19014
rect 2498 18912 2504 18964
rect 2556 18912 2562 18964
rect 3418 18912 3424 18964
rect 3476 18912 3482 18964
rect 4433 18955 4491 18961
rect 4433 18921 4445 18955
rect 4479 18952 4491 18955
rect 4614 18952 4620 18964
rect 4479 18924 4620 18952
rect 4479 18921 4491 18924
rect 4433 18915 4491 18921
rect 4614 18912 4620 18924
rect 4672 18912 4678 18964
rect 5721 18955 5779 18961
rect 5721 18921 5733 18955
rect 5767 18952 5779 18955
rect 6270 18952 6276 18964
rect 5767 18924 6276 18952
rect 5767 18921 5779 18924
rect 5721 18915 5779 18921
rect 6270 18912 6276 18924
rect 6328 18912 6334 18964
rect 7190 18912 7196 18964
rect 7248 18952 7254 18964
rect 9769 18955 9827 18961
rect 7248 18924 9352 18952
rect 7248 18912 7254 18924
rect 2866 18844 2872 18896
rect 2924 18884 2930 18896
rect 3053 18887 3111 18893
rect 3053 18884 3065 18887
rect 2924 18856 3065 18884
rect 2924 18844 2930 18856
rect 3053 18853 3065 18856
rect 3099 18884 3111 18887
rect 4062 18884 4068 18896
rect 3099 18856 4068 18884
rect 3099 18853 3111 18856
rect 3053 18847 3111 18853
rect 4062 18844 4068 18856
rect 4120 18844 4126 18896
rect 4801 18887 4859 18893
rect 4801 18853 4813 18887
rect 4847 18884 4859 18887
rect 6362 18884 6368 18896
rect 4847 18856 6368 18884
rect 4847 18853 4859 18856
rect 4801 18847 4859 18853
rect 4816 18816 4844 18847
rect 6362 18844 6368 18856
rect 6420 18844 6426 18896
rect 6546 18844 6552 18896
rect 6604 18884 6610 18896
rect 7837 18887 7895 18893
rect 6604 18856 7748 18884
rect 6604 18844 6610 18856
rect 6178 18816 6184 18828
rect 4724 18788 4844 18816
rect 5644 18788 6184 18816
rect 3234 18708 3240 18760
rect 3292 18708 3298 18760
rect 3418 18708 3424 18760
rect 3476 18748 3482 18760
rect 3605 18751 3663 18757
rect 3605 18748 3617 18751
rect 3476 18720 3617 18748
rect 3476 18708 3482 18720
rect 3605 18717 3617 18720
rect 3651 18717 3663 18751
rect 3605 18711 3663 18717
rect 3878 18708 3884 18760
rect 3936 18708 3942 18760
rect 3970 18708 3976 18760
rect 4028 18748 4034 18760
rect 4065 18751 4123 18757
rect 4065 18748 4077 18751
rect 4028 18720 4077 18748
rect 4028 18708 4034 18720
rect 4065 18717 4077 18720
rect 4111 18717 4123 18751
rect 4065 18711 4123 18717
rect 4301 18751 4359 18757
rect 4301 18717 4313 18751
rect 4347 18748 4359 18751
rect 4724 18748 4752 18788
rect 4347 18720 4752 18748
rect 4347 18717 4359 18720
rect 4301 18711 4359 18717
rect 4798 18708 4804 18760
rect 4856 18748 4862 18760
rect 5169 18751 5227 18757
rect 5169 18748 5181 18751
rect 4856 18720 5181 18748
rect 4856 18708 4862 18720
rect 5169 18717 5181 18720
rect 5215 18717 5227 18751
rect 5169 18711 5227 18717
rect 5258 18708 5264 18760
rect 5316 18748 5322 18760
rect 5644 18757 5672 18788
rect 6178 18776 6184 18788
rect 6236 18776 6242 18828
rect 7098 18776 7104 18828
rect 7156 18776 7162 18828
rect 5589 18751 5672 18757
rect 5589 18748 5601 18751
rect 5316 18720 5601 18748
rect 5316 18708 5322 18720
rect 5589 18717 5601 18720
rect 5635 18720 5672 18751
rect 6089 18751 6147 18757
rect 5635 18717 5647 18720
rect 5589 18711 5647 18717
rect 6089 18717 6101 18751
rect 6135 18748 6147 18751
rect 6270 18748 6276 18760
rect 6135 18720 6276 18748
rect 6135 18717 6147 18720
rect 6089 18711 6147 18717
rect 6270 18708 6276 18720
rect 6328 18708 6334 18760
rect 6454 18708 6460 18760
rect 6512 18708 6518 18760
rect 6641 18751 6699 18757
rect 6641 18717 6653 18751
rect 6687 18748 6699 18751
rect 7558 18748 7564 18760
rect 6687 18720 7564 18748
rect 6687 18717 6699 18720
rect 6641 18711 6699 18717
rect 2406 18640 2412 18692
rect 2464 18640 2470 18692
rect 3326 18640 3332 18692
rect 3384 18680 3390 18692
rect 4157 18683 4215 18689
rect 4157 18680 4169 18683
rect 3384 18652 4169 18680
rect 3384 18640 3390 18652
rect 4157 18649 4169 18652
rect 4203 18680 4215 18683
rect 4706 18680 4712 18692
rect 4203 18652 4712 18680
rect 4203 18649 4215 18652
rect 4157 18643 4215 18649
rect 4706 18640 4712 18652
rect 4764 18640 4770 18692
rect 4985 18683 5043 18689
rect 4985 18649 4997 18683
rect 5031 18680 5043 18683
rect 5074 18680 5080 18692
rect 5031 18652 5080 18680
rect 5031 18649 5043 18652
rect 4985 18643 5043 18649
rect 5074 18640 5080 18652
rect 5132 18640 5138 18692
rect 5353 18683 5411 18689
rect 5353 18649 5365 18683
rect 5399 18649 5411 18683
rect 5353 18643 5411 18649
rect 5445 18683 5503 18689
rect 5445 18649 5457 18683
rect 5491 18680 5503 18683
rect 5810 18680 5816 18692
rect 5491 18652 5816 18680
rect 5491 18649 5503 18652
rect 5445 18643 5503 18649
rect 5368 18612 5396 18643
rect 5810 18640 5816 18652
rect 5868 18640 5874 18692
rect 5902 18612 5908 18624
rect 5368 18584 5908 18612
rect 5902 18572 5908 18584
rect 5960 18572 5966 18624
rect 6086 18572 6092 18624
rect 6144 18612 6150 18624
rect 6656 18612 6684 18711
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 7720 18680 7748 18856
rect 7837 18853 7849 18887
rect 7883 18884 7895 18887
rect 8202 18884 8208 18896
rect 7883 18856 8208 18884
rect 7883 18853 7895 18856
rect 7837 18847 7895 18853
rect 8202 18844 8208 18856
rect 8260 18844 8266 18896
rect 8665 18887 8723 18893
rect 8665 18853 8677 18887
rect 8711 18884 8723 18887
rect 9214 18884 9220 18896
rect 8711 18856 9220 18884
rect 8711 18853 8723 18856
rect 8665 18847 8723 18853
rect 9214 18844 9220 18856
rect 9272 18844 9278 18896
rect 7926 18776 7932 18828
rect 7984 18816 7990 18828
rect 7984 18788 8156 18816
rect 7984 18776 7990 18788
rect 8018 18708 8024 18760
rect 8076 18708 8082 18760
rect 8128 18757 8156 18788
rect 8220 18788 9260 18816
rect 8113 18751 8171 18757
rect 8113 18717 8125 18751
rect 8159 18717 8171 18751
rect 8113 18711 8171 18717
rect 8220 18680 8248 18788
rect 8294 18708 8300 18760
rect 8352 18708 8358 18760
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 7720 18652 8248 18680
rect 6144 18584 6684 18612
rect 6144 18572 6150 18584
rect 8202 18572 8208 18624
rect 8260 18612 8266 18624
rect 8404 18612 8432 18711
rect 8478 18708 8484 18760
rect 8536 18757 8542 18760
rect 8536 18751 8591 18757
rect 8536 18717 8545 18751
rect 8579 18748 8591 18751
rect 8938 18748 8944 18760
rect 8579 18720 8944 18748
rect 8579 18717 8591 18720
rect 8536 18711 8591 18717
rect 8536 18708 8542 18711
rect 8938 18708 8944 18720
rect 8996 18708 9002 18760
rect 9232 18757 9260 18788
rect 9217 18751 9275 18757
rect 9217 18717 9229 18751
rect 9263 18717 9275 18751
rect 9324 18748 9352 18924
rect 9769 18921 9781 18955
rect 9815 18952 9827 18955
rect 9858 18952 9864 18964
rect 9815 18924 9864 18952
rect 9815 18921 9827 18924
rect 9769 18915 9827 18921
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 10502 18912 10508 18964
rect 10560 18912 10566 18964
rect 11241 18955 11299 18961
rect 11241 18921 11253 18955
rect 11287 18952 11299 18955
rect 11287 18924 16988 18952
rect 11287 18921 11299 18924
rect 11241 18915 11299 18921
rect 9950 18844 9956 18896
rect 10008 18884 10014 18896
rect 10008 18856 11468 18884
rect 10008 18844 10014 18856
rect 9674 18757 9680 18760
rect 9493 18751 9551 18757
rect 9493 18748 9505 18751
rect 9324 18720 9505 18748
rect 9217 18711 9275 18717
rect 9493 18717 9505 18720
rect 9539 18717 9551 18751
rect 9493 18711 9551 18717
rect 9637 18751 9680 18757
rect 9637 18717 9649 18751
rect 9637 18711 9680 18717
rect 9674 18708 9680 18711
rect 9732 18708 9738 18760
rect 9858 18708 9864 18760
rect 9916 18748 9922 18760
rect 9953 18751 10011 18757
rect 9953 18748 9965 18751
rect 9916 18720 9965 18748
rect 9916 18708 9922 18720
rect 9953 18717 9965 18720
rect 9999 18717 10011 18751
rect 10326 18751 10384 18757
rect 10326 18748 10338 18751
rect 9953 18711 10011 18717
rect 10060 18720 10338 18748
rect 9401 18683 9459 18689
rect 9401 18649 9413 18683
rect 9447 18649 9459 18683
rect 9692 18680 9720 18708
rect 10060 18680 10088 18720
rect 10326 18717 10338 18720
rect 10372 18717 10384 18751
rect 10326 18711 10384 18717
rect 9692 18652 10088 18680
rect 9401 18643 9459 18649
rect 8260 18584 8432 18612
rect 8260 18572 8266 18584
rect 9030 18572 9036 18624
rect 9088 18612 9094 18624
rect 9416 18612 9444 18643
rect 10134 18640 10140 18692
rect 10192 18640 10198 18692
rect 10226 18640 10232 18692
rect 10284 18640 10290 18692
rect 10341 18680 10369 18711
rect 10686 18708 10692 18760
rect 10744 18708 10750 18760
rect 11057 18751 11115 18757
rect 11057 18748 11069 18751
rect 10789 18720 11069 18748
rect 10789 18680 10817 18720
rect 11057 18717 11069 18720
rect 11103 18717 11115 18751
rect 11440 18748 11468 18856
rect 11974 18844 11980 18896
rect 12032 18884 12038 18896
rect 12032 18856 12572 18884
rect 12032 18844 12038 18856
rect 12434 18776 12440 18828
rect 12492 18776 12498 18828
rect 12158 18748 12164 18760
rect 11440 18720 12164 18748
rect 11057 18711 11115 18717
rect 12158 18708 12164 18720
rect 12216 18748 12222 18760
rect 12253 18751 12311 18757
rect 12253 18748 12265 18751
rect 12216 18720 12265 18748
rect 12216 18708 12222 18720
rect 12253 18717 12265 18720
rect 12299 18717 12311 18751
rect 12253 18711 12311 18717
rect 10341 18652 10817 18680
rect 10873 18683 10931 18689
rect 10873 18649 10885 18683
rect 10919 18649 10931 18683
rect 10873 18643 10931 18649
rect 10152 18612 10180 18640
rect 10888 18612 10916 18643
rect 10962 18640 10968 18692
rect 11020 18680 11026 18692
rect 12342 18680 12348 18692
rect 11020 18652 12348 18680
rect 11020 18640 11026 18652
rect 12342 18640 12348 18652
rect 12400 18640 12406 18692
rect 12469 18689 12497 18776
rect 12544 18757 12572 18856
rect 12802 18844 12808 18896
rect 12860 18844 12866 18896
rect 13354 18884 13360 18896
rect 12912 18856 13360 18884
rect 12710 18776 12716 18828
rect 12768 18816 12774 18828
rect 12912 18816 12940 18856
rect 13354 18844 13360 18856
rect 13412 18844 13418 18896
rect 13446 18844 13452 18896
rect 13504 18884 13510 18896
rect 13541 18887 13599 18893
rect 13541 18884 13553 18887
rect 13504 18856 13553 18884
rect 13504 18844 13510 18856
rect 13541 18853 13553 18856
rect 13587 18853 13599 18887
rect 13541 18847 13599 18853
rect 15013 18887 15071 18893
rect 15013 18853 15025 18887
rect 15059 18884 15071 18887
rect 15470 18884 15476 18896
rect 15059 18856 15476 18884
rect 15059 18853 15071 18856
rect 15013 18847 15071 18853
rect 15470 18844 15476 18856
rect 15528 18844 15534 18896
rect 16960 18884 16988 18924
rect 17034 18912 17040 18964
rect 17092 18912 17098 18964
rect 20622 18952 20628 18964
rect 19168 18924 20628 18952
rect 19168 18884 19196 18924
rect 20622 18912 20628 18924
rect 20680 18912 20686 18964
rect 21726 18912 21732 18964
rect 21784 18912 21790 18964
rect 23474 18912 23480 18964
rect 23532 18952 23538 18964
rect 25133 18955 25191 18961
rect 25133 18952 25145 18955
rect 23532 18924 25145 18952
rect 23532 18912 23538 18924
rect 25133 18921 25145 18924
rect 25179 18952 25191 18955
rect 27522 18952 27528 18964
rect 25179 18924 27528 18952
rect 25179 18921 25191 18924
rect 25133 18915 25191 18921
rect 27522 18912 27528 18924
rect 27580 18912 27586 18964
rect 27890 18912 27896 18964
rect 27948 18952 27954 18964
rect 27985 18955 28043 18961
rect 27985 18952 27997 18955
rect 27948 18924 27997 18952
rect 27948 18912 27954 18924
rect 27985 18921 27997 18924
rect 28031 18921 28043 18955
rect 28902 18952 28908 18964
rect 27985 18915 28043 18921
rect 28368 18924 28908 18952
rect 16960 18856 19196 18884
rect 19242 18844 19248 18896
rect 19300 18884 19306 18896
rect 21174 18884 21180 18896
rect 19300 18856 21180 18884
rect 19300 18844 19306 18856
rect 21174 18844 21180 18856
rect 21232 18844 21238 18896
rect 22094 18884 22100 18896
rect 21829 18856 22100 18884
rect 12768 18788 12940 18816
rect 12768 18776 12774 18788
rect 12529 18751 12587 18757
rect 12529 18717 12541 18751
rect 12575 18717 12587 18751
rect 12529 18711 12587 18717
rect 12626 18751 12684 18757
rect 12626 18717 12638 18751
rect 12672 18748 12684 18751
rect 12912 18748 12940 18788
rect 13262 18776 13268 18828
rect 13320 18816 13326 18828
rect 13320 18788 13400 18816
rect 13320 18776 13326 18788
rect 13372 18757 13400 18788
rect 14918 18776 14924 18828
rect 14976 18816 14982 18828
rect 21829 18816 21857 18856
rect 22094 18844 22100 18856
rect 22152 18844 22158 18896
rect 14976 18788 19288 18816
rect 14976 18776 14982 18788
rect 12672 18720 12940 18748
rect 12989 18751 13047 18757
rect 12672 18717 12684 18720
rect 12626 18711 12684 18717
rect 12989 18717 13001 18751
rect 13035 18717 13047 18751
rect 12989 18711 13047 18717
rect 13357 18751 13415 18757
rect 13357 18717 13369 18751
rect 13403 18748 13415 18751
rect 13630 18748 13636 18760
rect 13403 18720 13636 18748
rect 13403 18717 13415 18720
rect 13357 18711 13415 18717
rect 12437 18683 12497 18689
rect 12437 18649 12449 18683
rect 12483 18652 12497 18683
rect 12483 18649 12495 18652
rect 12437 18643 12495 18649
rect 12710 18640 12716 18692
rect 12768 18680 12774 18692
rect 13004 18680 13032 18711
rect 13630 18708 13636 18720
rect 13688 18708 13694 18760
rect 14458 18708 14464 18760
rect 14516 18708 14522 18760
rect 14642 18708 14648 18760
rect 14700 18708 14706 18760
rect 14826 18708 14832 18760
rect 14884 18708 14890 18760
rect 16761 18751 16819 18757
rect 16761 18748 16773 18751
rect 16132 18720 16773 18748
rect 12768 18652 13032 18680
rect 12768 18640 12774 18652
rect 13170 18640 13176 18692
rect 13228 18640 13234 18692
rect 13265 18683 13323 18689
rect 13265 18649 13277 18683
rect 13311 18649 13323 18683
rect 13265 18643 13323 18649
rect 9088 18584 10916 18612
rect 9088 18572 9094 18584
rect 11882 18572 11888 18624
rect 11940 18612 11946 18624
rect 12158 18612 12164 18624
rect 11940 18584 12164 18612
rect 11940 18572 11946 18584
rect 12158 18572 12164 18584
rect 12216 18612 12222 18624
rect 13280 18612 13308 18643
rect 14366 18640 14372 18692
rect 14424 18680 14430 18692
rect 14737 18683 14795 18689
rect 14737 18680 14749 18683
rect 14424 18652 14749 18680
rect 14424 18640 14430 18652
rect 14737 18649 14749 18652
rect 14783 18649 14795 18683
rect 14737 18643 14795 18649
rect 12216 18584 13308 18612
rect 12216 18572 12222 18584
rect 13446 18572 13452 18624
rect 13504 18612 13510 18624
rect 16132 18612 16160 18720
rect 16761 18717 16773 18720
rect 16807 18717 16819 18751
rect 16761 18711 16819 18717
rect 16853 18751 16911 18757
rect 16853 18717 16865 18751
rect 16899 18748 16911 18751
rect 16942 18748 16948 18760
rect 16899 18720 16948 18748
rect 16899 18717 16911 18720
rect 16853 18711 16911 18717
rect 16776 18680 16804 18711
rect 16942 18708 16948 18720
rect 17000 18708 17006 18760
rect 17037 18751 17095 18757
rect 17037 18717 17049 18751
rect 17083 18748 17095 18751
rect 17218 18748 17224 18760
rect 17083 18720 17224 18748
rect 17083 18717 17095 18720
rect 17037 18711 17095 18717
rect 17218 18708 17224 18720
rect 17276 18748 17282 18760
rect 19150 18748 19156 18760
rect 17276 18720 19156 18748
rect 17276 18708 17282 18720
rect 19150 18708 19156 18720
rect 19208 18708 19214 18760
rect 19260 18757 19288 18788
rect 21744 18788 21857 18816
rect 19245 18751 19303 18757
rect 19245 18717 19257 18751
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 19429 18751 19487 18757
rect 19429 18717 19441 18751
rect 19475 18748 19487 18751
rect 19978 18748 19984 18760
rect 19475 18720 19984 18748
rect 19475 18717 19487 18720
rect 19429 18711 19487 18717
rect 19978 18708 19984 18720
rect 20036 18708 20042 18760
rect 21542 18708 21548 18760
rect 21600 18708 21606 18760
rect 21744 18757 21772 18788
rect 21910 18776 21916 18828
rect 21968 18816 21974 18828
rect 23474 18816 23480 18828
rect 21968 18788 23480 18816
rect 21968 18776 21974 18788
rect 23474 18776 23480 18788
rect 23532 18776 23538 18828
rect 24854 18776 24860 18828
rect 24912 18816 24918 18828
rect 25041 18819 25099 18825
rect 25041 18816 25053 18819
rect 24912 18788 25053 18816
rect 24912 18776 24918 18788
rect 25041 18785 25053 18788
rect 25087 18785 25099 18819
rect 25041 18779 25099 18785
rect 28169 18819 28227 18825
rect 28169 18785 28181 18819
rect 28215 18816 28227 18819
rect 28368 18816 28396 18924
rect 28902 18912 28908 18924
rect 28960 18912 28966 18964
rect 29365 18955 29423 18961
rect 29365 18921 29377 18955
rect 29411 18952 29423 18955
rect 30098 18952 30104 18964
rect 29411 18924 30104 18952
rect 29411 18921 29423 18924
rect 29365 18915 29423 18921
rect 30098 18912 30104 18924
rect 30156 18912 30162 18964
rect 31665 18955 31723 18961
rect 31665 18921 31677 18955
rect 31711 18952 31723 18955
rect 31846 18952 31852 18964
rect 31711 18924 31852 18952
rect 31711 18921 31723 18924
rect 31665 18915 31723 18921
rect 31846 18912 31852 18924
rect 31904 18912 31910 18964
rect 37458 18912 37464 18964
rect 37516 18952 37522 18964
rect 38473 18955 38531 18961
rect 37516 18924 38240 18952
rect 37516 18912 37522 18924
rect 28445 18887 28503 18893
rect 28445 18853 28457 18887
rect 28491 18884 28503 18887
rect 36538 18884 36544 18896
rect 28491 18856 36544 18884
rect 28491 18853 28503 18856
rect 28445 18847 28503 18853
rect 36538 18844 36544 18856
rect 36596 18844 36602 18896
rect 38212 18893 38240 18924
rect 38473 18921 38485 18955
rect 38519 18952 38531 18955
rect 38654 18952 38660 18964
rect 38519 18924 38660 18952
rect 38519 18921 38531 18924
rect 38473 18915 38531 18921
rect 38654 18912 38660 18924
rect 38712 18912 38718 18964
rect 41782 18952 41788 18964
rect 40144 18924 41788 18952
rect 38197 18887 38255 18893
rect 38197 18853 38209 18887
rect 38243 18853 38255 18887
rect 38197 18847 38255 18853
rect 40034 18844 40040 18896
rect 40092 18844 40098 18896
rect 40144 18893 40172 18924
rect 41782 18912 41788 18924
rect 41840 18912 41846 18964
rect 40129 18887 40187 18893
rect 40129 18853 40141 18887
rect 40175 18853 40187 18887
rect 40129 18847 40187 18853
rect 42429 18887 42487 18893
rect 42429 18853 42441 18887
rect 42475 18884 42487 18887
rect 42475 18856 43208 18884
rect 42475 18853 42487 18856
rect 42429 18847 42487 18853
rect 29546 18816 29552 18828
rect 28215 18788 28396 18816
rect 29012 18788 29552 18816
rect 28215 18785 28227 18788
rect 28169 18779 28227 18785
rect 21729 18751 21787 18757
rect 21729 18726 21741 18751
rect 21652 18717 21741 18726
rect 21775 18717 21787 18751
rect 21652 18711 21787 18717
rect 21652 18698 21772 18711
rect 21818 18708 21824 18760
rect 21876 18708 21882 18760
rect 24026 18708 24032 18760
rect 24084 18748 24090 18760
rect 24949 18751 25007 18757
rect 24949 18748 24961 18751
rect 24084 18720 24961 18748
rect 24084 18708 24090 18720
rect 24949 18717 24961 18720
rect 24995 18717 25007 18751
rect 25056 18748 25084 18779
rect 27985 18751 28043 18757
rect 27985 18748 27997 18751
rect 25056 18720 27997 18748
rect 24949 18711 25007 18717
rect 27985 18717 27997 18720
rect 28031 18717 28043 18751
rect 27985 18711 28043 18717
rect 28258 18708 28264 18760
rect 28316 18708 28322 18760
rect 28534 18708 28540 18760
rect 28592 18748 28598 18760
rect 28810 18748 28816 18760
rect 28592 18720 28816 18748
rect 28592 18708 28598 18720
rect 28810 18708 28816 18720
rect 28868 18708 28874 18760
rect 28902 18708 28908 18760
rect 28960 18748 28966 18760
rect 29012 18748 29040 18788
rect 29546 18776 29552 18788
rect 29604 18776 29610 18828
rect 31018 18776 31024 18828
rect 31076 18816 31082 18828
rect 31481 18819 31539 18825
rect 31481 18816 31493 18819
rect 31076 18788 31493 18816
rect 31076 18776 31082 18788
rect 31481 18785 31493 18788
rect 31527 18816 31539 18819
rect 31754 18816 31760 18828
rect 31527 18788 31760 18816
rect 31527 18785 31539 18788
rect 31481 18779 31539 18785
rect 31754 18776 31760 18788
rect 31812 18776 31818 18828
rect 37274 18776 37280 18828
rect 37332 18816 37338 18828
rect 37553 18819 37611 18825
rect 37553 18816 37565 18819
rect 37332 18788 37565 18816
rect 37332 18776 37338 18788
rect 37553 18785 37565 18788
rect 37599 18785 37611 18819
rect 40052 18816 40080 18844
rect 37553 18779 37611 18785
rect 38028 18788 40080 18816
rect 28960 18720 29040 18748
rect 28960 18708 28966 18720
rect 29086 18708 29092 18760
rect 29144 18708 29150 18760
rect 29178 18708 29184 18760
rect 29236 18708 29242 18760
rect 30742 18708 30748 18760
rect 30800 18748 30806 18760
rect 31389 18751 31447 18757
rect 31389 18748 31401 18751
rect 30800 18720 31401 18748
rect 30800 18708 30806 18720
rect 31389 18717 31401 18720
rect 31435 18717 31447 18751
rect 31665 18751 31723 18757
rect 31665 18748 31677 18751
rect 31389 18711 31447 18717
rect 31496 18720 31677 18748
rect 20714 18680 20720 18692
rect 16776 18652 20720 18680
rect 20714 18640 20720 18652
rect 20772 18640 20778 18692
rect 20898 18640 20904 18692
rect 20956 18680 20962 18692
rect 21652 18680 21680 18698
rect 31496 18692 31524 18720
rect 31665 18717 31677 18720
rect 31711 18717 31723 18751
rect 31665 18711 31723 18717
rect 32582 18708 32588 18760
rect 32640 18748 32646 18760
rect 36998 18748 37004 18760
rect 32640 18720 37004 18748
rect 32640 18708 32646 18720
rect 36998 18708 37004 18720
rect 37056 18708 37062 18760
rect 37090 18708 37096 18760
rect 37148 18748 37154 18760
rect 38028 18757 38056 18788
rect 41046 18776 41052 18828
rect 41104 18776 41110 18828
rect 43180 18760 43208 18856
rect 43806 18776 43812 18828
rect 43864 18776 43870 18828
rect 37461 18751 37519 18757
rect 37461 18748 37473 18751
rect 37148 18720 37473 18748
rect 37148 18708 37154 18720
rect 37461 18717 37473 18720
rect 37507 18717 37519 18751
rect 37461 18711 37519 18717
rect 38013 18751 38071 18757
rect 38013 18717 38025 18751
rect 38059 18717 38071 18751
rect 38013 18711 38071 18717
rect 38102 18708 38108 18760
rect 38160 18708 38166 18760
rect 38286 18708 38292 18760
rect 38344 18708 38350 18760
rect 38930 18708 38936 18760
rect 38988 18748 38994 18760
rect 40037 18751 40095 18757
rect 40037 18748 40049 18751
rect 38988 18720 40049 18748
rect 38988 18708 38994 18720
rect 40037 18717 40049 18720
rect 40083 18717 40095 18751
rect 40037 18711 40095 18717
rect 40221 18751 40279 18757
rect 40221 18717 40233 18751
rect 40267 18717 40279 18751
rect 40221 18711 40279 18717
rect 20956 18652 21680 18680
rect 20956 18640 20962 18652
rect 22094 18640 22100 18692
rect 22152 18680 22158 18692
rect 22152 18652 28994 18680
rect 22152 18640 22158 18652
rect 13504 18584 16160 18612
rect 13504 18572 13510 18584
rect 16574 18572 16580 18624
rect 16632 18572 16638 18624
rect 17218 18572 17224 18624
rect 17276 18612 17282 18624
rect 17494 18612 17500 18624
rect 17276 18584 17500 18612
rect 17276 18572 17282 18584
rect 17494 18572 17500 18584
rect 17552 18572 17558 18624
rect 17770 18572 17776 18624
rect 17828 18612 17834 18624
rect 19518 18612 19524 18624
rect 17828 18584 19524 18612
rect 17828 18572 17834 18584
rect 19518 18572 19524 18584
rect 19576 18572 19582 18624
rect 19613 18615 19671 18621
rect 19613 18581 19625 18615
rect 19659 18612 19671 18615
rect 21542 18612 21548 18624
rect 19659 18584 21548 18612
rect 19659 18581 19671 18584
rect 19613 18575 19671 18581
rect 21542 18572 21548 18584
rect 21600 18572 21606 18624
rect 22005 18615 22063 18621
rect 22005 18581 22017 18615
rect 22051 18612 22063 18615
rect 22370 18612 22376 18624
rect 22051 18584 22376 18612
rect 22051 18581 22063 18584
rect 22005 18575 22063 18581
rect 22370 18572 22376 18584
rect 22428 18572 22434 18624
rect 25317 18615 25375 18621
rect 25317 18581 25329 18615
rect 25363 18612 25375 18615
rect 28534 18612 28540 18624
rect 25363 18584 28540 18612
rect 25363 18581 25375 18584
rect 25317 18575 25375 18581
rect 28534 18572 28540 18584
rect 28592 18572 28598 18624
rect 28718 18572 28724 18624
rect 28776 18572 28782 18624
rect 28966 18612 28994 18652
rect 29362 18640 29368 18692
rect 29420 18680 29426 18692
rect 30650 18680 30656 18692
rect 29420 18652 30656 18680
rect 29420 18640 29426 18652
rect 30650 18640 30656 18652
rect 30708 18640 30714 18692
rect 31478 18640 31484 18692
rect 31536 18640 31542 18692
rect 34974 18680 34980 18692
rect 31726 18652 34980 18680
rect 31726 18612 31754 18652
rect 34974 18640 34980 18652
rect 35032 18640 35038 18692
rect 38746 18640 38752 18692
rect 38804 18680 38810 18692
rect 40236 18680 40264 18711
rect 40310 18708 40316 18760
rect 40368 18708 40374 18760
rect 40497 18751 40555 18757
rect 40497 18717 40509 18751
rect 40543 18748 40555 18751
rect 40862 18748 40868 18760
rect 40543 18720 40868 18748
rect 40543 18717 40555 18720
rect 40497 18711 40555 18717
rect 40862 18708 40868 18720
rect 40920 18708 40926 18760
rect 43162 18708 43168 18760
rect 43220 18708 43226 18760
rect 44269 18751 44327 18757
rect 44269 18717 44281 18751
rect 44315 18717 44327 18751
rect 44269 18711 44327 18717
rect 38804 18652 40264 18680
rect 40328 18680 40356 18708
rect 41138 18680 41144 18692
rect 40328 18652 41144 18680
rect 38804 18640 38810 18652
rect 41138 18640 41144 18652
rect 41196 18640 41202 18692
rect 41316 18683 41374 18689
rect 41316 18649 41328 18683
rect 41362 18680 41374 18683
rect 41598 18680 41604 18692
rect 41362 18652 41604 18680
rect 41362 18649 41374 18652
rect 41316 18643 41374 18649
rect 41598 18640 41604 18652
rect 41656 18640 41662 18692
rect 41690 18640 41696 18692
rect 41748 18680 41754 18692
rect 44284 18680 44312 18711
rect 41748 18652 44312 18680
rect 41748 18640 41754 18652
rect 28966 18584 31754 18612
rect 31849 18615 31907 18621
rect 31849 18581 31861 18615
rect 31895 18612 31907 18615
rect 32306 18612 32312 18624
rect 31895 18584 32312 18612
rect 31895 18581 31907 18584
rect 31849 18575 31907 18581
rect 32306 18572 32312 18584
rect 32364 18572 32370 18624
rect 34054 18572 34060 18624
rect 34112 18612 34118 18624
rect 37182 18612 37188 18624
rect 34112 18584 37188 18612
rect 34112 18572 34118 18584
rect 37182 18572 37188 18584
rect 37240 18572 37246 18624
rect 37829 18615 37887 18621
rect 37829 18581 37841 18615
rect 37875 18612 37887 18615
rect 39574 18612 39580 18624
rect 37875 18584 39580 18612
rect 37875 18581 37887 18584
rect 37829 18575 37887 18581
rect 39574 18572 39580 18584
rect 39632 18572 39638 18624
rect 39853 18615 39911 18621
rect 39853 18581 39865 18615
rect 39899 18612 39911 18615
rect 40126 18612 40132 18624
rect 39899 18584 40132 18612
rect 39899 18581 39911 18584
rect 39853 18575 39911 18581
rect 40126 18572 40132 18584
rect 40184 18572 40190 18624
rect 42518 18572 42524 18624
rect 42576 18572 42582 18624
rect 43254 18572 43260 18624
rect 43312 18572 43318 18624
rect 44450 18572 44456 18624
rect 44508 18572 44514 18624
rect 1104 18522 44896 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 44896 18522
rect 1104 18448 44896 18470
rect 3421 18411 3479 18417
rect 3421 18377 3433 18411
rect 3467 18408 3479 18411
rect 3602 18408 3608 18420
rect 3467 18380 3608 18408
rect 3467 18377 3479 18380
rect 3421 18371 3479 18377
rect 3602 18368 3608 18380
rect 3660 18368 3666 18420
rect 4798 18368 4804 18420
rect 4856 18408 4862 18420
rect 4856 18380 6684 18408
rect 4856 18368 4862 18380
rect 5276 18349 5304 18380
rect 4065 18343 4123 18349
rect 4065 18309 4077 18343
rect 4111 18340 4123 18343
rect 5261 18343 5319 18349
rect 4111 18312 5120 18340
rect 4111 18309 4123 18312
rect 4065 18303 4123 18309
rect 2130 18232 2136 18284
rect 2188 18272 2194 18284
rect 2498 18272 2504 18284
rect 2188 18244 2504 18272
rect 2188 18232 2194 18244
rect 2498 18232 2504 18244
rect 2556 18232 2562 18284
rect 2866 18232 2872 18284
rect 2924 18232 2930 18284
rect 3418 18232 3424 18284
rect 3476 18272 3482 18284
rect 3697 18275 3755 18281
rect 3697 18272 3709 18275
rect 3476 18244 3709 18272
rect 3476 18232 3482 18244
rect 3697 18241 3709 18244
rect 3743 18241 3755 18275
rect 3697 18235 3755 18241
rect 2590 18164 2596 18216
rect 2648 18164 2654 18216
rect 3050 18164 3056 18216
rect 3108 18164 3114 18216
rect 2608 18136 2636 18164
rect 4080 18136 4108 18303
rect 4249 18275 4307 18281
rect 4249 18241 4261 18275
rect 4295 18272 4307 18275
rect 4614 18272 4620 18284
rect 4295 18244 4620 18272
rect 4295 18241 4307 18244
rect 4249 18235 4307 18241
rect 4614 18232 4620 18244
rect 4672 18232 4678 18284
rect 5092 18272 5120 18312
rect 5261 18309 5273 18343
rect 5307 18309 5319 18343
rect 5261 18303 5319 18309
rect 5353 18343 5411 18349
rect 5353 18309 5365 18343
rect 5399 18340 5411 18343
rect 5902 18340 5908 18352
rect 5399 18312 5908 18340
rect 5399 18309 5411 18312
rect 5353 18303 5411 18309
rect 5902 18300 5908 18312
rect 5960 18300 5966 18352
rect 6656 18349 6684 18380
rect 6822 18368 6828 18420
rect 6880 18408 6886 18420
rect 10134 18408 10140 18420
rect 6880 18380 10140 18408
rect 6880 18368 6886 18380
rect 10134 18368 10140 18380
rect 10192 18368 10198 18420
rect 10226 18368 10232 18420
rect 10284 18408 10290 18420
rect 11882 18408 11888 18420
rect 10284 18380 11888 18408
rect 10284 18368 10290 18380
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 12342 18368 12348 18420
rect 12400 18408 12406 18420
rect 13262 18408 13268 18420
rect 12400 18380 13268 18408
rect 12400 18368 12406 18380
rect 13262 18368 13268 18380
rect 13320 18368 13326 18420
rect 13354 18368 13360 18420
rect 13412 18408 13418 18420
rect 15289 18411 15347 18417
rect 13412 18380 15056 18408
rect 13412 18368 13418 18380
rect 6641 18343 6699 18349
rect 6641 18309 6653 18343
rect 6687 18340 6699 18343
rect 8202 18340 8208 18352
rect 6687 18312 8208 18340
rect 6687 18309 6699 18312
rect 6641 18303 6699 18309
rect 8202 18300 8208 18312
rect 8260 18300 8266 18352
rect 8294 18300 8300 18352
rect 8352 18300 8358 18352
rect 8386 18300 8392 18352
rect 8444 18300 8450 18352
rect 9125 18343 9183 18349
rect 9125 18309 9137 18343
rect 9171 18340 9183 18343
rect 9674 18340 9680 18352
rect 9171 18312 9680 18340
rect 9171 18309 9183 18312
rect 9125 18303 9183 18309
rect 9674 18300 9680 18312
rect 9732 18340 9738 18352
rect 10686 18340 10692 18352
rect 9732 18312 10692 18340
rect 9732 18300 9738 18312
rect 10686 18300 10692 18312
rect 10744 18300 10750 18352
rect 12454 18343 12512 18349
rect 12454 18309 12466 18343
rect 12500 18340 12512 18343
rect 13446 18340 13452 18352
rect 12500 18312 13452 18340
rect 12500 18309 12512 18312
rect 12454 18303 12512 18309
rect 13446 18300 13452 18312
rect 13504 18300 13510 18352
rect 13906 18300 13912 18352
rect 13964 18300 13970 18352
rect 15028 18349 15056 18380
rect 15289 18377 15301 18411
rect 15335 18408 15347 18411
rect 16022 18408 16028 18420
rect 15335 18380 16028 18408
rect 15335 18377 15347 18380
rect 15289 18371 15347 18377
rect 16022 18368 16028 18380
rect 16080 18408 16086 18420
rect 16942 18408 16948 18420
rect 16080 18380 16948 18408
rect 16080 18368 16086 18380
rect 16942 18368 16948 18380
rect 17000 18368 17006 18420
rect 18138 18368 18144 18420
rect 18196 18368 18202 18420
rect 19610 18368 19616 18420
rect 19668 18408 19674 18420
rect 19797 18411 19855 18417
rect 19797 18408 19809 18411
rect 19668 18380 19809 18408
rect 19668 18368 19674 18380
rect 19797 18377 19809 18380
rect 19843 18408 19855 18411
rect 20898 18408 20904 18420
rect 19843 18380 20904 18408
rect 19843 18377 19855 18380
rect 19797 18371 19855 18377
rect 20898 18368 20904 18380
rect 20956 18368 20962 18420
rect 21560 18380 23060 18408
rect 15013 18343 15071 18349
rect 15013 18309 15025 18343
rect 15059 18340 15071 18343
rect 15378 18340 15384 18352
rect 15059 18312 15384 18340
rect 15059 18309 15071 18312
rect 15013 18303 15071 18309
rect 15378 18300 15384 18312
rect 15436 18300 15442 18352
rect 17862 18340 17868 18352
rect 17236 18312 17868 18340
rect 5166 18281 5172 18284
rect 5164 18272 5172 18281
rect 5092 18244 5172 18272
rect 5164 18235 5172 18244
rect 5166 18232 5172 18235
rect 5224 18232 5230 18284
rect 5537 18275 5595 18281
rect 5537 18241 5549 18275
rect 5583 18241 5595 18275
rect 5537 18235 5595 18241
rect 5552 18204 5580 18235
rect 5718 18232 5724 18284
rect 5776 18232 5782 18284
rect 6089 18275 6147 18281
rect 6089 18241 6101 18275
rect 6135 18241 6147 18275
rect 6089 18235 6147 18241
rect 5810 18204 5816 18216
rect 5552 18176 5816 18204
rect 5810 18164 5816 18176
rect 5868 18204 5874 18216
rect 6104 18204 6132 18235
rect 6362 18232 6368 18284
rect 6420 18272 6426 18284
rect 6457 18275 6515 18281
rect 6457 18272 6469 18275
rect 6420 18244 6469 18272
rect 6420 18232 6426 18244
rect 6457 18241 6469 18244
rect 6503 18241 6515 18275
rect 6457 18235 6515 18241
rect 6733 18275 6791 18281
rect 6733 18241 6745 18275
rect 6779 18241 6791 18275
rect 6733 18235 6791 18241
rect 6748 18204 6776 18235
rect 6822 18232 6828 18284
rect 6880 18281 6886 18284
rect 6880 18272 6888 18281
rect 6880 18244 6925 18272
rect 6880 18235 6888 18244
rect 6880 18232 6886 18235
rect 7558 18232 7564 18284
rect 7616 18272 7622 18284
rect 7926 18272 7932 18284
rect 7616 18244 7932 18272
rect 7616 18232 7622 18244
rect 7926 18232 7932 18244
rect 7984 18272 7990 18284
rect 8113 18275 8171 18281
rect 8113 18272 8125 18275
rect 7984 18244 8125 18272
rect 7984 18232 7990 18244
rect 8113 18241 8125 18244
rect 8159 18241 8171 18275
rect 8478 18272 8484 18284
rect 8536 18281 8542 18284
rect 8444 18244 8484 18272
rect 8113 18235 8171 18241
rect 8478 18232 8484 18244
rect 8536 18235 8544 18281
rect 8849 18275 8907 18281
rect 8849 18241 8861 18275
rect 8895 18241 8907 18275
rect 8849 18235 8907 18241
rect 8536 18232 8542 18235
rect 7834 18204 7840 18216
rect 5868 18176 7840 18204
rect 5868 18164 5874 18176
rect 7834 18164 7840 18176
rect 7892 18164 7898 18216
rect 8682 18207 8740 18213
rect 8682 18204 8694 18207
rect 8496 18176 8694 18204
rect 8496 18148 8524 18176
rect 8682 18173 8694 18176
rect 8728 18173 8740 18207
rect 8864 18204 8892 18235
rect 9030 18232 9036 18284
rect 9088 18232 9094 18284
rect 9214 18272 9220 18284
rect 9272 18281 9278 18284
rect 9180 18244 9220 18272
rect 9214 18232 9220 18244
rect 9272 18235 9280 18281
rect 10318 18272 10324 18284
rect 9329 18244 10324 18272
rect 9272 18232 9278 18235
rect 8938 18204 8944 18216
rect 8864 18176 8944 18204
rect 8682 18167 8740 18173
rect 8938 18164 8944 18176
rect 8996 18204 9002 18216
rect 9329 18204 9357 18244
rect 10318 18232 10324 18244
rect 10376 18232 10382 18284
rect 11885 18275 11943 18281
rect 11885 18241 11897 18275
rect 11931 18241 11943 18275
rect 11885 18235 11943 18241
rect 8996 18176 9357 18204
rect 9418 18207 9476 18213
rect 8996 18164 9002 18176
rect 9418 18173 9430 18207
rect 9464 18204 9476 18207
rect 9950 18204 9956 18216
rect 9464 18176 9956 18204
rect 9464 18173 9476 18176
rect 9418 18167 9476 18173
rect 9950 18164 9956 18176
rect 10008 18164 10014 18216
rect 10134 18164 10140 18216
rect 10192 18204 10198 18216
rect 11900 18204 11928 18235
rect 11974 18232 11980 18284
rect 12032 18272 12038 18284
rect 12069 18275 12127 18281
rect 12069 18272 12081 18275
rect 12032 18244 12081 18272
rect 12032 18232 12038 18244
rect 12069 18241 12081 18244
rect 12115 18241 12127 18275
rect 12069 18235 12127 18241
rect 12158 18232 12164 18284
rect 12216 18232 12222 18284
rect 12258 18275 12316 18281
rect 12258 18241 12270 18275
rect 12304 18272 12316 18275
rect 12618 18272 12624 18284
rect 12304 18244 12624 18272
rect 12304 18241 12316 18244
rect 12258 18235 12316 18241
rect 12618 18232 12624 18244
rect 12676 18232 12682 18284
rect 13170 18272 13176 18284
rect 12728 18244 13176 18272
rect 12728 18204 12756 18244
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 13354 18232 13360 18284
rect 13412 18272 13418 18284
rect 13725 18275 13783 18281
rect 13725 18272 13737 18275
rect 13412 18244 13737 18272
rect 13412 18232 13418 18244
rect 13725 18241 13737 18244
rect 13771 18241 13783 18275
rect 13725 18235 13783 18241
rect 14001 18275 14059 18281
rect 14001 18241 14013 18275
rect 14047 18241 14059 18275
rect 14001 18235 14059 18241
rect 10192 18176 12756 18204
rect 10192 18164 10198 18176
rect 12802 18164 12808 18216
rect 12860 18164 12866 18216
rect 12986 18164 12992 18216
rect 13044 18204 13050 18216
rect 13081 18207 13139 18213
rect 13081 18204 13093 18207
rect 13044 18176 13093 18204
rect 13044 18164 13050 18176
rect 13081 18173 13093 18176
rect 13127 18173 13139 18207
rect 13081 18167 13139 18173
rect 2608 18108 4108 18136
rect 4985 18139 5043 18145
rect 4985 18105 4997 18139
rect 5031 18136 5043 18139
rect 5442 18136 5448 18148
rect 5031 18108 5448 18136
rect 5031 18105 5043 18108
rect 4985 18099 5043 18105
rect 5442 18096 5448 18108
rect 5500 18096 5506 18148
rect 6822 18136 6828 18148
rect 6288 18108 6828 18136
rect 3970 18028 3976 18080
rect 4028 18068 4034 18080
rect 4525 18071 4583 18077
rect 4525 18068 4537 18071
rect 4028 18040 4537 18068
rect 4028 18028 4034 18040
rect 4525 18037 4537 18040
rect 4571 18068 4583 18071
rect 6288 18068 6316 18108
rect 6822 18096 6828 18108
rect 6880 18096 6886 18148
rect 7006 18096 7012 18148
rect 7064 18096 7070 18148
rect 8478 18096 8484 18148
rect 8536 18096 8542 18148
rect 10410 18096 10416 18148
rect 10468 18136 10474 18148
rect 14016 18136 14044 18235
rect 14090 18232 14096 18284
rect 14148 18232 14154 18284
rect 14734 18232 14740 18284
rect 14792 18232 14798 18284
rect 14918 18232 14924 18284
rect 14976 18232 14982 18284
rect 15102 18232 15108 18284
rect 15160 18232 15166 18284
rect 17236 18281 17264 18312
rect 17862 18300 17868 18312
rect 17920 18300 17926 18352
rect 18506 18300 18512 18352
rect 18564 18340 18570 18352
rect 21450 18340 21456 18352
rect 18564 18312 21456 18340
rect 18564 18300 18570 18312
rect 21450 18300 21456 18312
rect 21508 18300 21514 18352
rect 17037 18275 17095 18281
rect 17037 18241 17049 18275
rect 17083 18241 17095 18275
rect 17037 18235 17095 18241
rect 17221 18275 17279 18281
rect 17221 18241 17233 18275
rect 17267 18241 17279 18275
rect 17221 18235 17279 18241
rect 16666 18164 16672 18216
rect 16724 18204 16730 18216
rect 17052 18204 17080 18235
rect 17310 18232 17316 18284
rect 17368 18272 17374 18284
rect 17586 18272 17592 18284
rect 17368 18244 17592 18272
rect 17368 18232 17374 18244
rect 17586 18232 17592 18244
rect 17644 18232 17650 18284
rect 17678 18232 17684 18284
rect 17736 18232 17742 18284
rect 17957 18275 18015 18281
rect 17957 18241 17969 18275
rect 18003 18272 18015 18275
rect 18230 18272 18236 18284
rect 18003 18244 18236 18272
rect 18003 18241 18015 18244
rect 17957 18235 18015 18241
rect 18230 18232 18236 18244
rect 18288 18232 18294 18284
rect 19242 18232 19248 18284
rect 19300 18272 19306 18284
rect 19337 18275 19395 18281
rect 19337 18272 19349 18275
rect 19300 18244 19349 18272
rect 19300 18232 19306 18244
rect 19337 18241 19349 18244
rect 19383 18241 19395 18275
rect 19337 18235 19395 18241
rect 19610 18232 19616 18284
rect 19668 18232 19674 18284
rect 19794 18232 19800 18284
rect 19852 18272 19858 18284
rect 21560 18272 21588 18380
rect 19852 18244 21588 18272
rect 21652 18312 22508 18340
rect 19852 18232 19858 18244
rect 16724 18176 17080 18204
rect 16724 18164 16730 18176
rect 17126 18164 17132 18216
rect 17184 18204 17190 18216
rect 17770 18204 17776 18216
rect 17184 18176 17776 18204
rect 17184 18164 17190 18176
rect 17770 18164 17776 18176
rect 17828 18164 17834 18216
rect 19153 18207 19211 18213
rect 19153 18173 19165 18207
rect 19199 18204 19211 18207
rect 19429 18207 19487 18213
rect 19429 18204 19441 18207
rect 19199 18176 19441 18204
rect 19199 18173 19211 18176
rect 19153 18167 19211 18173
rect 19429 18173 19441 18176
rect 19475 18204 19487 18207
rect 19978 18204 19984 18216
rect 19475 18176 19984 18204
rect 19475 18173 19487 18176
rect 19429 18167 19487 18173
rect 19978 18164 19984 18176
rect 20036 18204 20042 18216
rect 20162 18204 20168 18216
rect 20036 18176 20168 18204
rect 20036 18164 20042 18176
rect 20162 18164 20168 18176
rect 20220 18164 20226 18216
rect 21542 18164 21548 18216
rect 21600 18204 21606 18216
rect 21652 18204 21680 18312
rect 22480 18284 22508 18312
rect 22922 18300 22928 18352
rect 22980 18300 22986 18352
rect 23032 18340 23060 18380
rect 23290 18368 23296 18420
rect 23348 18368 23354 18420
rect 24026 18368 24032 18420
rect 24084 18368 24090 18420
rect 24854 18368 24860 18420
rect 24912 18408 24918 18420
rect 25590 18408 25596 18420
rect 24912 18380 25596 18408
rect 24912 18368 24918 18380
rect 25590 18368 25596 18380
rect 25648 18408 25654 18420
rect 25648 18380 27108 18408
rect 25648 18368 25654 18380
rect 23032 18312 25360 18340
rect 22186 18232 22192 18284
rect 22244 18232 22250 18284
rect 22370 18232 22376 18284
rect 22428 18232 22434 18284
rect 22462 18232 22468 18284
rect 22520 18232 22526 18284
rect 22830 18232 22836 18284
rect 22888 18232 22894 18284
rect 22940 18272 22968 18300
rect 23109 18275 23167 18281
rect 23109 18272 23121 18275
rect 22940 18244 23121 18272
rect 23109 18241 23121 18244
rect 23155 18241 23167 18275
rect 23109 18235 23167 18241
rect 23566 18232 23572 18284
rect 23624 18232 23630 18284
rect 23845 18275 23903 18281
rect 23845 18241 23857 18275
rect 23891 18272 23903 18275
rect 24026 18272 24032 18284
rect 23891 18244 24032 18272
rect 23891 18241 23903 18244
rect 23845 18235 23903 18241
rect 24026 18232 24032 18244
rect 24084 18232 24090 18284
rect 25332 18281 25360 18312
rect 26234 18300 26240 18352
rect 26292 18340 26298 18352
rect 26292 18312 26648 18340
rect 26292 18300 26298 18312
rect 25317 18275 25375 18281
rect 25317 18241 25329 18275
rect 25363 18241 25375 18275
rect 25317 18235 25375 18241
rect 25406 18232 25412 18284
rect 25464 18232 25470 18284
rect 26142 18232 26148 18284
rect 26200 18272 26206 18284
rect 26510 18272 26516 18284
rect 26200 18244 26516 18272
rect 26200 18232 26206 18244
rect 26510 18232 26516 18244
rect 26568 18232 26574 18284
rect 26620 18272 26648 18312
rect 26970 18300 26976 18352
rect 27028 18300 27034 18352
rect 27080 18340 27108 18380
rect 27890 18368 27896 18420
rect 27948 18408 27954 18420
rect 28994 18408 29000 18420
rect 27948 18380 29000 18408
rect 27948 18368 27954 18380
rect 28994 18368 29000 18380
rect 29052 18368 29058 18420
rect 29733 18411 29791 18417
rect 29196 18380 29408 18408
rect 27080 18312 28396 18340
rect 27249 18275 27307 18281
rect 27249 18272 27261 18275
rect 26620 18244 27261 18272
rect 27249 18241 27261 18244
rect 27295 18272 27307 18275
rect 28258 18272 28264 18284
rect 27295 18244 28264 18272
rect 27295 18241 27307 18244
rect 27249 18235 27307 18241
rect 28258 18232 28264 18244
rect 28316 18232 28322 18284
rect 28368 18272 28396 18312
rect 28534 18300 28540 18352
rect 28592 18340 28598 18352
rect 29196 18340 29224 18380
rect 28592 18312 29224 18340
rect 28592 18300 28598 18312
rect 29270 18300 29276 18352
rect 29328 18349 29334 18352
rect 29328 18303 29338 18349
rect 29380 18340 29408 18380
rect 29733 18377 29745 18411
rect 29779 18408 29791 18411
rect 30742 18408 30748 18420
rect 29779 18380 30748 18408
rect 29779 18377 29791 18380
rect 29733 18371 29791 18377
rect 30742 18368 30748 18380
rect 30800 18368 30806 18420
rect 31665 18411 31723 18417
rect 31665 18377 31677 18411
rect 31711 18377 31723 18411
rect 31665 18371 31723 18377
rect 31680 18340 31708 18371
rect 32582 18368 32588 18420
rect 32640 18368 32646 18420
rect 34348 18380 34560 18408
rect 32125 18343 32183 18349
rect 32125 18340 32137 18343
rect 29380 18312 31616 18340
rect 31680 18312 32137 18340
rect 29328 18300 29334 18303
rect 28368 18262 29040 18272
rect 29104 18262 29500 18272
rect 28368 18244 29500 18262
rect 29012 18234 29132 18244
rect 21600 18176 21680 18204
rect 21600 18164 21606 18176
rect 22922 18164 22928 18216
rect 22980 18164 22986 18216
rect 23382 18164 23388 18216
rect 23440 18204 23446 18216
rect 23661 18207 23719 18213
rect 23661 18204 23673 18207
rect 23440 18176 23673 18204
rect 23440 18164 23446 18176
rect 23661 18173 23673 18176
rect 23707 18173 23719 18207
rect 23661 18167 23719 18173
rect 27062 18164 27068 18216
rect 27120 18164 27126 18216
rect 28442 18204 28448 18216
rect 27264 18176 28448 18204
rect 27264 18148 27292 18176
rect 28442 18164 28448 18176
rect 28500 18164 28506 18216
rect 29362 18164 29368 18216
rect 29420 18164 29426 18216
rect 29472 18204 29500 18244
rect 29546 18232 29552 18284
rect 29604 18232 29610 18284
rect 31202 18232 31208 18284
rect 31260 18232 31266 18284
rect 31386 18232 31392 18284
rect 31444 18272 31450 18284
rect 31481 18275 31539 18281
rect 31481 18272 31493 18275
rect 31444 18244 31493 18272
rect 31444 18232 31450 18244
rect 31481 18241 31493 18244
rect 31527 18241 31539 18275
rect 31588 18272 31616 18312
rect 32125 18309 32137 18312
rect 32171 18309 32183 18343
rect 32125 18303 32183 18309
rect 32950 18300 32956 18352
rect 33008 18340 33014 18352
rect 34348 18340 34376 18380
rect 33008 18312 34376 18340
rect 33008 18300 33014 18312
rect 34532 18303 34560 18380
rect 37090 18368 37096 18420
rect 37148 18368 37154 18420
rect 40862 18368 40868 18420
rect 40920 18368 40926 18420
rect 41598 18368 41604 18420
rect 41656 18368 41662 18420
rect 34517 18297 34575 18303
rect 36630 18300 36636 18352
rect 36688 18300 36694 18352
rect 41322 18300 41328 18352
rect 41380 18340 41386 18352
rect 41380 18312 42196 18340
rect 41380 18300 41386 18312
rect 31662 18272 31668 18284
rect 31588 18244 31668 18272
rect 31481 18235 31539 18241
rect 31662 18232 31668 18244
rect 31720 18232 31726 18284
rect 32306 18232 32312 18284
rect 32364 18232 32370 18284
rect 32401 18275 32459 18281
rect 32401 18241 32413 18275
rect 32447 18272 32459 18275
rect 32766 18272 32772 18284
rect 32447 18244 32772 18272
rect 32447 18241 32459 18244
rect 32401 18235 32459 18241
rect 32766 18232 32772 18244
rect 32824 18232 32830 18284
rect 32876 18244 33456 18272
rect 31297 18207 31355 18213
rect 31297 18204 31309 18207
rect 29472 18176 31309 18204
rect 31297 18173 31309 18176
rect 31343 18173 31355 18207
rect 31297 18167 31355 18173
rect 10468 18108 14044 18136
rect 14277 18139 14335 18145
rect 10468 18096 10474 18108
rect 14277 18105 14289 18139
rect 14323 18136 14335 18139
rect 14323 18108 22600 18136
rect 14323 18105 14335 18108
rect 14277 18099 14335 18105
rect 4571 18040 6316 18068
rect 4571 18037 4583 18040
rect 4525 18031 4583 18037
rect 6362 18028 6368 18080
rect 6420 18068 6426 18080
rect 12158 18068 12164 18080
rect 6420 18040 12164 18068
rect 6420 18028 6426 18040
rect 12158 18028 12164 18040
rect 12216 18028 12222 18080
rect 12986 18028 12992 18080
rect 13044 18068 13050 18080
rect 14090 18068 14096 18080
rect 13044 18040 14096 18068
rect 13044 18028 13050 18040
rect 14090 18028 14096 18040
rect 14148 18028 14154 18080
rect 16850 18028 16856 18080
rect 16908 18068 16914 18080
rect 17037 18071 17095 18077
rect 17037 18068 17049 18071
rect 16908 18040 17049 18068
rect 16908 18028 16914 18040
rect 17037 18037 17049 18040
rect 17083 18037 17095 18071
rect 17037 18031 17095 18037
rect 17218 18028 17224 18080
rect 17276 18068 17282 18080
rect 17497 18071 17555 18077
rect 17497 18068 17509 18071
rect 17276 18040 17509 18068
rect 17276 18028 17282 18040
rect 17497 18037 17509 18040
rect 17543 18037 17555 18071
rect 17497 18031 17555 18037
rect 17586 18028 17592 18080
rect 17644 18068 17650 18080
rect 17681 18071 17739 18077
rect 17681 18068 17693 18071
rect 17644 18040 17693 18068
rect 17644 18028 17650 18040
rect 17681 18037 17693 18040
rect 17727 18037 17739 18071
rect 17681 18031 17739 18037
rect 19334 18028 19340 18080
rect 19392 18068 19398 18080
rect 19886 18068 19892 18080
rect 19392 18040 19892 18068
rect 19392 18028 19398 18040
rect 19886 18028 19892 18040
rect 19944 18028 19950 18080
rect 22370 18028 22376 18080
rect 22428 18028 22434 18080
rect 22572 18068 22600 18108
rect 22646 18096 22652 18148
rect 22704 18096 22710 18148
rect 27246 18096 27252 18148
rect 27304 18096 27310 18148
rect 27614 18096 27620 18148
rect 27672 18136 27678 18148
rect 28718 18136 28724 18148
rect 27672 18108 28724 18136
rect 27672 18096 27678 18108
rect 28718 18096 28724 18108
rect 28776 18136 28782 18148
rect 29089 18139 29147 18145
rect 29089 18136 29101 18139
rect 28776 18108 29101 18136
rect 28776 18096 28782 18108
rect 29089 18105 29101 18108
rect 29135 18136 29147 18139
rect 29380 18136 29408 18164
rect 32876 18136 32904 18244
rect 33134 18164 33140 18216
rect 33192 18204 33198 18216
rect 33318 18204 33324 18216
rect 33192 18176 33324 18204
rect 33192 18164 33198 18176
rect 33318 18164 33324 18176
rect 33376 18164 33382 18216
rect 33428 18204 33456 18244
rect 34054 18232 34060 18284
rect 34112 18272 34118 18284
rect 34149 18275 34207 18281
rect 34149 18272 34161 18275
rect 34112 18244 34161 18272
rect 34112 18232 34118 18244
rect 34149 18241 34161 18244
rect 34195 18241 34207 18275
rect 34149 18235 34207 18241
rect 34238 18232 34244 18284
rect 34296 18232 34302 18284
rect 34425 18275 34483 18281
rect 34425 18241 34437 18275
rect 34471 18241 34483 18275
rect 34517 18263 34529 18297
rect 34563 18263 34575 18297
rect 34517 18257 34575 18263
rect 34425 18235 34483 18241
rect 33428 18176 34192 18204
rect 29135 18108 29408 18136
rect 31312 18108 32904 18136
rect 29135 18105 29147 18108
rect 29089 18099 29147 18105
rect 23014 18068 23020 18080
rect 22572 18040 23020 18068
rect 23014 18028 23020 18040
rect 23072 18028 23078 18080
rect 23109 18071 23167 18077
rect 23109 18037 23121 18071
rect 23155 18068 23167 18071
rect 23474 18068 23480 18080
rect 23155 18040 23480 18068
rect 23155 18037 23167 18040
rect 23109 18031 23167 18037
rect 23474 18028 23480 18040
rect 23532 18028 23538 18080
rect 23750 18028 23756 18080
rect 23808 18028 23814 18080
rect 25406 18028 25412 18080
rect 25464 18028 25470 18080
rect 25682 18028 25688 18080
rect 25740 18028 25746 18080
rect 26878 18028 26884 18080
rect 26936 18068 26942 18080
rect 26973 18071 27031 18077
rect 26973 18068 26985 18071
rect 26936 18040 26985 18068
rect 26936 18028 26942 18040
rect 26973 18037 26985 18040
rect 27019 18037 27031 18071
rect 26973 18031 27031 18037
rect 27433 18071 27491 18077
rect 27433 18037 27445 18071
rect 27479 18068 27491 18071
rect 27706 18068 27712 18080
rect 27479 18040 27712 18068
rect 27479 18037 27491 18040
rect 27433 18031 27491 18037
rect 27706 18028 27712 18040
rect 27764 18028 27770 18080
rect 29178 18028 29184 18080
rect 29236 18068 29242 18080
rect 31312 18077 31340 18108
rect 33042 18096 33048 18148
rect 33100 18136 33106 18148
rect 34054 18136 34060 18148
rect 33100 18108 34060 18136
rect 33100 18096 33106 18108
rect 34054 18096 34060 18108
rect 34112 18096 34118 18148
rect 34164 18136 34192 18176
rect 34440 18136 34468 18235
rect 34698 18232 34704 18284
rect 34756 18232 34762 18284
rect 36906 18232 36912 18284
rect 36964 18232 36970 18284
rect 37366 18232 37372 18284
rect 37424 18232 37430 18284
rect 37458 18232 37464 18284
rect 37516 18272 37522 18284
rect 37645 18275 37703 18281
rect 37645 18272 37657 18275
rect 37516 18244 37657 18272
rect 37516 18232 37522 18244
rect 37645 18241 37657 18244
rect 37691 18241 37703 18275
rect 37645 18235 37703 18241
rect 41509 18275 41567 18281
rect 41509 18241 41521 18275
rect 41555 18272 41567 18275
rect 41690 18272 41696 18284
rect 41555 18244 41696 18272
rect 41555 18241 41567 18244
rect 41509 18235 41567 18241
rect 41690 18232 41696 18244
rect 41748 18232 41754 18284
rect 41782 18232 41788 18284
rect 41840 18232 41846 18284
rect 41874 18232 41880 18284
rect 41932 18232 41938 18284
rect 42168 18281 42196 18312
rect 42153 18275 42211 18281
rect 42153 18241 42165 18275
rect 42199 18241 42211 18275
rect 42153 18235 42211 18241
rect 43162 18232 43168 18284
rect 43220 18272 43226 18284
rect 44269 18275 44327 18281
rect 44269 18272 44281 18275
rect 43220 18244 44281 18272
rect 43220 18232 43226 18244
rect 44269 18241 44281 18244
rect 44315 18241 44327 18275
rect 44269 18235 44327 18241
rect 34882 18164 34888 18216
rect 34940 18204 34946 18216
rect 36725 18207 36783 18213
rect 36725 18204 36737 18207
rect 34940 18176 36737 18204
rect 34940 18164 34946 18176
rect 36725 18173 36737 18176
rect 36771 18173 36783 18207
rect 36725 18167 36783 18173
rect 37274 18164 37280 18216
rect 37332 18204 37338 18216
rect 37737 18207 37795 18213
rect 37737 18204 37749 18207
rect 37332 18176 37749 18204
rect 37332 18164 37338 18176
rect 37737 18173 37749 18176
rect 37783 18173 37795 18207
rect 37737 18167 37795 18173
rect 40310 18164 40316 18216
rect 40368 18164 40374 18216
rect 42061 18207 42119 18213
rect 42061 18173 42073 18207
rect 42107 18204 42119 18207
rect 42518 18204 42524 18216
rect 42107 18176 42524 18204
rect 42107 18173 42119 18176
rect 42061 18167 42119 18173
rect 42518 18164 42524 18176
rect 42576 18164 42582 18216
rect 35342 18136 35348 18148
rect 34164 18108 35348 18136
rect 35342 18096 35348 18108
rect 35400 18096 35406 18148
rect 37369 18139 37427 18145
rect 37369 18105 37381 18139
rect 37415 18136 37427 18139
rect 38194 18136 38200 18148
rect 37415 18108 38200 18136
rect 37415 18105 37427 18108
rect 37369 18099 37427 18105
rect 38194 18096 38200 18108
rect 38252 18096 38258 18148
rect 29273 18071 29331 18077
rect 29273 18068 29285 18071
rect 29236 18040 29285 18068
rect 29236 18028 29242 18040
rect 29273 18037 29285 18040
rect 29319 18037 29331 18071
rect 29273 18031 29331 18037
rect 31297 18071 31355 18077
rect 31297 18037 31309 18071
rect 31343 18037 31355 18071
rect 31297 18031 31355 18037
rect 31662 18028 31668 18080
rect 31720 18068 31726 18080
rect 32125 18071 32183 18077
rect 32125 18068 32137 18071
rect 31720 18040 32137 18068
rect 31720 18028 31726 18040
rect 32125 18037 32137 18040
rect 32171 18037 32183 18071
rect 32125 18031 32183 18037
rect 32306 18028 32312 18080
rect 32364 18068 32370 18080
rect 33778 18068 33784 18080
rect 32364 18040 33784 18068
rect 32364 18028 32370 18040
rect 33778 18028 33784 18040
rect 33836 18028 33842 18080
rect 33962 18028 33968 18080
rect 34020 18028 34026 18080
rect 34146 18028 34152 18080
rect 34204 18028 34210 18080
rect 34514 18028 34520 18080
rect 34572 18028 34578 18080
rect 34698 18028 34704 18080
rect 34756 18068 34762 18080
rect 34882 18068 34888 18080
rect 34756 18040 34888 18068
rect 34756 18028 34762 18040
rect 34882 18028 34888 18040
rect 34940 18028 34946 18080
rect 34974 18028 34980 18080
rect 35032 18068 35038 18080
rect 36633 18071 36691 18077
rect 36633 18068 36645 18071
rect 35032 18040 36645 18068
rect 35032 18028 35038 18040
rect 36633 18037 36645 18040
rect 36679 18037 36691 18071
rect 36633 18031 36691 18037
rect 37458 18028 37464 18080
rect 37516 18068 37522 18080
rect 37553 18071 37611 18077
rect 37553 18068 37565 18071
rect 37516 18040 37565 18068
rect 37516 18028 37522 18040
rect 37553 18037 37565 18040
rect 37599 18068 37611 18071
rect 38102 18068 38108 18080
rect 37599 18040 38108 18068
rect 37599 18037 37611 18040
rect 37553 18031 37611 18037
rect 38102 18028 38108 18040
rect 38160 18028 38166 18080
rect 38654 18028 38660 18080
rect 38712 18068 38718 18080
rect 39669 18071 39727 18077
rect 39669 18068 39681 18071
rect 38712 18040 39681 18068
rect 38712 18028 38718 18040
rect 39669 18037 39681 18040
rect 39715 18037 39727 18071
rect 39669 18031 39727 18037
rect 41782 18028 41788 18080
rect 41840 18068 41846 18080
rect 42518 18068 42524 18080
rect 41840 18040 42524 18068
rect 41840 18028 41846 18040
rect 42518 18028 42524 18040
rect 42576 18028 42582 18080
rect 44082 18028 44088 18080
rect 44140 18068 44146 18080
rect 44453 18071 44511 18077
rect 44453 18068 44465 18071
rect 44140 18040 44465 18068
rect 44140 18028 44146 18040
rect 44453 18037 44465 18040
rect 44499 18037 44511 18071
rect 44453 18031 44511 18037
rect 1104 17978 44896 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 44896 17978
rect 1104 17904 44896 17926
rect 2406 17824 2412 17876
rect 2464 17824 2470 17876
rect 2498 17824 2504 17876
rect 2556 17864 2562 17876
rect 2556 17836 2774 17864
rect 2556 17824 2562 17836
rect 2590 17620 2596 17672
rect 2648 17620 2654 17672
rect 2746 17524 2774 17836
rect 3050 17824 3056 17876
rect 3108 17864 3114 17876
rect 3145 17867 3203 17873
rect 3145 17864 3157 17867
rect 3108 17836 3157 17864
rect 3108 17824 3114 17836
rect 3145 17833 3157 17836
rect 3191 17864 3203 17867
rect 3191 17836 4752 17864
rect 3191 17833 3203 17836
rect 3145 17827 3203 17833
rect 4433 17799 4491 17805
rect 4433 17765 4445 17799
rect 4479 17765 4491 17799
rect 4724 17796 4752 17836
rect 4798 17824 4804 17876
rect 4856 17864 4862 17876
rect 5353 17867 5411 17873
rect 5353 17864 5365 17867
rect 4856 17836 5365 17864
rect 4856 17824 4862 17836
rect 5353 17833 5365 17836
rect 5399 17833 5411 17867
rect 5353 17827 5411 17833
rect 6270 17824 6276 17876
rect 6328 17864 6334 17876
rect 6328 17836 7236 17864
rect 6328 17824 6334 17836
rect 6546 17796 6552 17808
rect 4724 17768 6552 17796
rect 4433 17759 4491 17765
rect 4448 17728 4476 17759
rect 6546 17756 6552 17768
rect 6604 17756 6610 17808
rect 6733 17799 6791 17805
rect 6733 17765 6745 17799
rect 6779 17796 6791 17799
rect 6914 17796 6920 17808
rect 6779 17768 6920 17796
rect 6779 17765 6791 17768
rect 6733 17759 6791 17765
rect 6914 17756 6920 17768
rect 6972 17756 6978 17808
rect 7208 17796 7236 17836
rect 7282 17824 7288 17876
rect 7340 17864 7346 17876
rect 7742 17864 7748 17876
rect 7340 17836 7748 17864
rect 7340 17824 7346 17836
rect 7742 17824 7748 17836
rect 7800 17824 7806 17876
rect 8018 17824 8024 17876
rect 8076 17864 8082 17876
rect 8113 17867 8171 17873
rect 8113 17864 8125 17867
rect 8076 17836 8125 17864
rect 8076 17824 8082 17836
rect 8113 17833 8125 17836
rect 8159 17833 8171 17867
rect 8113 17827 8171 17833
rect 8202 17824 8208 17876
rect 8260 17864 8266 17876
rect 9674 17864 9680 17876
rect 8260 17836 9680 17864
rect 8260 17824 8266 17836
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 9950 17824 9956 17876
rect 10008 17824 10014 17876
rect 10318 17824 10324 17876
rect 10376 17864 10382 17876
rect 10962 17864 10968 17876
rect 10376 17836 10968 17864
rect 10376 17824 10382 17836
rect 10962 17824 10968 17836
rect 11020 17824 11026 17876
rect 11698 17824 11704 17876
rect 11756 17864 11762 17876
rect 12618 17864 12624 17876
rect 11756 17836 12624 17864
rect 11756 17824 11762 17836
rect 12618 17824 12624 17836
rect 12676 17864 12682 17876
rect 13538 17864 13544 17876
rect 12676 17836 13544 17864
rect 12676 17824 12682 17836
rect 13538 17824 13544 17836
rect 13596 17824 13602 17876
rect 15194 17824 15200 17876
rect 15252 17824 15258 17876
rect 16298 17824 16304 17876
rect 16356 17864 16362 17876
rect 16669 17867 16727 17873
rect 16669 17864 16681 17867
rect 16356 17836 16681 17864
rect 16356 17824 16362 17836
rect 16669 17833 16681 17836
rect 16715 17833 16727 17867
rect 16669 17827 16727 17833
rect 17129 17867 17187 17873
rect 17129 17833 17141 17867
rect 17175 17864 17187 17867
rect 22830 17864 22836 17876
rect 17175 17836 22836 17864
rect 17175 17833 17187 17836
rect 17129 17827 17187 17833
rect 22830 17824 22836 17836
rect 22888 17824 22894 17876
rect 22925 17867 22983 17873
rect 22925 17833 22937 17867
rect 22971 17833 22983 17867
rect 22925 17827 22983 17833
rect 23385 17867 23443 17873
rect 23385 17833 23397 17867
rect 23431 17864 23443 17867
rect 23566 17864 23572 17876
rect 23431 17836 23572 17864
rect 23431 17833 23443 17836
rect 23385 17827 23443 17833
rect 8386 17796 8392 17808
rect 7208 17768 8392 17796
rect 8386 17756 8392 17768
rect 8444 17796 8450 17808
rect 12253 17799 12311 17805
rect 8444 17768 12112 17796
rect 8444 17756 8450 17768
rect 12084 17728 12112 17768
rect 12253 17765 12265 17799
rect 12299 17796 12311 17799
rect 13722 17796 13728 17808
rect 12299 17768 13728 17796
rect 12299 17765 12311 17768
rect 12253 17759 12311 17765
rect 13722 17756 13728 17768
rect 13780 17756 13786 17808
rect 17770 17756 17776 17808
rect 17828 17796 17834 17808
rect 22940 17796 22968 17827
rect 23566 17824 23572 17836
rect 23624 17824 23630 17876
rect 24026 17824 24032 17876
rect 24084 17864 24090 17876
rect 24084 17836 25820 17864
rect 24084 17824 24090 17836
rect 24946 17796 24952 17808
rect 17828 17768 24952 17796
rect 17828 17756 17834 17768
rect 24946 17756 24952 17768
rect 25004 17756 25010 17808
rect 25792 17796 25820 17836
rect 25958 17824 25964 17876
rect 26016 17824 26022 17876
rect 26234 17824 26240 17876
rect 26292 17824 26298 17876
rect 26970 17824 26976 17876
rect 27028 17824 27034 17876
rect 27522 17824 27528 17876
rect 27580 17864 27586 17876
rect 27709 17867 27767 17873
rect 27709 17864 27721 17867
rect 27580 17836 27721 17864
rect 27580 17824 27586 17836
rect 27709 17833 27721 17836
rect 27755 17833 27767 17867
rect 28166 17864 28172 17876
rect 27709 17827 27767 17833
rect 27908 17836 28172 17864
rect 27246 17796 27252 17808
rect 25792 17768 27252 17796
rect 4448 17700 11100 17728
rect 2866 17620 2872 17672
rect 2924 17660 2930 17672
rect 2961 17663 3019 17669
rect 2961 17660 2973 17663
rect 2924 17632 2973 17660
rect 2924 17620 2930 17632
rect 2961 17629 2973 17632
rect 3007 17629 3019 17663
rect 2961 17623 3019 17629
rect 3326 17620 3332 17672
rect 3384 17620 3390 17672
rect 4249 17663 4307 17669
rect 4249 17629 4261 17663
rect 4295 17660 4307 17663
rect 4614 17660 4620 17672
rect 4295 17632 4620 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 4614 17620 4620 17632
rect 4672 17620 4678 17672
rect 4706 17620 4712 17672
rect 4764 17660 4770 17672
rect 4890 17660 4896 17672
rect 4764 17632 4896 17660
rect 4764 17620 4770 17632
rect 4890 17620 4896 17632
rect 4948 17620 4954 17672
rect 5537 17663 5595 17669
rect 5537 17629 5549 17663
rect 5583 17660 5595 17663
rect 5994 17660 6000 17672
rect 5583 17632 6000 17660
rect 5583 17629 5595 17632
rect 5537 17623 5595 17629
rect 5994 17620 6000 17632
rect 6052 17620 6058 17672
rect 6178 17620 6184 17672
rect 6236 17620 6242 17672
rect 6454 17660 6460 17672
rect 6288 17632 6460 17660
rect 3234 17552 3240 17604
rect 3292 17592 3298 17604
rect 5721 17595 5779 17601
rect 5721 17592 5733 17595
rect 3292 17564 5733 17592
rect 3292 17552 3298 17564
rect 5721 17561 5733 17564
rect 5767 17561 5779 17595
rect 5721 17555 5779 17561
rect 5902 17552 5908 17604
rect 5960 17592 5966 17604
rect 6288 17592 6316 17632
rect 6454 17620 6460 17632
rect 6512 17620 6518 17672
rect 6601 17663 6659 17669
rect 6601 17629 6613 17663
rect 6647 17660 6659 17663
rect 6730 17660 6736 17672
rect 6647 17632 6736 17660
rect 6647 17629 6659 17632
rect 6601 17623 6659 17629
rect 6730 17620 6736 17632
rect 6788 17620 6794 17672
rect 7469 17663 7527 17669
rect 7469 17629 7481 17663
rect 7515 17660 7527 17663
rect 7650 17660 7656 17672
rect 7515 17632 7656 17660
rect 7515 17629 7527 17632
rect 7469 17623 7527 17629
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 7745 17663 7803 17669
rect 7745 17629 7757 17663
rect 7791 17660 7803 17663
rect 8202 17660 8208 17672
rect 7791 17632 8208 17660
rect 7791 17629 7803 17632
rect 7745 17623 7803 17629
rect 8202 17620 8208 17632
rect 8260 17620 8266 17672
rect 9401 17663 9459 17669
rect 9401 17660 9413 17663
rect 8404 17632 9413 17660
rect 5960 17564 6316 17592
rect 5960 17552 5966 17564
rect 6362 17552 6368 17604
rect 6420 17552 6426 17604
rect 7834 17552 7840 17604
rect 7892 17552 7898 17604
rect 7954 17595 8012 17601
rect 7954 17561 7966 17595
rect 8000 17592 8012 17595
rect 8294 17592 8300 17604
rect 8000 17564 8300 17592
rect 8000 17561 8012 17564
rect 7954 17555 8012 17561
rect 8294 17552 8300 17564
rect 8352 17552 8358 17604
rect 3513 17527 3571 17533
rect 3513 17524 3525 17527
rect 2746 17496 3525 17524
rect 3513 17493 3525 17496
rect 3559 17524 3571 17527
rect 7190 17524 7196 17536
rect 3559 17496 7196 17524
rect 3559 17493 3571 17496
rect 3513 17487 3571 17493
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 7282 17484 7288 17536
rect 7340 17524 7346 17536
rect 8404 17524 8432 17632
rect 7340 17496 8432 17524
rect 9140 17524 9168 17632
rect 9401 17629 9413 17632
rect 9447 17629 9459 17663
rect 9401 17623 9459 17629
rect 9766 17620 9772 17672
rect 9824 17669 9830 17672
rect 9824 17660 9832 17669
rect 11072 17660 11100 17700
rect 12084 17700 12848 17728
rect 9824 17632 9869 17660
rect 11072 17632 11652 17660
rect 9824 17623 9832 17632
rect 9824 17620 9830 17623
rect 9214 17552 9220 17604
rect 9272 17592 9278 17604
rect 9490 17592 9496 17604
rect 9272 17564 9496 17592
rect 9272 17552 9278 17564
rect 9490 17552 9496 17564
rect 9548 17592 9554 17604
rect 9585 17595 9643 17601
rect 9585 17592 9597 17595
rect 9548 17564 9597 17592
rect 9548 17552 9554 17564
rect 9585 17561 9597 17564
rect 9631 17561 9643 17595
rect 9585 17555 9643 17561
rect 9677 17595 9735 17601
rect 9677 17561 9689 17595
rect 9723 17592 9735 17595
rect 11330 17592 11336 17604
rect 9723 17564 11336 17592
rect 9723 17561 9735 17564
rect 9677 17555 9735 17561
rect 11330 17552 11336 17564
rect 11388 17592 11394 17604
rect 11514 17592 11520 17604
rect 11388 17564 11520 17592
rect 11388 17552 11394 17564
rect 11514 17552 11520 17564
rect 11572 17552 11578 17604
rect 9950 17524 9956 17536
rect 9140 17496 9956 17524
rect 7340 17484 7346 17496
rect 9950 17484 9956 17496
rect 10008 17484 10014 17536
rect 11624 17524 11652 17632
rect 11698 17620 11704 17672
rect 11756 17620 11762 17672
rect 11974 17620 11980 17672
rect 12032 17620 12038 17672
rect 12084 17669 12112 17700
rect 12074 17663 12132 17669
rect 12074 17629 12086 17663
rect 12120 17629 12132 17663
rect 12074 17623 12132 17629
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17629 12495 17663
rect 12437 17623 12495 17629
rect 12713 17663 12771 17669
rect 12713 17629 12725 17663
rect 12759 17629 12771 17663
rect 12713 17623 12771 17629
rect 11882 17552 11888 17604
rect 11940 17552 11946 17604
rect 12452 17592 12480 17623
rect 11992 17564 12480 17592
rect 11992 17524 12020 17564
rect 11624 17496 12020 17524
rect 12158 17484 12164 17536
rect 12216 17524 12222 17536
rect 12728 17524 12756 17623
rect 12820 17592 12848 17700
rect 12894 17688 12900 17740
rect 12952 17728 12958 17740
rect 16761 17731 16819 17737
rect 16761 17728 16773 17731
rect 12952 17700 16773 17728
rect 12952 17688 12958 17700
rect 16761 17697 16773 17700
rect 16807 17697 16819 17731
rect 16761 17691 16819 17697
rect 17034 17688 17040 17740
rect 17092 17728 17098 17740
rect 17092 17700 19748 17728
rect 17092 17688 17098 17700
rect 12986 17620 12992 17672
rect 13044 17660 13050 17672
rect 13044 17632 15240 17660
rect 13044 17620 13050 17632
rect 13354 17592 13360 17604
rect 12820 17564 13360 17592
rect 13354 17552 13360 17564
rect 13412 17552 13418 17604
rect 14918 17552 14924 17604
rect 14976 17552 14982 17604
rect 15102 17552 15108 17604
rect 15160 17552 15166 17604
rect 15212 17592 15240 17632
rect 15286 17620 15292 17672
rect 15344 17660 15350 17672
rect 16114 17660 16120 17672
rect 15344 17632 16120 17660
rect 15344 17620 15350 17632
rect 16114 17620 16120 17632
rect 16172 17620 16178 17672
rect 16574 17620 16580 17672
rect 16632 17660 16638 17672
rect 16669 17663 16727 17669
rect 16669 17660 16681 17663
rect 16632 17632 16681 17660
rect 16632 17620 16638 17632
rect 16669 17629 16681 17632
rect 16715 17629 16727 17663
rect 16669 17623 16727 17629
rect 16850 17620 16856 17672
rect 16908 17660 16914 17672
rect 16945 17663 17003 17669
rect 16945 17660 16957 17663
rect 16908 17632 16957 17660
rect 16908 17620 16914 17632
rect 16945 17629 16957 17632
rect 16991 17629 17003 17663
rect 16945 17623 17003 17629
rect 19610 17620 19616 17672
rect 19668 17620 19674 17672
rect 19720 17660 19748 17700
rect 19794 17688 19800 17740
rect 19852 17688 19858 17740
rect 23014 17688 23020 17740
rect 23072 17688 23078 17740
rect 26142 17728 26148 17740
rect 23124 17700 26148 17728
rect 20254 17660 20260 17672
rect 19720 17632 20260 17660
rect 20254 17620 20260 17632
rect 20312 17620 20318 17672
rect 22186 17620 22192 17672
rect 22244 17620 22250 17672
rect 22370 17620 22376 17672
rect 22428 17660 22434 17672
rect 22554 17660 22560 17672
rect 22428 17632 22560 17660
rect 22428 17620 22434 17632
rect 22554 17620 22560 17632
rect 22612 17660 22618 17672
rect 23124 17660 23152 17700
rect 26142 17688 26148 17700
rect 26200 17688 26206 17740
rect 22612 17632 23152 17660
rect 22612 17620 22618 17632
rect 23198 17620 23204 17672
rect 23256 17620 23262 17672
rect 25222 17620 25228 17672
rect 25280 17660 25286 17672
rect 25593 17663 25651 17669
rect 25593 17660 25605 17663
rect 25280 17632 25605 17660
rect 25280 17620 25286 17632
rect 25593 17629 25605 17632
rect 25639 17629 25651 17663
rect 25593 17623 25651 17629
rect 25682 17620 25688 17672
rect 25740 17660 25746 17672
rect 26237 17663 26295 17669
rect 26237 17660 26249 17663
rect 25740 17632 26249 17660
rect 25740 17620 25746 17632
rect 26237 17629 26249 17632
rect 26283 17629 26295 17663
rect 26237 17623 26295 17629
rect 26326 17620 26332 17672
rect 26384 17660 26390 17672
rect 26528 17669 26556 17768
rect 27246 17756 27252 17768
rect 27304 17756 27310 17808
rect 27614 17728 27620 17740
rect 27172 17700 27620 17728
rect 27172 17669 27200 17700
rect 27614 17688 27620 17700
rect 27672 17688 27678 17740
rect 27908 17737 27936 17836
rect 28166 17824 28172 17836
rect 28224 17864 28230 17876
rect 29730 17864 29736 17876
rect 28224 17836 29736 17864
rect 28224 17824 28230 17836
rect 29730 17824 29736 17836
rect 29788 17824 29794 17876
rect 29822 17824 29828 17876
rect 29880 17824 29886 17876
rect 31386 17824 31392 17876
rect 31444 17824 31450 17876
rect 31941 17867 31999 17873
rect 31941 17833 31953 17867
rect 31987 17864 31999 17867
rect 32306 17864 32312 17876
rect 31987 17836 32312 17864
rect 31987 17833 31999 17836
rect 31941 17827 31999 17833
rect 32306 17824 32312 17836
rect 32364 17824 32370 17876
rect 32493 17867 32551 17873
rect 32493 17833 32505 17867
rect 32539 17864 32551 17867
rect 32950 17864 32956 17876
rect 32539 17836 32956 17864
rect 32539 17833 32551 17836
rect 32493 17827 32551 17833
rect 32950 17824 32956 17836
rect 33008 17824 33014 17876
rect 33229 17867 33287 17873
rect 33229 17833 33241 17867
rect 33275 17833 33287 17867
rect 33229 17827 33287 17833
rect 27982 17756 27988 17808
rect 28040 17796 28046 17808
rect 33244 17796 33272 17827
rect 33410 17824 33416 17876
rect 33468 17864 33474 17876
rect 33870 17864 33876 17876
rect 33468 17836 33876 17864
rect 33468 17824 33474 17836
rect 33870 17824 33876 17836
rect 33928 17824 33934 17876
rect 34054 17824 34060 17876
rect 34112 17824 34118 17876
rect 34238 17824 34244 17876
rect 34296 17864 34302 17876
rect 35345 17867 35403 17873
rect 35345 17864 35357 17867
rect 34296 17836 35357 17864
rect 34296 17824 34302 17836
rect 35345 17833 35357 17836
rect 35391 17833 35403 17867
rect 35345 17827 35403 17833
rect 35713 17867 35771 17873
rect 35713 17833 35725 17867
rect 35759 17864 35771 17867
rect 36173 17867 36231 17873
rect 36173 17864 36185 17867
rect 35759 17836 36185 17864
rect 35759 17833 35771 17836
rect 35713 17827 35771 17833
rect 36173 17833 36185 17836
rect 36219 17833 36231 17867
rect 36173 17827 36231 17833
rect 36262 17824 36268 17876
rect 36320 17824 36326 17876
rect 37182 17824 37188 17876
rect 37240 17864 37246 17876
rect 37277 17867 37335 17873
rect 37277 17864 37289 17867
rect 37240 17836 37289 17864
rect 37240 17824 37246 17836
rect 37277 17833 37289 17836
rect 37323 17833 37335 17867
rect 37277 17827 37335 17833
rect 37737 17867 37795 17873
rect 37737 17833 37749 17867
rect 37783 17864 37795 17867
rect 38746 17864 38752 17876
rect 37783 17836 38752 17864
rect 37783 17833 37795 17836
rect 37737 17827 37795 17833
rect 38746 17824 38752 17836
rect 38804 17824 38810 17876
rect 40034 17864 40040 17876
rect 38856 17836 40040 17864
rect 34333 17799 34391 17805
rect 34333 17796 34345 17799
rect 28040 17768 33088 17796
rect 33244 17768 34345 17796
rect 28040 17756 28046 17768
rect 27893 17731 27951 17737
rect 27893 17697 27905 17731
rect 27939 17697 27951 17731
rect 27893 17691 27951 17697
rect 28166 17688 28172 17740
rect 28224 17728 28230 17740
rect 28626 17728 28632 17740
rect 28224 17700 28632 17728
rect 28224 17688 28230 17700
rect 28626 17688 28632 17700
rect 28684 17728 28690 17740
rect 31202 17728 31208 17740
rect 28684 17700 31208 17728
rect 28684 17688 28690 17700
rect 31202 17688 31208 17700
rect 31260 17688 31266 17740
rect 31754 17688 31760 17740
rect 31812 17688 31818 17740
rect 32398 17688 32404 17740
rect 32456 17688 32462 17740
rect 26421 17663 26479 17669
rect 26421 17660 26433 17663
rect 26384 17632 26433 17660
rect 26384 17620 26390 17632
rect 26421 17629 26433 17632
rect 26467 17629 26479 17663
rect 26421 17623 26479 17629
rect 26513 17663 26571 17669
rect 26513 17629 26525 17663
rect 26559 17629 26571 17663
rect 26513 17623 26571 17629
rect 27157 17663 27215 17669
rect 27157 17629 27169 17663
rect 27203 17629 27215 17663
rect 27157 17623 27215 17629
rect 27249 17663 27307 17669
rect 27249 17629 27261 17663
rect 27295 17660 27307 17663
rect 27522 17660 27528 17672
rect 27295 17632 27528 17660
rect 27295 17629 27307 17632
rect 27249 17623 27307 17629
rect 19334 17592 19340 17604
rect 15212 17564 19340 17592
rect 19334 17552 19340 17564
rect 19392 17592 19398 17604
rect 19429 17595 19487 17601
rect 19429 17592 19441 17595
rect 19392 17564 19441 17592
rect 19392 17552 19398 17564
rect 19429 17561 19441 17564
rect 19475 17561 19487 17595
rect 22204 17592 22232 17620
rect 22925 17595 22983 17601
rect 22925 17592 22937 17595
rect 22204 17564 22937 17592
rect 19429 17555 19487 17561
rect 22925 17561 22937 17564
rect 22971 17592 22983 17595
rect 23014 17592 23020 17604
rect 22971 17564 23020 17592
rect 22971 17561 22983 17564
rect 22925 17555 22983 17561
rect 23014 17552 23020 17564
rect 23072 17552 23078 17604
rect 25240 17592 25268 17620
rect 23124 17564 25268 17592
rect 25777 17595 25835 17601
rect 13170 17524 13176 17536
rect 12216 17496 13176 17524
rect 12216 17484 12222 17496
rect 13170 17484 13176 17496
rect 13228 17484 13234 17536
rect 14458 17484 14464 17536
rect 14516 17524 14522 17536
rect 17126 17524 17132 17536
rect 14516 17496 17132 17524
rect 14516 17484 14522 17496
rect 17126 17484 17132 17496
rect 17184 17524 17190 17536
rect 17770 17524 17776 17536
rect 17184 17496 17776 17524
rect 17184 17484 17190 17496
rect 17770 17484 17776 17496
rect 17828 17484 17834 17536
rect 17862 17484 17868 17536
rect 17920 17524 17926 17536
rect 22094 17524 22100 17536
rect 17920 17496 22100 17524
rect 17920 17484 17926 17496
rect 22094 17484 22100 17496
rect 22152 17484 22158 17536
rect 22186 17484 22192 17536
rect 22244 17524 22250 17536
rect 23124 17524 23152 17564
rect 25777 17561 25789 17595
rect 25823 17561 25835 17595
rect 25777 17555 25835 17561
rect 22244 17496 23152 17524
rect 22244 17484 22250 17496
rect 24578 17484 24584 17536
rect 24636 17524 24642 17536
rect 25792 17524 25820 17555
rect 26786 17552 26792 17604
rect 26844 17592 26850 17604
rect 26973 17595 27031 17601
rect 26973 17592 26985 17595
rect 26844 17564 26985 17592
rect 26844 17552 26850 17564
rect 26973 17561 26985 17564
rect 27019 17561 27031 17595
rect 27172 17592 27200 17623
rect 27522 17620 27528 17632
rect 27580 17620 27586 17672
rect 27982 17620 27988 17672
rect 28040 17620 28046 17672
rect 28074 17620 28080 17672
rect 28132 17660 28138 17672
rect 29362 17660 29368 17672
rect 28132 17632 29368 17660
rect 28132 17620 28138 17632
rect 29362 17620 29368 17632
rect 29420 17620 29426 17672
rect 29730 17620 29736 17672
rect 29788 17620 29794 17672
rect 29825 17663 29883 17669
rect 29825 17629 29837 17663
rect 29871 17660 29883 17663
rect 30282 17660 30288 17672
rect 29871 17632 30288 17660
rect 29871 17629 29883 17632
rect 29825 17623 29883 17629
rect 30282 17620 30288 17632
rect 30340 17620 30346 17672
rect 31110 17620 31116 17672
rect 31168 17620 31174 17672
rect 31386 17620 31392 17672
rect 31444 17620 31450 17672
rect 31938 17620 31944 17672
rect 31996 17620 32002 17672
rect 32493 17663 32551 17669
rect 32493 17629 32505 17663
rect 32539 17660 32551 17663
rect 32582 17660 32588 17672
rect 32539 17632 32588 17660
rect 32539 17629 32551 17632
rect 32493 17623 32551 17629
rect 32582 17620 32588 17632
rect 32640 17620 32646 17672
rect 27709 17595 27767 17601
rect 27172 17564 27292 17592
rect 26973 17555 27031 17561
rect 27264 17536 27292 17564
rect 27709 17561 27721 17595
rect 27755 17561 27767 17595
rect 27709 17555 27767 17561
rect 26418 17524 26424 17536
rect 24636 17496 26424 17524
rect 24636 17484 24642 17496
rect 26418 17484 26424 17496
rect 26476 17484 26482 17536
rect 26694 17484 26700 17536
rect 26752 17484 26758 17536
rect 26881 17527 26939 17533
rect 26881 17493 26893 17527
rect 26927 17524 26939 17527
rect 27246 17524 27252 17536
rect 26927 17496 27252 17524
rect 26927 17493 26939 17496
rect 26881 17487 26939 17493
rect 27246 17484 27252 17496
rect 27304 17484 27310 17536
rect 27433 17527 27491 17533
rect 27433 17493 27445 17527
rect 27479 17524 27491 17527
rect 27724 17524 27752 17555
rect 29546 17552 29552 17604
rect 29604 17601 29610 17604
rect 29604 17592 29613 17601
rect 29604 17564 29649 17592
rect 29604 17555 29613 17564
rect 29604 17552 29610 17555
rect 31662 17552 31668 17604
rect 31720 17552 31726 17604
rect 32217 17595 32275 17601
rect 32217 17592 32229 17595
rect 31956 17564 32229 17592
rect 27479 17496 27752 17524
rect 28169 17527 28227 17533
rect 27479 17493 27491 17496
rect 27433 17487 27491 17493
rect 28169 17493 28181 17527
rect 28215 17524 28227 17527
rect 28442 17524 28448 17536
rect 28215 17496 28448 17524
rect 28215 17493 28227 17496
rect 28169 17487 28227 17493
rect 28442 17484 28448 17496
rect 28500 17484 28506 17536
rect 28810 17484 28816 17536
rect 28868 17524 28874 17536
rect 30009 17527 30067 17533
rect 30009 17524 30021 17527
rect 28868 17496 30021 17524
rect 28868 17484 28874 17496
rect 30009 17493 30021 17496
rect 30055 17524 30067 17527
rect 31018 17524 31024 17536
rect 30055 17496 31024 17524
rect 30055 17493 30067 17496
rect 30009 17487 30067 17493
rect 31018 17484 31024 17496
rect 31076 17484 31082 17536
rect 31573 17527 31631 17533
rect 31573 17493 31585 17527
rect 31619 17524 31631 17527
rect 31956 17524 31984 17564
rect 32217 17561 32229 17564
rect 32263 17561 32275 17595
rect 32217 17555 32275 17561
rect 32953 17595 33011 17601
rect 32953 17561 32965 17595
rect 32999 17561 33011 17595
rect 33060 17592 33088 17768
rect 34333 17765 34345 17768
rect 34379 17765 34391 17799
rect 34333 17759 34391 17765
rect 35253 17799 35311 17805
rect 35253 17765 35265 17799
rect 35299 17796 35311 17799
rect 36280 17796 36308 17824
rect 35299 17768 36308 17796
rect 35299 17765 35311 17768
rect 35253 17759 35311 17765
rect 36538 17756 36544 17808
rect 36596 17796 36602 17808
rect 36596 17768 37780 17796
rect 36596 17756 36602 17768
rect 33134 17688 33140 17740
rect 33192 17688 33198 17740
rect 35158 17728 35164 17740
rect 33428 17700 35164 17728
rect 33226 17620 33232 17672
rect 33284 17620 33290 17672
rect 33428 17592 33456 17700
rect 35158 17688 35164 17700
rect 35216 17688 35222 17740
rect 35437 17731 35495 17737
rect 35437 17728 35449 17731
rect 35268 17700 35449 17728
rect 33778 17670 33784 17672
rect 33505 17663 33563 17669
rect 33505 17629 33517 17663
rect 33551 17660 33563 17663
rect 33612 17660 33784 17670
rect 33551 17642 33784 17660
rect 33551 17632 33640 17642
rect 33551 17629 33563 17632
rect 33505 17623 33563 17629
rect 33778 17620 33784 17642
rect 33836 17620 33842 17672
rect 33962 17620 33968 17672
rect 34020 17620 34026 17672
rect 34057 17663 34115 17669
rect 34057 17629 34069 17663
rect 34103 17629 34115 17663
rect 34057 17623 34115 17629
rect 33060 17564 33456 17592
rect 32953 17555 33011 17561
rect 31619 17496 31984 17524
rect 31619 17493 31631 17496
rect 31573 17487 31631 17493
rect 32122 17484 32128 17536
rect 32180 17484 32186 17536
rect 32677 17527 32735 17533
rect 32677 17493 32689 17527
rect 32723 17524 32735 17527
rect 32968 17524 32996 17555
rect 33594 17552 33600 17604
rect 33652 17592 33658 17604
rect 33689 17595 33747 17601
rect 33689 17592 33701 17595
rect 33652 17564 33701 17592
rect 33652 17552 33658 17564
rect 33689 17561 33701 17564
rect 33735 17561 33747 17595
rect 33689 17555 33747 17561
rect 33870 17552 33876 17604
rect 33928 17592 33934 17604
rect 34072 17592 34100 17623
rect 34422 17620 34428 17672
rect 34480 17660 34486 17672
rect 35268 17660 35296 17700
rect 35437 17697 35449 17700
rect 35483 17697 35495 17731
rect 35437 17691 35495 17697
rect 36357 17731 36415 17737
rect 36357 17697 36369 17731
rect 36403 17728 36415 17731
rect 36722 17728 36728 17740
rect 36403 17700 36728 17728
rect 36403 17697 36415 17700
rect 36357 17691 36415 17697
rect 36722 17688 36728 17700
rect 36780 17688 36786 17740
rect 37752 17728 37780 17768
rect 37826 17756 37832 17808
rect 37884 17796 37890 17808
rect 38381 17799 38439 17805
rect 38381 17796 38393 17799
rect 37884 17768 38393 17796
rect 37884 17756 37890 17768
rect 38381 17765 38393 17768
rect 38427 17765 38439 17799
rect 38381 17759 38439 17765
rect 38470 17756 38476 17808
rect 38528 17796 38534 17808
rect 38856 17796 38884 17836
rect 40034 17824 40040 17836
rect 40092 17824 40098 17876
rect 41509 17867 41567 17873
rect 41509 17833 41521 17867
rect 41555 17864 41567 17867
rect 43254 17864 43260 17876
rect 41555 17836 43260 17864
rect 41555 17833 41567 17836
rect 41509 17827 41567 17833
rect 43254 17824 43260 17836
rect 43312 17824 43318 17876
rect 38528 17768 38884 17796
rect 41233 17799 41291 17805
rect 38528 17756 38534 17768
rect 41233 17765 41245 17799
rect 41279 17796 41291 17799
rect 41690 17796 41696 17808
rect 41279 17768 41696 17796
rect 41279 17765 41291 17768
rect 41233 17759 41291 17765
rect 41690 17756 41696 17768
rect 41748 17756 41754 17808
rect 41969 17799 42027 17805
rect 41969 17765 41981 17799
rect 42015 17796 42027 17799
rect 42702 17796 42708 17808
rect 42015 17768 42708 17796
rect 42015 17765 42027 17768
rect 41969 17759 42027 17765
rect 42702 17756 42708 17768
rect 42760 17756 42766 17808
rect 38930 17728 38936 17740
rect 37752 17700 38936 17728
rect 38930 17688 38936 17700
rect 38988 17688 38994 17740
rect 42153 17731 42211 17737
rect 41432 17700 42104 17728
rect 34480 17632 35296 17660
rect 34480 17620 34486 17632
rect 35342 17620 35348 17672
rect 35400 17620 35406 17672
rect 36446 17620 36452 17672
rect 36504 17620 36510 17672
rect 37093 17663 37151 17669
rect 37093 17660 37105 17663
rect 36556 17632 37105 17660
rect 33928 17564 34100 17592
rect 34885 17595 34943 17601
rect 33928 17552 33934 17564
rect 34885 17561 34897 17595
rect 34931 17561 34943 17595
rect 34885 17555 34943 17561
rect 32723 17496 32996 17524
rect 33413 17527 33471 17533
rect 32723 17493 32735 17496
rect 32677 17487 32735 17493
rect 33413 17493 33425 17527
rect 33459 17524 33471 17527
rect 34146 17524 34152 17536
rect 33459 17496 34152 17524
rect 33459 17493 33471 17496
rect 33413 17487 33471 17493
rect 34146 17484 34152 17496
rect 34204 17484 34210 17536
rect 34900 17524 34928 17555
rect 35066 17552 35072 17604
rect 35124 17552 35130 17604
rect 35158 17552 35164 17604
rect 35216 17592 35222 17604
rect 35216 17564 35480 17592
rect 35216 17552 35222 17564
rect 35342 17524 35348 17536
rect 34900 17496 35348 17524
rect 35342 17484 35348 17496
rect 35400 17484 35406 17536
rect 35452 17524 35480 17564
rect 36078 17552 36084 17604
rect 36136 17592 36142 17604
rect 36173 17595 36231 17601
rect 36173 17592 36185 17595
rect 36136 17564 36185 17592
rect 36136 17552 36142 17564
rect 36173 17561 36185 17564
rect 36219 17561 36231 17595
rect 36173 17555 36231 17561
rect 36556 17524 36584 17632
rect 37093 17629 37105 17632
rect 37139 17660 37151 17663
rect 37461 17663 37519 17669
rect 37461 17660 37473 17663
rect 37139 17632 37473 17660
rect 37139 17629 37151 17632
rect 37093 17623 37151 17629
rect 37461 17629 37473 17632
rect 37507 17629 37519 17663
rect 37461 17623 37519 17629
rect 37550 17620 37556 17672
rect 37608 17620 37614 17672
rect 38194 17620 38200 17672
rect 38252 17620 38258 17672
rect 38838 17620 38844 17672
rect 38896 17620 38902 17672
rect 39850 17620 39856 17672
rect 39908 17620 39914 17672
rect 40126 17669 40132 17672
rect 40120 17660 40132 17669
rect 40087 17632 40132 17660
rect 40120 17623 40132 17632
rect 40126 17620 40132 17623
rect 40184 17620 40190 17672
rect 41322 17620 41328 17672
rect 41380 17660 41386 17672
rect 41432 17669 41460 17700
rect 41417 17663 41475 17669
rect 41417 17660 41429 17663
rect 41380 17632 41429 17660
rect 41380 17620 41386 17632
rect 41417 17629 41429 17632
rect 41463 17629 41475 17663
rect 41417 17623 41475 17629
rect 41693 17663 41751 17669
rect 41693 17629 41705 17663
rect 41739 17629 41751 17663
rect 41693 17623 41751 17629
rect 37277 17595 37335 17601
rect 37277 17592 37289 17595
rect 36648 17564 37289 17592
rect 36648 17533 36676 17564
rect 37277 17561 37289 17564
rect 37323 17561 37335 17595
rect 37277 17555 37335 17561
rect 38657 17595 38715 17601
rect 38657 17561 38669 17595
rect 38703 17592 38715 17595
rect 38746 17592 38752 17604
rect 38703 17564 38752 17592
rect 38703 17561 38715 17564
rect 38657 17555 38715 17561
rect 38746 17552 38752 17564
rect 38804 17552 38810 17604
rect 39022 17552 39028 17604
rect 39080 17552 39086 17604
rect 39574 17552 39580 17604
rect 39632 17592 39638 17604
rect 41708 17592 41736 17623
rect 41782 17620 41788 17672
rect 41840 17620 41846 17672
rect 42076 17669 42104 17700
rect 42153 17697 42165 17731
rect 42199 17728 42211 17731
rect 43073 17731 43131 17737
rect 43073 17728 43085 17731
rect 42199 17700 43085 17728
rect 42199 17697 42211 17700
rect 42153 17691 42211 17697
rect 43073 17697 43085 17700
rect 43119 17697 43131 17731
rect 43073 17691 43131 17697
rect 42061 17663 42119 17669
rect 42061 17629 42073 17663
rect 42107 17629 42119 17663
rect 42277 17663 42335 17669
rect 42277 17660 42289 17663
rect 42061 17623 42119 17629
rect 42260 17629 42289 17660
rect 42323 17629 42335 17663
rect 42260 17623 42335 17629
rect 42429 17663 42487 17669
rect 42429 17629 42441 17663
rect 42475 17660 42487 17663
rect 42518 17660 42524 17672
rect 42475 17632 42524 17660
rect 42475 17629 42487 17632
rect 42429 17623 42487 17629
rect 39632 17564 41736 17592
rect 39632 17552 39638 17564
rect 35452 17496 36584 17524
rect 36633 17527 36691 17533
rect 36633 17493 36645 17527
rect 36679 17493 36691 17527
rect 36633 17487 36691 17493
rect 36998 17484 37004 17536
rect 37056 17524 37062 17536
rect 42260 17524 42288 17623
rect 42518 17620 42524 17632
rect 42576 17620 42582 17672
rect 43717 17663 43775 17669
rect 43717 17629 43729 17663
rect 43763 17660 43775 17663
rect 43806 17660 43812 17672
rect 43763 17632 43812 17660
rect 43763 17629 43775 17632
rect 43717 17623 43775 17629
rect 43806 17620 43812 17632
rect 43864 17620 43870 17672
rect 37056 17496 42288 17524
rect 42613 17527 42671 17533
rect 37056 17484 37062 17496
rect 42613 17493 42625 17527
rect 42659 17524 42671 17527
rect 42702 17524 42708 17536
rect 42659 17496 42708 17524
rect 42659 17493 42671 17496
rect 42613 17487 42671 17493
rect 42702 17484 42708 17496
rect 42760 17484 42766 17536
rect 1104 17434 44896 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 44896 17434
rect 1104 17360 44896 17382
rect 3786 17280 3792 17332
rect 3844 17320 3850 17332
rect 3970 17320 3976 17332
rect 3844 17292 3976 17320
rect 3844 17280 3850 17292
rect 3970 17280 3976 17292
rect 4028 17280 4034 17332
rect 5166 17280 5172 17332
rect 5224 17320 5230 17332
rect 5442 17320 5448 17332
rect 5224 17292 5448 17320
rect 5224 17280 5230 17292
rect 5442 17280 5448 17292
rect 5500 17280 5506 17332
rect 8389 17323 8447 17329
rect 8389 17289 8401 17323
rect 8435 17320 8447 17323
rect 8570 17320 8576 17332
rect 8435 17292 8576 17320
rect 8435 17289 8447 17292
rect 8389 17283 8447 17289
rect 8570 17280 8576 17292
rect 8628 17280 8634 17332
rect 8941 17323 8999 17329
rect 8941 17289 8953 17323
rect 8987 17320 8999 17323
rect 9030 17320 9036 17332
rect 8987 17292 9036 17320
rect 8987 17289 8999 17292
rect 8941 17283 8999 17289
rect 9030 17280 9036 17292
rect 9088 17280 9094 17332
rect 9306 17280 9312 17332
rect 9364 17280 9370 17332
rect 10689 17323 10747 17329
rect 10689 17289 10701 17323
rect 10735 17289 10747 17323
rect 10689 17283 10747 17289
rect 4706 17212 4712 17264
rect 4764 17252 4770 17264
rect 4982 17252 4988 17264
rect 4764 17224 4988 17252
rect 4764 17212 4770 17224
rect 4982 17212 4988 17224
rect 5040 17212 5046 17264
rect 7101 17255 7159 17261
rect 7101 17221 7113 17255
rect 7147 17252 7159 17255
rect 7653 17255 7711 17261
rect 7653 17252 7665 17255
rect 7147 17224 7665 17252
rect 7147 17221 7159 17224
rect 7101 17215 7159 17221
rect 7653 17221 7665 17224
rect 7699 17252 7711 17255
rect 7834 17252 7840 17264
rect 7699 17224 7840 17252
rect 7699 17221 7711 17224
rect 7653 17215 7711 17221
rect 7834 17212 7840 17224
rect 7892 17212 7898 17264
rect 8113 17255 8171 17261
rect 8113 17221 8125 17255
rect 8159 17252 8171 17255
rect 8202 17252 8208 17264
rect 8159 17224 8208 17252
rect 8159 17221 8171 17224
rect 8113 17215 8171 17221
rect 8202 17212 8208 17224
rect 8260 17212 8266 17264
rect 10704 17252 10732 17283
rect 11698 17280 11704 17332
rect 11756 17280 11762 17332
rect 14921 17323 14979 17329
rect 12268 17292 14688 17320
rect 12268 17252 12296 17292
rect 9508 17224 12296 17252
rect 9508 17196 9536 17224
rect 2222 17144 2228 17196
rect 2280 17144 2286 17196
rect 3602 17144 3608 17196
rect 3660 17144 3666 17196
rect 4249 17187 4307 17193
rect 4249 17153 4261 17187
rect 4295 17153 4307 17187
rect 4249 17147 4307 17153
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17184 4491 17187
rect 5442 17184 5448 17196
rect 4479 17156 5448 17184
rect 4479 17153 4491 17156
rect 4433 17147 4491 17153
rect 4264 17116 4292 17147
rect 5442 17144 5448 17156
rect 5500 17144 5506 17196
rect 6089 17187 6147 17193
rect 6089 17153 6101 17187
rect 6135 17184 6147 17187
rect 6822 17184 6828 17196
rect 6135 17156 6828 17184
rect 6135 17153 6147 17156
rect 6089 17147 6147 17153
rect 6822 17144 6828 17156
rect 6880 17144 6886 17196
rect 6917 17187 6975 17193
rect 6917 17153 6929 17187
rect 6963 17184 6975 17187
rect 7285 17187 7343 17193
rect 6963 17156 7052 17184
rect 6963 17153 6975 17156
rect 6917 17147 6975 17153
rect 4706 17116 4712 17128
rect 4264 17088 4712 17116
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 5074 17076 5080 17128
rect 5132 17116 5138 17128
rect 7024 17116 7052 17156
rect 7285 17153 7297 17187
rect 7331 17184 7343 17187
rect 7926 17184 7932 17196
rect 7331 17156 7932 17184
rect 7331 17153 7343 17156
rect 7285 17147 7343 17153
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 8754 17144 8760 17196
rect 8812 17144 8818 17196
rect 9122 17144 9128 17196
rect 9180 17144 9186 17196
rect 9490 17144 9496 17196
rect 9548 17144 9554 17196
rect 9677 17187 9735 17193
rect 9677 17153 9689 17187
rect 9723 17153 9735 17187
rect 9677 17147 9735 17153
rect 7558 17116 7564 17128
rect 5132 17088 7564 17116
rect 5132 17076 5138 17088
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 7742 17076 7748 17128
rect 7800 17116 7806 17128
rect 8205 17119 8263 17125
rect 8205 17116 8217 17119
rect 7800 17088 8217 17116
rect 7800 17076 7806 17088
rect 8205 17085 8217 17088
rect 8251 17085 8263 17119
rect 9692 17116 9720 17147
rect 9766 17144 9772 17196
rect 9824 17144 9830 17196
rect 9858 17144 9864 17196
rect 9916 17193 9922 17196
rect 9916 17184 9924 17193
rect 9916 17156 9961 17184
rect 9916 17147 9924 17156
rect 9916 17144 9922 17147
rect 10134 17144 10140 17196
rect 10192 17184 10198 17196
rect 10502 17184 10508 17196
rect 10192 17156 10508 17184
rect 10192 17144 10198 17156
rect 10502 17144 10508 17156
rect 10560 17144 10566 17196
rect 10686 17144 10692 17196
rect 10744 17184 10750 17196
rect 10781 17187 10839 17193
rect 10781 17184 10793 17187
rect 10744 17156 10793 17184
rect 10744 17144 10750 17156
rect 10781 17153 10793 17156
rect 10827 17153 10839 17187
rect 10781 17147 10839 17153
rect 11422 17144 11428 17196
rect 11480 17184 11486 17196
rect 11977 17187 12035 17193
rect 11977 17184 11989 17187
rect 11480 17156 11989 17184
rect 11480 17144 11486 17156
rect 11977 17153 11989 17156
rect 12023 17153 12035 17187
rect 11977 17147 12035 17153
rect 12161 17187 12219 17193
rect 12161 17153 12173 17187
rect 12207 17184 12219 17187
rect 12268 17184 12296 17224
rect 12529 17255 12587 17261
rect 12529 17221 12541 17255
rect 12575 17252 12587 17255
rect 12618 17252 12624 17264
rect 12575 17224 12624 17252
rect 12575 17221 12587 17224
rect 12529 17215 12587 17221
rect 12618 17212 12624 17224
rect 12676 17252 12682 17264
rect 14001 17255 14059 17261
rect 12676 17224 13400 17252
rect 12676 17212 12682 17224
rect 12207 17156 12296 17184
rect 12345 17187 12403 17193
rect 12207 17153 12219 17156
rect 12161 17147 12219 17153
rect 12345 17153 12357 17187
rect 12391 17153 12403 17187
rect 12345 17147 12403 17153
rect 10226 17116 10232 17128
rect 9692 17088 10232 17116
rect 8205 17079 8263 17085
rect 10226 17076 10232 17088
rect 10284 17076 10290 17128
rect 11054 17076 11060 17128
rect 11112 17116 11118 17128
rect 11609 17119 11667 17125
rect 11609 17116 11621 17119
rect 11112 17088 11621 17116
rect 11112 17076 11118 17088
rect 11609 17085 11621 17088
rect 11655 17085 11667 17119
rect 11609 17079 11667 17085
rect 11882 17076 11888 17128
rect 11940 17116 11946 17128
rect 12176 17116 12204 17147
rect 11940 17088 12204 17116
rect 11940 17076 11946 17088
rect 3694 17008 3700 17060
rect 3752 17048 3758 17060
rect 3752 17020 5396 17048
rect 3752 17008 3758 17020
rect 5368 16992 5396 17020
rect 5534 17008 5540 17060
rect 5592 17048 5598 17060
rect 5905 17051 5963 17057
rect 5905 17048 5917 17051
rect 5592 17020 5917 17048
rect 5592 17008 5598 17020
rect 5905 17017 5917 17020
rect 5951 17048 5963 17051
rect 6270 17048 6276 17060
rect 5951 17020 6276 17048
rect 5951 17017 5963 17020
rect 5905 17011 5963 17017
rect 6270 17008 6276 17020
rect 6328 17008 6334 17060
rect 7469 17051 7527 17057
rect 7469 17017 7481 17051
rect 7515 17048 7527 17051
rect 7653 17051 7711 17057
rect 7653 17048 7665 17051
rect 7515 17020 7665 17048
rect 7515 17017 7527 17020
rect 7469 17011 7527 17017
rect 7653 17017 7665 17020
rect 7699 17048 7711 17051
rect 8294 17048 8300 17060
rect 7699 17020 8300 17048
rect 7699 17017 7711 17020
rect 7653 17011 7711 17017
rect 8294 17008 8300 17020
rect 8352 17008 8358 17060
rect 10045 17051 10103 17057
rect 10045 17017 10057 17051
rect 10091 17048 10103 17051
rect 10962 17048 10968 17060
rect 10091 17020 10968 17048
rect 10091 17017 10103 17020
rect 10045 17011 10103 17017
rect 10962 17008 10968 17020
rect 11020 17008 11026 17060
rect 2314 16940 2320 16992
rect 2372 16940 2378 16992
rect 3878 16940 3884 16992
rect 3936 16980 3942 16992
rect 4065 16983 4123 16989
rect 4065 16980 4077 16983
rect 3936 16952 4077 16980
rect 3936 16940 3942 16952
rect 4065 16949 4077 16952
rect 4111 16949 4123 16983
rect 4065 16943 4123 16949
rect 4709 16983 4767 16989
rect 4709 16949 4721 16983
rect 4755 16980 4767 16983
rect 4890 16980 4896 16992
rect 4755 16952 4896 16980
rect 4755 16949 4767 16952
rect 4709 16943 4767 16949
rect 4890 16940 4896 16952
rect 4948 16940 4954 16992
rect 5350 16940 5356 16992
rect 5408 16980 5414 16992
rect 12360 16980 12388 17147
rect 12986 17144 12992 17196
rect 13044 17144 13050 17196
rect 13170 17144 13176 17196
rect 13228 17144 13234 17196
rect 13262 17144 13268 17196
rect 13320 17144 13326 17196
rect 13372 17193 13400 17224
rect 14001 17221 14013 17255
rect 14047 17252 14059 17255
rect 14458 17252 14464 17264
rect 14047 17224 14464 17252
rect 14047 17221 14059 17224
rect 14001 17215 14059 17221
rect 14458 17212 14464 17224
rect 14516 17212 14522 17264
rect 13362 17187 13420 17193
rect 13362 17153 13374 17187
rect 13408 17184 13420 17187
rect 13408 17156 13492 17184
rect 13408 17153 13420 17156
rect 13362 17147 13420 17153
rect 13464 17116 13492 17156
rect 13722 17144 13728 17196
rect 13780 17144 13786 17196
rect 13906 17144 13912 17196
rect 13964 17144 13970 17196
rect 14090 17144 14096 17196
rect 14148 17193 14154 17196
rect 14660 17193 14688 17292
rect 14921 17289 14933 17323
rect 14967 17289 14979 17323
rect 14921 17283 14979 17289
rect 19078 17323 19136 17329
rect 19078 17289 19090 17323
rect 19124 17320 19136 17323
rect 19610 17320 19616 17332
rect 19124 17292 19616 17320
rect 19124 17289 19136 17292
rect 19078 17283 19136 17289
rect 14148 17184 14156 17193
rect 14645 17187 14703 17193
rect 14148 17156 14193 17184
rect 14148 17147 14156 17156
rect 14645 17153 14657 17187
rect 14691 17153 14703 17187
rect 14645 17147 14703 17153
rect 14148 17144 14154 17147
rect 14461 17119 14519 17125
rect 14461 17116 14473 17119
rect 13464 17088 14473 17116
rect 14461 17085 14473 17088
rect 14507 17085 14519 17119
rect 14461 17079 14519 17085
rect 13538 17008 13544 17060
rect 13596 17008 13602 17060
rect 14182 17008 14188 17060
rect 14240 17048 14246 17060
rect 14277 17051 14335 17057
rect 14277 17048 14289 17051
rect 14240 17020 14289 17048
rect 14240 17008 14246 17020
rect 14277 17017 14289 17020
rect 14323 17017 14335 17051
rect 14936 17048 14964 17283
rect 19610 17280 19616 17292
rect 19668 17280 19674 17332
rect 22094 17280 22100 17332
rect 22152 17320 22158 17332
rect 23106 17320 23112 17332
rect 22152 17292 23112 17320
rect 22152 17280 22158 17292
rect 23106 17280 23112 17292
rect 23164 17280 23170 17332
rect 23385 17323 23443 17329
rect 23385 17289 23397 17323
rect 23431 17289 23443 17323
rect 23385 17283 23443 17289
rect 16850 17212 16856 17264
rect 16908 17252 16914 17264
rect 23198 17252 23204 17264
rect 16908 17224 23204 17252
rect 16908 17212 16914 17224
rect 23198 17212 23204 17224
rect 23256 17212 23262 17264
rect 23400 17252 23428 17283
rect 24394 17280 24400 17332
rect 24452 17320 24458 17332
rect 24762 17320 24768 17332
rect 24452 17292 24768 17320
rect 24452 17280 24458 17292
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 26786 17280 26792 17332
rect 26844 17320 26850 17332
rect 27154 17320 27160 17332
rect 26844 17292 27160 17320
rect 26844 17280 26850 17292
rect 27154 17280 27160 17292
rect 27212 17280 27218 17332
rect 27341 17323 27399 17329
rect 27341 17289 27353 17323
rect 27387 17320 27399 17323
rect 31662 17320 31668 17332
rect 27387 17292 31668 17320
rect 27387 17289 27399 17292
rect 27341 17283 27399 17289
rect 31662 17280 31668 17292
rect 31720 17320 31726 17332
rect 31938 17320 31944 17332
rect 31720 17292 31944 17320
rect 31720 17280 31726 17292
rect 31938 17280 31944 17292
rect 31996 17280 32002 17332
rect 34054 17280 34060 17332
rect 34112 17320 34118 17332
rect 34112 17292 35664 17320
rect 34112 17280 34118 17292
rect 26234 17252 26240 17264
rect 23400 17224 26240 17252
rect 26234 17212 26240 17224
rect 26292 17252 26298 17264
rect 26292 17224 26464 17252
rect 26292 17212 26298 17224
rect 15010 17144 15016 17196
rect 15068 17144 15074 17196
rect 17770 17144 17776 17196
rect 17828 17184 17834 17196
rect 18509 17187 18567 17193
rect 18509 17184 18521 17187
rect 17828 17156 18521 17184
rect 17828 17144 17834 17156
rect 18509 17153 18521 17156
rect 18555 17153 18567 17187
rect 18509 17147 18567 17153
rect 18690 17144 18696 17196
rect 18748 17144 18754 17196
rect 18782 17144 18788 17196
rect 18840 17144 18846 17196
rect 18882 17187 18940 17193
rect 18882 17153 18894 17187
rect 18928 17153 18940 17187
rect 18882 17147 18940 17153
rect 15838 17076 15844 17128
rect 15896 17116 15902 17128
rect 17954 17116 17960 17128
rect 15896 17088 17960 17116
rect 15896 17076 15902 17088
rect 17954 17076 17960 17088
rect 18012 17116 18018 17128
rect 18897 17116 18925 17147
rect 19150 17144 19156 17196
rect 19208 17184 19214 17196
rect 19245 17187 19303 17193
rect 19245 17184 19257 17187
rect 19208 17156 19257 17184
rect 19208 17144 19214 17156
rect 19245 17153 19257 17156
rect 19291 17153 19303 17187
rect 19245 17147 19303 17153
rect 19429 17187 19487 17193
rect 19429 17153 19441 17187
rect 19475 17184 19487 17187
rect 20254 17184 20260 17196
rect 19475 17156 20260 17184
rect 19475 17153 19487 17156
rect 19429 17147 19487 17153
rect 20254 17144 20260 17156
rect 20312 17144 20318 17196
rect 22738 17144 22744 17196
rect 22796 17184 22802 17196
rect 23017 17187 23075 17193
rect 23017 17184 23029 17187
rect 22796 17156 23029 17184
rect 22796 17144 22802 17156
rect 23017 17153 23029 17156
rect 23063 17153 23075 17187
rect 23017 17147 23075 17153
rect 24762 17144 24768 17196
rect 24820 17144 24826 17196
rect 25041 17187 25099 17193
rect 25041 17153 25053 17187
rect 25087 17184 25099 17187
rect 26326 17184 26332 17196
rect 25087 17156 26332 17184
rect 25087 17153 25099 17156
rect 25041 17147 25099 17153
rect 26326 17144 26332 17156
rect 26384 17144 26390 17196
rect 18012 17088 18925 17116
rect 18012 17076 18018 17088
rect 19058 17076 19064 17128
rect 19116 17116 19122 17128
rect 24302 17116 24308 17128
rect 19116 17088 24308 17116
rect 19116 17076 19122 17088
rect 24302 17076 24308 17088
rect 24360 17076 24366 17128
rect 24854 17076 24860 17128
rect 24912 17076 24918 17128
rect 25314 17116 25320 17128
rect 24964 17088 25320 17116
rect 24026 17048 24032 17060
rect 14936 17020 24032 17048
rect 14277 17011 14335 17017
rect 24026 17008 24032 17020
rect 24084 17008 24090 17060
rect 5408 16952 12388 16980
rect 5408 16940 5414 16952
rect 12894 16940 12900 16992
rect 12952 16980 12958 16992
rect 14090 16980 14096 16992
rect 12952 16952 14096 16980
rect 12952 16940 12958 16952
rect 14090 16940 14096 16952
rect 14148 16940 14154 16992
rect 14366 16940 14372 16992
rect 14424 16980 14430 16992
rect 18782 16980 18788 16992
rect 14424 16952 18788 16980
rect 14424 16940 14430 16952
rect 18782 16940 18788 16952
rect 18840 16980 18846 16992
rect 19150 16980 19156 16992
rect 18840 16952 19156 16980
rect 18840 16940 18846 16952
rect 19150 16940 19156 16952
rect 19208 16940 19214 16992
rect 19334 16940 19340 16992
rect 19392 16940 19398 16992
rect 19426 16940 19432 16992
rect 19484 16980 19490 16992
rect 19613 16983 19671 16989
rect 19613 16980 19625 16983
rect 19484 16952 19625 16980
rect 19484 16940 19490 16952
rect 19613 16949 19625 16952
rect 19659 16949 19671 16983
rect 19613 16943 19671 16949
rect 19794 16940 19800 16992
rect 19852 16980 19858 16992
rect 24578 16980 24584 16992
rect 19852 16952 24584 16980
rect 19852 16940 19858 16952
rect 24578 16940 24584 16952
rect 24636 16940 24642 16992
rect 24964 16989 24992 17088
rect 25314 17076 25320 17088
rect 25372 17076 25378 17128
rect 26436 17116 26464 17224
rect 26694 17212 26700 17264
rect 26752 17252 26758 17264
rect 26752 17224 27292 17252
rect 26752 17212 26758 17224
rect 26510 17144 26516 17196
rect 26568 17184 26574 17196
rect 26973 17187 27031 17193
rect 26973 17184 26985 17187
rect 26568 17156 26985 17184
rect 26568 17144 26574 17156
rect 26973 17153 26985 17156
rect 27019 17153 27031 17187
rect 27264 17184 27292 17224
rect 27706 17212 27712 17264
rect 27764 17212 27770 17264
rect 28966 17224 30696 17252
rect 27893 17187 27951 17193
rect 27893 17184 27905 17187
rect 27264 17156 27905 17184
rect 26973 17147 27031 17153
rect 27893 17153 27905 17156
rect 27939 17153 27951 17187
rect 27893 17147 27951 17153
rect 27985 17187 28043 17193
rect 27985 17153 27997 17187
rect 28031 17184 28043 17187
rect 28074 17184 28080 17196
rect 28031 17156 28080 17184
rect 28031 17153 28043 17156
rect 27985 17147 28043 17153
rect 28074 17144 28080 17156
rect 28132 17144 28138 17196
rect 27065 17119 27123 17125
rect 27065 17116 27077 17119
rect 26436 17088 27077 17116
rect 27065 17085 27077 17088
rect 27111 17085 27123 17119
rect 27065 17079 27123 17085
rect 27154 17076 27160 17128
rect 27212 17116 27218 17128
rect 28966 17116 28994 17224
rect 29457 17187 29515 17193
rect 29457 17153 29469 17187
rect 29503 17184 29515 17187
rect 29638 17184 29644 17196
rect 29503 17156 29644 17184
rect 29503 17153 29515 17156
rect 29457 17147 29515 17153
rect 29638 17144 29644 17156
rect 29696 17144 29702 17196
rect 30668 17184 30696 17224
rect 32122 17212 32128 17264
rect 32180 17212 32186 17264
rect 32306 17212 32312 17264
rect 32364 17212 32370 17264
rect 35636 17261 35664 17292
rect 36078 17280 36084 17332
rect 36136 17280 36142 17332
rect 36817 17323 36875 17329
rect 36817 17289 36829 17323
rect 36863 17320 36875 17323
rect 37274 17320 37280 17332
rect 36863 17292 37280 17320
rect 36863 17289 36875 17292
rect 36817 17283 36875 17289
rect 37274 17280 37280 17292
rect 37332 17280 37338 17332
rect 38289 17323 38347 17329
rect 38289 17289 38301 17323
rect 38335 17320 38347 17323
rect 38470 17320 38476 17332
rect 38335 17292 38476 17320
rect 38335 17289 38347 17292
rect 38289 17283 38347 17289
rect 35621 17255 35679 17261
rect 35621 17221 35633 17255
rect 35667 17221 35679 17255
rect 35621 17215 35679 17221
rect 35710 17212 35716 17264
rect 35768 17252 35774 17264
rect 36354 17252 36360 17264
rect 35768 17224 36360 17252
rect 35768 17212 35774 17224
rect 36354 17212 36360 17224
rect 36412 17212 36418 17264
rect 36906 17212 36912 17264
rect 36964 17252 36970 17264
rect 38304 17252 38332 17283
rect 38470 17280 38476 17292
rect 38528 17280 38534 17332
rect 40218 17320 40224 17332
rect 38764 17292 40224 17320
rect 36964 17224 38332 17252
rect 36964 17212 36970 17224
rect 31386 17184 31392 17196
rect 30668 17156 31392 17184
rect 31386 17144 31392 17156
rect 31444 17184 31450 17196
rect 31561 17193 31619 17199
rect 31561 17184 31573 17193
rect 31444 17159 31573 17184
rect 31607 17159 31619 17193
rect 31444 17156 31619 17159
rect 31444 17144 31450 17156
rect 31561 17153 31619 17156
rect 31757 17187 31815 17193
rect 31757 17153 31769 17187
rect 31803 17153 31815 17187
rect 35526 17184 35532 17196
rect 31757 17147 31815 17153
rect 31956 17156 35532 17184
rect 27212 17088 28994 17116
rect 27212 17076 27218 17088
rect 29546 17076 29552 17128
rect 29604 17116 29610 17128
rect 30282 17116 30288 17128
rect 29604 17088 30288 17116
rect 29604 17076 29610 17088
rect 30282 17076 30288 17088
rect 30340 17076 30346 17128
rect 31772 17116 31800 17147
rect 31726 17088 31800 17116
rect 29825 17051 29883 17057
rect 29825 17048 29837 17051
rect 28092 17020 29837 17048
rect 24949 16983 25007 16989
rect 24949 16949 24961 16983
rect 24995 16949 25007 16983
rect 24949 16943 25007 16949
rect 25038 16940 25044 16992
rect 25096 16980 25102 16992
rect 25225 16983 25283 16989
rect 25225 16980 25237 16983
rect 25096 16952 25237 16980
rect 25096 16940 25102 16952
rect 25225 16949 25237 16952
rect 25271 16949 25283 16983
rect 25225 16943 25283 16949
rect 26878 16940 26884 16992
rect 26936 16980 26942 16992
rect 27154 16980 27160 16992
rect 26936 16952 27160 16980
rect 26936 16940 26942 16952
rect 27154 16940 27160 16952
rect 27212 16940 27218 16992
rect 27801 16983 27859 16989
rect 27801 16949 27813 16983
rect 27847 16980 27859 16983
rect 27982 16980 27988 16992
rect 27847 16952 27988 16980
rect 27847 16949 27859 16952
rect 27801 16943 27859 16949
rect 27982 16940 27988 16952
rect 28040 16980 28046 16992
rect 28092 16980 28120 17020
rect 29825 17017 29837 17020
rect 29871 17048 29883 17051
rect 30190 17048 30196 17060
rect 29871 17020 30196 17048
rect 29871 17017 29883 17020
rect 29825 17011 29883 17017
rect 30190 17008 30196 17020
rect 30248 17008 30254 17060
rect 31478 17008 31484 17060
rect 31536 17048 31542 17060
rect 31726 17048 31754 17088
rect 31956 17057 31984 17156
rect 35526 17144 35532 17156
rect 35584 17144 35590 17196
rect 35894 17144 35900 17196
rect 35952 17144 35958 17196
rect 36630 17144 36636 17196
rect 36688 17144 36694 17196
rect 37642 17144 37648 17196
rect 37700 17144 37706 17196
rect 37844 17193 37872 17224
rect 37829 17187 37887 17193
rect 37829 17153 37841 17187
rect 37875 17153 37887 17187
rect 37829 17147 37887 17153
rect 38378 17144 38384 17196
rect 38436 17144 38442 17196
rect 38565 17187 38623 17193
rect 38565 17153 38577 17187
rect 38611 17184 38623 17187
rect 38654 17184 38660 17196
rect 38611 17156 38660 17184
rect 38611 17153 38623 17156
rect 38565 17147 38623 17153
rect 38654 17144 38660 17156
rect 38712 17144 38718 17196
rect 38764 17193 38792 17292
rect 40218 17280 40224 17292
rect 40276 17280 40282 17332
rect 40310 17280 40316 17332
rect 40368 17320 40374 17332
rect 40681 17323 40739 17329
rect 40681 17320 40693 17323
rect 40368 17292 40693 17320
rect 40368 17280 40374 17292
rect 40681 17289 40693 17292
rect 40727 17289 40739 17323
rect 40681 17283 40739 17289
rect 41230 17280 41236 17332
rect 41288 17320 41294 17332
rect 41782 17320 41788 17332
rect 41288 17292 41788 17320
rect 41288 17280 41294 17292
rect 41782 17280 41788 17292
rect 41840 17280 41846 17332
rect 43806 17280 43812 17332
rect 43864 17280 43870 17332
rect 38838 17212 38844 17264
rect 38896 17252 38902 17264
rect 39850 17252 39856 17264
rect 38896 17224 39856 17252
rect 38896 17212 38902 17224
rect 38749 17187 38807 17193
rect 38749 17153 38761 17187
rect 38795 17153 38807 17187
rect 38749 17147 38807 17153
rect 38930 17144 38936 17196
rect 38988 17184 38994 17196
rect 39316 17193 39344 17224
rect 39850 17212 39856 17224
rect 39908 17212 39914 17264
rect 39025 17187 39083 17193
rect 39025 17184 39037 17187
rect 38988 17156 39037 17184
rect 38988 17144 38994 17156
rect 39025 17153 39037 17156
rect 39071 17153 39083 17187
rect 39025 17147 39083 17153
rect 39301 17187 39359 17193
rect 39301 17153 39313 17187
rect 39347 17153 39359 17187
rect 39557 17187 39615 17193
rect 39557 17184 39569 17187
rect 39301 17147 39359 17153
rect 39408 17156 39569 17184
rect 35434 17076 35440 17128
rect 35492 17116 35498 17128
rect 35710 17116 35716 17128
rect 35492 17088 35716 17116
rect 35492 17076 35498 17088
rect 35710 17076 35716 17088
rect 35768 17076 35774 17128
rect 36446 17076 36452 17128
rect 36504 17076 36510 17128
rect 36538 17076 36544 17128
rect 36596 17116 36602 17128
rect 38841 17119 38899 17125
rect 38841 17116 38853 17119
rect 36596 17088 38853 17116
rect 36596 17076 36602 17088
rect 38841 17085 38853 17088
rect 38887 17085 38899 17119
rect 38841 17079 38899 17085
rect 39209 17119 39267 17125
rect 39209 17085 39221 17119
rect 39255 17116 39267 17119
rect 39408 17116 39436 17156
rect 39557 17153 39569 17156
rect 39603 17153 39615 17187
rect 39557 17147 39615 17153
rect 42426 17144 42432 17196
rect 42484 17144 42490 17196
rect 42702 17193 42708 17196
rect 42696 17184 42708 17193
rect 42663 17156 42708 17184
rect 42696 17147 42708 17156
rect 42702 17144 42708 17147
rect 42760 17144 42766 17196
rect 43824 17184 43852 17280
rect 44269 17187 44327 17193
rect 44269 17184 44281 17187
rect 43824 17156 44281 17184
rect 44269 17153 44281 17156
rect 44315 17153 44327 17187
rect 44269 17147 44327 17153
rect 39255 17088 39436 17116
rect 39255 17085 39267 17088
rect 39209 17079 39267 17085
rect 31536 17020 31754 17048
rect 31941 17051 31999 17057
rect 31536 17008 31542 17020
rect 31941 17017 31953 17051
rect 31987 17017 31999 17051
rect 31941 17011 31999 17017
rect 32493 17051 32551 17057
rect 32493 17017 32505 17051
rect 32539 17048 32551 17051
rect 36722 17048 36728 17060
rect 32539 17020 36728 17048
rect 32539 17017 32551 17020
rect 32493 17011 32551 17017
rect 36722 17008 36728 17020
rect 36780 17008 36786 17060
rect 37734 17008 37740 17060
rect 37792 17048 37798 17060
rect 38013 17051 38071 17057
rect 38013 17048 38025 17051
rect 37792 17020 38025 17048
rect 37792 17008 37798 17020
rect 38013 17017 38025 17020
rect 38059 17048 38071 17051
rect 38933 17051 38991 17057
rect 38059 17020 38608 17048
rect 38059 17017 38071 17020
rect 38013 17011 38071 17017
rect 28040 16952 28120 16980
rect 28169 16983 28227 16989
rect 28040 16940 28046 16952
rect 28169 16949 28181 16983
rect 28215 16980 28227 16983
rect 29362 16980 29368 16992
rect 28215 16952 29368 16980
rect 28215 16949 28227 16952
rect 28169 16943 28227 16949
rect 29362 16940 29368 16952
rect 29420 16940 29426 16992
rect 29454 16940 29460 16992
rect 29512 16980 29518 16992
rect 29730 16980 29736 16992
rect 29512 16952 29736 16980
rect 29512 16940 29518 16952
rect 29730 16940 29736 16952
rect 29788 16940 29794 16992
rect 31662 16940 31668 16992
rect 31720 16940 31726 16992
rect 33134 16940 33140 16992
rect 33192 16980 33198 16992
rect 35621 16983 35679 16989
rect 35621 16980 35633 16983
rect 33192 16952 35633 16980
rect 33192 16940 33198 16952
rect 35621 16949 35633 16952
rect 35667 16949 35679 16983
rect 35621 16943 35679 16949
rect 35710 16940 35716 16992
rect 35768 16980 35774 16992
rect 36357 16983 36415 16989
rect 36357 16980 36369 16983
rect 35768 16952 36369 16980
rect 35768 16940 35774 16952
rect 36357 16949 36369 16952
rect 36403 16949 36415 16983
rect 36357 16943 36415 16949
rect 37182 16940 37188 16992
rect 37240 16980 37246 16992
rect 37369 16983 37427 16989
rect 37369 16980 37381 16983
rect 37240 16952 37381 16980
rect 37240 16940 37246 16952
rect 37369 16949 37381 16952
rect 37415 16949 37427 16983
rect 37369 16943 37427 16949
rect 37642 16940 37648 16992
rect 37700 16980 37706 16992
rect 38286 16980 38292 16992
rect 37700 16952 38292 16980
rect 37700 16940 37706 16952
rect 38286 16940 38292 16952
rect 38344 16980 38350 16992
rect 38470 16980 38476 16992
rect 38344 16952 38476 16980
rect 38344 16940 38350 16952
rect 38470 16940 38476 16952
rect 38528 16940 38534 16992
rect 38580 16980 38608 17020
rect 38933 17017 38945 17051
rect 38979 17017 38991 17051
rect 38933 17011 38991 17017
rect 38948 16980 38976 17011
rect 44450 17008 44456 17060
rect 44508 17008 44514 17060
rect 41230 16980 41236 16992
rect 38580 16952 41236 16980
rect 41230 16940 41236 16952
rect 41288 16940 41294 16992
rect 1104 16890 44896 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 44896 16890
rect 1104 16816 44896 16838
rect 2501 16779 2559 16785
rect 2501 16745 2513 16779
rect 2547 16776 2559 16779
rect 3234 16776 3240 16788
rect 2547 16748 3240 16776
rect 2547 16745 2559 16748
rect 2501 16739 2559 16745
rect 3234 16736 3240 16748
rect 3292 16736 3298 16788
rect 3605 16779 3663 16785
rect 3605 16745 3617 16779
rect 3651 16776 3663 16779
rect 3694 16776 3700 16788
rect 3651 16748 3700 16776
rect 3651 16745 3663 16748
rect 3605 16739 3663 16745
rect 3694 16736 3700 16748
rect 3752 16736 3758 16788
rect 4341 16779 4399 16785
rect 4341 16745 4353 16779
rect 4387 16776 4399 16779
rect 4614 16776 4620 16788
rect 4387 16748 4620 16776
rect 4387 16745 4399 16748
rect 4341 16739 4399 16745
rect 4614 16736 4620 16748
rect 4672 16736 4678 16788
rect 7024 16748 8708 16776
rect 1765 16711 1823 16717
rect 1765 16677 1777 16711
rect 1811 16708 1823 16711
rect 2130 16708 2136 16720
rect 1811 16680 2136 16708
rect 1811 16677 1823 16680
rect 1765 16671 1823 16677
rect 2130 16668 2136 16680
rect 2188 16668 2194 16720
rect 2869 16711 2927 16717
rect 2869 16677 2881 16711
rect 2915 16708 2927 16711
rect 3053 16711 3111 16717
rect 3053 16708 3065 16711
rect 2915 16680 3065 16708
rect 2915 16677 2927 16680
rect 2869 16671 2927 16677
rect 3053 16677 3065 16680
rect 3099 16708 3111 16711
rect 3970 16708 3976 16720
rect 3099 16680 3976 16708
rect 3099 16677 3111 16680
rect 3053 16671 3111 16677
rect 3970 16668 3976 16680
rect 4028 16668 4034 16720
rect 4154 16708 4160 16720
rect 4080 16680 4160 16708
rect 2314 16600 2320 16652
rect 2372 16640 2378 16652
rect 4080 16649 4108 16680
rect 4154 16668 4160 16680
rect 4212 16708 4218 16720
rect 5074 16708 5080 16720
rect 4212 16680 5080 16708
rect 4212 16668 4218 16680
rect 5074 16668 5080 16680
rect 5132 16668 5138 16720
rect 5258 16668 5264 16720
rect 5316 16668 5322 16720
rect 5442 16668 5448 16720
rect 5500 16708 5506 16720
rect 5500 16680 5948 16708
rect 5500 16668 5506 16680
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 2372 16612 4077 16640
rect 2372 16600 2378 16612
rect 842 16532 848 16584
rect 900 16572 906 16584
rect 3252 16581 3280 16612
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 4709 16643 4767 16649
rect 4709 16609 4721 16643
rect 4755 16640 4767 16643
rect 5276 16640 5304 16668
rect 5920 16640 5948 16680
rect 5994 16668 6000 16720
rect 6052 16708 6058 16720
rect 6178 16708 6184 16720
rect 6052 16680 6184 16708
rect 6052 16668 6058 16680
rect 6178 16668 6184 16680
rect 6236 16668 6242 16720
rect 7024 16640 7052 16748
rect 7466 16668 7472 16720
rect 7524 16668 7530 16720
rect 8021 16711 8079 16717
rect 8021 16677 8033 16711
rect 8067 16708 8079 16711
rect 8294 16708 8300 16720
rect 8067 16680 8300 16708
rect 8067 16677 8079 16680
rect 8021 16671 8079 16677
rect 8294 16668 8300 16680
rect 8352 16668 8358 16720
rect 8570 16668 8576 16720
rect 8628 16668 8634 16720
rect 8680 16708 8708 16748
rect 8754 16736 8760 16788
rect 8812 16736 8818 16788
rect 10134 16776 10140 16788
rect 8864 16748 10140 16776
rect 8864 16708 8892 16748
rect 10134 16736 10140 16748
rect 10192 16736 10198 16788
rect 19794 16776 19800 16788
rect 17420 16748 19800 16776
rect 17420 16720 17448 16748
rect 19794 16736 19800 16748
rect 19852 16736 19858 16788
rect 21082 16736 21088 16788
rect 21140 16736 21146 16788
rect 21821 16779 21879 16785
rect 21821 16745 21833 16779
rect 21867 16776 21879 16779
rect 22278 16776 22284 16788
rect 21867 16748 22284 16776
rect 21867 16745 21879 16748
rect 21821 16739 21879 16745
rect 22278 16736 22284 16748
rect 22336 16736 22342 16788
rect 22465 16779 22523 16785
rect 22465 16745 22477 16779
rect 22511 16776 22523 16779
rect 22554 16776 22560 16788
rect 22511 16748 22560 16776
rect 22511 16745 22523 16748
rect 22465 16739 22523 16745
rect 22554 16736 22560 16748
rect 22612 16736 22618 16788
rect 22833 16779 22891 16785
rect 22833 16745 22845 16779
rect 22879 16776 22891 16779
rect 23106 16776 23112 16788
rect 22879 16748 23112 16776
rect 22879 16745 22891 16748
rect 22833 16739 22891 16745
rect 23106 16736 23112 16748
rect 23164 16736 23170 16788
rect 24302 16736 24308 16788
rect 24360 16776 24366 16788
rect 24673 16779 24731 16785
rect 24673 16776 24685 16779
rect 24360 16748 24685 16776
rect 24360 16736 24366 16748
rect 24673 16745 24685 16748
rect 24719 16745 24731 16779
rect 24673 16739 24731 16745
rect 24857 16779 24915 16785
rect 24857 16745 24869 16779
rect 24903 16745 24915 16779
rect 24857 16739 24915 16745
rect 9858 16708 9864 16720
rect 8680 16680 8892 16708
rect 9232 16680 9864 16708
rect 4755 16612 5856 16640
rect 5920 16612 7052 16640
rect 7101 16643 7159 16649
rect 4755 16609 4767 16612
rect 4709 16603 4767 16609
rect 1397 16575 1455 16581
rect 1397 16572 1409 16575
rect 900 16544 1409 16572
rect 900 16532 906 16544
rect 1397 16541 1409 16544
rect 1443 16541 1455 16575
rect 2685 16575 2743 16581
rect 2685 16572 2697 16575
rect 1397 16535 1455 16541
rect 1596 16544 2697 16572
rect 1596 16445 1624 16544
rect 2685 16541 2697 16544
rect 2731 16541 2743 16575
rect 2685 16535 2743 16541
rect 3237 16575 3295 16581
rect 3237 16541 3249 16575
rect 3283 16541 3295 16575
rect 3237 16535 3295 16541
rect 3510 16532 3516 16584
rect 3568 16572 3574 16584
rect 3881 16575 3939 16581
rect 3881 16572 3893 16575
rect 3568 16544 3893 16572
rect 3568 16532 3574 16544
rect 3881 16541 3893 16544
rect 3927 16541 3939 16575
rect 3881 16535 3939 16541
rect 3970 16532 3976 16584
rect 4028 16532 4034 16584
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16541 4215 16575
rect 4157 16535 4215 16541
rect 4893 16575 4951 16581
rect 4893 16541 4905 16575
rect 4939 16541 4951 16575
rect 4893 16535 4951 16541
rect 1762 16464 1768 16516
rect 1820 16464 1826 16516
rect 2225 16507 2283 16513
rect 2225 16473 2237 16507
rect 2271 16504 2283 16507
rect 2958 16504 2964 16516
rect 2271 16476 2964 16504
rect 2271 16473 2283 16476
rect 2225 16467 2283 16473
rect 2958 16464 2964 16476
rect 3016 16464 3022 16516
rect 3050 16464 3056 16516
rect 3108 16504 3114 16516
rect 3421 16507 3479 16513
rect 3421 16504 3433 16507
rect 3108 16476 3433 16504
rect 3108 16464 3114 16476
rect 3421 16473 3433 16476
rect 3467 16504 3479 16507
rect 4172 16504 4200 16535
rect 3467 16476 4200 16504
rect 4908 16504 4936 16535
rect 4982 16532 4988 16584
rect 5040 16572 5046 16584
rect 5261 16575 5319 16581
rect 5261 16572 5273 16575
rect 5040 16544 5273 16572
rect 5040 16532 5046 16544
rect 5261 16541 5273 16544
rect 5307 16572 5319 16575
rect 5350 16572 5356 16584
rect 5307 16544 5356 16572
rect 5307 16541 5319 16544
rect 5261 16535 5319 16541
rect 5350 16532 5356 16544
rect 5408 16532 5414 16584
rect 5445 16575 5503 16581
rect 5445 16541 5457 16575
rect 5491 16572 5503 16575
rect 5534 16572 5540 16584
rect 5491 16544 5540 16572
rect 5491 16541 5503 16544
rect 5445 16535 5503 16541
rect 5534 16532 5540 16544
rect 5592 16532 5598 16584
rect 5828 16581 5856 16612
rect 7101 16609 7113 16643
rect 7147 16640 7159 16643
rect 7484 16640 7512 16668
rect 8588 16640 8616 16668
rect 7147 16612 8616 16640
rect 7147 16609 7159 16612
rect 7101 16603 7159 16609
rect 5813 16575 5871 16581
rect 5813 16541 5825 16575
rect 5859 16541 5871 16575
rect 5813 16535 5871 16541
rect 5902 16532 5908 16584
rect 5960 16572 5966 16584
rect 6089 16575 6147 16581
rect 6089 16572 6101 16575
rect 5960 16544 6101 16572
rect 5960 16532 5966 16544
rect 6089 16541 6101 16544
rect 6135 16541 6147 16575
rect 6089 16535 6147 16541
rect 6454 16532 6460 16584
rect 6512 16532 6518 16584
rect 7009 16575 7067 16581
rect 7009 16541 7021 16575
rect 7055 16572 7067 16575
rect 7374 16572 7380 16584
rect 7055 16544 7380 16572
rect 7055 16541 7067 16544
rect 7009 16535 7067 16541
rect 7374 16532 7380 16544
rect 7432 16532 7438 16584
rect 7466 16532 7472 16584
rect 7524 16572 7530 16584
rect 7653 16575 7711 16581
rect 7653 16572 7665 16575
rect 7524 16544 7665 16572
rect 7524 16532 7530 16544
rect 7653 16541 7665 16544
rect 7699 16541 7711 16575
rect 7653 16535 7711 16541
rect 7834 16532 7840 16584
rect 7892 16572 7898 16584
rect 8573 16575 8631 16581
rect 8573 16572 8585 16575
rect 7892 16544 8585 16572
rect 7892 16532 7898 16544
rect 8573 16541 8585 16544
rect 8619 16541 8631 16575
rect 8573 16535 8631 16541
rect 8938 16532 8944 16584
rect 8996 16572 9002 16584
rect 9125 16575 9183 16581
rect 9125 16572 9137 16575
rect 8996 16544 9137 16572
rect 8996 16532 9002 16544
rect 9125 16541 9137 16544
rect 9171 16541 9183 16575
rect 9232 16572 9260 16680
rect 9858 16668 9864 16680
rect 9916 16668 9922 16720
rect 11606 16708 11612 16720
rect 9968 16680 11612 16708
rect 9306 16600 9312 16652
rect 9364 16640 9370 16652
rect 9364 16612 9541 16640
rect 9364 16600 9370 16612
rect 9513 16581 9541 16612
rect 9968 16581 9996 16680
rect 10594 16600 10600 16652
rect 10652 16600 10658 16652
rect 10962 16600 10968 16652
rect 11020 16600 11026 16652
rect 11440 16640 11468 16680
rect 11606 16668 11612 16680
rect 11664 16668 11670 16720
rect 11698 16668 11704 16720
rect 11756 16708 11762 16720
rect 17034 16708 17040 16720
rect 11756 16680 17040 16708
rect 11756 16668 11762 16680
rect 17034 16668 17040 16680
rect 17092 16668 17098 16720
rect 17402 16668 17408 16720
rect 17460 16668 17466 16720
rect 17862 16668 17868 16720
rect 17920 16668 17926 16720
rect 21361 16711 21419 16717
rect 21361 16677 21373 16711
rect 21407 16708 21419 16711
rect 24872 16708 24900 16739
rect 25498 16736 25504 16788
rect 25556 16736 25562 16788
rect 26786 16736 26792 16788
rect 26844 16776 26850 16788
rect 28166 16776 28172 16788
rect 26844 16748 28172 16776
rect 26844 16736 26850 16748
rect 28166 16736 28172 16748
rect 28224 16736 28230 16788
rect 28442 16736 28448 16788
rect 28500 16736 28506 16788
rect 31662 16776 31668 16788
rect 28966 16748 31668 16776
rect 21407 16680 24900 16708
rect 21407 16677 21419 16680
rect 21361 16671 21419 16677
rect 25130 16668 25136 16720
rect 25188 16708 25194 16720
rect 25188 16680 25452 16708
rect 25188 16668 25194 16680
rect 25424 16652 25452 16680
rect 25866 16668 25872 16720
rect 25924 16668 25930 16720
rect 26878 16668 26884 16720
rect 26936 16708 26942 16720
rect 27338 16708 27344 16720
rect 26936 16680 27344 16708
rect 26936 16668 26942 16680
rect 27338 16668 27344 16680
rect 27396 16668 27402 16720
rect 28966 16708 28994 16748
rect 31662 16736 31668 16748
rect 31720 16736 31726 16788
rect 31938 16736 31944 16788
rect 31996 16776 32002 16788
rect 32125 16779 32183 16785
rect 32125 16776 32137 16779
rect 31996 16748 32137 16776
rect 31996 16736 32002 16748
rect 32125 16745 32137 16748
rect 32171 16745 32183 16779
rect 32125 16739 32183 16745
rect 32490 16736 32496 16788
rect 32548 16736 32554 16788
rect 33410 16736 33416 16788
rect 33468 16776 33474 16788
rect 34054 16776 34060 16788
rect 33468 16748 34060 16776
rect 33468 16736 33474 16748
rect 34054 16736 34060 16748
rect 34112 16776 34118 16788
rect 35894 16776 35900 16788
rect 34112 16748 35900 16776
rect 34112 16736 34118 16748
rect 35894 16736 35900 16748
rect 35952 16776 35958 16788
rect 37182 16776 37188 16788
rect 35952 16748 37188 16776
rect 35952 16736 35958 16748
rect 37182 16736 37188 16748
rect 37240 16736 37246 16788
rect 37458 16736 37464 16788
rect 37516 16776 37522 16788
rect 37516 16748 37688 16776
rect 37516 16736 37522 16748
rect 27448 16680 28994 16708
rect 12710 16640 12716 16652
rect 11072 16612 11376 16640
rect 11440 16612 12716 16640
rect 9498 16575 9556 16581
rect 9232 16544 9444 16572
rect 9125 16535 9183 16541
rect 5629 16507 5687 16513
rect 5629 16504 5641 16507
rect 4908 16476 5641 16504
rect 3467 16473 3479 16476
rect 3421 16467 3479 16473
rect 1581 16439 1639 16445
rect 1581 16405 1593 16439
rect 1627 16405 1639 16439
rect 1581 16399 1639 16405
rect 3234 16396 3240 16448
rect 3292 16436 3298 16448
rect 3329 16439 3387 16445
rect 3329 16436 3341 16439
rect 3292 16408 3341 16436
rect 3292 16396 3298 16408
rect 3329 16405 3341 16408
rect 3375 16436 3387 16439
rect 3510 16436 3516 16448
rect 3375 16408 3516 16436
rect 3375 16405 3387 16408
rect 3329 16399 3387 16405
rect 3510 16396 3516 16408
rect 3568 16396 3574 16448
rect 4062 16396 4068 16448
rect 4120 16436 4126 16448
rect 4908 16436 4936 16476
rect 5629 16473 5641 16476
rect 5675 16473 5687 16507
rect 5629 16467 5687 16473
rect 5721 16507 5779 16513
rect 5721 16473 5733 16507
rect 5767 16504 5779 16507
rect 7558 16504 7564 16516
rect 5767 16476 5948 16504
rect 5767 16473 5779 16476
rect 5721 16467 5779 16473
rect 5920 16448 5948 16476
rect 6012 16476 7564 16504
rect 4120 16408 4936 16436
rect 5169 16439 5227 16445
rect 4120 16396 4126 16408
rect 5169 16405 5181 16439
rect 5215 16436 5227 16439
rect 5534 16436 5540 16448
rect 5215 16408 5540 16436
rect 5215 16405 5227 16408
rect 5169 16399 5227 16405
rect 5534 16396 5540 16408
rect 5592 16396 5598 16448
rect 5902 16396 5908 16448
rect 5960 16396 5966 16448
rect 6012 16445 6040 16476
rect 7558 16464 7564 16476
rect 7616 16464 7622 16516
rect 7742 16464 7748 16516
rect 7800 16504 7806 16516
rect 8021 16507 8079 16513
rect 8021 16504 8033 16507
rect 7800 16476 8033 16504
rect 7800 16464 7806 16476
rect 8021 16473 8033 16476
rect 8067 16473 8079 16507
rect 8021 16467 8079 16473
rect 9030 16464 9036 16516
rect 9088 16504 9094 16516
rect 9416 16513 9444 16544
rect 9498 16541 9510 16575
rect 9544 16541 9556 16575
rect 9498 16535 9556 16541
rect 9953 16575 10011 16581
rect 9953 16541 9965 16575
rect 9999 16541 10011 16575
rect 9953 16535 10011 16541
rect 10045 16575 10103 16581
rect 10045 16541 10057 16575
rect 10091 16541 10103 16575
rect 10045 16535 10103 16541
rect 9309 16507 9367 16513
rect 9309 16504 9321 16507
rect 9088 16476 9321 16504
rect 9088 16464 9094 16476
rect 9309 16473 9321 16476
rect 9355 16473 9367 16507
rect 9309 16467 9367 16473
rect 9401 16507 9459 16513
rect 9401 16473 9413 16507
rect 9447 16473 9459 16507
rect 10060 16504 10088 16535
rect 10134 16532 10140 16584
rect 10192 16572 10198 16584
rect 10413 16575 10471 16581
rect 10413 16572 10425 16575
rect 10192 16544 10425 16572
rect 10192 16532 10198 16544
rect 10413 16541 10425 16544
rect 10459 16541 10471 16575
rect 11072 16572 11100 16612
rect 10413 16535 10471 16541
rect 10520 16544 11100 16572
rect 10520 16504 10548 16544
rect 11238 16532 11244 16584
rect 11296 16532 11302 16584
rect 11348 16572 11376 16612
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 15286 16640 15292 16652
rect 12820 16612 15292 16640
rect 11614 16575 11672 16581
rect 11614 16572 11626 16575
rect 11348 16544 11626 16572
rect 11614 16541 11626 16544
rect 11660 16541 11672 16575
rect 11614 16535 11672 16541
rect 9401 16467 9459 16473
rect 9508 16476 10548 16504
rect 9508 16448 9536 16476
rect 10594 16464 10600 16516
rect 10652 16504 10658 16516
rect 11422 16504 11428 16516
rect 10652 16476 11428 16504
rect 10652 16464 10658 16476
rect 11422 16464 11428 16476
rect 11480 16464 11486 16516
rect 11517 16507 11575 16513
rect 11517 16473 11529 16507
rect 11563 16504 11575 16507
rect 12820 16504 12848 16612
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 15838 16640 15844 16652
rect 15764 16612 15844 16640
rect 15764 16581 15792 16612
rect 15838 16600 15844 16612
rect 15896 16600 15902 16652
rect 16040 16612 16252 16640
rect 15749 16575 15807 16581
rect 15749 16541 15761 16575
rect 15795 16541 15807 16575
rect 16040 16572 16068 16612
rect 15749 16535 15807 16541
rect 15856 16544 16068 16572
rect 11563 16476 12848 16504
rect 11563 16473 11575 16476
rect 11517 16467 11575 16473
rect 12986 16464 12992 16516
rect 13044 16504 13050 16516
rect 15856 16504 15884 16544
rect 16114 16532 16120 16584
rect 16172 16532 16178 16584
rect 16224 16572 16252 16612
rect 16960 16612 17908 16640
rect 16960 16572 16988 16612
rect 17880 16572 17908 16612
rect 19518 16600 19524 16652
rect 19576 16640 19582 16652
rect 20993 16643 21051 16649
rect 20993 16640 21005 16643
rect 19576 16612 21005 16640
rect 19576 16600 19582 16612
rect 20993 16609 21005 16612
rect 21039 16609 21051 16643
rect 20993 16603 21051 16609
rect 22278 16600 22284 16652
rect 22336 16640 22342 16652
rect 22336 16612 22876 16640
rect 22336 16600 22342 16612
rect 16224 16544 16988 16572
rect 17052 16544 17816 16572
rect 17880 16544 21128 16572
rect 13044 16476 15884 16504
rect 13044 16464 13050 16476
rect 15930 16464 15936 16516
rect 15988 16464 15994 16516
rect 16022 16464 16028 16516
rect 16080 16464 16086 16516
rect 17052 16513 17080 16544
rect 17037 16507 17095 16513
rect 17037 16504 17049 16507
rect 16132 16476 17049 16504
rect 5997 16439 6055 16445
rect 5997 16405 6009 16439
rect 6043 16405 6055 16439
rect 5997 16399 6055 16405
rect 6454 16396 6460 16448
rect 6512 16436 6518 16448
rect 7374 16436 7380 16448
rect 6512 16408 7380 16436
rect 6512 16396 6518 16408
rect 7374 16396 7380 16408
rect 7432 16396 7438 16448
rect 8202 16396 8208 16448
rect 8260 16436 8266 16448
rect 8481 16439 8539 16445
rect 8481 16436 8493 16439
rect 8260 16408 8493 16436
rect 8260 16396 8266 16408
rect 8481 16405 8493 16408
rect 8527 16405 8539 16439
rect 8481 16399 8539 16405
rect 9490 16396 9496 16448
rect 9548 16396 9554 16448
rect 9694 16439 9752 16445
rect 9694 16405 9706 16439
rect 9740 16436 9752 16439
rect 10962 16436 10968 16448
rect 9740 16408 10968 16436
rect 9740 16405 9752 16408
rect 9694 16399 9752 16405
rect 10962 16396 10968 16408
rect 11020 16396 11026 16448
rect 11146 16396 11152 16448
rect 11204 16436 11210 16448
rect 11801 16439 11859 16445
rect 11801 16436 11813 16439
rect 11204 16408 11813 16436
rect 11204 16396 11210 16408
rect 11801 16405 11813 16408
rect 11847 16405 11859 16439
rect 11801 16399 11859 16405
rect 15102 16396 15108 16448
rect 15160 16436 15166 16448
rect 16132 16436 16160 16476
rect 17037 16473 17049 16476
rect 17083 16473 17095 16507
rect 17218 16504 17224 16516
rect 17037 16467 17095 16473
rect 17144 16476 17224 16504
rect 15160 16408 16160 16436
rect 16301 16439 16359 16445
rect 15160 16396 15166 16408
rect 16301 16405 16313 16439
rect 16347 16436 16359 16439
rect 17144 16436 17172 16476
rect 17218 16464 17224 16476
rect 17276 16504 17282 16516
rect 17497 16507 17555 16513
rect 17276 16476 17448 16504
rect 17276 16464 17282 16476
rect 16347 16408 17172 16436
rect 17420 16436 17448 16476
rect 17497 16473 17509 16507
rect 17543 16504 17555 16507
rect 17586 16504 17592 16516
rect 17543 16476 17592 16504
rect 17543 16473 17555 16476
rect 17497 16467 17555 16473
rect 17586 16464 17592 16476
rect 17644 16464 17650 16516
rect 17681 16507 17739 16513
rect 17681 16473 17693 16507
rect 17727 16473 17739 16507
rect 17681 16467 17739 16473
rect 17696 16436 17724 16467
rect 17420 16408 17724 16436
rect 17788 16436 17816 16544
rect 20530 16464 20536 16516
rect 20588 16504 20594 16516
rect 20901 16507 20959 16513
rect 20901 16504 20913 16507
rect 20588 16476 20913 16504
rect 20588 16464 20594 16476
rect 20901 16473 20913 16476
rect 20947 16473 20959 16507
rect 21100 16504 21128 16544
rect 21174 16532 21180 16584
rect 21232 16532 21238 16584
rect 22186 16572 22192 16584
rect 21560 16544 22192 16572
rect 21453 16507 21511 16513
rect 21453 16504 21465 16507
rect 21100 16476 21465 16504
rect 20901 16467 20959 16473
rect 21453 16473 21465 16476
rect 21499 16504 21511 16507
rect 21560 16504 21588 16544
rect 22186 16532 22192 16544
rect 22244 16532 22250 16584
rect 22646 16532 22652 16584
rect 22704 16532 22710 16584
rect 22848 16581 22876 16612
rect 24302 16600 24308 16652
rect 24360 16640 24366 16652
rect 24360 16612 24900 16640
rect 24360 16600 24366 16612
rect 24872 16581 24900 16612
rect 25038 16600 25044 16652
rect 25096 16600 25102 16652
rect 25406 16600 25412 16652
rect 25464 16640 25470 16652
rect 25501 16643 25559 16649
rect 25501 16640 25513 16643
rect 25464 16612 25513 16640
rect 25464 16600 25470 16612
rect 25501 16609 25513 16612
rect 25547 16609 25559 16643
rect 25501 16603 25559 16609
rect 26326 16600 26332 16652
rect 26384 16640 26390 16652
rect 27448 16640 27476 16680
rect 29362 16668 29368 16720
rect 29420 16708 29426 16720
rect 31386 16708 31392 16720
rect 29420 16680 31392 16708
rect 29420 16668 29426 16680
rect 31386 16668 31392 16680
rect 31444 16668 31450 16720
rect 32030 16668 32036 16720
rect 32088 16668 32094 16720
rect 32398 16708 32404 16720
rect 32140 16680 32404 16708
rect 26384 16612 27476 16640
rect 26384 16600 26390 16612
rect 28534 16600 28540 16652
rect 28592 16600 28598 16652
rect 30834 16600 30840 16652
rect 30892 16640 30898 16652
rect 30892 16612 31432 16640
rect 30892 16600 30898 16612
rect 22833 16575 22891 16581
rect 22833 16541 22845 16575
rect 22879 16541 22891 16575
rect 22833 16535 22891 16541
rect 24857 16575 24915 16581
rect 24857 16541 24869 16575
rect 24903 16541 24915 16575
rect 24857 16535 24915 16541
rect 25130 16532 25136 16584
rect 25188 16532 25194 16584
rect 25685 16575 25743 16581
rect 25685 16541 25697 16575
rect 25731 16572 25743 16575
rect 25774 16572 25780 16584
rect 25731 16544 25780 16572
rect 25731 16541 25743 16544
rect 25685 16535 25743 16541
rect 25774 16532 25780 16544
rect 25832 16532 25838 16584
rect 28761 16575 28819 16581
rect 28761 16541 28773 16575
rect 28807 16572 28819 16575
rect 28994 16572 29000 16584
rect 28807 16544 29000 16572
rect 28807 16541 28819 16544
rect 28761 16535 28819 16541
rect 28994 16532 29000 16544
rect 29052 16532 29058 16584
rect 31294 16572 31300 16584
rect 29104 16544 31300 16572
rect 21499 16476 21588 16504
rect 21637 16507 21695 16513
rect 21499 16473 21511 16476
rect 21453 16467 21511 16473
rect 21637 16473 21649 16507
rect 21683 16473 21695 16507
rect 21637 16467 21695 16473
rect 21652 16436 21680 16467
rect 22278 16464 22284 16516
rect 22336 16504 22342 16516
rect 24118 16504 24124 16516
rect 22336 16476 24124 16504
rect 22336 16464 22342 16476
rect 24118 16464 24124 16476
rect 24176 16464 24182 16516
rect 24946 16464 24952 16516
rect 25004 16504 25010 16516
rect 25409 16507 25467 16513
rect 25409 16504 25421 16507
rect 25004 16476 25421 16504
rect 25004 16464 25010 16476
rect 25409 16473 25421 16476
rect 25455 16473 25467 16507
rect 25409 16467 25467 16473
rect 25958 16464 25964 16516
rect 26016 16464 26022 16516
rect 26142 16464 26148 16516
rect 26200 16504 26206 16516
rect 26878 16504 26884 16516
rect 26200 16476 26884 16504
rect 26200 16464 26206 16476
rect 26878 16464 26884 16476
rect 26936 16464 26942 16516
rect 28258 16464 28264 16516
rect 28316 16504 28322 16516
rect 28445 16507 28503 16513
rect 28445 16504 28457 16507
rect 28316 16476 28457 16504
rect 28316 16464 28322 16476
rect 28445 16473 28457 16476
rect 28491 16473 28503 16507
rect 29104 16504 29132 16544
rect 31294 16532 31300 16544
rect 31352 16532 31358 16584
rect 31404 16572 31432 16612
rect 31754 16600 31760 16652
rect 31812 16640 31818 16652
rect 32140 16640 32168 16680
rect 32398 16668 32404 16680
rect 32456 16668 32462 16720
rect 37660 16717 37688 16748
rect 38470 16736 38476 16788
rect 38528 16776 38534 16788
rect 38565 16779 38623 16785
rect 38565 16776 38577 16779
rect 38528 16748 38577 16776
rect 38528 16736 38534 16748
rect 38565 16745 38577 16748
rect 38611 16745 38623 16779
rect 38565 16739 38623 16745
rect 37645 16711 37703 16717
rect 37645 16677 37657 16711
rect 37691 16677 37703 16711
rect 37645 16671 37703 16677
rect 38378 16668 38384 16720
rect 38436 16708 38442 16720
rect 39298 16708 39304 16720
rect 38436 16680 39304 16708
rect 38436 16668 38442 16680
rect 39298 16668 39304 16680
rect 39356 16668 39362 16720
rect 31812 16612 32168 16640
rect 32217 16643 32275 16649
rect 31812 16600 31818 16612
rect 32217 16609 32229 16643
rect 32263 16640 32275 16643
rect 32306 16640 32312 16652
rect 32263 16612 32312 16640
rect 32263 16609 32275 16612
rect 32217 16603 32275 16609
rect 32306 16600 32312 16612
rect 32364 16600 32370 16652
rect 37734 16600 37740 16652
rect 37792 16600 37798 16652
rect 37829 16643 37887 16649
rect 37829 16609 37841 16643
rect 37875 16640 37887 16643
rect 38746 16640 38752 16652
rect 37875 16612 38752 16640
rect 37875 16609 37887 16612
rect 37829 16603 37887 16609
rect 38746 16600 38752 16612
rect 38804 16600 38810 16652
rect 31665 16575 31723 16581
rect 31665 16572 31677 16575
rect 31404 16544 31677 16572
rect 31665 16541 31677 16544
rect 31711 16541 31723 16575
rect 31665 16535 31723 16541
rect 32030 16532 32036 16584
rect 32088 16572 32094 16584
rect 32125 16575 32183 16581
rect 32125 16572 32137 16575
rect 32088 16544 32137 16572
rect 32088 16532 32094 16544
rect 32125 16541 32137 16544
rect 32171 16572 32183 16575
rect 33226 16572 33232 16584
rect 32171 16544 33232 16572
rect 32171 16541 32183 16544
rect 32125 16535 32183 16541
rect 33226 16532 33232 16544
rect 33284 16532 33290 16584
rect 33410 16532 33416 16584
rect 33468 16572 33474 16584
rect 37553 16575 37611 16581
rect 37553 16572 37565 16575
rect 33468 16544 37565 16572
rect 33468 16532 33474 16544
rect 37553 16541 37565 16544
rect 37599 16541 37611 16575
rect 37553 16535 37611 16541
rect 38013 16575 38071 16581
rect 38013 16541 38025 16575
rect 38059 16572 38071 16575
rect 38657 16575 38715 16581
rect 38657 16572 38669 16575
rect 38059 16544 38669 16572
rect 38059 16541 38071 16544
rect 38013 16535 38071 16541
rect 38657 16541 38669 16544
rect 38703 16572 38715 16575
rect 40218 16572 40224 16584
rect 38703 16544 40224 16572
rect 38703 16541 38715 16544
rect 38657 16535 38715 16541
rect 40218 16532 40224 16544
rect 40276 16532 40282 16584
rect 40310 16532 40316 16584
rect 40368 16572 40374 16584
rect 44269 16575 44327 16581
rect 44269 16572 44281 16575
rect 40368 16544 44281 16572
rect 40368 16532 40374 16544
rect 44269 16541 44281 16544
rect 44315 16541 44327 16575
rect 44269 16535 44327 16541
rect 28445 16467 28503 16473
rect 28828 16476 29132 16504
rect 17788 16408 21680 16436
rect 16347 16405 16359 16408
rect 16301 16399 16359 16405
rect 22186 16396 22192 16448
rect 22244 16436 22250 16448
rect 22738 16436 22744 16448
rect 22244 16408 22744 16436
rect 22244 16396 22250 16408
rect 22738 16396 22744 16408
rect 22796 16396 22802 16448
rect 25317 16439 25375 16445
rect 25317 16405 25329 16439
rect 25363 16436 25375 16439
rect 28828 16436 28856 16476
rect 29362 16464 29368 16516
rect 29420 16504 29426 16516
rect 29914 16504 29920 16516
rect 29420 16476 29920 16504
rect 29420 16464 29426 16476
rect 29914 16464 29920 16476
rect 29972 16464 29978 16516
rect 36814 16504 36820 16516
rect 31956 16476 32260 16504
rect 25363 16408 28856 16436
rect 25363 16405 25375 16408
rect 25317 16399 25375 16405
rect 28902 16396 28908 16448
rect 28960 16396 28966 16448
rect 29178 16396 29184 16448
rect 29236 16436 29242 16448
rect 31956 16436 31984 16476
rect 29236 16408 31984 16436
rect 32232 16436 32260 16476
rect 35912 16476 36820 16504
rect 35912 16436 35940 16476
rect 36814 16464 36820 16476
rect 36872 16464 36878 16516
rect 37826 16464 37832 16516
rect 37884 16504 37890 16516
rect 38197 16507 38255 16513
rect 38197 16504 38209 16507
rect 37884 16476 38209 16504
rect 37884 16464 37890 16476
rect 38197 16473 38209 16476
rect 38243 16473 38255 16507
rect 38197 16467 38255 16473
rect 38562 16464 38568 16516
rect 38620 16504 38626 16516
rect 42426 16504 42432 16516
rect 38620 16476 42432 16504
rect 38620 16464 38626 16476
rect 42426 16464 42432 16476
rect 42484 16464 42490 16516
rect 32232 16408 35940 16436
rect 29236 16396 29242 16408
rect 35986 16396 35992 16448
rect 36044 16436 36050 16448
rect 36906 16436 36912 16448
rect 36044 16408 36912 16436
rect 36044 16396 36050 16408
rect 36906 16396 36912 16408
rect 36964 16396 36970 16448
rect 37366 16396 37372 16448
rect 37424 16396 37430 16448
rect 44450 16396 44456 16448
rect 44508 16396 44514 16448
rect 1104 16346 44896 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 44896 16346
rect 1104 16272 44896 16294
rect 1581 16235 1639 16241
rect 1581 16201 1593 16235
rect 1627 16232 1639 16235
rect 2222 16232 2228 16244
rect 1627 16204 2228 16232
rect 1627 16201 1639 16204
rect 1581 16195 1639 16201
rect 2222 16192 2228 16204
rect 2280 16192 2286 16244
rect 5445 16235 5503 16241
rect 4448 16204 5396 16232
rect 2958 16164 2964 16176
rect 2056 16136 2964 16164
rect 842 16056 848 16108
rect 900 16096 906 16108
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 900 16068 1409 16096
rect 900 16056 906 16068
rect 1397 16065 1409 16068
rect 1443 16065 1455 16099
rect 1397 16059 1455 16065
rect 1762 16056 1768 16108
rect 1820 16096 1826 16108
rect 2056 16105 2084 16136
rect 2958 16124 2964 16136
rect 3016 16124 3022 16176
rect 1949 16099 2007 16105
rect 1949 16096 1961 16099
rect 1820 16068 1961 16096
rect 1820 16056 1826 16068
rect 1872 15960 1900 16068
rect 1949 16065 1961 16068
rect 1995 16065 2007 16099
rect 1949 16059 2007 16065
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16065 2099 16099
rect 2041 16059 2099 16065
rect 2133 16099 2191 16105
rect 2133 16065 2145 16099
rect 2179 16096 2191 16099
rect 2314 16096 2320 16108
rect 2179 16068 2320 16096
rect 2179 16065 2191 16068
rect 2133 16059 2191 16065
rect 2314 16056 2320 16068
rect 2372 16056 2378 16108
rect 2774 16056 2780 16108
rect 2832 16056 2838 16108
rect 3513 16099 3571 16105
rect 3513 16065 3525 16099
rect 3559 16065 3571 16099
rect 3513 16059 3571 16065
rect 2222 15988 2228 16040
rect 2280 15988 2286 16040
rect 2409 16031 2467 16037
rect 2409 15997 2421 16031
rect 2455 16028 2467 16031
rect 3418 16028 3424 16040
rect 2455 16000 3424 16028
rect 2455 15997 2467 16000
rect 2409 15991 2467 15997
rect 3418 15988 3424 16000
rect 3476 15988 3482 16040
rect 1872 15932 2912 15960
rect 2884 15901 2912 15932
rect 2869 15895 2927 15901
rect 2869 15861 2881 15895
rect 2915 15892 2927 15895
rect 3050 15892 3056 15904
rect 2915 15864 3056 15892
rect 2915 15861 2927 15864
rect 2869 15855 2927 15861
rect 3050 15852 3056 15864
rect 3108 15892 3114 15904
rect 3418 15892 3424 15904
rect 3108 15864 3424 15892
rect 3108 15852 3114 15864
rect 3418 15852 3424 15864
rect 3476 15852 3482 15904
rect 3528 15892 3556 16059
rect 3878 16056 3884 16108
rect 3936 16096 3942 16108
rect 4448 16096 4476 16204
rect 4525 16167 4583 16173
rect 4525 16133 4537 16167
rect 4571 16164 4583 16167
rect 5258 16164 5264 16176
rect 4571 16136 5264 16164
rect 4571 16133 4583 16136
rect 4525 16127 4583 16133
rect 5258 16124 5264 16136
rect 5316 16124 5322 16176
rect 3936 16068 4476 16096
rect 3936 16056 3942 16068
rect 4614 16056 4620 16108
rect 4672 16056 4678 16108
rect 5368 16096 5396 16204
rect 5445 16201 5457 16235
rect 5491 16232 5503 16235
rect 6362 16232 6368 16244
rect 5491 16204 6368 16232
rect 5491 16201 5503 16204
rect 5445 16195 5503 16201
rect 6362 16192 6368 16204
rect 6420 16192 6426 16244
rect 6638 16192 6644 16244
rect 6696 16192 6702 16244
rect 6914 16192 6920 16244
rect 6972 16232 6978 16244
rect 8573 16235 8631 16241
rect 6972 16204 8156 16232
rect 6972 16192 6978 16204
rect 5537 16167 5595 16173
rect 5537 16133 5549 16167
rect 5583 16164 5595 16167
rect 5994 16164 6000 16176
rect 5583 16136 6000 16164
rect 5583 16133 5595 16136
rect 5537 16127 5595 16133
rect 5994 16124 6000 16136
rect 6052 16124 6058 16176
rect 6181 16167 6239 16173
rect 6181 16133 6193 16167
rect 6227 16164 6239 16167
rect 6730 16164 6736 16176
rect 6227 16136 6736 16164
rect 6227 16133 6239 16136
rect 6181 16127 6239 16133
rect 6730 16124 6736 16136
rect 6788 16164 6794 16176
rect 8128 16164 8156 16204
rect 8573 16201 8585 16235
rect 8619 16232 8631 16235
rect 9122 16232 9128 16244
rect 8619 16204 9128 16232
rect 8619 16201 8631 16204
rect 8573 16195 8631 16201
rect 9122 16192 9128 16204
rect 9180 16192 9186 16244
rect 9490 16192 9496 16244
rect 9548 16232 9554 16244
rect 9548 16204 10732 16232
rect 9548 16192 9554 16204
rect 8846 16164 8852 16176
rect 6788 16136 8064 16164
rect 8128 16136 8852 16164
rect 6788 16124 6794 16136
rect 5368 16068 5764 16096
rect 3605 16031 3663 16037
rect 3605 15997 3617 16031
rect 3651 16028 3663 16031
rect 3694 16028 3700 16040
rect 3651 16000 3700 16028
rect 3651 15997 3663 16000
rect 3605 15991 3663 15997
rect 3694 15988 3700 16000
rect 3752 15988 3758 16040
rect 3786 15988 3792 16040
rect 3844 16028 3850 16040
rect 4065 16031 4123 16037
rect 4065 16028 4077 16031
rect 3844 16000 4077 16028
rect 3844 15988 3850 16000
rect 4065 15997 4077 16000
rect 4111 16028 4123 16031
rect 5736 16028 5764 16068
rect 5810 16056 5816 16108
rect 5868 16056 5874 16108
rect 6362 16056 6368 16108
rect 6420 16096 6426 16108
rect 7009 16099 7067 16105
rect 7009 16096 7021 16099
rect 6420 16068 7021 16096
rect 6420 16056 6426 16068
rect 7009 16065 7021 16068
rect 7055 16065 7067 16099
rect 7009 16059 7067 16065
rect 6914 16028 6920 16040
rect 4111 16000 4936 16028
rect 5736 16000 6920 16028
rect 4111 15997 4123 16000
rect 4065 15991 4123 15997
rect 4908 15960 4936 16000
rect 6914 15988 6920 16000
rect 6972 15988 6978 16040
rect 7024 16028 7052 16059
rect 7282 16056 7288 16108
rect 7340 16096 7346 16108
rect 7576 16105 7604 16136
rect 7377 16099 7435 16105
rect 7377 16096 7389 16099
rect 7340 16068 7389 16096
rect 7340 16056 7346 16068
rect 7377 16065 7389 16068
rect 7423 16065 7435 16099
rect 7377 16059 7435 16065
rect 7561 16099 7619 16105
rect 7561 16065 7573 16099
rect 7607 16065 7619 16099
rect 7561 16059 7619 16065
rect 7834 16056 7840 16108
rect 7892 16096 7898 16108
rect 7929 16099 7987 16105
rect 7929 16096 7941 16099
rect 7892 16068 7941 16096
rect 7892 16056 7898 16068
rect 7929 16065 7941 16068
rect 7975 16065 7987 16099
rect 8036 16096 8064 16136
rect 8846 16124 8852 16136
rect 8904 16124 8910 16176
rect 9398 16164 9404 16176
rect 9324 16136 9404 16164
rect 8036 16068 8725 16096
rect 7929 16059 7987 16065
rect 7024 16000 7420 16028
rect 7282 15960 7288 15972
rect 4908 15932 7288 15960
rect 7282 15920 7288 15932
rect 7340 15920 7346 15972
rect 4798 15892 4804 15904
rect 3528 15864 4804 15892
rect 4798 15852 4804 15864
rect 4856 15892 4862 15904
rect 6362 15892 6368 15904
rect 4856 15864 6368 15892
rect 4856 15852 4862 15864
rect 6362 15852 6368 15864
rect 6420 15852 6426 15904
rect 7392 15892 7420 16000
rect 8018 15988 8024 16040
rect 8076 16028 8082 16040
rect 8202 16028 8208 16040
rect 8076 16000 8208 16028
rect 8076 15988 8082 16000
rect 8202 15988 8208 16000
rect 8260 15988 8266 16040
rect 8297 16031 8355 16037
rect 8297 15997 8309 16031
rect 8343 15997 8355 16031
rect 8297 15991 8355 15997
rect 7742 15920 7748 15972
rect 7800 15960 7806 15972
rect 8312 15960 8340 15991
rect 8386 15988 8392 16040
rect 8444 16037 8450 16040
rect 8444 16031 8472 16037
rect 8460 15997 8472 16031
rect 8697 16028 8725 16068
rect 8754 16056 8760 16108
rect 8812 16056 8818 16108
rect 9030 16056 9036 16108
rect 9088 16096 9094 16108
rect 9217 16099 9275 16105
rect 9217 16096 9229 16099
rect 9088 16068 9229 16096
rect 9088 16056 9094 16068
rect 9217 16065 9229 16068
rect 9263 16065 9275 16099
rect 9217 16059 9275 16065
rect 9122 16028 9128 16040
rect 8697 16000 9128 16028
rect 8444 15991 8472 15997
rect 8444 15988 8450 15991
rect 9122 15988 9128 16000
rect 9180 16028 9186 16040
rect 9324 16037 9352 16136
rect 9398 16124 9404 16136
rect 9456 16124 9462 16176
rect 10502 16124 10508 16176
rect 10560 16124 10566 16176
rect 9585 16100 9643 16105
rect 9585 16099 9653 16100
rect 9585 16065 9597 16099
rect 9631 16065 9653 16099
rect 9585 16059 9653 16065
rect 9309 16031 9367 16037
rect 9309 16028 9321 16031
rect 9180 16000 9321 16028
rect 9180 15988 9186 16000
rect 9309 15997 9321 16000
rect 9355 15997 9367 16031
rect 9309 15991 9367 15997
rect 9493 16031 9551 16037
rect 9493 15997 9505 16031
rect 9539 15997 9551 16031
rect 9493 15991 9551 15997
rect 7800 15932 8340 15960
rect 8941 15963 8999 15969
rect 7800 15920 7806 15932
rect 8941 15929 8953 15963
rect 8987 15960 8999 15963
rect 9030 15960 9036 15972
rect 8987 15932 9036 15960
rect 8987 15929 8999 15932
rect 8941 15923 8999 15929
rect 9030 15920 9036 15932
rect 9088 15920 9094 15972
rect 9398 15920 9404 15972
rect 9456 15960 9462 15972
rect 9508 15960 9536 15991
rect 9456 15932 9536 15960
rect 9625 15960 9653 16059
rect 10318 16056 10324 16108
rect 10376 16056 10382 16108
rect 10594 16056 10600 16108
rect 10652 16056 10658 16108
rect 10704 16105 10732 16204
rect 10778 16192 10784 16244
rect 10836 16232 10842 16244
rect 10873 16235 10931 16241
rect 10873 16232 10885 16235
rect 10836 16204 10885 16232
rect 10836 16192 10842 16204
rect 10873 16201 10885 16204
rect 10919 16232 10931 16235
rect 11146 16232 11152 16244
rect 10919 16204 11152 16232
rect 10919 16201 10931 16204
rect 10873 16195 10931 16201
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 11422 16192 11428 16244
rect 11480 16232 11486 16244
rect 11606 16232 11612 16244
rect 11480 16204 11612 16232
rect 11480 16192 11486 16204
rect 11606 16192 11612 16204
rect 11664 16232 11670 16244
rect 15289 16235 15347 16241
rect 11664 16204 12388 16232
rect 11664 16192 11670 16204
rect 11054 16124 11060 16176
rect 11112 16164 11118 16176
rect 11793 16167 11851 16173
rect 11793 16164 11805 16167
rect 11112 16136 11805 16164
rect 11112 16124 11118 16136
rect 11793 16133 11805 16136
rect 11839 16164 11851 16167
rect 12158 16164 12164 16176
rect 11839 16136 12164 16164
rect 11839 16133 11851 16136
rect 11793 16127 11851 16133
rect 12158 16124 12164 16136
rect 12216 16124 12222 16176
rect 12360 16108 12388 16204
rect 15289 16201 15301 16235
rect 15335 16232 15347 16235
rect 15378 16232 15384 16244
rect 15335 16204 15384 16232
rect 15335 16201 15347 16204
rect 15289 16195 15347 16201
rect 15378 16192 15384 16204
rect 15436 16232 15442 16244
rect 15838 16232 15844 16244
rect 15436 16204 15844 16232
rect 15436 16192 15442 16204
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 16758 16192 16764 16244
rect 16816 16232 16822 16244
rect 17497 16235 17555 16241
rect 17497 16232 17509 16235
rect 16816 16204 17509 16232
rect 16816 16192 16822 16204
rect 17497 16201 17509 16204
rect 17543 16201 17555 16235
rect 17497 16195 17555 16201
rect 17770 16192 17776 16244
rect 17828 16232 17834 16244
rect 20070 16232 20076 16244
rect 17828 16204 20076 16232
rect 17828 16192 17834 16204
rect 20070 16192 20076 16204
rect 20128 16192 20134 16244
rect 20530 16192 20536 16244
rect 20588 16192 20594 16244
rect 22002 16192 22008 16244
rect 22060 16232 22066 16244
rect 22189 16235 22247 16241
rect 22189 16232 22201 16235
rect 22060 16204 22201 16232
rect 22060 16192 22066 16204
rect 22189 16201 22201 16204
rect 22235 16201 22247 16235
rect 22189 16195 22247 16201
rect 22738 16192 22744 16244
rect 22796 16232 22802 16244
rect 22796 16204 23520 16232
rect 22796 16192 22802 16204
rect 15194 16124 15200 16176
rect 15252 16124 15258 16176
rect 17586 16164 17592 16176
rect 15304 16136 17592 16164
rect 10689 16099 10747 16105
rect 10689 16065 10701 16099
rect 10735 16065 10747 16099
rect 10689 16059 10747 16065
rect 11606 16056 11612 16108
rect 11664 16056 11670 16108
rect 11882 16056 11888 16108
rect 11940 16056 11946 16108
rect 12066 16105 12072 16108
rect 12029 16099 12072 16105
rect 12029 16065 12041 16099
rect 12029 16059 12072 16065
rect 12066 16056 12072 16059
rect 12124 16056 12130 16108
rect 12342 16056 12348 16108
rect 12400 16056 12406 16108
rect 12618 16056 12624 16108
rect 12676 16096 12682 16108
rect 12713 16099 12771 16105
rect 12713 16096 12725 16099
rect 12676 16068 12725 16096
rect 12676 16056 12682 16068
rect 12713 16065 12725 16068
rect 12759 16065 12771 16099
rect 12713 16059 12771 16065
rect 12986 16056 12992 16108
rect 13044 16056 13050 16108
rect 10778 15988 10784 16040
rect 10836 16028 10842 16040
rect 13081 16031 13139 16037
rect 13081 16028 13093 16031
rect 10836 16000 13093 16028
rect 10836 15988 10842 16000
rect 13081 15997 13093 16000
rect 13127 16028 13139 16031
rect 15102 16028 15108 16040
rect 13127 16000 15108 16028
rect 13127 15997 13139 16000
rect 13081 15991 13139 15997
rect 15102 15988 15108 16000
rect 15160 15988 15166 16040
rect 10226 15960 10232 15972
rect 9625 15932 10232 15960
rect 9456 15920 9462 15932
rect 9214 15892 9220 15904
rect 7392 15864 9220 15892
rect 9214 15852 9220 15864
rect 9272 15892 9278 15904
rect 9625 15892 9653 15932
rect 10226 15920 10232 15932
rect 10284 15920 10290 15972
rect 11330 15920 11336 15972
rect 11388 15960 11394 15972
rect 12161 15963 12219 15969
rect 12161 15960 12173 15963
rect 11388 15932 12173 15960
rect 11388 15920 11394 15932
rect 12161 15929 12173 15932
rect 12207 15960 12219 15963
rect 12986 15960 12992 15972
rect 12207 15932 12992 15960
rect 12207 15929 12219 15932
rect 12161 15923 12219 15929
rect 12986 15920 12992 15932
rect 13044 15920 13050 15972
rect 15304 15960 15332 16136
rect 17586 16124 17592 16136
rect 17644 16164 17650 16176
rect 18601 16167 18659 16173
rect 18601 16164 18613 16167
rect 17644 16136 18613 16164
rect 17644 16124 17650 16136
rect 18601 16133 18613 16136
rect 18647 16133 18659 16167
rect 22278 16164 22284 16176
rect 18601 16127 18659 16133
rect 18708 16136 22284 16164
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16065 15715 16099
rect 15657 16059 15715 16065
rect 13188 15932 15332 15960
rect 15672 15960 15700 16059
rect 15838 16056 15844 16108
rect 15896 16056 15902 16108
rect 15930 16056 15936 16108
rect 15988 16056 15994 16108
rect 16077 16099 16135 16105
rect 16077 16065 16089 16099
rect 16123 16096 16135 16099
rect 16390 16096 16396 16108
rect 16123 16068 16396 16096
rect 16123 16065 16135 16068
rect 16077 16059 16135 16065
rect 16390 16056 16396 16068
rect 16448 16056 16454 16108
rect 16666 16056 16672 16108
rect 16724 16096 16730 16108
rect 17037 16099 17095 16105
rect 17037 16096 17049 16099
rect 16724 16068 17049 16096
rect 16724 16056 16730 16068
rect 17037 16065 17049 16068
rect 17083 16096 17095 16099
rect 17083 16068 17264 16096
rect 17083 16065 17095 16068
rect 17037 16059 17095 16065
rect 16942 15988 16948 16040
rect 17000 16028 17006 16040
rect 17129 16031 17187 16037
rect 17129 16028 17141 16031
rect 17000 16000 17141 16028
rect 17000 15988 17006 16000
rect 17129 15997 17141 16000
rect 17175 15997 17187 16031
rect 17236 16028 17264 16068
rect 17310 16056 17316 16108
rect 17368 16056 17374 16108
rect 18708 16096 18736 16136
rect 22278 16124 22284 16136
rect 22336 16124 22342 16176
rect 22462 16124 22468 16176
rect 22520 16164 22526 16176
rect 22520 16136 22968 16164
rect 22520 16124 22526 16136
rect 17420 16068 18736 16096
rect 17420 16028 17448 16068
rect 18874 16056 18880 16108
rect 18932 16056 18938 16108
rect 20070 16056 20076 16108
rect 20128 16056 20134 16108
rect 20346 16056 20352 16108
rect 20404 16056 20410 16108
rect 22370 16056 22376 16108
rect 22428 16056 22434 16108
rect 22646 16056 22652 16108
rect 22704 16056 22710 16108
rect 22940 16105 22968 16136
rect 22741 16099 22799 16105
rect 22741 16065 22753 16099
rect 22787 16065 22799 16099
rect 22741 16059 22799 16065
rect 22925 16099 22983 16105
rect 22925 16065 22937 16099
rect 22971 16065 22983 16099
rect 22925 16059 22983 16065
rect 23017 16099 23075 16105
rect 23017 16065 23029 16099
rect 23063 16096 23075 16099
rect 23382 16096 23388 16108
rect 23063 16068 23388 16096
rect 23063 16065 23075 16068
rect 23017 16059 23075 16065
rect 17236 16000 17448 16028
rect 17129 15991 17187 15997
rect 18598 15988 18604 16040
rect 18656 16028 18662 16040
rect 18693 16031 18751 16037
rect 18693 16028 18705 16031
rect 18656 16000 18705 16028
rect 18656 15988 18662 16000
rect 18693 15997 18705 16000
rect 18739 15997 18751 16031
rect 18693 15991 18751 15997
rect 20165 16031 20223 16037
rect 20165 15997 20177 16031
rect 20211 15997 20223 16031
rect 20165 15991 20223 15997
rect 15746 15960 15752 15972
rect 15672 15932 15752 15960
rect 9272 15864 9653 15892
rect 9272 15852 9278 15864
rect 9950 15852 9956 15904
rect 10008 15852 10014 15904
rect 10318 15852 10324 15904
rect 10376 15892 10382 15904
rect 10870 15892 10876 15904
rect 10376 15864 10876 15892
rect 10376 15852 10382 15864
rect 10870 15852 10876 15864
rect 10928 15852 10934 15904
rect 11146 15852 11152 15904
rect 11204 15892 11210 15904
rect 13188 15901 13216 15932
rect 15746 15920 15752 15932
rect 15804 15960 15810 15972
rect 16114 15960 16120 15972
rect 15804 15932 16120 15960
rect 15804 15920 15810 15932
rect 16114 15920 16120 15932
rect 16172 15920 16178 15972
rect 16206 15920 16212 15972
rect 16264 15920 16270 15972
rect 18322 15920 18328 15972
rect 18380 15960 18386 15972
rect 18380 15932 20116 15960
rect 18380 15920 18386 15932
rect 13173 15895 13231 15901
rect 13173 15892 13185 15895
rect 11204 15864 13185 15892
rect 11204 15852 11210 15864
rect 13173 15861 13185 15864
rect 13219 15861 13231 15895
rect 13173 15855 13231 15861
rect 13262 15852 13268 15904
rect 13320 15892 13326 15904
rect 13357 15895 13415 15901
rect 13357 15892 13369 15895
rect 13320 15864 13369 15892
rect 13320 15852 13326 15864
rect 13357 15861 13369 15864
rect 13403 15861 13415 15895
rect 13357 15855 13415 15861
rect 13722 15852 13728 15904
rect 13780 15892 13786 15904
rect 17034 15892 17040 15904
rect 13780 15864 17040 15892
rect 13780 15852 13786 15864
rect 17034 15852 17040 15864
rect 17092 15852 17098 15904
rect 17218 15852 17224 15904
rect 17276 15852 17282 15904
rect 18782 15852 18788 15904
rect 18840 15852 18846 15904
rect 19058 15852 19064 15904
rect 19116 15852 19122 15904
rect 20088 15901 20116 15932
rect 20180 15904 20208 15991
rect 21634 15988 21640 16040
rect 21692 16028 21698 16040
rect 22465 16031 22523 16037
rect 22465 16028 22477 16031
rect 21692 16000 22477 16028
rect 21692 15988 21698 16000
rect 22465 15997 22477 16000
rect 22511 15997 22523 16031
rect 22465 15991 22523 15997
rect 22554 15988 22560 16040
rect 22612 16028 22618 16040
rect 22763 16028 22791 16059
rect 23382 16056 23388 16068
rect 23440 16056 23446 16108
rect 23492 16096 23520 16204
rect 25130 16192 25136 16244
rect 25188 16232 25194 16244
rect 25409 16235 25467 16241
rect 25409 16232 25421 16235
rect 25188 16204 25421 16232
rect 25188 16192 25194 16204
rect 25409 16201 25421 16204
rect 25455 16232 25467 16235
rect 26145 16235 26203 16241
rect 25455 16204 26004 16232
rect 25455 16201 25467 16204
rect 25409 16195 25467 16201
rect 24946 16124 24952 16176
rect 25004 16164 25010 16176
rect 25976 16173 26004 16204
rect 26145 16201 26157 16235
rect 26191 16232 26203 16235
rect 26602 16232 26608 16244
rect 26191 16204 26608 16232
rect 26191 16201 26203 16204
rect 26145 16195 26203 16201
rect 26602 16192 26608 16204
rect 26660 16232 26666 16244
rect 28074 16232 28080 16244
rect 26660 16204 28080 16232
rect 26660 16192 26666 16204
rect 28074 16192 28080 16204
rect 28132 16192 28138 16244
rect 28994 16192 29000 16244
rect 29052 16192 29058 16244
rect 30834 16232 30840 16244
rect 30484 16204 30840 16232
rect 25041 16167 25099 16173
rect 25041 16164 25053 16167
rect 25004 16136 25053 16164
rect 25004 16124 25010 16136
rect 25041 16133 25053 16136
rect 25087 16133 25099 16167
rect 25777 16167 25835 16173
rect 25777 16164 25789 16167
rect 25041 16127 25099 16133
rect 25148 16136 25789 16164
rect 25148 16096 25176 16136
rect 25777 16133 25789 16136
rect 25823 16133 25835 16167
rect 25777 16127 25835 16133
rect 25961 16167 26019 16173
rect 25961 16133 25973 16167
rect 26007 16133 26019 16167
rect 25961 16127 26019 16133
rect 26326 16124 26332 16176
rect 26384 16164 26390 16176
rect 30484 16164 30512 16204
rect 30834 16192 30840 16204
rect 30892 16192 30898 16244
rect 32398 16192 32404 16244
rect 32456 16192 32462 16244
rect 32582 16192 32588 16244
rect 32640 16232 32646 16244
rect 32640 16204 32904 16232
rect 32640 16192 32646 16204
rect 26384 16136 30512 16164
rect 26384 16124 26390 16136
rect 30742 16124 30748 16176
rect 30800 16164 30806 16176
rect 30800 16136 32812 16164
rect 30800 16124 30806 16136
rect 23492 16068 25176 16096
rect 25225 16099 25283 16105
rect 25225 16065 25237 16099
rect 25271 16096 25283 16099
rect 25498 16096 25504 16108
rect 25271 16068 25504 16096
rect 25271 16065 25283 16068
rect 25225 16059 25283 16065
rect 25498 16056 25504 16068
rect 25556 16056 25562 16108
rect 25590 16056 25596 16108
rect 25648 16096 25654 16108
rect 27522 16096 27528 16108
rect 25648 16068 27528 16096
rect 25648 16056 25654 16068
rect 27522 16056 27528 16068
rect 27580 16096 27586 16108
rect 29181 16099 29239 16105
rect 29181 16096 29193 16099
rect 27580 16068 29193 16096
rect 27580 16056 27586 16068
rect 29181 16065 29193 16068
rect 29227 16065 29239 16099
rect 29181 16059 29239 16065
rect 29457 16099 29515 16105
rect 29457 16065 29469 16099
rect 29503 16065 29515 16099
rect 29457 16059 29515 16065
rect 29549 16099 29607 16105
rect 29549 16065 29561 16099
rect 29595 16096 29607 16099
rect 29638 16096 29644 16108
rect 29595 16068 29644 16096
rect 29595 16065 29607 16068
rect 29549 16059 29607 16065
rect 22612 16000 22791 16028
rect 22612 15988 22618 16000
rect 29362 15988 29368 16040
rect 29420 15988 29426 16040
rect 29472 16028 29500 16059
rect 29638 16056 29644 16068
rect 29696 16056 29702 16108
rect 29733 16099 29791 16105
rect 29733 16065 29745 16099
rect 29779 16096 29791 16099
rect 29822 16096 29828 16108
rect 29779 16068 29828 16096
rect 29779 16065 29791 16068
rect 29733 16059 29791 16065
rect 29822 16056 29828 16068
rect 29880 16056 29886 16108
rect 32582 16056 32588 16108
rect 32640 16056 32646 16108
rect 30098 16028 30104 16040
rect 29472 16000 30104 16028
rect 30098 15988 30104 16000
rect 30156 15988 30162 16040
rect 32398 15988 32404 16040
rect 32456 16028 32462 16040
rect 32677 16031 32735 16037
rect 32677 16028 32689 16031
rect 32456 16000 32689 16028
rect 32456 15988 32462 16000
rect 32677 15997 32689 16000
rect 32723 15997 32735 16031
rect 32784 16028 32812 16136
rect 32876 16096 32904 16204
rect 32950 16192 32956 16244
rect 33008 16192 33014 16244
rect 36538 16192 36544 16244
rect 36596 16232 36602 16244
rect 36596 16204 38654 16232
rect 36596 16192 36602 16204
rect 33686 16124 33692 16176
rect 33744 16164 33750 16176
rect 37277 16167 37335 16173
rect 37277 16164 37289 16167
rect 33744 16136 36032 16164
rect 33744 16124 33750 16136
rect 33045 16099 33103 16105
rect 33045 16096 33057 16099
rect 32876 16068 33057 16096
rect 33045 16065 33057 16068
rect 33091 16065 33103 16099
rect 33045 16059 33103 16065
rect 34882 16056 34888 16108
rect 34940 16096 34946 16108
rect 35069 16099 35127 16105
rect 35069 16096 35081 16099
rect 34940 16068 35081 16096
rect 34940 16056 34946 16068
rect 35069 16065 35081 16068
rect 35115 16065 35127 16099
rect 35069 16059 35127 16065
rect 35342 16056 35348 16108
rect 35400 16056 35406 16108
rect 35802 16056 35808 16108
rect 35860 16056 35866 16108
rect 36004 16105 36032 16136
rect 36280 16136 37289 16164
rect 36280 16105 36308 16136
rect 37277 16133 37289 16136
rect 37323 16133 37335 16167
rect 38626 16164 38654 16204
rect 38746 16192 38752 16244
rect 38804 16192 38810 16244
rect 42794 16164 42800 16176
rect 38626 16136 42800 16164
rect 37277 16127 37335 16133
rect 42794 16124 42800 16136
rect 42852 16124 42858 16176
rect 35989 16099 36047 16105
rect 35989 16065 36001 16099
rect 36035 16065 36047 16099
rect 35989 16059 36047 16065
rect 36265 16099 36323 16105
rect 36265 16065 36277 16099
rect 36311 16065 36323 16099
rect 36265 16059 36323 16065
rect 36357 16099 36415 16105
rect 36357 16065 36369 16099
rect 36403 16096 36415 16099
rect 36817 16099 36875 16105
rect 36403 16068 36768 16096
rect 36403 16065 36415 16068
rect 36357 16059 36415 16065
rect 34330 16028 34336 16040
rect 32784 16000 34336 16028
rect 32677 15991 32735 15997
rect 34330 15988 34336 16000
rect 34388 15988 34394 16040
rect 34790 15988 34796 16040
rect 34848 16028 34854 16040
rect 35161 16031 35219 16037
rect 35161 16028 35173 16031
rect 34848 16000 35173 16028
rect 34848 15988 34854 16000
rect 35161 15997 35173 16000
rect 35207 15997 35219 16031
rect 35161 15991 35219 15997
rect 36081 16031 36139 16037
rect 36081 15997 36093 16031
rect 36127 16028 36139 16031
rect 36538 16028 36544 16040
rect 36127 16000 36544 16028
rect 36127 15997 36139 16000
rect 36081 15991 36139 15997
rect 36538 15988 36544 16000
rect 36596 15988 36602 16040
rect 36630 15988 36636 16040
rect 36688 15988 36694 16040
rect 36740 16028 36768 16068
rect 36817 16065 36829 16099
rect 36863 16096 36875 16099
rect 36906 16096 36912 16108
rect 36863 16068 36912 16096
rect 36863 16065 36875 16068
rect 36817 16059 36875 16065
rect 36906 16056 36912 16068
rect 36964 16056 36970 16108
rect 39022 16056 39028 16108
rect 39080 16096 39086 16108
rect 39393 16099 39451 16105
rect 39393 16096 39405 16099
rect 39080 16068 39405 16096
rect 39080 16056 39086 16068
rect 39393 16065 39405 16068
rect 39439 16096 39451 16099
rect 44269 16099 44327 16105
rect 44269 16096 44281 16099
rect 39439 16068 44281 16096
rect 39439 16065 39451 16068
rect 39393 16059 39451 16065
rect 44269 16065 44281 16068
rect 44315 16065 44327 16099
rect 44269 16059 44327 16065
rect 36740 16000 36860 16028
rect 22646 15960 22652 15972
rect 20364 15932 22652 15960
rect 20073 15895 20131 15901
rect 20073 15861 20085 15895
rect 20119 15861 20131 15895
rect 20073 15855 20131 15861
rect 20162 15852 20168 15904
rect 20220 15892 20226 15904
rect 20364 15892 20392 15932
rect 22646 15920 22652 15932
rect 22704 15920 22710 15972
rect 22738 15920 22744 15972
rect 22796 15960 22802 15972
rect 25222 15960 25228 15972
rect 22796 15932 25228 15960
rect 22796 15920 22802 15932
rect 25222 15920 25228 15932
rect 25280 15920 25286 15972
rect 25866 15920 25872 15972
rect 25924 15960 25930 15972
rect 35434 15960 35440 15972
rect 25924 15932 35440 15960
rect 25924 15920 25930 15932
rect 20220 15864 20392 15892
rect 20220 15852 20226 15864
rect 22094 15852 22100 15904
rect 22152 15892 22158 15904
rect 22373 15895 22431 15901
rect 22373 15892 22385 15895
rect 22152 15864 22385 15892
rect 22152 15852 22158 15864
rect 22373 15861 22385 15864
rect 22419 15861 22431 15895
rect 22373 15855 22431 15861
rect 23014 15852 23020 15904
rect 23072 15852 23078 15904
rect 23198 15852 23204 15904
rect 23256 15852 23262 15904
rect 24118 15852 24124 15904
rect 24176 15892 24182 15904
rect 26326 15892 26332 15904
rect 24176 15864 26332 15892
rect 24176 15852 24182 15864
rect 26326 15852 26332 15864
rect 26384 15852 26390 15904
rect 26510 15852 26516 15904
rect 26568 15892 26574 15904
rect 29181 15895 29239 15901
rect 29181 15892 29193 15895
rect 26568 15864 29193 15892
rect 26568 15852 26574 15864
rect 29181 15861 29193 15864
rect 29227 15861 29239 15895
rect 29181 15855 29239 15861
rect 29730 15852 29736 15904
rect 29788 15852 29794 15904
rect 29917 15895 29975 15901
rect 29917 15861 29929 15895
rect 29963 15892 29975 15895
rect 30098 15892 30104 15904
rect 29963 15864 30104 15892
rect 29963 15861 29975 15864
rect 29917 15855 29975 15861
rect 30098 15852 30104 15864
rect 30156 15892 30162 15904
rect 32306 15892 32312 15904
rect 30156 15864 32312 15892
rect 30156 15852 30162 15864
rect 32306 15852 32312 15864
rect 32364 15852 32370 15904
rect 32582 15852 32588 15904
rect 32640 15852 32646 15904
rect 32766 15852 32772 15904
rect 32824 15892 32830 15904
rect 33594 15892 33600 15904
rect 32824 15864 33600 15892
rect 32824 15852 32830 15864
rect 33594 15852 33600 15864
rect 33652 15852 33658 15904
rect 35084 15901 35112 15932
rect 35434 15920 35440 15932
rect 35492 15920 35498 15972
rect 35529 15963 35587 15969
rect 35529 15929 35541 15963
rect 35575 15960 35587 15963
rect 35897 15963 35955 15969
rect 35897 15960 35909 15963
rect 35575 15932 35909 15960
rect 35575 15929 35587 15932
rect 35529 15923 35587 15929
rect 35897 15929 35909 15932
rect 35943 15929 35955 15963
rect 35897 15923 35955 15929
rect 36722 15920 36728 15972
rect 36780 15920 36786 15972
rect 36832 15960 36860 16000
rect 36998 15988 37004 16040
rect 37056 16028 37062 16040
rect 37921 16031 37979 16037
rect 37921 16028 37933 16031
rect 37056 16000 37933 16028
rect 37056 15988 37062 16000
rect 37921 15997 37933 16000
rect 37967 16028 37979 16031
rect 37967 16000 38608 16028
rect 37967 15997 37979 16000
rect 37921 15991 37979 15997
rect 38013 15963 38071 15969
rect 38013 15960 38025 15963
rect 36832 15932 38025 15960
rect 38013 15929 38025 15932
rect 38059 15929 38071 15963
rect 38580 15960 38608 16000
rect 38654 15988 38660 16040
rect 38712 15988 38718 16040
rect 44266 15960 44272 15972
rect 38580 15932 44272 15960
rect 38013 15923 38071 15929
rect 44266 15920 44272 15932
rect 44324 15920 44330 15972
rect 35069 15895 35127 15901
rect 35069 15861 35081 15895
rect 35115 15861 35127 15895
rect 35069 15855 35127 15861
rect 35621 15895 35679 15901
rect 35621 15861 35633 15895
rect 35667 15892 35679 15895
rect 35802 15892 35808 15904
rect 35667 15864 35808 15892
rect 35667 15861 35679 15864
rect 35621 15855 35679 15861
rect 35802 15852 35808 15864
rect 35860 15852 35866 15904
rect 37001 15895 37059 15901
rect 37001 15861 37013 15895
rect 37047 15892 37059 15895
rect 37182 15892 37188 15904
rect 37047 15864 37188 15892
rect 37047 15861 37059 15864
rect 37001 15855 37059 15861
rect 37182 15852 37188 15864
rect 37240 15852 37246 15904
rect 44450 15852 44456 15904
rect 44508 15852 44514 15904
rect 1104 15802 44896 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 44896 15802
rect 1104 15728 44896 15750
rect 1581 15691 1639 15697
rect 1581 15657 1593 15691
rect 1627 15688 1639 15691
rect 2774 15688 2780 15700
rect 1627 15660 2780 15688
rect 1627 15657 1639 15660
rect 1581 15651 1639 15657
rect 2774 15648 2780 15660
rect 2832 15648 2838 15700
rect 5353 15691 5411 15697
rect 5353 15657 5365 15691
rect 5399 15688 5411 15691
rect 5718 15688 5724 15700
rect 5399 15660 5724 15688
rect 5399 15657 5411 15660
rect 5353 15651 5411 15657
rect 5718 15648 5724 15660
rect 5776 15648 5782 15700
rect 5902 15648 5908 15700
rect 5960 15648 5966 15700
rect 6638 15648 6644 15700
rect 6696 15648 6702 15700
rect 6748 15660 7052 15688
rect 2869 15623 2927 15629
rect 2869 15589 2881 15623
rect 2915 15620 2927 15623
rect 2958 15620 2964 15632
rect 2915 15592 2964 15620
rect 2915 15589 2927 15592
rect 2869 15583 2927 15589
rect 2958 15580 2964 15592
rect 3016 15620 3022 15632
rect 3970 15620 3976 15632
rect 3016 15592 3976 15620
rect 3016 15580 3022 15592
rect 3970 15580 3976 15592
rect 4028 15580 4034 15632
rect 5442 15580 5448 15632
rect 5500 15580 5506 15632
rect 5629 15623 5687 15629
rect 5629 15589 5641 15623
rect 5675 15620 5687 15623
rect 6748 15620 6776 15660
rect 5675 15592 6776 15620
rect 5675 15589 5687 15592
rect 5629 15583 5687 15589
rect 3605 15555 3663 15561
rect 3605 15521 3617 15555
rect 3651 15552 3663 15555
rect 5460 15552 5488 15580
rect 3651 15524 5488 15552
rect 3651 15521 3663 15524
rect 3605 15515 3663 15521
rect 6270 15512 6276 15564
rect 6328 15512 6334 15564
rect 6638 15512 6644 15564
rect 6696 15552 6702 15564
rect 7024 15552 7052 15660
rect 7190 15648 7196 15700
rect 7248 15688 7254 15700
rect 7558 15688 7564 15700
rect 7248 15660 7564 15688
rect 7248 15648 7254 15660
rect 7558 15648 7564 15660
rect 7616 15648 7622 15700
rect 8481 15691 8539 15697
rect 8481 15657 8493 15691
rect 8527 15688 8539 15691
rect 8754 15688 8760 15700
rect 8527 15660 8760 15688
rect 8527 15657 8539 15660
rect 8481 15651 8539 15657
rect 8754 15648 8760 15660
rect 8812 15648 8818 15700
rect 8846 15648 8852 15700
rect 8904 15688 8910 15700
rect 8904 15660 10548 15688
rect 8904 15648 8910 15660
rect 7098 15580 7104 15632
rect 7156 15620 7162 15632
rect 7377 15623 7435 15629
rect 7377 15620 7389 15623
rect 7156 15592 7389 15620
rect 7156 15580 7162 15592
rect 7377 15589 7389 15592
rect 7423 15589 7435 15623
rect 9674 15620 9680 15632
rect 7377 15583 7435 15589
rect 9416 15592 9680 15620
rect 6696 15524 6960 15552
rect 7024 15524 7604 15552
rect 6696 15512 6702 15524
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 2406 15444 2412 15496
rect 2464 15444 2470 15496
rect 2682 15444 2688 15496
rect 2740 15484 2746 15496
rect 3421 15487 3479 15493
rect 3421 15484 3433 15487
rect 2740 15456 3433 15484
rect 2740 15444 2746 15456
rect 3421 15453 3433 15456
rect 3467 15484 3479 15487
rect 4062 15484 4068 15496
rect 3467 15456 4068 15484
rect 3467 15453 3479 15456
rect 3421 15447 3479 15453
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 5169 15487 5227 15493
rect 5169 15453 5181 15487
rect 5215 15484 5227 15487
rect 5445 15487 5503 15493
rect 5445 15484 5457 15487
rect 5215 15456 5457 15484
rect 5215 15453 5227 15456
rect 5169 15447 5227 15453
rect 5445 15453 5457 15456
rect 5491 15453 5503 15487
rect 5445 15447 5503 15453
rect 5721 15487 5779 15493
rect 5721 15453 5733 15487
rect 5767 15453 5779 15487
rect 5721 15447 5779 15453
rect 2869 15419 2927 15425
rect 2869 15385 2881 15419
rect 2915 15385 2927 15419
rect 5460 15416 5488 15447
rect 5626 15416 5632 15428
rect 5460 15388 5632 15416
rect 2869 15379 2927 15385
rect 2222 15308 2228 15360
rect 2280 15348 2286 15360
rect 2593 15351 2651 15357
rect 2593 15348 2605 15351
rect 2280 15320 2605 15348
rect 2280 15308 2286 15320
rect 2593 15317 2605 15320
rect 2639 15348 2651 15351
rect 2774 15348 2780 15360
rect 2639 15320 2780 15348
rect 2639 15317 2651 15320
rect 2593 15311 2651 15317
rect 2774 15308 2780 15320
rect 2832 15348 2838 15360
rect 2884 15348 2912 15379
rect 5626 15376 5632 15388
rect 5684 15376 5690 15428
rect 3234 15348 3240 15360
rect 2832 15320 3240 15348
rect 2832 15308 2838 15320
rect 3234 15308 3240 15320
rect 3292 15308 3298 15360
rect 3329 15351 3387 15357
rect 3329 15317 3341 15351
rect 3375 15348 3387 15351
rect 3510 15348 3516 15360
rect 3375 15320 3516 15348
rect 3375 15317 3387 15320
rect 3329 15311 3387 15317
rect 3510 15308 3516 15320
rect 3568 15308 3574 15360
rect 5736 15348 5764 15447
rect 5902 15444 5908 15496
rect 5960 15484 5966 15496
rect 6089 15487 6147 15493
rect 6089 15484 6101 15487
rect 5960 15456 6101 15484
rect 5960 15444 5966 15456
rect 6089 15453 6101 15456
rect 6135 15453 6147 15487
rect 6288 15484 6316 15512
rect 6932 15496 6960 15524
rect 6365 15487 6423 15493
rect 6365 15484 6377 15487
rect 6288 15456 6377 15484
rect 6089 15447 6147 15453
rect 6365 15453 6377 15456
rect 6411 15453 6423 15487
rect 6365 15447 6423 15453
rect 6509 15487 6567 15493
rect 6509 15453 6521 15487
rect 6555 15484 6567 15487
rect 6730 15484 6736 15496
rect 6555 15456 6736 15484
rect 6555 15453 6567 15456
rect 6509 15447 6567 15453
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 6825 15487 6883 15493
rect 6825 15453 6837 15487
rect 6871 15462 6883 15487
rect 6914 15462 6920 15496
rect 6871 15453 6920 15462
rect 6825 15447 6920 15453
rect 6840 15444 6920 15447
rect 6972 15444 6978 15496
rect 7245 15487 7303 15493
rect 7245 15453 7257 15487
rect 7291 15484 7303 15487
rect 7374 15484 7380 15496
rect 7291 15456 7380 15484
rect 7291 15453 7303 15456
rect 7245 15447 7303 15453
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 7576 15493 7604 15524
rect 7650 15512 7656 15564
rect 7708 15552 7714 15564
rect 7708 15524 8248 15552
rect 7708 15512 7714 15524
rect 7561 15487 7619 15493
rect 7561 15453 7573 15487
rect 7607 15453 7619 15487
rect 7926 15484 7932 15496
rect 7561 15447 7619 15453
rect 7668 15456 7932 15484
rect 6840 15434 6960 15444
rect 6270 15376 6276 15428
rect 6328 15376 6334 15428
rect 7006 15376 7012 15428
rect 7064 15376 7070 15428
rect 7098 15376 7104 15428
rect 7156 15376 7162 15428
rect 5902 15348 5908 15360
rect 5736 15320 5908 15348
rect 5902 15308 5908 15320
rect 5960 15308 5966 15360
rect 6730 15308 6736 15360
rect 6788 15348 6794 15360
rect 7668 15348 7696 15456
rect 7926 15444 7932 15456
rect 7984 15484 7990 15496
rect 8021 15487 8079 15493
rect 8021 15484 8033 15487
rect 7984 15456 8033 15484
rect 7984 15444 7990 15456
rect 8021 15453 8033 15456
rect 8067 15453 8079 15487
rect 8021 15447 8079 15453
rect 8110 15444 8116 15496
rect 8168 15444 8174 15496
rect 8220 15493 8248 15524
rect 8205 15487 8263 15493
rect 8205 15453 8217 15487
rect 8251 15453 8263 15487
rect 8205 15447 8263 15453
rect 8389 15487 8447 15493
rect 8389 15453 8401 15487
rect 8435 15484 8447 15487
rect 8481 15487 8539 15493
rect 8481 15484 8493 15487
rect 8435 15456 8493 15484
rect 8435 15453 8447 15456
rect 8389 15447 8447 15453
rect 8481 15453 8493 15456
rect 8527 15453 8539 15487
rect 8481 15447 8539 15453
rect 8570 15444 8576 15496
rect 8628 15484 8634 15496
rect 9416 15493 9444 15592
rect 9674 15580 9680 15592
rect 9732 15580 9738 15632
rect 10520 15620 10548 15660
rect 10594 15648 10600 15700
rect 10652 15688 10658 15700
rect 10652 15660 11744 15688
rect 10652 15648 10658 15660
rect 10870 15620 10876 15632
rect 10520 15592 10876 15620
rect 10870 15580 10876 15592
rect 10928 15580 10934 15632
rect 11606 15620 11612 15632
rect 11072 15592 11612 15620
rect 9490 15512 9496 15564
rect 9548 15512 9554 15564
rect 9953 15555 10011 15561
rect 9953 15521 9965 15555
rect 9999 15552 10011 15555
rect 10318 15552 10324 15564
rect 9999 15524 10324 15552
rect 9999 15521 10011 15524
rect 9953 15515 10011 15521
rect 10318 15512 10324 15524
rect 10376 15512 10382 15564
rect 10410 15512 10416 15564
rect 10468 15512 10474 15564
rect 11072 15561 11100 15592
rect 11606 15580 11612 15592
rect 11664 15580 11670 15632
rect 11057 15555 11115 15561
rect 11057 15521 11069 15555
rect 11103 15521 11115 15555
rect 11716 15552 11744 15660
rect 12618 15648 12624 15700
rect 12676 15688 12682 15700
rect 14645 15691 14703 15697
rect 12676 15660 13308 15688
rect 12676 15648 12682 15660
rect 12710 15580 12716 15632
rect 12768 15620 12774 15632
rect 12894 15620 12900 15632
rect 12768 15592 12900 15620
rect 12768 15580 12774 15592
rect 12894 15580 12900 15592
rect 12952 15580 12958 15632
rect 12986 15580 12992 15632
rect 13044 15620 13050 15632
rect 13081 15623 13139 15629
rect 13081 15620 13093 15623
rect 13044 15592 13093 15620
rect 13044 15580 13050 15592
rect 13081 15589 13093 15592
rect 13127 15589 13139 15623
rect 13081 15583 13139 15589
rect 12802 15552 12808 15564
rect 11716 15524 12808 15552
rect 11057 15515 11115 15521
rect 8665 15487 8723 15493
rect 8665 15484 8677 15487
rect 8628 15456 8677 15484
rect 8628 15444 8634 15456
rect 8665 15453 8677 15456
rect 8711 15453 8723 15487
rect 8665 15447 8723 15453
rect 8941 15487 8999 15493
rect 8941 15453 8953 15487
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 9401 15487 9459 15493
rect 9401 15453 9413 15487
rect 9447 15453 9459 15487
rect 9401 15447 9459 15453
rect 8956 15416 8984 15447
rect 7760 15388 8984 15416
rect 9508 15416 9536 15512
rect 9766 15444 9772 15496
rect 9824 15484 9830 15496
rect 11072 15484 11100 15515
rect 12802 15512 12808 15524
rect 12860 15552 12866 15564
rect 13280 15552 13308 15660
rect 14645 15657 14657 15691
rect 14691 15688 14703 15691
rect 14918 15688 14924 15700
rect 14691 15660 14924 15688
rect 14691 15657 14703 15660
rect 14645 15651 14703 15657
rect 14918 15648 14924 15660
rect 14976 15688 14982 15700
rect 16485 15691 16543 15697
rect 14976 15660 16252 15688
rect 14976 15648 14982 15660
rect 13909 15623 13967 15629
rect 13909 15589 13921 15623
rect 13955 15620 13967 15623
rect 14366 15620 14372 15632
rect 13955 15592 14372 15620
rect 13955 15589 13967 15592
rect 13909 15583 13967 15589
rect 14366 15580 14372 15592
rect 14424 15580 14430 15632
rect 15930 15580 15936 15632
rect 15988 15620 15994 15632
rect 16114 15620 16120 15632
rect 15988 15592 16120 15620
rect 15988 15580 15994 15592
rect 16114 15580 16120 15592
rect 16172 15580 16178 15632
rect 16224 15620 16252 15660
rect 16485 15657 16497 15691
rect 16531 15688 16543 15691
rect 20162 15688 20168 15700
rect 16531 15660 20168 15688
rect 16531 15657 16543 15660
rect 16485 15651 16543 15657
rect 20162 15648 20168 15660
rect 20220 15648 20226 15700
rect 22278 15648 22284 15700
rect 22336 15648 22342 15700
rect 22554 15648 22560 15700
rect 22612 15688 22618 15700
rect 22741 15691 22799 15697
rect 22741 15688 22753 15691
rect 22612 15660 22753 15688
rect 22612 15648 22618 15660
rect 22741 15657 22753 15660
rect 22787 15657 22799 15691
rect 22741 15651 22799 15657
rect 23842 15648 23848 15700
rect 23900 15648 23906 15700
rect 25590 15648 25596 15700
rect 25648 15688 25654 15700
rect 25648 15660 25728 15688
rect 25648 15648 25654 15660
rect 17770 15620 17776 15632
rect 16224 15592 17776 15620
rect 17770 15580 17776 15592
rect 17828 15580 17834 15632
rect 17954 15580 17960 15632
rect 18012 15620 18018 15632
rect 18012 15592 18460 15620
rect 18012 15580 18018 15592
rect 14829 15555 14887 15561
rect 14829 15552 14841 15555
rect 12860 15524 13124 15552
rect 13280 15524 14841 15552
rect 12860 15512 12866 15524
rect 9824 15456 11100 15484
rect 9824 15444 9830 15456
rect 11146 15444 11152 15496
rect 11204 15444 11210 15496
rect 11517 15487 11575 15493
rect 11517 15453 11529 15487
rect 11563 15453 11575 15487
rect 11517 15447 11575 15453
rect 11532 15416 11560 15447
rect 11698 15444 11704 15496
rect 11756 15444 11762 15496
rect 12529 15487 12587 15493
rect 12529 15484 12541 15487
rect 11808 15456 12541 15484
rect 11808 15416 11836 15456
rect 12529 15453 12541 15456
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 12710 15444 12716 15496
rect 12768 15444 12774 15496
rect 12894 15444 12900 15496
rect 12952 15493 12958 15496
rect 12952 15484 12960 15493
rect 13096 15484 13124 15524
rect 14829 15521 14841 15524
rect 14875 15521 14887 15555
rect 14829 15515 14887 15521
rect 15102 15512 15108 15564
rect 15160 15552 15166 15564
rect 16022 15552 16028 15564
rect 15160 15524 16028 15552
rect 15160 15512 15166 15524
rect 16022 15512 16028 15524
rect 16080 15512 16086 15564
rect 14090 15484 14096 15496
rect 12952 15456 12997 15484
rect 13096 15456 14096 15484
rect 12952 15447 12960 15456
rect 12952 15444 12958 15447
rect 14090 15444 14096 15456
rect 14148 15444 14154 15496
rect 14182 15444 14188 15496
rect 14240 15484 14246 15496
rect 14461 15487 14519 15493
rect 14461 15484 14473 15487
rect 14240 15456 14473 15484
rect 14240 15444 14246 15456
rect 14461 15453 14473 15456
rect 14507 15453 14519 15487
rect 14461 15447 14519 15453
rect 14734 15444 14740 15496
rect 14792 15484 14798 15496
rect 15930 15484 15936 15496
rect 14792 15456 15936 15484
rect 14792 15444 14798 15456
rect 15930 15444 15936 15456
rect 15988 15444 15994 15496
rect 16390 15493 16396 15496
rect 16353 15487 16396 15493
rect 16353 15453 16365 15487
rect 16353 15447 16396 15453
rect 16390 15444 16396 15447
rect 16448 15444 16454 15496
rect 16758 15444 16764 15496
rect 16816 15484 16822 15496
rect 17681 15487 17739 15493
rect 17681 15484 17693 15487
rect 16816 15456 17693 15484
rect 16816 15444 16822 15456
rect 17681 15453 17693 15456
rect 17727 15453 17739 15487
rect 17681 15447 17739 15453
rect 17954 15444 17960 15496
rect 18012 15444 18018 15496
rect 18046 15444 18052 15496
rect 18104 15493 18110 15496
rect 18432 15493 18460 15592
rect 19058 15580 19064 15632
rect 19116 15620 19122 15632
rect 25700 15620 25728 15660
rect 28074 15648 28080 15700
rect 28132 15648 28138 15700
rect 28258 15648 28264 15700
rect 28316 15648 28322 15700
rect 29086 15648 29092 15700
rect 29144 15688 29150 15700
rect 29549 15691 29607 15697
rect 29549 15688 29561 15691
rect 29144 15660 29561 15688
rect 29144 15648 29150 15660
rect 29549 15657 29561 15660
rect 29595 15657 29607 15691
rect 29549 15651 29607 15657
rect 29914 15648 29920 15700
rect 29972 15648 29978 15700
rect 31846 15648 31852 15700
rect 31904 15688 31910 15700
rect 32401 15691 32459 15697
rect 32401 15688 32413 15691
rect 31904 15660 32413 15688
rect 31904 15648 31910 15660
rect 32401 15657 32413 15660
rect 32447 15657 32459 15691
rect 32401 15651 32459 15657
rect 31754 15620 31760 15632
rect 19116 15592 24992 15620
rect 25700 15592 31760 15620
rect 19116 15580 19122 15592
rect 22462 15512 22468 15564
rect 22520 15552 22526 15564
rect 24964 15552 24992 15592
rect 31754 15580 31760 15592
rect 31812 15580 31818 15632
rect 27893 15555 27951 15561
rect 27893 15552 27905 15555
rect 22520 15524 24900 15552
rect 24964 15524 27905 15552
rect 22520 15512 22526 15524
rect 18104 15484 18112 15493
rect 18250 15487 18308 15493
rect 18250 15484 18262 15487
rect 18104 15456 18149 15484
rect 18104 15447 18112 15456
rect 18248 15453 18262 15484
rect 18296 15453 18308 15487
rect 18248 15447 18308 15453
rect 18417 15487 18475 15493
rect 18417 15453 18429 15487
rect 18463 15484 18475 15487
rect 18506 15484 18512 15496
rect 18463 15456 18512 15484
rect 18463 15453 18475 15456
rect 18417 15447 18475 15453
rect 18104 15444 18110 15447
rect 12161 15419 12219 15425
rect 12161 15416 12173 15419
rect 9508 15388 11836 15416
rect 11900 15388 12173 15416
rect 7760 15357 7788 15388
rect 6788 15320 7696 15348
rect 7745 15351 7803 15357
rect 6788 15308 6794 15320
rect 7745 15317 7757 15351
rect 7791 15317 7803 15351
rect 7745 15311 7803 15317
rect 8478 15308 8484 15360
rect 8536 15348 8542 15360
rect 9030 15348 9036 15360
rect 8536 15320 9036 15348
rect 8536 15308 8542 15320
rect 9030 15308 9036 15320
rect 9088 15308 9094 15360
rect 9125 15351 9183 15357
rect 9125 15317 9137 15351
rect 9171 15348 9183 15351
rect 10042 15348 10048 15360
rect 9171 15320 10048 15348
rect 9171 15317 9183 15320
rect 9125 15311 9183 15317
rect 10042 15308 10048 15320
rect 10100 15308 10106 15360
rect 10778 15308 10784 15360
rect 10836 15308 10842 15360
rect 10870 15308 10876 15360
rect 10928 15348 10934 15360
rect 11900 15348 11928 15388
rect 12161 15385 12173 15388
rect 12207 15385 12219 15419
rect 12161 15379 12219 15385
rect 12342 15376 12348 15428
rect 12400 15416 12406 15428
rect 12802 15416 12808 15428
rect 12400 15388 12808 15416
rect 12400 15376 12406 15388
rect 12802 15376 12808 15388
rect 12860 15376 12866 15428
rect 13722 15376 13728 15428
rect 13780 15376 13786 15428
rect 13906 15376 13912 15428
rect 13964 15416 13970 15428
rect 14277 15419 14335 15425
rect 14277 15416 14289 15419
rect 13964 15388 14289 15416
rect 13964 15376 13970 15388
rect 14277 15385 14289 15388
rect 14323 15385 14335 15419
rect 14277 15379 14335 15385
rect 14366 15376 14372 15428
rect 14424 15376 14430 15428
rect 16117 15419 16175 15425
rect 16117 15385 16129 15419
rect 16163 15385 16175 15419
rect 16117 15379 16175 15385
rect 10928 15320 11928 15348
rect 10928 15308 10934 15320
rect 11974 15308 11980 15360
rect 12032 15348 12038 15360
rect 12069 15351 12127 15357
rect 12069 15348 12081 15351
rect 12032 15320 12081 15348
rect 12032 15308 12038 15320
rect 12069 15317 12081 15320
rect 12115 15317 12127 15351
rect 12069 15311 12127 15317
rect 14734 15308 14740 15360
rect 14792 15348 14798 15360
rect 15838 15348 15844 15360
rect 14792 15320 15844 15348
rect 14792 15308 14798 15320
rect 15838 15308 15844 15320
rect 15896 15348 15902 15360
rect 16132 15348 16160 15379
rect 16206 15376 16212 15428
rect 16264 15376 16270 15428
rect 17865 15419 17923 15425
rect 17865 15385 17877 15419
rect 17911 15385 17923 15419
rect 17865 15379 17923 15385
rect 15896 15320 16160 15348
rect 15896 15308 15902 15320
rect 16298 15308 16304 15360
rect 16356 15348 16362 15360
rect 16482 15348 16488 15360
rect 16356 15320 16488 15348
rect 16356 15308 16362 15320
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 17494 15308 17500 15360
rect 17552 15348 17558 15360
rect 17880 15348 17908 15379
rect 18138 15376 18144 15428
rect 18196 15416 18202 15428
rect 18248 15416 18276 15447
rect 18506 15444 18512 15456
rect 18564 15444 18570 15496
rect 18690 15444 18696 15496
rect 18748 15444 18754 15496
rect 18874 15493 18880 15496
rect 18837 15487 18880 15493
rect 18837 15453 18849 15487
rect 18837 15447 18880 15453
rect 18874 15444 18880 15447
rect 18932 15444 18938 15496
rect 22370 15444 22376 15496
rect 22428 15484 22434 15496
rect 22557 15487 22615 15493
rect 22557 15484 22569 15487
rect 22428 15456 22569 15484
rect 22428 15444 22434 15456
rect 22557 15453 22569 15456
rect 22603 15453 22615 15487
rect 22557 15447 22615 15453
rect 23198 15444 23204 15496
rect 23256 15484 23262 15496
rect 23845 15487 23903 15493
rect 23845 15484 23857 15487
rect 23256 15456 23857 15484
rect 23256 15444 23262 15456
rect 23845 15453 23857 15456
rect 23891 15453 23903 15487
rect 23845 15447 23903 15453
rect 23937 15487 23995 15493
rect 23937 15453 23949 15487
rect 23983 15453 23995 15487
rect 24872 15484 24900 15524
rect 27893 15521 27905 15524
rect 27939 15521 27951 15555
rect 29178 15552 29184 15564
rect 27893 15515 27951 15521
rect 28000 15524 29184 15552
rect 25409 15487 25467 15493
rect 25409 15484 25421 15487
rect 24872 15456 25421 15484
rect 23937 15447 23995 15453
rect 25409 15453 25421 15456
rect 25455 15453 25467 15487
rect 25409 15447 25467 15453
rect 25501 15487 25559 15493
rect 25501 15453 25513 15487
rect 25547 15453 25559 15487
rect 25501 15447 25559 15453
rect 25685 15487 25743 15493
rect 25685 15453 25697 15487
rect 25731 15484 25743 15487
rect 26326 15484 26332 15496
rect 25731 15456 26332 15484
rect 25731 15453 25743 15456
rect 25685 15447 25743 15453
rect 18196 15388 18276 15416
rect 18601 15419 18659 15425
rect 18196 15376 18202 15388
rect 18601 15385 18613 15419
rect 18647 15385 18659 15419
rect 18601 15379 18659 15385
rect 18616 15348 18644 15379
rect 19426 15376 19432 15428
rect 19484 15416 19490 15428
rect 22278 15416 22284 15428
rect 19484 15388 22284 15416
rect 19484 15376 19490 15388
rect 22278 15376 22284 15388
rect 22336 15376 22342 15428
rect 23290 15376 23296 15428
rect 23348 15416 23354 15428
rect 23952 15416 23980 15447
rect 25516 15416 25544 15447
rect 26326 15444 26332 15456
rect 26384 15444 26390 15496
rect 26694 15444 26700 15496
rect 26752 15484 26758 15496
rect 28000 15484 28028 15524
rect 29178 15512 29184 15524
rect 29236 15512 29242 15564
rect 32416 15552 32444 15651
rect 32582 15648 32588 15700
rect 32640 15648 32646 15700
rect 32858 15648 32864 15700
rect 32916 15648 32922 15700
rect 33318 15648 33324 15700
rect 33376 15648 33382 15700
rect 33502 15648 33508 15700
rect 33560 15648 33566 15700
rect 34241 15691 34299 15697
rect 34241 15657 34253 15691
rect 34287 15688 34299 15691
rect 34330 15688 34336 15700
rect 34287 15660 34336 15688
rect 34287 15657 34299 15660
rect 34241 15651 34299 15657
rect 34330 15648 34336 15660
rect 34388 15648 34394 15700
rect 34425 15691 34483 15697
rect 34425 15657 34437 15691
rect 34471 15688 34483 15691
rect 34790 15688 34796 15700
rect 34471 15660 34796 15688
rect 34471 15657 34483 15660
rect 34425 15651 34483 15657
rect 34790 15648 34796 15660
rect 34848 15648 34854 15700
rect 35161 15691 35219 15697
rect 35161 15657 35173 15691
rect 35207 15688 35219 15691
rect 35207 15660 36584 15688
rect 35207 15657 35219 15660
rect 35161 15651 35219 15657
rect 32674 15580 32680 15632
rect 32732 15620 32738 15632
rect 33042 15620 33048 15632
rect 32732 15592 33048 15620
rect 32732 15580 32738 15592
rect 33042 15580 33048 15592
rect 33100 15580 33106 15632
rect 33226 15620 33232 15632
rect 33152 15592 33232 15620
rect 33152 15561 33180 15592
rect 33226 15580 33232 15592
rect 33284 15580 33290 15632
rect 36556 15620 36584 15660
rect 36998 15648 37004 15700
rect 37056 15648 37062 15700
rect 37274 15688 37280 15700
rect 37108 15660 37280 15688
rect 37108 15620 37136 15660
rect 37274 15648 37280 15660
rect 37332 15648 37338 15700
rect 36556 15592 37136 15620
rect 32861 15555 32919 15561
rect 32861 15552 32873 15555
rect 32416 15524 32873 15552
rect 32861 15521 32873 15524
rect 32907 15521 32919 15555
rect 32861 15515 32919 15521
rect 33137 15555 33195 15561
rect 33137 15521 33149 15555
rect 33183 15521 33195 15555
rect 33137 15515 33195 15521
rect 34698 15512 34704 15564
rect 34756 15512 34762 15564
rect 34790 15512 34796 15564
rect 34848 15512 34854 15564
rect 40957 15555 41015 15561
rect 40957 15521 40969 15555
rect 41003 15552 41015 15555
rect 41414 15552 41420 15564
rect 41003 15524 41420 15552
rect 41003 15521 41015 15524
rect 40957 15515 41015 15521
rect 41414 15512 41420 15524
rect 41472 15512 41478 15564
rect 26752 15456 28028 15484
rect 28077 15487 28135 15493
rect 26752 15444 26758 15456
rect 28077 15453 28089 15487
rect 28123 15453 28135 15487
rect 28077 15447 28135 15453
rect 23348 15388 23980 15416
rect 24136 15388 25544 15416
rect 23348 15376 23354 15388
rect 17552 15320 18644 15348
rect 18986 15351 19044 15357
rect 17552 15308 17558 15320
rect 18986 15317 18998 15351
rect 19032 15348 19044 15351
rect 23750 15348 23756 15360
rect 19032 15320 23756 15348
rect 19032 15317 19044 15320
rect 18986 15311 19044 15317
rect 23750 15308 23756 15320
rect 23808 15348 23814 15360
rect 24136 15348 24164 15388
rect 26234 15376 26240 15428
rect 26292 15416 26298 15428
rect 26881 15419 26939 15425
rect 26881 15416 26893 15419
rect 26292 15388 26893 15416
rect 26292 15376 26298 15388
rect 26881 15385 26893 15388
rect 26927 15416 26939 15419
rect 26970 15416 26976 15428
rect 26927 15388 26976 15416
rect 26927 15385 26939 15388
rect 26881 15379 26939 15385
rect 26970 15376 26976 15388
rect 27028 15376 27034 15428
rect 27798 15376 27804 15428
rect 27856 15376 27862 15428
rect 28092 15416 28120 15447
rect 29546 15444 29552 15496
rect 29604 15444 29610 15496
rect 29638 15444 29644 15496
rect 29696 15484 29702 15496
rect 32766 15484 32772 15496
rect 29696 15456 32772 15484
rect 29696 15444 29702 15456
rect 32766 15444 32772 15456
rect 32824 15444 32830 15496
rect 32950 15444 32956 15496
rect 33008 15444 33014 15496
rect 33042 15444 33048 15496
rect 33100 15444 33106 15496
rect 33318 15444 33324 15496
rect 33376 15444 33382 15496
rect 33594 15444 33600 15496
rect 33652 15444 33658 15496
rect 34057 15487 34115 15493
rect 34057 15484 34069 15487
rect 33888 15456 34069 15484
rect 32214 15416 32220 15428
rect 28092 15388 32220 15416
rect 32214 15376 32220 15388
rect 32272 15416 32278 15428
rect 32858 15416 32864 15428
rect 32272 15388 32864 15416
rect 32272 15376 32278 15388
rect 32858 15376 32864 15388
rect 32916 15376 32922 15428
rect 33778 15376 33784 15428
rect 33836 15376 33842 15428
rect 23808 15320 24164 15348
rect 23808 15308 23814 15320
rect 24210 15308 24216 15360
rect 24268 15308 24274 15360
rect 25222 15308 25228 15360
rect 25280 15308 25286 15360
rect 25682 15308 25688 15360
rect 25740 15348 25746 15360
rect 26142 15348 26148 15360
rect 25740 15320 26148 15348
rect 25740 15308 25746 15320
rect 26142 15308 26148 15320
rect 26200 15308 26206 15360
rect 27062 15308 27068 15360
rect 27120 15308 27126 15360
rect 27522 15308 27528 15360
rect 27580 15348 27586 15360
rect 30742 15348 30748 15360
rect 27580 15320 30748 15348
rect 27580 15308 27586 15320
rect 30742 15308 30748 15320
rect 30800 15308 30806 15360
rect 31202 15308 31208 15360
rect 31260 15348 31266 15360
rect 33888 15348 33916 15456
rect 34057 15453 34069 15456
rect 34103 15453 34115 15487
rect 34057 15447 34115 15453
rect 34238 15444 34244 15496
rect 34296 15444 34302 15496
rect 34716 15484 34744 15512
rect 34977 15487 35035 15493
rect 34977 15484 34989 15487
rect 34716 15456 34989 15484
rect 34977 15453 34989 15456
rect 35023 15453 35035 15487
rect 34977 15447 35035 15453
rect 35621 15487 35679 15493
rect 35621 15453 35633 15487
rect 35667 15453 35679 15487
rect 35621 15447 35679 15453
rect 35888 15487 35946 15493
rect 35888 15453 35900 15487
rect 35934 15453 35946 15487
rect 37093 15487 37151 15493
rect 37093 15484 37105 15487
rect 35888 15447 35946 15453
rect 37016 15456 37105 15484
rect 33965 15419 34023 15425
rect 33965 15385 33977 15419
rect 34011 15416 34023 15419
rect 34701 15419 34759 15425
rect 34701 15416 34713 15419
rect 34011 15388 34713 15416
rect 34011 15385 34023 15388
rect 33965 15379 34023 15385
rect 34701 15385 34713 15388
rect 34747 15385 34759 15419
rect 34701 15379 34759 15385
rect 31260 15320 33916 15348
rect 35636 15348 35664 15447
rect 35802 15376 35808 15428
rect 35860 15416 35866 15428
rect 35912 15416 35940 15447
rect 35860 15388 35940 15416
rect 35860 15376 35866 15388
rect 37016 15348 37044 15456
rect 37093 15453 37105 15456
rect 37139 15484 37151 15487
rect 37642 15484 37648 15496
rect 37139 15456 37648 15484
rect 37139 15453 37151 15456
rect 37093 15447 37151 15453
rect 37642 15444 37648 15456
rect 37700 15484 37706 15496
rect 38562 15484 38568 15496
rect 37700 15456 38568 15484
rect 37700 15444 37706 15456
rect 38562 15444 38568 15456
rect 38620 15444 38626 15496
rect 40218 15444 40224 15496
rect 40276 15484 40282 15496
rect 40865 15487 40923 15493
rect 40865 15484 40877 15487
rect 40276 15456 40877 15484
rect 40276 15444 40282 15456
rect 40865 15453 40877 15456
rect 40911 15453 40923 15487
rect 40865 15447 40923 15453
rect 41141 15487 41199 15493
rect 41141 15453 41153 15487
rect 41187 15453 41199 15487
rect 41141 15447 41199 15453
rect 37182 15376 37188 15428
rect 37240 15416 37246 15428
rect 37338 15419 37396 15425
rect 37338 15416 37350 15419
rect 37240 15388 37350 15416
rect 37240 15376 37246 15388
rect 37338 15385 37350 15388
rect 37384 15385 37396 15419
rect 41156 15416 41184 15447
rect 41230 15444 41236 15496
rect 41288 15444 41294 15496
rect 41509 15487 41567 15493
rect 41509 15453 41521 15487
rect 41555 15484 41567 15487
rect 42334 15484 42340 15496
rect 41555 15456 42340 15484
rect 41555 15453 41567 15456
rect 41509 15447 41567 15453
rect 42334 15444 42340 15456
rect 42392 15444 42398 15496
rect 44269 15487 44327 15493
rect 44269 15453 44281 15487
rect 44315 15453 44327 15487
rect 44269 15447 44327 15453
rect 37338 15379 37396 15385
rect 38396 15388 41184 15416
rect 41417 15419 41475 15425
rect 35636 15320 37044 15348
rect 31260 15308 31266 15320
rect 37090 15308 37096 15360
rect 37148 15348 37154 15360
rect 38396 15348 38424 15388
rect 41417 15385 41429 15419
rect 41463 15416 41475 15419
rect 41754 15419 41812 15425
rect 41754 15416 41766 15419
rect 41463 15388 41766 15416
rect 41463 15385 41475 15388
rect 41417 15379 41475 15385
rect 41754 15385 41766 15388
rect 41800 15385 41812 15419
rect 44284 15416 44312 15447
rect 41754 15379 41812 15385
rect 41892 15388 44312 15416
rect 37148 15320 38424 15348
rect 38473 15351 38531 15357
rect 37148 15308 37154 15320
rect 38473 15317 38485 15351
rect 38519 15348 38531 15351
rect 38654 15348 38660 15360
rect 38519 15320 38660 15348
rect 38519 15317 38531 15320
rect 38473 15311 38531 15317
rect 38654 15308 38660 15320
rect 38712 15348 38718 15360
rect 41892 15348 41920 15388
rect 38712 15320 41920 15348
rect 42889 15351 42947 15357
rect 38712 15308 38718 15320
rect 42889 15317 42901 15351
rect 42935 15348 42947 15351
rect 43070 15348 43076 15360
rect 42935 15320 43076 15348
rect 42935 15317 42947 15320
rect 42889 15311 42947 15317
rect 43070 15308 43076 15320
rect 43128 15308 43134 15360
rect 44082 15308 44088 15360
rect 44140 15348 44146 15360
rect 44453 15351 44511 15357
rect 44453 15348 44465 15351
rect 44140 15320 44465 15348
rect 44140 15308 44146 15320
rect 44453 15317 44465 15320
rect 44499 15317 44511 15351
rect 44453 15311 44511 15317
rect 1104 15258 44896 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 44896 15258
rect 1104 15184 44896 15206
rect 2590 15104 2596 15156
rect 2648 15144 2654 15156
rect 3145 15147 3203 15153
rect 3145 15144 3157 15147
rect 2648 15116 3157 15144
rect 2648 15104 2654 15116
rect 3145 15113 3157 15116
rect 3191 15113 3203 15147
rect 3145 15107 3203 15113
rect 3234 15104 3240 15156
rect 3292 15144 3298 15156
rect 8110 15144 8116 15156
rect 3292 15116 8116 15144
rect 3292 15104 3298 15116
rect 3053 15079 3111 15085
rect 3053 15045 3065 15079
rect 3099 15076 3111 15079
rect 3602 15076 3608 15088
rect 3099 15048 3608 15076
rect 3099 15045 3111 15048
rect 3053 15039 3111 15045
rect 3602 15036 3608 15048
rect 3660 15036 3666 15088
rect 6472 15085 6500 15116
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 8386 15104 8392 15156
rect 8444 15144 8450 15156
rect 8846 15144 8852 15156
rect 8444 15116 8852 15144
rect 8444 15104 8450 15116
rect 8846 15104 8852 15116
rect 8904 15104 8910 15156
rect 9033 15147 9091 15153
rect 9033 15113 9045 15147
rect 9079 15144 9091 15147
rect 10686 15144 10692 15156
rect 9079 15116 10692 15144
rect 9079 15113 9091 15116
rect 9033 15107 9091 15113
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 11054 15104 11060 15156
rect 11112 15104 11118 15156
rect 11606 15104 11612 15156
rect 11664 15144 11670 15156
rect 11974 15144 11980 15156
rect 11664 15116 11980 15144
rect 11664 15104 11670 15116
rect 11974 15104 11980 15116
rect 12032 15104 12038 15156
rect 12158 15104 12164 15156
rect 12216 15144 12222 15156
rect 12529 15147 12587 15153
rect 12216 15116 12480 15144
rect 12216 15104 12222 15116
rect 6457 15079 6515 15085
rect 6457 15045 6469 15079
rect 6503 15045 6515 15079
rect 6457 15039 6515 15045
rect 6914 15036 6920 15088
rect 6972 15076 6978 15088
rect 6972 15048 7420 15076
rect 6972 15036 6978 15048
rect 2498 14968 2504 15020
rect 2556 15008 2562 15020
rect 3329 15011 3387 15017
rect 3329 15008 3341 15011
rect 2556 14980 3341 15008
rect 2556 14968 2562 14980
rect 3329 14977 3341 14980
rect 3375 14977 3387 15011
rect 3329 14971 3387 14977
rect 3510 14968 3516 15020
rect 3568 15008 3574 15020
rect 5997 15011 6055 15017
rect 5997 15008 6009 15011
rect 3568 14980 6009 15008
rect 3568 14968 3574 14980
rect 5997 14977 6009 14980
rect 6043 14977 6055 15011
rect 5997 14971 6055 14977
rect 2593 14943 2651 14949
rect 2593 14909 2605 14943
rect 2639 14909 2651 14943
rect 2593 14903 2651 14909
rect 2608 14804 2636 14903
rect 2682 14900 2688 14952
rect 2740 14900 2746 14952
rect 2774 14900 2780 14952
rect 2832 14900 2838 14952
rect 2869 14943 2927 14949
rect 2869 14909 2881 14943
rect 2915 14940 2927 14943
rect 3528 14940 3556 14968
rect 2915 14912 3556 14940
rect 6012 14940 6040 14971
rect 7098 14968 7104 15020
rect 7156 15008 7162 15020
rect 7285 15011 7343 15017
rect 7285 15008 7297 15011
rect 7156 14980 7297 15008
rect 7156 14968 7162 14980
rect 7285 14977 7297 14980
rect 7331 14977 7343 15011
rect 7392 15008 7420 15048
rect 7742 15036 7748 15088
rect 7800 15076 7806 15088
rect 8297 15079 8355 15085
rect 8297 15076 8309 15079
rect 7800 15048 8309 15076
rect 7800 15036 7806 15048
rect 8297 15045 8309 15048
rect 8343 15045 8355 15079
rect 8297 15039 8355 15045
rect 8757 15079 8815 15085
rect 8757 15045 8769 15079
rect 8803 15076 8815 15079
rect 9214 15076 9220 15088
rect 8803 15048 9220 15076
rect 8803 15045 8815 15048
rect 8757 15039 8815 15045
rect 7926 15008 7932 15020
rect 7392 14980 7932 15008
rect 7285 14971 7343 14977
rect 7926 14968 7932 14980
rect 7984 14968 7990 15020
rect 8018 14968 8024 15020
rect 8076 15008 8082 15020
rect 8772 15008 8800 15039
rect 9214 15036 9220 15048
rect 9272 15076 9278 15088
rect 9493 15079 9551 15085
rect 9493 15076 9505 15079
rect 9272 15048 9505 15076
rect 9272 15036 9278 15048
rect 9493 15045 9505 15048
rect 9539 15045 9551 15079
rect 9493 15039 9551 15045
rect 10042 15036 10048 15088
rect 10100 15076 10106 15088
rect 12452 15076 12480 15116
rect 12529 15113 12541 15147
rect 12575 15144 12587 15147
rect 13722 15144 13728 15156
rect 12575 15116 13728 15144
rect 12575 15113 12587 15116
rect 12529 15107 12587 15113
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 15102 15144 15108 15156
rect 14844 15116 15108 15144
rect 13078 15076 13084 15088
rect 10100 15048 12388 15076
rect 12452 15048 13084 15076
rect 10100 15036 10106 15048
rect 8076 14980 8800 15008
rect 8076 14968 8082 14980
rect 8846 14968 8852 15020
rect 8904 15008 8910 15020
rect 9125 15011 9183 15017
rect 9125 15008 9137 15011
rect 8904 14980 9137 15008
rect 8904 14968 8910 14980
rect 9125 14977 9137 14980
rect 9171 15008 9183 15011
rect 9306 15008 9312 15020
rect 9171 14980 9312 15008
rect 9171 14977 9183 14980
rect 9125 14971 9183 14977
rect 9306 14968 9312 14980
rect 9364 14968 9370 15020
rect 9858 14968 9864 15020
rect 9916 15008 9922 15020
rect 10321 15011 10379 15017
rect 10321 15008 10333 15011
rect 9916 14980 10333 15008
rect 9916 14968 9922 14980
rect 10321 14977 10333 14980
rect 10367 15008 10379 15011
rect 10502 15008 10508 15020
rect 10367 14980 10508 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 10502 14968 10508 14980
rect 10560 14968 10566 15020
rect 10689 15011 10747 15017
rect 10689 14977 10701 15011
rect 10735 14977 10747 15011
rect 10689 14971 10747 14977
rect 8478 14940 8484 14952
rect 6012 14912 8484 14940
rect 2915 14909 2927 14912
rect 2869 14903 2927 14909
rect 8478 14900 8484 14912
rect 8536 14900 8542 14952
rect 9401 14943 9459 14949
rect 9401 14940 9413 14943
rect 8680 14912 9413 14940
rect 6641 14875 6699 14881
rect 6641 14841 6653 14875
rect 6687 14872 6699 14875
rect 6914 14872 6920 14884
rect 6687 14844 6920 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 6914 14832 6920 14844
rect 6972 14832 6978 14884
rect 7834 14832 7840 14884
rect 7892 14872 7898 14884
rect 8297 14875 8355 14881
rect 8297 14872 8309 14875
rect 7892 14844 8309 14872
rect 7892 14832 7898 14844
rect 8297 14841 8309 14844
rect 8343 14872 8355 14875
rect 8680 14872 8708 14912
rect 9401 14909 9413 14912
rect 9447 14909 9459 14943
rect 9401 14903 9459 14909
rect 9490 14900 9496 14952
rect 9548 14940 9554 14952
rect 9610 14943 9668 14949
rect 9610 14940 9622 14943
rect 9548 14912 9622 14940
rect 9548 14900 9554 14912
rect 9610 14909 9622 14912
rect 9656 14909 9668 14943
rect 9610 14903 9668 14909
rect 9950 14900 9956 14952
rect 10008 14940 10014 14952
rect 10413 14943 10471 14949
rect 10413 14940 10425 14943
rect 10008 14912 10425 14940
rect 10008 14900 10014 14912
rect 10413 14909 10425 14912
rect 10459 14909 10471 14943
rect 10413 14903 10471 14909
rect 10594 14900 10600 14952
rect 10652 14900 10658 14952
rect 10704 14940 10732 14971
rect 10870 14968 10876 15020
rect 10928 15008 10934 15020
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 10928 14980 11713 15008
rect 10928 14968 10934 14980
rect 11701 14977 11713 14980
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 11882 14968 11888 15020
rect 11940 14968 11946 15020
rect 11974 14968 11980 15020
rect 12032 15008 12038 15020
rect 12360 15017 12388 15048
rect 13078 15036 13084 15048
rect 13136 15036 13142 15088
rect 13998 15036 14004 15088
rect 14056 15076 14062 15088
rect 14844 15085 14872 15116
rect 15102 15104 15108 15116
rect 15160 15104 15166 15156
rect 15194 15104 15200 15156
rect 15252 15144 15258 15156
rect 18414 15144 18420 15156
rect 15252 15116 18420 15144
rect 15252 15104 15258 15116
rect 18414 15104 18420 15116
rect 18472 15104 18478 15156
rect 18690 15104 18696 15156
rect 18748 15144 18754 15156
rect 18748 15116 18920 15144
rect 18748 15104 18754 15116
rect 14829 15079 14887 15085
rect 14056 15048 14780 15076
rect 14056 15036 14062 15048
rect 12069 15011 12127 15017
rect 12069 15008 12081 15011
rect 12032 14980 12081 15008
rect 12032 14968 12038 14980
rect 12069 14977 12081 14980
rect 12115 14977 12127 15011
rect 12069 14971 12127 14977
rect 12345 15011 12403 15017
rect 12345 14977 12357 15011
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 14550 14968 14556 15020
rect 14608 15008 14614 15020
rect 14645 15011 14703 15017
rect 14645 15008 14657 15011
rect 14608 14980 14657 15008
rect 14608 14968 14614 14980
rect 14645 14977 14657 14980
rect 14691 14977 14703 15011
rect 14752 15008 14780 15048
rect 14829 15045 14841 15079
rect 14875 15045 14887 15079
rect 14829 15039 14887 15045
rect 18506 15036 18512 15088
rect 18564 15076 18570 15088
rect 18892 15085 18920 15116
rect 21174 15104 21180 15156
rect 21232 15144 21238 15156
rect 23750 15144 23756 15156
rect 21232 15116 23756 15144
rect 21232 15104 21238 15116
rect 23750 15104 23756 15116
rect 23808 15104 23814 15156
rect 23842 15104 23848 15156
rect 23900 15104 23906 15156
rect 26234 15144 26240 15156
rect 23952 15116 26240 15144
rect 18877 15079 18935 15085
rect 18564 15048 18828 15076
rect 18564 15036 18570 15048
rect 14918 15008 14924 15020
rect 14752 14980 14924 15008
rect 14645 14971 14703 14977
rect 14918 14968 14924 14980
rect 14976 14968 14982 15020
rect 15065 15011 15123 15017
rect 15065 14977 15077 15011
rect 15111 15008 15123 15011
rect 15378 15008 15384 15020
rect 15111 14980 15384 15008
rect 15111 14977 15123 14980
rect 15065 14971 15123 14977
rect 15378 14968 15384 14980
rect 15436 14968 15442 15020
rect 15838 14968 15844 15020
rect 15896 15008 15902 15020
rect 18693 15011 18751 15017
rect 15896 14980 18644 15008
rect 15896 14968 15902 14980
rect 11606 14940 11612 14952
rect 10704 14912 11612 14940
rect 11606 14900 11612 14912
rect 11664 14900 11670 14952
rect 11900 14940 11928 14968
rect 16758 14940 16764 14952
rect 11900 14912 16764 14940
rect 16758 14900 16764 14912
rect 16816 14900 16822 14952
rect 11146 14872 11152 14884
rect 8343 14844 8708 14872
rect 8956 14844 11152 14872
rect 8343 14841 8355 14844
rect 8297 14835 8355 14841
rect 3970 14804 3976 14816
rect 2608 14776 3976 14804
rect 3970 14764 3976 14776
rect 4028 14764 4034 14816
rect 6086 14764 6092 14816
rect 6144 14764 6150 14816
rect 6270 14764 6276 14816
rect 6328 14804 6334 14816
rect 7006 14804 7012 14816
rect 6328 14776 7012 14804
rect 6328 14764 6334 14776
rect 7006 14764 7012 14776
rect 7064 14804 7070 14816
rect 7190 14804 7196 14816
rect 7064 14776 7196 14804
rect 7064 14764 7070 14776
rect 7190 14764 7196 14776
rect 7248 14764 7254 14816
rect 7469 14807 7527 14813
rect 7469 14773 7481 14807
rect 7515 14804 7527 14807
rect 8956 14804 8984 14844
rect 11146 14832 11152 14844
rect 11204 14832 11210 14884
rect 11698 14832 11704 14884
rect 11756 14872 11762 14884
rect 11885 14875 11943 14881
rect 11885 14872 11897 14875
rect 11756 14844 11897 14872
rect 11756 14832 11762 14844
rect 11885 14841 11897 14844
rect 11931 14872 11943 14875
rect 11931 14844 14504 14872
rect 11931 14841 11943 14844
rect 11885 14835 11943 14841
rect 7515 14776 8984 14804
rect 7515 14773 7527 14776
rect 7469 14767 7527 14773
rect 9766 14764 9772 14816
rect 9824 14764 9830 14816
rect 10502 14764 10508 14816
rect 10560 14804 10566 14816
rect 11514 14804 11520 14816
rect 10560 14776 11520 14804
rect 10560 14764 10566 14776
rect 11514 14764 11520 14776
rect 11572 14804 11578 14816
rect 12066 14804 12072 14816
rect 11572 14776 12072 14804
rect 11572 14764 11578 14776
rect 12066 14764 12072 14776
rect 12124 14764 12130 14816
rect 14476 14804 14504 14844
rect 14826 14832 14832 14884
rect 14884 14872 14890 14884
rect 15102 14872 15108 14884
rect 14884 14844 15108 14872
rect 14884 14832 14890 14844
rect 15102 14832 15108 14844
rect 15160 14832 15166 14884
rect 15197 14875 15255 14881
rect 15197 14841 15209 14875
rect 15243 14872 15255 14875
rect 16666 14872 16672 14884
rect 15243 14844 16672 14872
rect 15243 14841 15255 14844
rect 15197 14835 15255 14841
rect 16666 14832 16672 14844
rect 16724 14832 16730 14884
rect 18616 14872 18644 14980
rect 18693 14977 18705 15011
rect 18739 14977 18751 15011
rect 18800 15008 18828 15048
rect 18877 15045 18889 15079
rect 18923 15045 18935 15079
rect 18877 15039 18935 15045
rect 18969 15079 19027 15085
rect 18969 15045 18981 15079
rect 19015 15076 19027 15079
rect 19886 15076 19892 15088
rect 19015 15048 19892 15076
rect 19015 15045 19027 15048
rect 18969 15039 19027 15045
rect 19886 15036 19892 15048
rect 19944 15036 19950 15088
rect 23952 15076 23980 15116
rect 26234 15104 26240 15116
rect 26292 15104 26298 15156
rect 26605 15147 26663 15153
rect 26605 15113 26617 15147
rect 26651 15113 26663 15147
rect 26605 15107 26663 15113
rect 22066 15048 23980 15076
rect 24044 15048 26556 15076
rect 19066 15011 19124 15017
rect 19066 15008 19078 15011
rect 18800 14980 19078 15008
rect 18693 14971 18751 14977
rect 19066 14977 19078 14980
rect 19112 14977 19124 15011
rect 19066 14971 19124 14977
rect 18708 14940 18736 14971
rect 19242 14968 19248 15020
rect 19300 15008 19306 15020
rect 22066 15008 22094 15048
rect 23014 15008 23020 15020
rect 19300 14980 22094 15008
rect 22480 14980 23020 15008
rect 19300 14968 19306 14980
rect 19518 14940 19524 14952
rect 18708 14912 19524 14940
rect 19518 14900 19524 14912
rect 19576 14900 19582 14952
rect 22480 14940 22508 14980
rect 23014 14968 23020 14980
rect 23072 15008 23078 15020
rect 23566 15008 23572 15020
rect 23072 14980 23572 15008
rect 23072 14968 23078 14980
rect 23566 14968 23572 14980
rect 23624 14968 23630 15020
rect 23658 14968 23664 15020
rect 23716 15008 23722 15020
rect 24044 15017 24072 15048
rect 24029 15011 24087 15017
rect 24029 15008 24041 15011
rect 23716 14980 24041 15008
rect 23716 14968 23722 14980
rect 24029 14977 24041 14980
rect 24075 14977 24087 15011
rect 24029 14971 24087 14977
rect 24302 14968 24308 15020
rect 24360 14968 24366 15020
rect 26142 14968 26148 15020
rect 26200 14968 26206 15020
rect 26418 14968 26424 15020
rect 26476 14968 26482 15020
rect 19628 14912 22508 14940
rect 19245 14875 19303 14881
rect 18616 14844 18828 14872
rect 15746 14804 15752 14816
rect 14476 14776 15752 14804
rect 15746 14764 15752 14776
rect 15804 14764 15810 14816
rect 18800 14804 18828 14844
rect 19245 14841 19257 14875
rect 19291 14872 19303 14875
rect 19426 14872 19432 14884
rect 19291 14844 19432 14872
rect 19291 14841 19303 14844
rect 19245 14835 19303 14841
rect 19426 14832 19432 14844
rect 19484 14832 19490 14884
rect 19628 14804 19656 14912
rect 23750 14900 23756 14952
rect 23808 14940 23814 14952
rect 24121 14943 24179 14949
rect 24121 14940 24133 14943
rect 23808 14912 24133 14940
rect 23808 14900 23814 14912
rect 24121 14909 24133 14912
rect 24167 14909 24179 14943
rect 24121 14903 24179 14909
rect 25222 14900 25228 14952
rect 25280 14940 25286 14952
rect 26237 14943 26295 14949
rect 26237 14940 26249 14943
rect 25280 14912 26249 14940
rect 25280 14900 25286 14912
rect 26237 14909 26249 14912
rect 26283 14909 26295 14943
rect 26528 14940 26556 15048
rect 26620 15008 26648 15107
rect 27338 15104 27344 15156
rect 27396 15104 27402 15156
rect 27798 15104 27804 15156
rect 27856 15144 27862 15156
rect 27893 15147 27951 15153
rect 27893 15144 27905 15147
rect 27856 15116 27905 15144
rect 27856 15104 27862 15116
rect 27893 15113 27905 15116
rect 27939 15113 27951 15147
rect 31294 15144 31300 15156
rect 27893 15107 27951 15113
rect 30668 15116 31300 15144
rect 26878 15036 26884 15088
rect 26936 15076 26942 15088
rect 29454 15076 29460 15088
rect 26936 15048 29460 15076
rect 26936 15036 26942 15048
rect 29454 15036 29460 15048
rect 29512 15036 29518 15088
rect 29546 15036 29552 15088
rect 29604 15076 29610 15088
rect 30668 15085 30696 15116
rect 31294 15104 31300 15116
rect 31352 15104 31358 15156
rect 31570 15144 31576 15156
rect 31404 15116 31576 15144
rect 30653 15079 30711 15085
rect 30653 15076 30665 15079
rect 29604 15048 30665 15076
rect 29604 15036 29610 15048
rect 30653 15045 30665 15048
rect 30699 15045 30711 15079
rect 30653 15039 30711 15045
rect 26973 15011 27031 15017
rect 26973 15008 26985 15011
rect 26620 14980 26985 15008
rect 26973 14977 26985 14980
rect 27019 14977 27031 15011
rect 26973 14971 27031 14977
rect 27525 15011 27583 15017
rect 27525 14977 27537 15011
rect 27571 15008 27583 15011
rect 27706 15008 27712 15020
rect 27571 14980 27712 15008
rect 27571 14977 27583 14980
rect 27525 14971 27583 14977
rect 27706 14968 27712 14980
rect 27764 15008 27770 15020
rect 28718 15008 28724 15020
rect 27764 14980 28724 15008
rect 27764 14968 27770 14980
rect 28718 14968 28724 14980
rect 28776 14968 28782 15020
rect 30834 14968 30840 15020
rect 30892 14968 30898 15020
rect 30929 15011 30987 15017
rect 30929 14977 30941 15011
rect 30975 15008 30987 15011
rect 31110 15008 31116 15020
rect 30975 14980 31116 15008
rect 30975 14977 30987 14980
rect 30929 14971 30987 14977
rect 31110 14968 31116 14980
rect 31168 14968 31174 15020
rect 31202 14968 31208 15020
rect 31260 14968 31266 15020
rect 31404 15008 31432 15116
rect 31570 15104 31576 15116
rect 31628 15104 31634 15156
rect 31941 15147 31999 15153
rect 31941 15113 31953 15147
rect 31987 15144 31999 15147
rect 32950 15144 32956 15156
rect 31987 15116 32956 15144
rect 31987 15113 31999 15116
rect 31941 15107 31999 15113
rect 32950 15104 32956 15116
rect 33008 15144 33014 15156
rect 33778 15144 33784 15156
rect 33008 15116 33784 15144
rect 33008 15104 33014 15116
rect 33778 15104 33784 15116
rect 33836 15104 33842 15156
rect 33965 15147 34023 15153
rect 33965 15113 33977 15147
rect 34011 15144 34023 15147
rect 36170 15144 36176 15156
rect 34011 15116 36176 15144
rect 34011 15113 34023 15116
rect 33965 15107 34023 15113
rect 36170 15104 36176 15116
rect 36228 15104 36234 15156
rect 39022 15104 39028 15156
rect 39080 15104 39086 15156
rect 41414 15104 41420 15156
rect 41472 15144 41478 15156
rect 42429 15147 42487 15153
rect 42429 15144 42441 15147
rect 41472 15116 42441 15144
rect 41472 15104 41478 15116
rect 42429 15113 42441 15116
rect 42475 15113 42487 15147
rect 42429 15107 42487 15113
rect 33502 15036 33508 15088
rect 33560 15036 33566 15088
rect 37366 15036 37372 15088
rect 37424 15076 37430 15088
rect 37890 15079 37948 15085
rect 37890 15076 37902 15079
rect 37424 15048 37902 15076
rect 37424 15036 37430 15048
rect 37890 15045 37902 15048
rect 37936 15045 37948 15079
rect 37890 15039 37948 15045
rect 31481 15011 31539 15017
rect 31481 15008 31493 15011
rect 31404 14980 31493 15008
rect 31481 14977 31493 14980
rect 31527 14977 31539 15011
rect 31481 14971 31539 14977
rect 31570 14968 31576 15020
rect 31628 15008 31634 15020
rect 31665 15011 31723 15017
rect 31665 15008 31677 15011
rect 31628 14980 31677 15008
rect 31628 14968 31634 14980
rect 31665 14977 31677 14980
rect 31711 14977 31723 15011
rect 31665 14971 31723 14977
rect 31754 14968 31760 15020
rect 31812 15008 31818 15020
rect 33134 15008 33140 15020
rect 31812 14980 33140 15008
rect 31812 14968 31818 14980
rect 33134 14968 33140 14980
rect 33192 14968 33198 15020
rect 33686 14968 33692 15020
rect 33744 14968 33750 15020
rect 33781 15011 33839 15017
rect 33781 14977 33793 15011
rect 33827 14977 33839 15011
rect 33781 14971 33839 14977
rect 27065 14943 27123 14949
rect 27065 14940 27077 14943
rect 26528 14912 27077 14940
rect 26237 14903 26295 14909
rect 27065 14909 27077 14912
rect 27111 14909 27123 14943
rect 27065 14903 27123 14909
rect 27338 14900 27344 14952
rect 27396 14940 27402 14952
rect 27617 14943 27675 14949
rect 27617 14940 27629 14943
rect 27396 14912 27629 14940
rect 27396 14900 27402 14912
rect 27617 14909 27629 14912
rect 27663 14909 27675 14943
rect 27617 14903 27675 14909
rect 27798 14900 27804 14952
rect 27856 14940 27862 14952
rect 30650 14940 30656 14952
rect 27856 14912 30656 14940
rect 27856 14900 27862 14912
rect 30650 14900 30656 14912
rect 30708 14900 30714 14952
rect 31018 14900 31024 14952
rect 31076 14900 31082 14952
rect 31386 14900 31392 14952
rect 31444 14940 31450 14952
rect 33796 14940 33824 14971
rect 37642 14968 37648 15020
rect 37700 14968 37706 15020
rect 37734 14968 37740 15020
rect 37792 14968 37798 15020
rect 37752 14940 37780 14968
rect 31444 14912 37780 14940
rect 31444 14900 31450 14912
rect 43070 14900 43076 14952
rect 43128 14900 43134 14952
rect 19978 14832 19984 14884
rect 20036 14872 20042 14884
rect 20714 14872 20720 14884
rect 20036 14844 20720 14872
rect 20036 14832 20042 14844
rect 20714 14832 20720 14844
rect 20772 14872 20778 14884
rect 21634 14872 21640 14884
rect 20772 14844 21640 14872
rect 20772 14832 20778 14844
rect 21634 14832 21640 14844
rect 21692 14832 21698 14884
rect 30469 14875 30527 14881
rect 30469 14872 30481 14875
rect 24320 14844 30481 14872
rect 18800 14776 19656 14804
rect 20806 14764 20812 14816
rect 20864 14804 20870 14816
rect 23566 14804 23572 14816
rect 20864 14776 23572 14804
rect 20864 14764 20870 14776
rect 23566 14764 23572 14776
rect 23624 14764 23630 14816
rect 23658 14764 23664 14816
rect 23716 14804 23722 14816
rect 24118 14804 24124 14816
rect 23716 14776 24124 14804
rect 23716 14764 23722 14776
rect 24118 14764 24124 14776
rect 24176 14764 24182 14816
rect 24320 14813 24348 14844
rect 30469 14841 30481 14844
rect 30515 14872 30527 14875
rect 31202 14872 31208 14884
rect 30515 14844 31208 14872
rect 30515 14841 30527 14844
rect 30469 14835 30527 14841
rect 31202 14832 31208 14844
rect 31260 14832 31266 14884
rect 31294 14832 31300 14884
rect 31352 14872 31358 14884
rect 31352 14844 33548 14872
rect 31352 14832 31358 14844
rect 24305 14807 24363 14813
rect 24305 14773 24317 14807
rect 24351 14773 24363 14807
rect 24305 14767 24363 14773
rect 26326 14764 26332 14816
rect 26384 14804 26390 14816
rect 26878 14804 26884 14816
rect 26384 14776 26884 14804
rect 26384 14764 26390 14776
rect 26878 14764 26884 14776
rect 26936 14764 26942 14816
rect 27062 14764 27068 14816
rect 27120 14764 27126 14816
rect 27709 14807 27767 14813
rect 27709 14773 27721 14807
rect 27755 14804 27767 14807
rect 27798 14804 27804 14816
rect 27755 14776 27804 14804
rect 27755 14773 27767 14776
rect 27709 14767 27767 14773
rect 27798 14764 27804 14776
rect 27856 14764 27862 14816
rect 30926 14764 30932 14816
rect 30984 14764 30990 14816
rect 31389 14807 31447 14813
rect 31389 14773 31401 14807
rect 31435 14804 31447 14807
rect 31570 14804 31576 14816
rect 31435 14776 31576 14804
rect 31435 14773 31447 14776
rect 31389 14767 31447 14773
rect 31570 14764 31576 14776
rect 31628 14764 31634 14816
rect 31757 14807 31815 14813
rect 31757 14773 31769 14807
rect 31803 14804 31815 14807
rect 31846 14804 31852 14816
rect 31803 14776 31852 14804
rect 31803 14773 31815 14776
rect 31757 14767 31815 14773
rect 31846 14764 31852 14776
rect 31904 14764 31910 14816
rect 33520 14813 33548 14844
rect 33505 14807 33563 14813
rect 33505 14773 33517 14807
rect 33551 14773 33563 14807
rect 33505 14767 33563 14773
rect 1104 14714 44896 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 44896 14714
rect 1104 14640 44896 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 2406 14600 2412 14612
rect 1627 14572 2412 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 2406 14560 2412 14572
rect 2464 14560 2470 14612
rect 6089 14603 6147 14609
rect 6089 14569 6101 14603
rect 6135 14600 6147 14603
rect 7098 14600 7104 14612
rect 6135 14572 7104 14600
rect 6135 14569 6147 14572
rect 6089 14563 6147 14569
rect 7098 14560 7104 14572
rect 7156 14560 7162 14612
rect 7834 14560 7840 14612
rect 7892 14600 7898 14612
rect 7929 14603 7987 14609
rect 7929 14600 7941 14603
rect 7892 14572 7941 14600
rect 7892 14560 7898 14572
rect 7929 14569 7941 14572
rect 7975 14600 7987 14603
rect 8573 14603 8631 14609
rect 8573 14600 8585 14603
rect 7975 14572 8585 14600
rect 7975 14569 7987 14572
rect 7929 14563 7987 14569
rect 8573 14569 8585 14572
rect 8619 14600 8631 14603
rect 8619 14572 9469 14600
rect 8619 14569 8631 14572
rect 8573 14563 8631 14569
rect 6273 14535 6331 14541
rect 6273 14532 6285 14535
rect 5644 14504 6285 14532
rect 5644 14473 5672 14504
rect 6273 14501 6285 14504
rect 6319 14532 6331 14535
rect 7650 14532 7656 14544
rect 6319 14504 7656 14532
rect 6319 14501 6331 14504
rect 6273 14495 6331 14501
rect 7650 14492 7656 14504
rect 7708 14492 7714 14544
rect 8202 14532 8208 14544
rect 7852 14504 8208 14532
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14433 5687 14467
rect 5629 14427 5687 14433
rect 5905 14467 5963 14473
rect 5905 14433 5917 14467
rect 5951 14464 5963 14467
rect 6086 14464 6092 14476
rect 5951 14436 6092 14464
rect 5951 14433 5963 14436
rect 5905 14427 5963 14433
rect 6086 14424 6092 14436
rect 6144 14464 6150 14476
rect 6733 14467 6791 14473
rect 6733 14464 6745 14467
rect 6144 14436 6745 14464
rect 6144 14424 6150 14436
rect 6733 14433 6745 14436
rect 6779 14464 6791 14467
rect 7742 14464 7748 14476
rect 6779 14436 7748 14464
rect 6779 14433 6791 14436
rect 6733 14427 6791 14433
rect 7742 14424 7748 14436
rect 7800 14424 7806 14476
rect 7852 14473 7880 14504
rect 8202 14492 8208 14504
rect 8260 14492 8266 14544
rect 8757 14535 8815 14541
rect 8757 14501 8769 14535
rect 8803 14532 8815 14535
rect 9122 14532 9128 14544
rect 8803 14504 9128 14532
rect 8803 14501 8815 14504
rect 8757 14495 8815 14501
rect 9122 14492 9128 14504
rect 9180 14492 9186 14544
rect 7837 14467 7895 14473
rect 7837 14433 7849 14467
rect 7883 14433 7895 14467
rect 7837 14427 7895 14433
rect 8018 14424 8024 14476
rect 8076 14424 8082 14476
rect 8941 14467 8999 14473
rect 8588 14436 8892 14464
rect 842 14356 848 14408
rect 900 14396 906 14408
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 900 14368 1409 14396
rect 900 14356 906 14368
rect 1397 14365 1409 14368
rect 1443 14365 1455 14399
rect 5077 14399 5135 14405
rect 5077 14396 5089 14399
rect 1397 14359 1455 14365
rect 2332 14368 5089 14396
rect 2332 14340 2360 14368
rect 5077 14365 5089 14368
rect 5123 14365 5135 14399
rect 5077 14359 5135 14365
rect 5721 14399 5779 14405
rect 5721 14365 5733 14399
rect 5767 14365 5779 14399
rect 5721 14359 5779 14365
rect 5813 14399 5871 14405
rect 5813 14365 5825 14399
rect 5859 14396 5871 14399
rect 6914 14396 6920 14408
rect 5859 14368 6920 14396
rect 5859 14365 5871 14368
rect 5813 14359 5871 14365
rect 2314 14288 2320 14340
rect 2372 14288 2378 14340
rect 3970 14288 3976 14340
rect 4028 14328 4034 14340
rect 5736 14328 5764 14359
rect 6288 14337 6316 14368
rect 6914 14356 6920 14368
rect 6972 14396 6978 14408
rect 8036 14396 8064 14424
rect 6972 14368 8064 14396
rect 6972 14356 6978 14368
rect 8386 14356 8392 14408
rect 8444 14396 8450 14408
rect 8588 14405 8616 14436
rect 8481 14399 8539 14405
rect 8481 14396 8493 14399
rect 8444 14368 8493 14396
rect 8444 14356 8450 14368
rect 8481 14365 8493 14368
rect 8527 14365 8539 14399
rect 8481 14359 8539 14365
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14365 8631 14399
rect 8754 14396 8760 14408
rect 8573 14359 8631 14365
rect 8680 14368 8760 14396
rect 4028 14300 5764 14328
rect 4028 14288 4034 14300
rect 2225 14263 2283 14269
rect 2225 14229 2237 14263
rect 2271 14260 2283 14263
rect 2774 14260 2780 14272
rect 2271 14232 2780 14260
rect 2271 14229 2283 14232
rect 2225 14223 2283 14229
rect 2774 14220 2780 14232
rect 2832 14220 2838 14272
rect 4798 14220 4804 14272
rect 4856 14260 4862 14272
rect 5261 14263 5319 14269
rect 5261 14260 5273 14263
rect 4856 14232 5273 14260
rect 4856 14220 4862 14232
rect 5261 14229 5273 14232
rect 5307 14229 5319 14263
rect 5736 14260 5764 14300
rect 6273 14331 6331 14337
rect 6273 14297 6285 14331
rect 6319 14297 6331 14331
rect 6273 14291 6331 14297
rect 7742 14288 7748 14340
rect 7800 14328 7806 14340
rect 8205 14331 8263 14337
rect 8205 14328 8217 14331
rect 7800 14300 8217 14328
rect 7800 14288 7806 14300
rect 8205 14297 8217 14300
rect 8251 14297 8263 14331
rect 8205 14291 8263 14297
rect 8297 14331 8355 14337
rect 8297 14297 8309 14331
rect 8343 14328 8355 14331
rect 8680 14328 8708 14368
rect 8754 14356 8760 14368
rect 8812 14356 8818 14408
rect 8864 14396 8892 14436
rect 8941 14433 8953 14467
rect 8987 14464 8999 14467
rect 9214 14464 9220 14476
rect 8987 14436 9220 14464
rect 8987 14433 8999 14436
rect 8941 14427 8999 14433
rect 9214 14424 9220 14436
rect 9272 14424 9278 14476
rect 9441 14473 9469 14572
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 12618 14600 12624 14612
rect 9824 14572 12624 14600
rect 9824 14560 9830 14572
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 16574 14560 16580 14612
rect 16632 14600 16638 14612
rect 16632 14572 19932 14600
rect 16632 14560 16638 14572
rect 9582 14492 9588 14544
rect 9640 14532 9646 14544
rect 16485 14535 16543 14541
rect 9640 14504 15608 14532
rect 9640 14492 9646 14504
rect 9426 14467 9484 14473
rect 9426 14433 9438 14467
rect 9472 14433 9484 14467
rect 9426 14427 9484 14433
rect 11698 14424 11704 14476
rect 11756 14464 11762 14476
rect 13354 14464 13360 14476
rect 11756 14436 13360 14464
rect 11756 14424 11762 14436
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 13906 14424 13912 14476
rect 13964 14464 13970 14476
rect 14645 14467 14703 14473
rect 13964 14436 14320 14464
rect 13964 14424 13970 14436
rect 9306 14396 9312 14408
rect 8864 14368 9312 14396
rect 9306 14356 9312 14368
rect 9364 14356 9370 14408
rect 9674 14356 9680 14408
rect 9732 14356 9738 14408
rect 14093 14399 14151 14405
rect 14093 14365 14105 14399
rect 14139 14396 14151 14399
rect 14182 14396 14188 14408
rect 14139 14368 14188 14396
rect 14139 14365 14151 14368
rect 14093 14359 14151 14365
rect 14182 14356 14188 14368
rect 14240 14356 14246 14408
rect 14292 14405 14320 14436
rect 14645 14433 14657 14467
rect 14691 14464 14703 14467
rect 15010 14464 15016 14476
rect 14691 14436 15016 14464
rect 14691 14433 14703 14436
rect 14645 14427 14703 14433
rect 15010 14424 15016 14436
rect 15068 14424 15074 14476
rect 15580 14405 15608 14504
rect 16485 14501 16497 14535
rect 16531 14532 16543 14535
rect 16666 14532 16672 14544
rect 16531 14504 16672 14532
rect 16531 14501 16543 14504
rect 16485 14495 16543 14501
rect 16666 14492 16672 14504
rect 16724 14492 16730 14544
rect 18598 14492 18604 14544
rect 18656 14532 18662 14544
rect 19242 14532 19248 14544
rect 18656 14504 19248 14532
rect 18656 14492 18662 14504
rect 19242 14492 19248 14504
rect 19300 14492 19306 14544
rect 19904 14541 19932 14572
rect 19978 14560 19984 14612
rect 20036 14600 20042 14612
rect 20073 14603 20131 14609
rect 20073 14600 20085 14603
rect 20036 14572 20085 14600
rect 20036 14560 20042 14572
rect 20073 14569 20085 14572
rect 20119 14569 20131 14603
rect 21821 14603 21879 14609
rect 21821 14600 21833 14603
rect 20073 14563 20131 14569
rect 20180 14572 21833 14600
rect 19889 14535 19947 14541
rect 19889 14501 19901 14535
rect 19935 14532 19947 14535
rect 20180 14532 20208 14572
rect 21821 14569 21833 14572
rect 21867 14600 21879 14603
rect 22741 14603 22799 14609
rect 21867 14572 22416 14600
rect 21867 14569 21879 14572
rect 21821 14563 21879 14569
rect 19935 14504 20208 14532
rect 19935 14501 19947 14504
rect 19889 14495 19947 14501
rect 20254 14492 20260 14544
rect 20312 14532 20318 14544
rect 22094 14532 22100 14544
rect 20312 14504 22100 14532
rect 20312 14492 20318 14504
rect 22094 14492 22100 14504
rect 22152 14492 22158 14544
rect 15746 14424 15752 14476
rect 15804 14464 15810 14476
rect 15804 14436 16349 14464
rect 15804 14424 15810 14436
rect 14277 14399 14335 14405
rect 14277 14365 14289 14399
rect 14323 14365 14335 14399
rect 14277 14359 14335 14365
rect 15565 14399 15623 14405
rect 15565 14365 15577 14399
rect 15611 14365 15623 14399
rect 15565 14359 15623 14365
rect 15933 14399 15991 14405
rect 15933 14365 15945 14399
rect 15979 14396 15991 14399
rect 16022 14396 16028 14408
rect 15979 14368 16028 14396
rect 15979 14365 15991 14368
rect 15933 14359 15991 14365
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 16114 14356 16120 14408
rect 16172 14356 16178 14408
rect 16321 14405 16349 14436
rect 20346 14424 20352 14476
rect 20404 14424 20410 14476
rect 16306 14399 16364 14405
rect 16306 14365 16318 14399
rect 16352 14365 16364 14399
rect 16306 14359 16364 14365
rect 16758 14356 16764 14408
rect 16816 14396 16822 14408
rect 19610 14396 19616 14408
rect 16816 14368 19616 14396
rect 16816 14356 16822 14368
rect 19610 14356 19616 14368
rect 19668 14356 19674 14408
rect 19794 14356 19800 14408
rect 19852 14396 19858 14408
rect 20070 14396 20076 14408
rect 19852 14368 20076 14396
rect 19852 14356 19858 14368
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 20162 14356 20168 14408
rect 20220 14396 20226 14408
rect 20364 14396 20392 14424
rect 20220 14368 20392 14396
rect 20220 14356 20226 14368
rect 20530 14356 20536 14408
rect 20588 14396 20594 14408
rect 21361 14399 21419 14405
rect 21361 14396 21373 14399
rect 20588 14368 21373 14396
rect 20588 14356 20594 14368
rect 21361 14365 21373 14368
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 21726 14356 21732 14408
rect 21784 14356 21790 14408
rect 21821 14399 21879 14405
rect 21821 14365 21833 14399
rect 21867 14365 21879 14399
rect 21821 14359 21879 14365
rect 9217 14331 9275 14337
rect 9217 14328 9229 14331
rect 8343 14300 8708 14328
rect 8772 14300 9229 14328
rect 8343 14297 8355 14300
rect 8297 14291 8355 14297
rect 6730 14260 6736 14272
rect 5736 14232 6736 14260
rect 5261 14223 5319 14229
rect 6730 14220 6736 14232
rect 6788 14260 6794 14272
rect 6825 14263 6883 14269
rect 6825 14260 6837 14263
rect 6788 14232 6837 14260
rect 6788 14220 6794 14232
rect 6825 14229 6837 14232
rect 6871 14229 6883 14263
rect 6825 14223 6883 14229
rect 7006 14220 7012 14272
rect 7064 14260 7070 14272
rect 7466 14260 7472 14272
rect 7064 14232 7472 14260
rect 7064 14220 7070 14232
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 7926 14220 7932 14272
rect 7984 14260 7990 14272
rect 8113 14263 8171 14269
rect 8113 14260 8125 14263
rect 7984 14232 8125 14260
rect 7984 14220 7990 14232
rect 8113 14229 8125 14232
rect 8159 14229 8171 14263
rect 8220 14260 8248 14291
rect 8772 14260 8800 14300
rect 9217 14297 9229 14300
rect 9263 14328 9275 14331
rect 9490 14328 9496 14340
rect 9263 14300 9496 14328
rect 9263 14297 9275 14300
rect 9217 14291 9275 14297
rect 9490 14288 9496 14300
rect 9548 14288 9554 14340
rect 15197 14331 15255 14337
rect 15197 14328 15209 14331
rect 12544 14300 15209 14328
rect 8220 14232 8800 14260
rect 9861 14263 9919 14269
rect 8113 14223 8171 14229
rect 9861 14229 9873 14263
rect 9907 14260 9919 14263
rect 12544 14260 12572 14300
rect 15197 14297 15209 14300
rect 15243 14297 15255 14331
rect 16209 14331 16267 14337
rect 16209 14328 16221 14331
rect 15197 14291 15255 14297
rect 15672 14300 16221 14328
rect 15672 14272 15700 14300
rect 16209 14297 16221 14300
rect 16255 14297 16267 14331
rect 16209 14291 16267 14297
rect 16850 14288 16856 14340
rect 16908 14328 16914 14340
rect 16908 14300 20300 14328
rect 16908 14288 16914 14300
rect 9907 14232 12572 14260
rect 14553 14263 14611 14269
rect 9907 14229 9919 14232
rect 9861 14223 9919 14229
rect 14553 14229 14565 14263
rect 14599 14260 14611 14263
rect 14826 14260 14832 14272
rect 14599 14232 14832 14260
rect 14599 14229 14611 14232
rect 14553 14223 14611 14229
rect 14826 14220 14832 14232
rect 14884 14220 14890 14272
rect 15102 14220 15108 14272
rect 15160 14260 15166 14272
rect 15289 14263 15347 14269
rect 15289 14260 15301 14263
rect 15160 14232 15301 14260
rect 15160 14220 15166 14232
rect 15289 14229 15301 14232
rect 15335 14229 15347 14263
rect 15289 14223 15347 14229
rect 15654 14220 15660 14272
rect 15712 14220 15718 14272
rect 17034 14220 17040 14272
rect 17092 14260 17098 14272
rect 19242 14260 19248 14272
rect 17092 14232 19248 14260
rect 17092 14220 17098 14232
rect 19242 14220 19248 14232
rect 19300 14220 19306 14272
rect 20272 14260 20300 14300
rect 20346 14288 20352 14340
rect 20404 14288 20410 14340
rect 21836 14260 21864 14359
rect 21910 14260 21916 14272
rect 20272 14232 21916 14260
rect 21910 14220 21916 14232
rect 21968 14220 21974 14272
rect 22002 14220 22008 14272
rect 22060 14220 22066 14272
rect 22388 14260 22416 14572
rect 22741 14569 22753 14603
rect 22787 14569 22799 14603
rect 22741 14563 22799 14569
rect 22554 14424 22560 14476
rect 22612 14424 22618 14476
rect 22756 14464 22784 14563
rect 22922 14560 22928 14612
rect 22980 14560 22986 14612
rect 23566 14560 23572 14612
rect 23624 14560 23630 14612
rect 24029 14603 24087 14609
rect 24029 14569 24041 14603
rect 24075 14600 24087 14603
rect 24302 14600 24308 14612
rect 24075 14572 24308 14600
rect 24075 14569 24087 14572
rect 24029 14563 24087 14569
rect 24302 14560 24308 14572
rect 24360 14560 24366 14612
rect 30926 14600 30932 14612
rect 28184 14572 30932 14600
rect 25590 14492 25596 14544
rect 25648 14532 25654 14544
rect 28184 14532 28212 14572
rect 30926 14560 30932 14572
rect 30984 14560 30990 14612
rect 31110 14560 31116 14612
rect 31168 14560 31174 14612
rect 31754 14532 31760 14544
rect 25648 14504 28212 14532
rect 30760 14504 31760 14532
rect 25648 14492 25654 14504
rect 23753 14467 23811 14473
rect 22756 14436 23704 14464
rect 22741 14399 22799 14405
rect 22741 14365 22753 14399
rect 22787 14396 22799 14399
rect 23014 14396 23020 14408
rect 22787 14368 23020 14396
rect 22787 14365 22799 14368
rect 22741 14359 22799 14365
rect 23014 14356 23020 14368
rect 23072 14396 23078 14408
rect 23569 14399 23627 14405
rect 23569 14396 23581 14399
rect 23072 14368 23581 14396
rect 23072 14356 23078 14368
rect 23569 14365 23581 14368
rect 23615 14365 23627 14399
rect 23569 14359 23627 14365
rect 22462 14288 22468 14340
rect 22520 14288 22526 14340
rect 23676 14328 23704 14436
rect 23753 14433 23765 14467
rect 23799 14464 23811 14467
rect 24026 14464 24032 14476
rect 23799 14436 24032 14464
rect 23799 14433 23811 14436
rect 23753 14427 23811 14433
rect 24026 14424 24032 14436
rect 24084 14424 24090 14476
rect 24118 14424 24124 14476
rect 24176 14464 24182 14476
rect 27338 14464 27344 14476
rect 24176 14436 27344 14464
rect 24176 14424 24182 14436
rect 27338 14424 27344 14436
rect 27396 14464 27402 14476
rect 30760 14464 30788 14504
rect 31754 14492 31760 14504
rect 31812 14492 31818 14544
rect 27396 14436 30788 14464
rect 27396 14424 27402 14436
rect 31570 14424 31576 14476
rect 31628 14464 31634 14476
rect 33686 14464 33692 14476
rect 31628 14436 33692 14464
rect 31628 14424 31634 14436
rect 33686 14424 33692 14436
rect 33744 14424 33750 14476
rect 23845 14399 23903 14405
rect 23845 14365 23857 14399
rect 23891 14396 23903 14399
rect 24670 14396 24676 14408
rect 23891 14368 24676 14396
rect 23891 14365 23903 14368
rect 23845 14359 23903 14365
rect 24670 14356 24676 14368
rect 24728 14356 24734 14408
rect 26418 14356 26424 14408
rect 26476 14396 26482 14408
rect 27430 14396 27436 14408
rect 26476 14368 27436 14396
rect 26476 14356 26482 14368
rect 27430 14356 27436 14368
rect 27488 14396 27494 14408
rect 30745 14399 30803 14405
rect 30745 14396 30757 14399
rect 27488 14368 30757 14396
rect 27488 14356 27494 14368
rect 30745 14365 30757 14368
rect 30791 14365 30803 14399
rect 30745 14359 30803 14365
rect 30834 14356 30840 14408
rect 30892 14356 30898 14408
rect 44266 14356 44272 14408
rect 44324 14356 44330 14408
rect 28810 14328 28816 14340
rect 23676 14300 28816 14328
rect 28810 14288 28816 14300
rect 28868 14288 28874 14340
rect 30282 14288 30288 14340
rect 30340 14328 30346 14340
rect 31846 14328 31852 14340
rect 30340 14300 31852 14328
rect 30340 14288 30346 14300
rect 31846 14288 31852 14300
rect 31904 14288 31910 14340
rect 30466 14260 30472 14272
rect 22388 14232 30472 14260
rect 30466 14220 30472 14232
rect 30524 14220 30530 14272
rect 44450 14220 44456 14272
rect 44508 14220 44514 14272
rect 1104 14170 44896 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 44896 14170
rect 1104 14096 44896 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 2314 14056 2320 14068
rect 1627 14028 2320 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 2314 14016 2320 14028
rect 2372 14016 2378 14068
rect 2498 14016 2504 14068
rect 2556 14016 2562 14068
rect 2774 14016 2780 14068
rect 2832 14056 2838 14068
rect 3237 14059 3295 14065
rect 2832 14028 3096 14056
rect 2832 14016 2838 14028
rect 2682 13948 2688 14000
rect 2740 13988 2746 14000
rect 3068 13997 3096 14028
rect 3237 14025 3249 14059
rect 3283 14056 3295 14059
rect 4614 14056 4620 14068
rect 3283 14028 4620 14056
rect 3283 14025 3295 14028
rect 3237 14019 3295 14025
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 4798 14016 4804 14068
rect 4856 14056 4862 14068
rect 5718 14056 5724 14068
rect 4856 14028 5724 14056
rect 4856 14016 4862 14028
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 5810 14016 5816 14068
rect 5868 14056 5874 14068
rect 5905 14059 5963 14065
rect 5905 14056 5917 14059
rect 5868 14028 5917 14056
rect 5868 14016 5874 14028
rect 5905 14025 5917 14028
rect 5951 14056 5963 14059
rect 10870 14056 10876 14068
rect 5951 14028 10876 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 10870 14016 10876 14028
rect 10928 14016 10934 14068
rect 11974 14056 11980 14068
rect 11532 14028 11980 14056
rect 2961 13991 3019 13997
rect 2961 13988 2973 13991
rect 2740 13960 2973 13988
rect 2740 13948 2746 13960
rect 2961 13957 2973 13960
rect 3007 13957 3019 13991
rect 3068 13991 3136 13997
rect 3068 13960 3090 13991
rect 2961 13951 3019 13957
rect 3078 13957 3090 13960
rect 3124 13957 3136 13991
rect 5169 13991 5227 13997
rect 5169 13988 5181 13991
rect 3078 13951 3136 13957
rect 4356 13960 5181 13988
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 2317 13923 2375 13929
rect 2317 13920 2329 13923
rect 1719 13892 2329 13920
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 2317 13889 2329 13892
rect 2363 13920 2375 13923
rect 3234 13920 3240 13932
rect 2363 13892 3240 13920
rect 2363 13889 2375 13892
rect 2317 13883 2375 13889
rect 3234 13880 3240 13892
rect 3292 13880 3298 13932
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13889 4215 13923
rect 4157 13883 4215 13889
rect 1857 13855 1915 13861
rect 1857 13821 1869 13855
rect 1903 13821 1915 13855
rect 1857 13815 1915 13821
rect 1949 13855 2007 13861
rect 1949 13821 1961 13855
rect 1995 13821 2007 13855
rect 1949 13815 2007 13821
rect 1578 13676 1584 13728
rect 1636 13716 1642 13728
rect 1872 13716 1900 13815
rect 1964 13784 1992 13815
rect 2038 13812 2044 13864
rect 2096 13812 2102 13864
rect 2130 13812 2136 13864
rect 2188 13852 2194 13864
rect 2593 13855 2651 13861
rect 2593 13852 2605 13855
rect 2188 13824 2605 13852
rect 2188 13812 2194 13824
rect 2593 13821 2605 13824
rect 2639 13821 2651 13855
rect 2593 13815 2651 13821
rect 2869 13855 2927 13861
rect 2869 13821 2881 13855
rect 2915 13821 2927 13855
rect 2869 13815 2927 13821
rect 2774 13784 2780 13796
rect 1964 13756 2780 13784
rect 2774 13744 2780 13756
rect 2832 13744 2838 13796
rect 2884 13716 2912 13815
rect 2958 13812 2964 13864
rect 3016 13852 3022 13864
rect 4172 13852 4200 13883
rect 3016 13824 4200 13852
rect 4356 13852 4384 13960
rect 5169 13957 5181 13960
rect 5215 13988 5227 13991
rect 5258 13988 5264 14000
rect 5215 13960 5264 13988
rect 5215 13957 5227 13960
rect 5169 13951 5227 13957
rect 5258 13948 5264 13960
rect 5316 13948 5322 14000
rect 7834 13948 7840 14000
rect 7892 13988 7898 14000
rect 11532 13988 11560 14028
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 12066 14016 12072 14068
rect 12124 14065 12130 14068
rect 12124 14056 12135 14065
rect 15565 14059 15623 14065
rect 12124 14028 12169 14056
rect 12124 14019 12135 14028
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 15838 14056 15844 14068
rect 15611 14028 15844 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 12124 14016 12130 14019
rect 15838 14016 15844 14028
rect 15896 14016 15902 14068
rect 16301 14059 16359 14065
rect 16301 14025 16313 14059
rect 16347 14056 16359 14059
rect 16850 14056 16856 14068
rect 16347 14028 16856 14056
rect 16347 14025 16359 14028
rect 16301 14019 16359 14025
rect 16850 14016 16856 14028
rect 16908 14016 16914 14068
rect 17126 14016 17132 14068
rect 17184 14056 17190 14068
rect 23017 14059 23075 14065
rect 17184 14028 18920 14056
rect 17184 14016 17190 14028
rect 12710 13988 12716 14000
rect 7892 13960 9076 13988
rect 7892 13948 7898 13960
rect 4433 13923 4491 13929
rect 4433 13889 4445 13923
rect 4479 13920 4491 13923
rect 5902 13920 5908 13932
rect 4479 13892 5908 13920
rect 4479 13889 4491 13892
rect 4433 13883 4491 13889
rect 5902 13880 5908 13892
rect 5960 13880 5966 13932
rect 8202 13880 8208 13932
rect 8260 13880 8266 13932
rect 8297 13923 8355 13929
rect 8297 13889 8309 13923
rect 8343 13889 8355 13923
rect 8297 13883 8355 13889
rect 4617 13855 4675 13861
rect 4617 13852 4629 13855
rect 4356 13824 4629 13852
rect 3016 13812 3022 13824
rect 4617 13821 4629 13824
rect 4663 13821 4675 13855
rect 4617 13815 4675 13821
rect 4709 13855 4767 13861
rect 4709 13821 4721 13855
rect 4755 13821 4767 13855
rect 4709 13815 4767 13821
rect 4341 13787 4399 13793
rect 4341 13753 4353 13787
rect 4387 13784 4399 13787
rect 4724 13784 4752 13815
rect 4798 13812 4804 13864
rect 4856 13812 4862 13864
rect 4890 13812 4896 13864
rect 4948 13852 4954 13864
rect 5442 13852 5448 13864
rect 4948 13824 5448 13852
rect 4948 13812 4954 13824
rect 5442 13812 5448 13824
rect 5500 13852 5506 13864
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5500 13824 5641 13852
rect 5500 13812 5506 13824
rect 5629 13821 5641 13824
rect 5675 13852 5687 13855
rect 5810 13852 5816 13864
rect 5675 13824 5816 13852
rect 5675 13821 5687 13824
rect 5629 13815 5687 13821
rect 5810 13812 5816 13824
rect 5868 13812 5874 13864
rect 6086 13812 6092 13864
rect 6144 13852 6150 13864
rect 6144 13824 8064 13852
rect 6144 13812 6150 13824
rect 5169 13787 5227 13793
rect 5169 13784 5181 13787
rect 4387 13756 5181 13784
rect 4387 13753 4399 13756
rect 4341 13747 4399 13753
rect 4632 13728 4660 13756
rect 5169 13753 5181 13756
rect 5215 13784 5227 13787
rect 5350 13784 5356 13796
rect 5215 13756 5356 13784
rect 5215 13753 5227 13756
rect 5169 13747 5227 13753
rect 5350 13744 5356 13756
rect 5408 13784 5414 13796
rect 6638 13784 6644 13796
rect 5408 13756 6644 13784
rect 5408 13744 5414 13756
rect 6638 13744 6644 13756
rect 6696 13744 6702 13796
rect 8036 13784 8064 13824
rect 8110 13812 8116 13864
rect 8168 13852 8174 13864
rect 8312 13852 8340 13883
rect 8570 13880 8576 13932
rect 8628 13880 8634 13932
rect 9048 13929 9076 13960
rect 9140 13960 11560 13988
rect 11716 13960 12716 13988
rect 9033 13923 9091 13929
rect 8680 13892 8892 13920
rect 8680 13852 8708 13892
rect 8168 13824 8340 13852
rect 8404 13824 8708 13852
rect 8168 13812 8174 13824
rect 8404 13784 8432 13824
rect 8754 13812 8760 13864
rect 8812 13812 8818 13864
rect 8864 13852 8892 13892
rect 9033 13889 9045 13923
rect 9079 13889 9091 13923
rect 9033 13883 9091 13889
rect 9140 13852 9168 13960
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13920 9459 13923
rect 9582 13920 9588 13932
rect 9447 13892 9588 13920
rect 9447 13889 9459 13892
rect 9401 13883 9459 13889
rect 9582 13880 9588 13892
rect 9640 13880 9646 13932
rect 10410 13880 10416 13932
rect 10468 13880 10474 13932
rect 11716 13929 11744 13960
rect 12710 13948 12716 13960
rect 12768 13948 12774 14000
rect 14660 13960 15148 13988
rect 11974 13929 11980 13932
rect 11149 13923 11207 13929
rect 11149 13920 11161 13923
rect 10520 13892 11161 13920
rect 8864 13824 9168 13852
rect 9214 13812 9220 13864
rect 9272 13852 9278 13864
rect 10520 13852 10548 13892
rect 11149 13889 11161 13892
rect 11195 13889 11207 13923
rect 11149 13883 11207 13889
rect 11517 13923 11575 13929
rect 11517 13889 11529 13923
rect 11563 13889 11575 13923
rect 11517 13883 11575 13889
rect 11701 13923 11759 13929
rect 11701 13889 11713 13923
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 11793 13923 11851 13929
rect 11793 13889 11805 13923
rect 11839 13889 11851 13923
rect 11793 13883 11851 13889
rect 11937 13923 11980 13929
rect 11937 13889 11949 13923
rect 12032 13920 12038 13932
rect 12894 13920 12900 13932
rect 12032 13892 12900 13920
rect 11937 13883 11980 13889
rect 9272 13824 10548 13852
rect 9272 13812 9278 13824
rect 10962 13812 10968 13864
rect 11020 13852 11026 13864
rect 11532 13852 11560 13883
rect 11020 13824 11560 13852
rect 11808 13852 11836 13883
rect 11974 13880 11980 13883
rect 12032 13880 12038 13892
rect 12894 13880 12900 13892
rect 12952 13880 12958 13932
rect 14550 13880 14556 13932
rect 14608 13880 14614 13932
rect 14660 13929 14688 13960
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13889 14703 13923
rect 14645 13883 14703 13889
rect 14918 13880 14924 13932
rect 14976 13920 14982 13932
rect 15013 13923 15071 13929
rect 15013 13920 15025 13923
rect 14976 13892 15025 13920
rect 14976 13880 14982 13892
rect 15013 13889 15025 13892
rect 15059 13889 15071 13923
rect 15120 13920 15148 13960
rect 15194 13948 15200 14000
rect 15252 13988 15258 14000
rect 17037 13991 17095 13997
rect 17037 13988 17049 13991
rect 15252 13960 17049 13988
rect 15252 13948 15258 13960
rect 17037 13957 17049 13960
rect 17083 13957 17095 13991
rect 17037 13951 17095 13957
rect 17144 13960 18736 13988
rect 15654 13920 15660 13932
rect 15120 13892 15660 13920
rect 15013 13883 15071 13889
rect 15654 13880 15660 13892
rect 15712 13880 15718 13932
rect 15749 13923 15807 13929
rect 15749 13889 15761 13923
rect 15795 13889 15807 13923
rect 15749 13883 15807 13889
rect 12158 13852 12164 13864
rect 11808 13824 12164 13852
rect 11020 13812 11026 13824
rect 8036 13756 8432 13784
rect 8570 13744 8576 13796
rect 8628 13744 8634 13796
rect 11532 13784 11560 13824
rect 12158 13812 12164 13824
rect 12216 13812 12222 13864
rect 15102 13812 15108 13864
rect 15160 13812 15166 13864
rect 15764 13852 15792 13883
rect 15930 13880 15936 13932
rect 15988 13880 15994 13932
rect 16022 13880 16028 13932
rect 16080 13880 16086 13932
rect 16117 13923 16175 13929
rect 16117 13889 16129 13923
rect 16163 13920 16175 13923
rect 16206 13920 16212 13932
rect 16163 13892 16212 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 16206 13880 16212 13892
rect 16264 13880 16270 13932
rect 17144 13852 17172 13960
rect 18708 13932 18736 13960
rect 17402 13880 17408 13932
rect 17460 13880 17466 13932
rect 17586 13880 17592 13932
rect 17644 13880 17650 13932
rect 17678 13880 17684 13932
rect 17736 13880 17742 13932
rect 17773 13923 17831 13929
rect 17773 13889 17785 13923
rect 17819 13920 17831 13923
rect 17954 13920 17960 13932
rect 17819 13892 17960 13920
rect 17819 13889 17831 13892
rect 17773 13883 17831 13889
rect 17954 13880 17960 13892
rect 18012 13880 18018 13932
rect 18690 13880 18696 13932
rect 18748 13880 18754 13932
rect 18892 13929 18920 14028
rect 21100 14028 22876 14056
rect 19610 13948 19616 14000
rect 19668 13988 19674 14000
rect 21100 13997 21128 14028
rect 22848 14000 22876 14028
rect 23017 14025 23029 14059
rect 23063 14056 23075 14059
rect 23106 14056 23112 14068
rect 23063 14028 23112 14056
rect 23063 14025 23075 14028
rect 23017 14019 23075 14025
rect 23106 14016 23112 14028
rect 23164 14016 23170 14068
rect 28074 14016 28080 14068
rect 28132 14016 28138 14068
rect 28353 14059 28411 14065
rect 28353 14025 28365 14059
rect 28399 14025 28411 14059
rect 28353 14019 28411 14025
rect 21085 13991 21143 13997
rect 21085 13988 21097 13991
rect 19668 13960 21097 13988
rect 19668 13948 19674 13960
rect 21085 13957 21097 13960
rect 21131 13957 21143 13991
rect 21085 13951 21143 13957
rect 22002 13948 22008 14000
rect 22060 13948 22066 14000
rect 22186 13948 22192 14000
rect 22244 13948 22250 14000
rect 22388 13960 22784 13988
rect 19150 13929 19156 13932
rect 18877 13923 18935 13929
rect 18877 13889 18889 13923
rect 18923 13889 18935 13923
rect 18877 13883 18935 13889
rect 18969 13923 19027 13929
rect 18969 13889 18981 13923
rect 19015 13889 19027 13923
rect 18969 13883 19027 13889
rect 19113 13923 19156 13929
rect 19113 13889 19125 13923
rect 19113 13883 19156 13889
rect 15764 13824 17172 13852
rect 17420 13852 17448 13880
rect 17862 13852 17868 13864
rect 17420 13824 17868 13852
rect 12342 13784 12348 13796
rect 11532 13756 12348 13784
rect 12342 13744 12348 13756
rect 12400 13744 12406 13796
rect 13814 13744 13820 13796
rect 13872 13784 13878 13796
rect 14182 13784 14188 13796
rect 13872 13756 14188 13784
rect 13872 13744 13878 13756
rect 14182 13744 14188 13756
rect 14240 13784 14246 13796
rect 15764 13784 15792 13824
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 18598 13852 18604 13864
rect 17972 13824 18604 13852
rect 14240 13756 15792 13784
rect 14240 13744 14246 13756
rect 16942 13744 16948 13796
rect 17000 13784 17006 13796
rect 17972 13793 18000 13824
rect 18598 13812 18604 13824
rect 18656 13812 18662 13864
rect 18782 13812 18788 13864
rect 18840 13852 18846 13864
rect 18984 13852 19012 13883
rect 19150 13880 19156 13883
rect 19208 13880 19214 13932
rect 19262 13923 19320 13929
rect 19262 13889 19274 13923
rect 19308 13920 19320 13923
rect 19702 13920 19708 13932
rect 19308 13892 19708 13920
rect 19308 13889 19320 13892
rect 19262 13883 19320 13889
rect 19702 13880 19708 13892
rect 19760 13920 19766 13932
rect 20901 13923 20959 13929
rect 20901 13920 20913 13923
rect 19760 13892 20913 13920
rect 19760 13880 19766 13892
rect 20901 13889 20913 13892
rect 20947 13920 20959 13923
rect 21821 13923 21879 13929
rect 21821 13920 21833 13923
rect 20947 13892 21833 13920
rect 20947 13889 20959 13892
rect 20901 13883 20959 13889
rect 21821 13889 21833 13892
rect 21867 13920 21879 13923
rect 22388 13920 22416 13960
rect 21867 13892 22416 13920
rect 21867 13889 21879 13892
rect 21821 13883 21879 13889
rect 22462 13880 22468 13932
rect 22520 13920 22526 13932
rect 22649 13923 22707 13929
rect 22649 13920 22661 13923
rect 22520 13892 22661 13920
rect 22520 13880 22526 13892
rect 22649 13889 22661 13892
rect 22695 13889 22707 13923
rect 22756 13920 22784 13960
rect 22830 13948 22836 14000
rect 22888 13948 22894 14000
rect 26142 13948 26148 14000
rect 26200 13988 26206 14000
rect 27617 13991 27675 13997
rect 27617 13988 27629 13991
rect 26200 13960 27629 13988
rect 26200 13948 26206 13960
rect 27617 13957 27629 13960
rect 27663 13957 27675 13991
rect 27617 13951 27675 13957
rect 27724 13960 28212 13988
rect 25590 13920 25596 13932
rect 22756 13892 25596 13920
rect 22649 13883 22707 13889
rect 25590 13880 25596 13892
rect 25648 13880 25654 13932
rect 25866 13880 25872 13932
rect 25924 13880 25930 13932
rect 26053 13923 26111 13929
rect 26053 13889 26065 13923
rect 26099 13920 26111 13923
rect 26234 13920 26240 13932
rect 26099 13892 26240 13920
rect 26099 13889 26111 13892
rect 26053 13883 26111 13889
rect 26234 13880 26240 13892
rect 26292 13880 26298 13932
rect 26421 13923 26479 13929
rect 26421 13889 26433 13923
rect 26467 13920 26479 13923
rect 26510 13920 26516 13932
rect 26467 13892 26516 13920
rect 26467 13889 26479 13892
rect 26421 13883 26479 13889
rect 26510 13880 26516 13892
rect 26568 13880 26574 13932
rect 26602 13880 26608 13932
rect 26660 13880 26666 13932
rect 26786 13880 26792 13932
rect 26844 13880 26850 13932
rect 26973 13923 27031 13929
rect 26973 13889 26985 13923
rect 27019 13889 27031 13923
rect 26973 13883 27031 13889
rect 18840 13824 19012 13852
rect 21269 13855 21327 13861
rect 18840 13812 18846 13824
rect 21269 13821 21281 13855
rect 21315 13852 21327 13855
rect 21726 13852 21732 13864
rect 21315 13824 21732 13852
rect 21315 13821 21327 13824
rect 21269 13815 21327 13821
rect 21726 13812 21732 13824
rect 21784 13852 21790 13864
rect 25314 13852 25320 13864
rect 21784 13824 25320 13852
rect 21784 13812 21790 13824
rect 25314 13812 25320 13824
rect 25372 13852 25378 13864
rect 26326 13852 26332 13864
rect 25372 13824 26332 13852
rect 25372 13812 25378 13824
rect 26326 13812 26332 13824
rect 26384 13812 26390 13864
rect 17957 13787 18015 13793
rect 17000 13756 17448 13784
rect 17000 13744 17006 13756
rect 1636 13688 2912 13716
rect 1636 13676 1642 13688
rect 4614 13676 4620 13728
rect 4672 13676 4678 13728
rect 5994 13676 6000 13728
rect 6052 13716 6058 13728
rect 8588 13716 8616 13744
rect 17420 13728 17448 13756
rect 17957 13753 17969 13787
rect 18003 13753 18015 13787
rect 17957 13747 18015 13753
rect 18064 13756 22094 13784
rect 6052 13688 8616 13716
rect 9217 13719 9275 13725
rect 6052 13676 6058 13688
rect 9217 13685 9229 13719
rect 9263 13716 9275 13719
rect 9582 13716 9588 13728
rect 9263 13688 9588 13716
rect 9263 13685 9275 13688
rect 9217 13679 9275 13685
rect 9582 13676 9588 13688
rect 9640 13676 9646 13728
rect 10594 13676 10600 13728
rect 10652 13676 10658 13728
rect 10870 13676 10876 13728
rect 10928 13716 10934 13728
rect 10965 13719 11023 13725
rect 10965 13716 10977 13719
rect 10928 13688 10977 13716
rect 10928 13676 10934 13688
rect 10965 13685 10977 13688
rect 11011 13685 11023 13719
rect 10965 13679 11023 13685
rect 17402 13676 17408 13728
rect 17460 13716 17466 13728
rect 18064 13716 18092 13756
rect 17460 13688 18092 13716
rect 22066 13716 22094 13756
rect 22278 13744 22284 13796
rect 22336 13784 22342 13796
rect 26988 13784 27016 13883
rect 27154 13880 27160 13932
rect 27212 13880 27218 13932
rect 27522 13880 27528 13932
rect 27580 13880 27586 13932
rect 27724 13864 27752 13960
rect 28184 13929 28212 13960
rect 27893 13923 27951 13929
rect 27893 13889 27905 13923
rect 27939 13889 27951 13923
rect 27893 13883 27951 13889
rect 28169 13923 28227 13929
rect 28169 13889 28181 13923
rect 28215 13889 28227 13923
rect 28368 13920 28396 14019
rect 28994 14016 29000 14068
rect 29052 14016 29058 14068
rect 32493 14059 32551 14065
rect 32493 14025 32505 14059
rect 32539 14056 32551 14059
rect 34606 14056 34612 14068
rect 32539 14028 34612 14056
rect 32539 14025 32551 14028
rect 32493 14019 32551 14025
rect 34606 14016 34612 14028
rect 34664 14016 34670 14068
rect 44082 14016 44088 14068
rect 44140 14056 44146 14068
rect 44453 14059 44511 14065
rect 44453 14056 44465 14059
rect 44140 14028 44465 14056
rect 44140 14016 44146 14028
rect 44453 14025 44465 14028
rect 44499 14025 44511 14059
rect 44453 14019 44511 14025
rect 28902 13948 28908 14000
rect 28960 13988 28966 14000
rect 28960 13948 28994 13988
rect 31662 13948 31668 14000
rect 31720 13988 31726 14000
rect 32125 13991 32183 13997
rect 32125 13988 32137 13991
rect 31720 13960 32137 13988
rect 31720 13948 31726 13960
rect 32125 13957 32137 13960
rect 32171 13957 32183 13991
rect 32125 13951 32183 13957
rect 32306 13948 32312 14000
rect 32364 13988 32370 14000
rect 33318 13988 33324 14000
rect 32364 13960 33324 13988
rect 32364 13948 32370 13960
rect 33318 13948 33324 13960
rect 33376 13948 33382 14000
rect 28534 13920 28540 13932
rect 28368 13892 28540 13920
rect 28169 13883 28227 13889
rect 27706 13812 27712 13864
rect 27764 13812 27770 13864
rect 27908 13852 27936 13883
rect 28534 13880 28540 13892
rect 28592 13920 28598 13932
rect 28813 13923 28871 13929
rect 28813 13920 28825 13923
rect 28592 13892 28825 13920
rect 28592 13880 28598 13892
rect 28813 13889 28825 13892
rect 28859 13889 28871 13923
rect 28966 13920 28994 13948
rect 33226 13920 33232 13932
rect 28966 13892 33232 13920
rect 28813 13883 28871 13889
rect 33226 13880 33232 13892
rect 33284 13880 33290 13932
rect 43070 13880 43076 13932
rect 43128 13920 43134 13932
rect 44269 13923 44327 13929
rect 44269 13920 44281 13923
rect 43128 13892 44281 13920
rect 43128 13880 43134 13892
rect 44269 13889 44281 13892
rect 44315 13889 44327 13923
rect 44269 13883 44327 13889
rect 34054 13852 34060 13864
rect 27908 13824 34060 13852
rect 34054 13812 34060 13824
rect 34112 13812 34118 13864
rect 28810 13784 28816 13796
rect 22336 13756 28816 13784
rect 22336 13744 22342 13756
rect 28810 13744 28816 13756
rect 28868 13744 28874 13796
rect 28902 13744 28908 13796
rect 28960 13784 28966 13796
rect 30282 13784 30288 13796
rect 28960 13756 30288 13784
rect 28960 13744 28966 13756
rect 30282 13744 30288 13756
rect 30340 13744 30346 13796
rect 32306 13784 32312 13796
rect 31726 13756 32312 13784
rect 25682 13716 25688 13728
rect 22066 13688 25688 13716
rect 17460 13676 17466 13688
rect 25682 13676 25688 13688
rect 25740 13716 25746 13728
rect 25869 13719 25927 13725
rect 25869 13716 25881 13719
rect 25740 13688 25881 13716
rect 25740 13676 25746 13688
rect 25869 13685 25881 13688
rect 25915 13685 25927 13719
rect 25869 13679 25927 13685
rect 26237 13719 26295 13725
rect 26237 13685 26249 13719
rect 26283 13716 26295 13719
rect 26418 13716 26424 13728
rect 26283 13688 26424 13716
rect 26283 13685 26295 13688
rect 26237 13679 26295 13685
rect 26418 13676 26424 13688
rect 26476 13676 26482 13728
rect 26694 13676 26700 13728
rect 26752 13716 26758 13728
rect 27893 13719 27951 13725
rect 27893 13716 27905 13719
rect 26752 13688 27905 13716
rect 26752 13676 26758 13688
rect 27893 13685 27905 13688
rect 27939 13716 27951 13719
rect 31726 13716 31754 13756
rect 32306 13744 32312 13756
rect 32364 13744 32370 13796
rect 27939 13688 31754 13716
rect 27939 13685 27951 13688
rect 27893 13679 27951 13685
rect 1104 13626 44896 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 44896 13626
rect 1104 13552 44896 13574
rect 2225 13515 2283 13521
rect 2225 13481 2237 13515
rect 2271 13512 2283 13515
rect 2866 13512 2872 13524
rect 2271 13484 2872 13512
rect 2271 13481 2283 13484
rect 2225 13475 2283 13481
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 4617 13515 4675 13521
rect 4617 13481 4629 13515
rect 4663 13512 4675 13515
rect 4706 13512 4712 13524
rect 4663 13484 4712 13512
rect 4663 13481 4675 13484
rect 4617 13475 4675 13481
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 4890 13472 4896 13524
rect 4948 13472 4954 13524
rect 5350 13472 5356 13524
rect 5408 13472 5414 13524
rect 5537 13515 5595 13521
rect 5537 13481 5549 13515
rect 5583 13512 5595 13515
rect 5718 13512 5724 13524
rect 5583 13484 5724 13512
rect 5583 13481 5595 13484
rect 5537 13475 5595 13481
rect 5718 13472 5724 13484
rect 5776 13512 5782 13524
rect 6546 13512 6552 13524
rect 5776 13484 6552 13512
rect 5776 13472 5782 13484
rect 6546 13472 6552 13484
rect 6604 13472 6610 13524
rect 6656 13484 6868 13512
rect 2409 13447 2467 13453
rect 2409 13413 2421 13447
rect 2455 13413 2467 13447
rect 2409 13407 2467 13413
rect 1578 13336 1584 13388
rect 1636 13336 1642 13388
rect 2038 13336 2044 13388
rect 2096 13385 2102 13388
rect 2096 13379 2124 13385
rect 2112 13376 2124 13379
rect 2424 13376 2452 13407
rect 2774 13404 2780 13456
rect 2832 13444 2838 13456
rect 3881 13447 3939 13453
rect 3881 13444 3893 13447
rect 2832 13416 3893 13444
rect 2832 13404 2838 13416
rect 3881 13413 3893 13416
rect 3927 13444 3939 13447
rect 4062 13444 4068 13456
rect 3927 13416 4068 13444
rect 3927 13413 3939 13416
rect 3881 13407 3939 13413
rect 4062 13404 4068 13416
rect 4120 13404 4126 13456
rect 5074 13404 5080 13456
rect 5132 13444 5138 13456
rect 5169 13447 5227 13453
rect 5169 13444 5181 13447
rect 5132 13416 5181 13444
rect 5132 13404 5138 13416
rect 5169 13413 5181 13416
rect 5215 13413 5227 13447
rect 5368 13444 5396 13472
rect 5368 13416 5488 13444
rect 5169 13407 5227 13413
rect 2682 13376 2688 13388
rect 2112 13348 2688 13376
rect 2112 13345 2124 13348
rect 2096 13339 2124 13345
rect 2096 13336 2102 13339
rect 2682 13336 2688 13348
rect 2740 13376 2746 13388
rect 3513 13379 3571 13385
rect 3513 13376 3525 13379
rect 2740 13348 3525 13376
rect 2740 13336 2746 13348
rect 3513 13345 3525 13348
rect 3559 13376 3571 13379
rect 4522 13376 4528 13388
rect 3559 13348 4528 13376
rect 3559 13345 3571 13348
rect 3513 13339 3571 13345
rect 4522 13336 4528 13348
rect 4580 13336 4586 13388
rect 5460 13376 5488 13416
rect 5810 13404 5816 13456
rect 5868 13404 5874 13456
rect 5902 13404 5908 13456
rect 5960 13444 5966 13456
rect 6656 13444 6684 13484
rect 5960 13416 6684 13444
rect 6840 13444 6868 13484
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 7377 13515 7435 13521
rect 7377 13512 7389 13515
rect 6972 13484 7389 13512
rect 6972 13472 6978 13484
rect 7377 13481 7389 13484
rect 7423 13481 7435 13515
rect 7377 13475 7435 13481
rect 7653 13515 7711 13521
rect 7653 13481 7665 13515
rect 7699 13512 7711 13515
rect 10410 13512 10416 13524
rect 7699 13484 10416 13512
rect 7699 13481 7711 13484
rect 7653 13475 7711 13481
rect 10410 13472 10416 13484
rect 10468 13472 10474 13524
rect 11241 13515 11299 13521
rect 11241 13481 11253 13515
rect 11287 13512 11299 13515
rect 11790 13512 11796 13524
rect 11287 13484 11796 13512
rect 11287 13481 11299 13484
rect 11241 13475 11299 13481
rect 11790 13472 11796 13484
rect 11848 13472 11854 13524
rect 11882 13472 11888 13524
rect 11940 13472 11946 13524
rect 12618 13512 12624 13524
rect 11992 13484 12624 13512
rect 11992 13456 12020 13484
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 13078 13472 13084 13524
rect 13136 13472 13142 13524
rect 13906 13472 13912 13524
rect 13964 13512 13970 13524
rect 13964 13484 17356 13512
rect 13964 13472 13970 13484
rect 8665 13447 8723 13453
rect 6840 13416 6873 13444
rect 5960 13404 5966 13416
rect 5441 13348 5488 13376
rect 5629 13379 5687 13385
rect 1949 13311 2007 13317
rect 1949 13277 1961 13311
rect 1995 13308 2007 13311
rect 2866 13308 2872 13320
rect 1995 13280 2872 13308
rect 1995 13277 2007 13280
rect 1949 13271 2007 13277
rect 2424 13249 2452 13280
rect 2866 13268 2872 13280
rect 2924 13268 2930 13320
rect 2961 13311 3019 13317
rect 2961 13277 2973 13311
rect 3007 13308 3019 13311
rect 4709 13311 4767 13317
rect 4709 13308 4721 13311
rect 3007 13280 3924 13308
rect 3007 13277 3019 13280
rect 2961 13271 3019 13277
rect 2409 13243 2467 13249
rect 2409 13209 2421 13243
rect 2455 13209 2467 13243
rect 2409 13203 2467 13209
rect 2774 13200 2780 13252
rect 2832 13240 2838 13252
rect 3896 13249 3924 13280
rect 4080 13280 4721 13308
rect 3329 13243 3387 13249
rect 3329 13240 3341 13243
rect 2832 13212 3341 13240
rect 2832 13200 2838 13212
rect 3329 13209 3341 13212
rect 3375 13240 3387 13243
rect 3881 13243 3939 13249
rect 3375 13212 3832 13240
rect 3375 13209 3387 13212
rect 3329 13203 3387 13209
rect 1857 13175 1915 13181
rect 1857 13141 1869 13175
rect 1903 13172 1915 13175
rect 2130 13172 2136 13184
rect 1903 13144 2136 13172
rect 1903 13141 1915 13144
rect 1857 13135 1915 13141
rect 2130 13132 2136 13144
rect 2188 13172 2194 13184
rect 2590 13172 2596 13184
rect 2188 13144 2596 13172
rect 2188 13132 2194 13144
rect 2590 13132 2596 13144
rect 2648 13172 2654 13184
rect 2869 13175 2927 13181
rect 2869 13172 2881 13175
rect 2648 13144 2881 13172
rect 2648 13132 2654 13144
rect 2869 13141 2881 13144
rect 2915 13141 2927 13175
rect 2869 13135 2927 13141
rect 3142 13132 3148 13184
rect 3200 13132 3206 13184
rect 3804 13172 3832 13212
rect 3881 13209 3893 13243
rect 3927 13240 3939 13243
rect 3970 13240 3976 13252
rect 3927 13212 3976 13240
rect 3927 13209 3939 13212
rect 3881 13203 3939 13209
rect 3970 13200 3976 13212
rect 4028 13200 4034 13252
rect 4080 13172 4108 13280
rect 4709 13277 4721 13280
rect 4755 13277 4767 13311
rect 4709 13271 4767 13277
rect 4798 13268 4804 13320
rect 4856 13308 4862 13320
rect 5441 13317 5469 13348
rect 5629 13345 5641 13379
rect 5675 13376 5687 13379
rect 5828 13376 5856 13404
rect 5675 13348 5948 13376
rect 5675 13345 5687 13348
rect 5629 13339 5687 13345
rect 4985 13311 5043 13317
rect 4985 13308 4997 13311
rect 4856 13280 4997 13308
rect 4856 13268 4862 13280
rect 4985 13277 4997 13280
rect 5031 13277 5043 13311
rect 4985 13271 5043 13277
rect 5408 13311 5469 13317
rect 5408 13277 5420 13311
rect 5454 13280 5469 13311
rect 5920 13308 5948 13348
rect 5994 13336 6000 13388
rect 6052 13336 6058 13388
rect 6380 13385 6408 13416
rect 6365 13379 6423 13385
rect 6365 13345 6377 13379
rect 6411 13345 6423 13379
rect 6365 13339 6423 13345
rect 6457 13379 6515 13385
rect 6457 13345 6469 13379
rect 6503 13376 6515 13379
rect 6638 13376 6644 13388
rect 6503 13348 6644 13376
rect 6503 13345 6515 13348
rect 6457 13339 6515 13345
rect 6638 13336 6644 13348
rect 6696 13336 6702 13388
rect 5920 13280 6291 13308
rect 5454 13277 5466 13280
rect 5408 13271 5466 13277
rect 4338 13200 4344 13252
rect 4396 13240 4402 13252
rect 4396 13212 4660 13240
rect 4396 13200 4402 13212
rect 3804 13144 4108 13172
rect 4433 13175 4491 13181
rect 4433 13141 4445 13175
rect 4479 13172 4491 13175
rect 4522 13172 4528 13184
rect 4479 13144 4528 13172
rect 4479 13141 4491 13144
rect 4433 13135 4491 13141
rect 4522 13132 4528 13144
rect 4580 13132 4586 13184
rect 4632 13172 4660 13212
rect 5258 13200 5264 13252
rect 5316 13240 5322 13252
rect 5902 13240 5908 13252
rect 5316 13212 5908 13240
rect 5316 13200 5322 13212
rect 5902 13200 5908 13212
rect 5960 13200 5966 13252
rect 6263 13249 6291 13280
rect 6546 13268 6552 13320
rect 6604 13308 6610 13320
rect 6733 13311 6791 13317
rect 6733 13308 6745 13311
rect 6604 13280 6745 13308
rect 6604 13268 6610 13280
rect 6733 13277 6745 13280
rect 6779 13277 6791 13311
rect 6845 13308 6873 13416
rect 8665 13413 8677 13447
rect 8711 13444 8723 13447
rect 8846 13444 8852 13456
rect 8711 13416 8852 13444
rect 8711 13413 8723 13416
rect 8665 13407 8723 13413
rect 8846 13404 8852 13416
rect 8904 13404 8910 13456
rect 9122 13404 9128 13456
rect 9180 13404 9186 13456
rect 9306 13404 9312 13456
rect 9364 13404 9370 13456
rect 9490 13404 9496 13456
rect 9548 13444 9554 13456
rect 10962 13444 10968 13456
rect 9548 13416 10968 13444
rect 9548 13404 9554 13416
rect 10962 13404 10968 13416
rect 11020 13404 11026 13456
rect 11514 13404 11520 13456
rect 11572 13444 11578 13456
rect 11974 13444 11980 13456
rect 11572 13416 11980 13444
rect 11572 13404 11578 13416
rect 11974 13404 11980 13416
rect 12032 13404 12038 13456
rect 13814 13444 13820 13456
rect 12544 13416 13820 13444
rect 8018 13336 8024 13388
rect 8076 13376 8082 13388
rect 9324 13376 9352 13404
rect 8076 13348 8432 13376
rect 9324 13348 9536 13376
rect 8076 13336 8082 13348
rect 7193 13311 7251 13317
rect 7193 13308 7205 13311
rect 6845 13280 7205 13308
rect 6733 13271 6791 13277
rect 7193 13277 7205 13280
rect 7239 13277 7251 13311
rect 7193 13271 7251 13277
rect 7466 13268 7472 13320
rect 7524 13268 7530 13320
rect 7558 13268 7564 13320
rect 7616 13308 7622 13320
rect 8404 13317 8432 13348
rect 7837 13311 7895 13317
rect 7837 13308 7849 13311
rect 7616 13280 7849 13308
rect 7616 13268 7622 13280
rect 7837 13277 7849 13280
rect 7883 13277 7895 13311
rect 7837 13271 7895 13277
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 8570 13268 8576 13320
rect 8628 13308 8634 13320
rect 9398 13317 9404 13320
rect 9257 13311 9315 13317
rect 9257 13308 9269 13311
rect 8628 13280 9269 13308
rect 8628 13268 8634 13280
rect 9257 13277 9269 13280
rect 9303 13277 9315 13311
rect 9257 13271 9315 13277
rect 9388 13311 9404 13317
rect 9388 13277 9400 13311
rect 9388 13271 9404 13277
rect 9398 13268 9404 13271
rect 9456 13268 9462 13320
rect 9508 13317 9536 13348
rect 9582 13336 9588 13388
rect 9640 13376 9646 13388
rect 12544 13376 12572 13416
rect 13814 13404 13820 13416
rect 13872 13404 13878 13456
rect 14182 13404 14188 13456
rect 14240 13444 14246 13456
rect 15470 13444 15476 13456
rect 14240 13416 15476 13444
rect 14240 13404 14246 13416
rect 15470 13404 15476 13416
rect 15528 13404 15534 13456
rect 17328 13444 17356 13484
rect 17402 13472 17408 13524
rect 17460 13472 17466 13524
rect 22278 13472 22284 13524
rect 22336 13472 22342 13524
rect 22462 13472 22468 13524
rect 22520 13472 22526 13524
rect 25317 13515 25375 13521
rect 25317 13481 25329 13515
rect 25363 13512 25375 13515
rect 26050 13512 26056 13524
rect 25363 13484 26056 13512
rect 25363 13481 25375 13484
rect 25317 13475 25375 13481
rect 26050 13472 26056 13484
rect 26108 13472 26114 13524
rect 26602 13472 26608 13524
rect 26660 13512 26666 13524
rect 26697 13515 26755 13521
rect 26697 13512 26709 13515
rect 26660 13484 26709 13512
rect 26660 13472 26666 13484
rect 26697 13481 26709 13484
rect 26743 13481 26755 13515
rect 27154 13512 27160 13524
rect 26697 13475 26755 13481
rect 26804 13484 27160 13512
rect 17770 13444 17776 13456
rect 17328 13416 17776 13444
rect 17770 13404 17776 13416
rect 17828 13444 17834 13456
rect 22094 13444 22100 13456
rect 17828 13416 22100 13444
rect 17828 13404 17834 13416
rect 22094 13404 22100 13416
rect 22152 13404 22158 13456
rect 26804 13444 26832 13484
rect 27154 13472 27160 13484
rect 27212 13472 27218 13524
rect 28905 13515 28963 13521
rect 28905 13481 28917 13515
rect 28951 13512 28963 13515
rect 28994 13512 29000 13524
rect 28951 13484 29000 13512
rect 28951 13481 28963 13484
rect 28905 13475 28963 13481
rect 28994 13472 29000 13484
rect 29052 13472 29058 13524
rect 29273 13515 29331 13521
rect 29273 13481 29285 13515
rect 29319 13512 29331 13515
rect 30006 13512 30012 13524
rect 29319 13484 30012 13512
rect 29319 13481 29331 13484
rect 29273 13475 29331 13481
rect 30006 13472 30012 13484
rect 30064 13472 30070 13524
rect 31389 13515 31447 13521
rect 31389 13481 31401 13515
rect 31435 13512 31447 13515
rect 36078 13512 36084 13524
rect 31435 13484 36084 13512
rect 31435 13481 31447 13484
rect 31389 13475 31447 13481
rect 36078 13472 36084 13484
rect 36136 13472 36142 13524
rect 22204 13416 26832 13444
rect 9640 13348 12572 13376
rect 9640 13336 9646 13348
rect 9692 13317 9720 13348
rect 9493 13311 9551 13317
rect 9493 13277 9505 13311
rect 9539 13277 9551 13311
rect 9493 13271 9551 13277
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 9950 13268 9956 13320
rect 10008 13268 10014 13320
rect 10042 13268 10048 13320
rect 10100 13308 10106 13320
rect 10704 13317 10732 13348
rect 10321 13311 10379 13317
rect 10321 13308 10333 13311
rect 10100 13280 10333 13308
rect 10100 13268 10106 13280
rect 10321 13277 10333 13280
rect 10367 13277 10379 13311
rect 10321 13271 10379 13277
rect 10689 13311 10747 13317
rect 10689 13277 10701 13311
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 10962 13268 10968 13320
rect 11020 13268 11026 13320
rect 11109 13311 11167 13317
rect 11109 13277 11121 13311
rect 11155 13308 11167 13311
rect 11514 13308 11520 13320
rect 11155 13280 11520 13308
rect 11155 13277 11167 13280
rect 11109 13271 11167 13277
rect 11514 13268 11520 13280
rect 11572 13268 11578 13320
rect 11698 13268 11704 13320
rect 11756 13268 11762 13320
rect 11974 13268 11980 13320
rect 12032 13317 12038 13320
rect 12032 13311 12075 13317
rect 12063 13277 12075 13311
rect 12032 13271 12075 13277
rect 12032 13268 12038 13271
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 12273 13308 12301 13348
rect 12216 13280 12301 13308
rect 12216 13268 12222 13280
rect 12342 13268 12348 13320
rect 12400 13308 12406 13320
rect 12544 13317 12572 13348
rect 12618 13336 12624 13388
rect 12676 13376 12682 13388
rect 15488 13376 15516 13404
rect 22204 13385 22232 13416
rect 22189 13379 22247 13385
rect 22189 13376 22201 13379
rect 12676 13348 13308 13376
rect 12676 13336 12682 13348
rect 12437 13311 12495 13317
rect 12437 13308 12449 13311
rect 12400 13280 12449 13308
rect 12400 13268 12406 13280
rect 12437 13277 12449 13280
rect 12483 13277 12495 13311
rect 12437 13271 12495 13277
rect 12529 13311 12587 13317
rect 12529 13277 12541 13311
rect 12575 13277 12587 13311
rect 12529 13271 12587 13277
rect 6248 13243 6306 13249
rect 6248 13209 6260 13243
rect 6294 13240 6306 13243
rect 6825 13243 6883 13249
rect 6825 13240 6837 13243
rect 6294 13212 6837 13240
rect 6294 13209 6306 13212
rect 6248 13203 6306 13209
rect 6825 13209 6837 13212
rect 6871 13209 6883 13243
rect 6825 13203 6883 13209
rect 6914 13200 6920 13252
rect 6972 13240 6978 13252
rect 7101 13243 7159 13249
rect 7101 13240 7113 13243
rect 6972 13212 7113 13240
rect 6972 13200 6978 13212
rect 7101 13209 7113 13212
rect 7147 13209 7159 13243
rect 7101 13203 7159 13209
rect 10870 13200 10876 13252
rect 10928 13240 10934 13252
rect 12253 13243 12311 13249
rect 12253 13240 12265 13243
rect 10928 13212 12265 13240
rect 10928 13200 10934 13212
rect 12253 13209 12265 13212
rect 12299 13209 12311 13243
rect 12452 13240 12480 13271
rect 12710 13268 12716 13320
rect 12768 13268 12774 13320
rect 12894 13268 12900 13320
rect 12952 13317 12958 13320
rect 13280 13317 13308 13348
rect 13372 13348 13768 13376
rect 15488 13348 19334 13376
rect 12952 13308 12960 13317
rect 13265 13311 13323 13317
rect 12952 13280 12997 13308
rect 12952 13271 12960 13280
rect 13265 13277 13277 13311
rect 13311 13277 13323 13311
rect 13265 13271 13323 13277
rect 12952 13268 12958 13271
rect 12805 13243 12863 13249
rect 12805 13240 12817 13243
rect 12452 13212 12817 13240
rect 12253 13203 12311 13209
rect 12805 13209 12817 13212
rect 12851 13240 12863 13243
rect 13372 13240 13400 13348
rect 13630 13268 13636 13320
rect 13688 13268 13694 13320
rect 12851 13212 13400 13240
rect 12851 13209 12863 13212
rect 12805 13203 12863 13209
rect 5350 13172 5356 13184
rect 4632 13144 5356 13172
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 6086 13132 6092 13184
rect 6144 13132 6150 13184
rect 6546 13132 6552 13184
rect 6604 13172 6610 13184
rect 7009 13175 7067 13181
rect 7009 13172 7021 13175
rect 6604 13144 7021 13172
rect 6604 13132 6610 13144
rect 7009 13141 7021 13144
rect 7055 13141 7067 13175
rect 7009 13135 7067 13141
rect 8110 13132 8116 13184
rect 8168 13172 8174 13184
rect 9858 13172 9864 13184
rect 8168 13144 9864 13172
rect 8168 13132 8174 13144
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 10137 13175 10195 13181
rect 10137 13141 10149 13175
rect 10183 13172 10195 13175
rect 10410 13172 10416 13184
rect 10183 13144 10416 13172
rect 10183 13141 10195 13144
rect 10137 13135 10195 13141
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 10505 13175 10563 13181
rect 10505 13141 10517 13175
rect 10551 13172 10563 13175
rect 11146 13172 11152 13184
rect 10551 13144 11152 13172
rect 10551 13141 10563 13144
rect 10505 13135 10563 13141
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 12268 13172 12296 13203
rect 13446 13200 13452 13252
rect 13504 13200 13510 13252
rect 13541 13243 13599 13249
rect 13541 13209 13553 13243
rect 13587 13209 13599 13243
rect 13740 13240 13768 13348
rect 14642 13268 14648 13320
rect 14700 13268 14706 13320
rect 15010 13268 15016 13320
rect 15068 13268 15074 13320
rect 15197 13311 15255 13317
rect 15197 13277 15209 13311
rect 15243 13308 15255 13311
rect 15654 13308 15660 13320
rect 15243 13280 15660 13308
rect 15243 13277 15255 13280
rect 15197 13271 15255 13277
rect 15654 13268 15660 13280
rect 15712 13308 15718 13320
rect 16853 13311 16911 13317
rect 15712 13280 16620 13308
rect 15712 13268 15718 13280
rect 16022 13240 16028 13252
rect 13740 13212 16028 13240
rect 13541 13203 13599 13209
rect 13556 13172 13584 13203
rect 16022 13200 16028 13212
rect 16080 13200 16086 13252
rect 12268 13144 13584 13172
rect 13817 13175 13875 13181
rect 13817 13141 13829 13175
rect 13863 13172 13875 13175
rect 13906 13172 13912 13184
rect 13863 13144 13912 13172
rect 13863 13141 13875 13144
rect 13817 13135 13875 13141
rect 13906 13132 13912 13144
rect 13964 13132 13970 13184
rect 14274 13132 14280 13184
rect 14332 13172 14338 13184
rect 14737 13175 14795 13181
rect 14737 13172 14749 13175
rect 14332 13144 14749 13172
rect 14332 13132 14338 13144
rect 14737 13141 14749 13144
rect 14783 13141 14795 13175
rect 16592 13172 16620 13280
rect 16853 13277 16865 13311
rect 16899 13308 16911 13311
rect 16942 13308 16948 13320
rect 16899 13280 16948 13308
rect 16899 13277 16911 13280
rect 16853 13271 16911 13277
rect 16942 13268 16948 13280
rect 17000 13268 17006 13320
rect 17226 13311 17284 13317
rect 17226 13277 17238 13311
rect 17272 13308 17284 13311
rect 17494 13308 17500 13320
rect 17272 13280 17500 13308
rect 17272 13277 17284 13280
rect 17226 13271 17284 13277
rect 17494 13268 17500 13280
rect 17552 13308 17558 13320
rect 17954 13308 17960 13320
rect 17552 13280 17960 13308
rect 17552 13268 17558 13280
rect 17954 13268 17960 13280
rect 18012 13268 18018 13320
rect 19306 13308 19334 13348
rect 19996 13348 22201 13376
rect 19996 13308 20024 13348
rect 22189 13345 22201 13348
rect 22235 13345 22247 13379
rect 26602 13376 26608 13388
rect 22189 13339 22247 13345
rect 25424 13348 26608 13376
rect 19306 13280 20024 13308
rect 22097 13311 22155 13317
rect 22097 13277 22109 13311
rect 22143 13308 22155 13311
rect 25424 13308 25452 13348
rect 26602 13336 26608 13348
rect 26660 13336 26666 13388
rect 26804 13385 26832 13416
rect 27065 13447 27123 13453
rect 27065 13413 27077 13447
rect 27111 13444 27123 13447
rect 27111 13416 31754 13444
rect 27111 13413 27123 13416
rect 27065 13407 27123 13413
rect 26789 13379 26847 13385
rect 26789 13345 26801 13379
rect 26835 13345 26847 13379
rect 28902 13376 28908 13388
rect 26789 13339 26847 13345
rect 26896 13348 28908 13376
rect 22143 13280 25452 13308
rect 25516 13280 26280 13308
rect 22143 13277 22155 13280
rect 22097 13271 22155 13277
rect 17034 13200 17040 13252
rect 17092 13200 17098 13252
rect 17126 13200 17132 13252
rect 17184 13240 17190 13252
rect 19150 13240 19156 13252
rect 17184 13212 19156 13240
rect 17184 13200 17190 13212
rect 19150 13200 19156 13212
rect 19208 13200 19214 13252
rect 20070 13200 20076 13252
rect 20128 13240 20134 13252
rect 22112 13240 22140 13271
rect 20128 13212 22140 13240
rect 20128 13200 20134 13212
rect 23474 13200 23480 13252
rect 23532 13240 23538 13252
rect 25516 13249 25544 13280
rect 25501 13243 25559 13249
rect 25501 13240 25513 13243
rect 23532 13212 25513 13240
rect 23532 13200 23538 13212
rect 25501 13209 25513 13212
rect 25547 13209 25559 13243
rect 25501 13203 25559 13209
rect 25685 13243 25743 13249
rect 25685 13209 25697 13243
rect 25731 13240 25743 13243
rect 25866 13240 25872 13252
rect 25731 13212 25872 13240
rect 25731 13209 25743 13212
rect 25685 13203 25743 13209
rect 18322 13172 18328 13184
rect 16592 13144 18328 13172
rect 14737 13135 14795 13141
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 22094 13132 22100 13184
rect 22152 13172 22158 13184
rect 25700 13172 25728 13203
rect 25866 13200 25872 13212
rect 25924 13200 25930 13252
rect 26252 13240 26280 13280
rect 26326 13268 26332 13320
rect 26384 13308 26390 13320
rect 26697 13311 26755 13317
rect 26697 13308 26709 13311
rect 26384 13280 26709 13308
rect 26384 13268 26390 13280
rect 26697 13277 26709 13280
rect 26743 13277 26755 13311
rect 26697 13271 26755 13277
rect 26896 13240 26924 13348
rect 28902 13336 28908 13348
rect 28960 13336 28966 13388
rect 29638 13376 29644 13388
rect 29012 13348 29644 13376
rect 28534 13268 28540 13320
rect 28592 13268 28598 13320
rect 28721 13311 28779 13317
rect 28721 13277 28733 13311
rect 28767 13308 28779 13311
rect 29012 13308 29040 13348
rect 29638 13336 29644 13348
rect 29696 13336 29702 13388
rect 31018 13336 31024 13388
rect 31076 13376 31082 13388
rect 31570 13376 31576 13388
rect 31076 13348 31576 13376
rect 31076 13336 31082 13348
rect 28767 13280 29040 13308
rect 29089 13311 29147 13317
rect 28767 13277 28779 13280
rect 28721 13271 28779 13277
rect 29089 13277 29101 13311
rect 29135 13308 29147 13311
rect 31386 13308 31392 13320
rect 29135 13280 31392 13308
rect 29135 13277 29147 13280
rect 29089 13271 29147 13277
rect 31386 13268 31392 13280
rect 31444 13268 31450 13320
rect 26252 13212 26924 13240
rect 28350 13200 28356 13252
rect 28408 13200 28414 13252
rect 28810 13200 28816 13252
rect 28868 13200 28874 13252
rect 29196 13212 29408 13240
rect 22152 13144 25728 13172
rect 28368 13172 28396 13200
rect 29196 13172 29224 13212
rect 28368 13144 29224 13172
rect 29380 13172 29408 13212
rect 29454 13200 29460 13252
rect 29512 13240 29518 13252
rect 30745 13243 30803 13249
rect 30745 13240 30757 13243
rect 29512 13212 30757 13240
rect 29512 13200 29518 13212
rect 30745 13209 30757 13212
rect 30791 13209 30803 13243
rect 30745 13203 30803 13209
rect 30926 13200 30932 13252
rect 30984 13200 30990 13252
rect 31110 13200 31116 13252
rect 31168 13200 31174 13252
rect 31496 13249 31524 13348
rect 31570 13336 31576 13348
rect 31628 13336 31634 13388
rect 31726 13376 31754 13416
rect 37918 13376 37924 13388
rect 31726 13348 37924 13376
rect 37918 13336 37924 13348
rect 37976 13336 37982 13388
rect 31481 13243 31539 13249
rect 31481 13209 31493 13243
rect 31527 13209 31539 13243
rect 31481 13203 31539 13209
rect 31662 13200 31668 13252
rect 31720 13200 31726 13252
rect 37550 13172 37556 13184
rect 29380 13144 37556 13172
rect 22152 13132 22158 13144
rect 37550 13132 37556 13144
rect 37608 13132 37614 13184
rect 1104 13082 44896 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 44896 13082
rect 1104 13008 44896 13030
rect 1578 12928 1584 12980
rect 1636 12968 1642 12980
rect 1673 12971 1731 12977
rect 1673 12968 1685 12971
rect 1636 12940 1685 12968
rect 1636 12928 1642 12940
rect 1673 12937 1685 12940
rect 1719 12937 1731 12971
rect 1673 12931 1731 12937
rect 2593 12971 2651 12977
rect 2593 12937 2605 12971
rect 2639 12968 2651 12971
rect 2682 12968 2688 12980
rect 2639 12940 2688 12968
rect 2639 12937 2651 12940
rect 2593 12931 2651 12937
rect 2682 12928 2688 12940
rect 2740 12928 2746 12980
rect 2777 12971 2835 12977
rect 2777 12937 2789 12971
rect 2823 12968 2835 12971
rect 3326 12968 3332 12980
rect 2823 12940 3332 12968
rect 2823 12937 2835 12940
rect 2777 12931 2835 12937
rect 3326 12928 3332 12940
rect 3384 12928 3390 12980
rect 3421 12971 3479 12977
rect 3421 12937 3433 12971
rect 3467 12968 3479 12971
rect 4798 12968 4804 12980
rect 3467 12940 4804 12968
rect 3467 12937 3479 12940
rect 3421 12931 3479 12937
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 5077 12971 5135 12977
rect 5077 12937 5089 12971
rect 5123 12968 5135 12971
rect 5534 12968 5540 12980
rect 5123 12940 5540 12968
rect 5123 12937 5135 12940
rect 5077 12931 5135 12937
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 6089 12971 6147 12977
rect 6089 12937 6101 12971
rect 6135 12968 6147 12971
rect 10042 12968 10048 12980
rect 6135 12940 10048 12968
rect 6135 12937 6147 12940
rect 6089 12931 6147 12937
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 10560 12940 11008 12968
rect 10560 12928 10566 12940
rect 2041 12903 2099 12909
rect 2041 12869 2053 12903
rect 2087 12900 2099 12903
rect 2498 12900 2504 12912
rect 2087 12872 2504 12900
rect 2087 12869 2099 12872
rect 2041 12863 2099 12869
rect 2498 12860 2504 12872
rect 2556 12860 2562 12912
rect 2746 12872 4016 12900
rect 1578 12792 1584 12844
rect 1636 12832 1642 12844
rect 1765 12835 1823 12841
rect 1765 12832 1777 12835
rect 1636 12804 1777 12832
rect 1636 12792 1642 12804
rect 1765 12801 1777 12804
rect 1811 12832 1823 12835
rect 2746 12832 2774 12872
rect 1811 12804 2774 12832
rect 1811 12801 1823 12804
rect 1765 12795 1823 12801
rect 2958 12792 2964 12844
rect 3016 12792 3022 12844
rect 3234 12792 3240 12844
rect 3292 12792 3298 12844
rect 3988 12841 4016 12872
rect 5350 12860 5356 12912
rect 5408 12900 5414 12912
rect 9582 12900 9588 12912
rect 5408 12872 6868 12900
rect 5408 12860 5414 12872
rect 3973 12835 4031 12841
rect 3973 12801 3985 12835
rect 4019 12801 4031 12835
rect 3973 12795 4031 12801
rect 4249 12835 4307 12841
rect 4249 12801 4261 12835
rect 4295 12832 4307 12835
rect 5258 12832 5264 12844
rect 4295 12804 5264 12832
rect 4295 12801 4307 12804
rect 4249 12795 4307 12801
rect 1670 12724 1676 12776
rect 1728 12764 1734 12776
rect 2498 12764 2504 12776
rect 1728 12736 2504 12764
rect 1728 12724 1734 12736
rect 2498 12724 2504 12736
rect 2556 12724 2562 12776
rect 2590 12724 2596 12776
rect 2648 12764 2654 12776
rect 3145 12767 3203 12773
rect 3145 12764 3157 12767
rect 2648 12736 3157 12764
rect 2648 12724 2654 12736
rect 3145 12733 3157 12736
rect 3191 12764 3203 12767
rect 4338 12764 4344 12776
rect 3191 12736 4344 12764
rect 3191 12733 3203 12736
rect 3145 12727 3203 12733
rect 4338 12724 4344 12736
rect 4396 12724 4402 12776
rect 2041 12699 2099 12705
rect 2041 12665 2053 12699
rect 2087 12696 2099 12699
rect 2866 12696 2872 12708
rect 2087 12668 2872 12696
rect 2087 12665 2099 12668
rect 2041 12659 2099 12665
rect 2866 12656 2872 12668
rect 2924 12656 2930 12708
rect 4157 12699 4215 12705
rect 4157 12665 4169 12699
rect 4203 12696 4215 12699
rect 4448 12696 4476 12804
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 5776 12804 5825 12832
rect 5776 12792 5782 12804
rect 5813 12801 5825 12804
rect 5859 12832 5871 12835
rect 6733 12835 6791 12841
rect 6733 12832 6745 12835
rect 5859 12804 6745 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 6733 12801 6745 12804
rect 6779 12801 6791 12835
rect 6733 12795 6791 12801
rect 4801 12767 4859 12773
rect 4801 12733 4813 12767
rect 4847 12764 4859 12767
rect 5442 12764 5448 12776
rect 4847 12736 5448 12764
rect 4847 12733 4859 12736
rect 4801 12727 4859 12733
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 5902 12724 5908 12776
rect 5960 12764 5966 12776
rect 6457 12767 6515 12773
rect 6457 12764 6469 12767
rect 5960 12736 6469 12764
rect 5960 12724 5966 12736
rect 6457 12733 6469 12736
rect 6503 12733 6515 12767
rect 6457 12727 6515 12733
rect 6546 12724 6552 12776
rect 6604 12724 6610 12776
rect 6641 12767 6699 12773
rect 6641 12733 6653 12767
rect 6687 12764 6699 12767
rect 6840 12764 6868 12872
rect 8404 12872 9588 12900
rect 7190 12792 7196 12844
rect 7248 12832 7254 12844
rect 8018 12832 8024 12844
rect 7248 12804 8024 12832
rect 7248 12792 7254 12804
rect 8018 12792 8024 12804
rect 8076 12832 8082 12844
rect 8404 12841 8432 12872
rect 9582 12860 9588 12872
rect 9640 12900 9646 12912
rect 10229 12903 10287 12909
rect 10229 12900 10241 12903
rect 9640 12872 10241 12900
rect 9640 12860 9646 12872
rect 10229 12869 10241 12872
rect 10275 12869 10287 12903
rect 10229 12863 10287 12869
rect 10318 12860 10324 12912
rect 10376 12900 10382 12912
rect 10980 12900 11008 12940
rect 11606 12928 11612 12980
rect 11664 12928 11670 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 13357 12971 13415 12977
rect 13357 12968 13369 12971
rect 12492 12940 13369 12968
rect 12492 12928 12498 12940
rect 13357 12937 13369 12940
rect 13403 12937 13415 12971
rect 14366 12968 14372 12980
rect 13357 12931 13415 12937
rect 14016 12940 14372 12968
rect 14016 12912 14044 12940
rect 14366 12928 14372 12940
rect 14424 12928 14430 12980
rect 14550 12928 14556 12980
rect 14608 12968 14614 12980
rect 15473 12971 15531 12977
rect 15473 12968 15485 12971
rect 14608 12940 15485 12968
rect 14608 12928 14614 12940
rect 15473 12937 15485 12940
rect 15519 12937 15531 12971
rect 17586 12968 17592 12980
rect 15473 12931 15531 12937
rect 17328 12940 17592 12968
rect 17328 12912 17356 12940
rect 17586 12928 17592 12940
rect 17644 12928 17650 12980
rect 18782 12968 18788 12980
rect 18064 12940 18788 12968
rect 12897 12903 12955 12909
rect 12897 12900 12909 12903
rect 10376 12872 10824 12900
rect 10980 12872 12909 12900
rect 10376 12860 10382 12872
rect 8389 12835 8447 12841
rect 8389 12832 8401 12835
rect 8076 12804 8401 12832
rect 8076 12792 8082 12804
rect 8389 12801 8401 12804
rect 8435 12801 8447 12835
rect 8389 12795 8447 12801
rect 8757 12835 8815 12841
rect 8757 12801 8769 12835
rect 8803 12832 8815 12835
rect 8846 12832 8852 12844
rect 8803 12804 8852 12832
rect 8803 12801 8815 12804
rect 8757 12795 8815 12801
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 8941 12835 8999 12841
rect 8941 12801 8953 12835
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 6687 12736 6868 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 7926 12724 7932 12776
rect 7984 12724 7990 12776
rect 8110 12724 8116 12776
rect 8168 12764 8174 12776
rect 8205 12767 8263 12773
rect 8205 12764 8217 12767
rect 8168 12736 8217 12764
rect 8168 12724 8174 12736
rect 8205 12733 8217 12736
rect 8251 12733 8263 12767
rect 8205 12727 8263 12733
rect 8956 12764 8984 12795
rect 9674 12792 9680 12844
rect 9732 12792 9738 12844
rect 9766 12792 9772 12844
rect 9824 12832 9830 12844
rect 10045 12835 10103 12841
rect 10045 12832 10057 12835
rect 9824 12804 10057 12832
rect 9824 12792 9830 12804
rect 10045 12801 10057 12804
rect 10091 12801 10103 12835
rect 10418 12835 10476 12841
rect 10418 12832 10430 12835
rect 10045 12795 10103 12801
rect 10341 12804 10430 12832
rect 10341 12764 10369 12804
rect 10418 12801 10430 12804
rect 10464 12832 10476 12835
rect 10686 12832 10692 12844
rect 10464 12804 10692 12832
rect 10464 12801 10476 12804
rect 10418 12795 10476 12801
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 10796 12841 10824 12872
rect 12897 12869 12909 12872
rect 12943 12869 12955 12903
rect 12897 12863 12955 12869
rect 13262 12860 13268 12912
rect 13320 12860 13326 12912
rect 13998 12860 14004 12912
rect 14056 12860 14062 12912
rect 14093 12903 14151 12909
rect 14093 12869 14105 12903
rect 14139 12900 14151 12903
rect 15010 12900 15016 12912
rect 14139 12872 15016 12900
rect 14139 12869 14151 12872
rect 14093 12863 14151 12869
rect 15010 12860 15016 12872
rect 15068 12860 15074 12912
rect 15212 12872 17264 12900
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 11146 12792 11152 12844
rect 11204 12792 11210 12844
rect 12158 12792 12164 12844
rect 12216 12792 12222 12844
rect 12434 12792 12440 12844
rect 12492 12832 12498 12844
rect 12529 12835 12587 12841
rect 12529 12832 12541 12835
rect 12492 12804 12541 12832
rect 12492 12792 12498 12804
rect 12529 12801 12541 12804
rect 12575 12801 12587 12835
rect 12529 12795 12587 12801
rect 12713 12835 12771 12841
rect 12713 12801 12725 12835
rect 12759 12832 12771 12835
rect 13081 12835 13139 12841
rect 13081 12832 13093 12835
rect 12759 12804 13093 12832
rect 12759 12801 12771 12804
rect 12713 12795 12771 12801
rect 13081 12801 13093 12804
rect 13127 12801 13139 12835
rect 13081 12795 13139 12801
rect 8956 12736 10369 12764
rect 10480 12736 11652 12764
rect 4203 12668 4476 12696
rect 4203 12665 4215 12668
rect 4157 12659 4215 12665
rect 4614 12656 4620 12708
rect 4672 12656 4678 12708
rect 4706 12656 4712 12708
rect 4764 12656 4770 12708
rect 5353 12699 5411 12705
rect 5353 12696 5365 12699
rect 4816 12668 5365 12696
rect 2498 12588 2504 12640
rect 2556 12628 2562 12640
rect 3970 12628 3976 12640
rect 2556 12600 3976 12628
rect 2556 12588 2562 12600
rect 3970 12588 3976 12600
rect 4028 12588 4034 12640
rect 4522 12588 4528 12640
rect 4580 12628 4586 12640
rect 4816 12628 4844 12668
rect 5353 12665 5365 12668
rect 5399 12665 5411 12699
rect 5353 12659 5411 12665
rect 4580 12600 4844 12628
rect 5368 12628 5396 12659
rect 5626 12656 5632 12708
rect 5684 12696 5690 12708
rect 6917 12699 6975 12705
rect 6917 12696 6929 12699
rect 5684 12668 6929 12696
rect 5684 12656 5690 12668
rect 6917 12665 6929 12668
rect 6963 12665 6975 12699
rect 6917 12659 6975 12665
rect 7374 12656 7380 12708
rect 7432 12696 7438 12708
rect 7742 12696 7748 12708
rect 7432 12668 7748 12696
rect 7432 12656 7438 12668
rect 7742 12656 7748 12668
rect 7800 12696 7806 12708
rect 8956 12696 8984 12736
rect 7800 12668 8984 12696
rect 7800 12656 7806 12668
rect 9490 12656 9496 12708
rect 9548 12656 9554 12708
rect 9582 12656 9588 12708
rect 9640 12696 9646 12708
rect 10480 12696 10508 12736
rect 9640 12668 10508 12696
rect 11624 12696 11652 12736
rect 12250 12724 12256 12776
rect 12308 12724 12314 12776
rect 13096 12764 13124 12795
rect 13814 12792 13820 12844
rect 13872 12792 13878 12844
rect 14237 12835 14295 12841
rect 14237 12801 14249 12835
rect 14283 12832 14295 12835
rect 14550 12832 14556 12844
rect 14283 12804 14556 12832
rect 14283 12801 14295 12804
rect 14237 12795 14295 12801
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 14734 12792 14740 12844
rect 14792 12792 14798 12844
rect 14826 12792 14832 12844
rect 14884 12792 14890 12844
rect 14926 12835 14984 12841
rect 14926 12801 14938 12835
rect 14972 12832 14984 12835
rect 15212 12832 15240 12872
rect 14972 12804 15240 12832
rect 14972 12801 14984 12804
rect 14926 12795 14984 12801
rect 14936 12764 14964 12795
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 15746 12832 15752 12844
rect 15344 12804 15752 12832
rect 15344 12792 15350 12804
rect 15746 12792 15752 12804
rect 15804 12792 15810 12844
rect 17126 12792 17132 12844
rect 17184 12792 17190 12844
rect 17236 12832 17264 12872
rect 17310 12860 17316 12912
rect 17368 12860 17374 12912
rect 17402 12860 17408 12912
rect 17460 12860 17466 12912
rect 17494 12832 17500 12844
rect 17552 12841 17558 12844
rect 18064 12841 18092 12940
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 18874 12928 18880 12980
rect 18932 12968 18938 12980
rect 18932 12940 20024 12968
rect 18932 12928 18938 12940
rect 18322 12860 18328 12912
rect 18380 12900 18386 12912
rect 19610 12900 19616 12912
rect 18380 12872 19616 12900
rect 18380 12860 18386 12872
rect 19610 12860 19616 12872
rect 19668 12900 19674 12912
rect 19797 12903 19855 12909
rect 19797 12900 19809 12903
rect 19668 12872 19809 12900
rect 19668 12860 19674 12872
rect 19797 12869 19809 12872
rect 19843 12869 19855 12903
rect 19797 12863 19855 12869
rect 18506 12841 18512 12844
rect 17236 12804 17500 12832
rect 17494 12792 17500 12804
rect 17552 12795 17560 12841
rect 18049 12835 18107 12841
rect 18049 12832 18061 12835
rect 17604 12804 18061 12832
rect 17552 12792 17558 12795
rect 13096 12736 14964 12764
rect 16022 12724 16028 12776
rect 16080 12764 16086 12776
rect 17604 12764 17632 12804
rect 18049 12801 18061 12804
rect 18095 12801 18107 12835
rect 18233 12835 18291 12841
rect 18233 12832 18245 12835
rect 18049 12795 18107 12801
rect 18156 12804 18245 12832
rect 16080 12736 17632 12764
rect 16080 12724 16086 12736
rect 17954 12724 17960 12776
rect 18012 12764 18018 12776
rect 18156 12764 18184 12804
rect 18233 12801 18245 12804
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 18469 12835 18512 12841
rect 18469 12801 18481 12835
rect 18469 12795 18512 12801
rect 18506 12792 18512 12795
rect 18564 12792 18570 12844
rect 18782 12792 18788 12844
rect 18840 12792 18846 12844
rect 19242 12841 19248 12844
rect 18969 12835 19027 12841
rect 18969 12801 18981 12835
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 19061 12835 19119 12841
rect 19061 12801 19073 12835
rect 19107 12801 19119 12835
rect 19061 12795 19119 12801
rect 19205 12835 19248 12841
rect 19205 12801 19217 12835
rect 19205 12795 19248 12801
rect 18984 12764 19012 12795
rect 18012 12736 18184 12764
rect 18248 12736 19012 12764
rect 18012 12724 18018 12736
rect 13446 12696 13452 12708
rect 11624 12668 13452 12696
rect 9640 12656 9646 12668
rect 13446 12656 13452 12668
rect 13504 12656 13510 12708
rect 14090 12656 14096 12708
rect 14148 12696 14154 12708
rect 15105 12699 15163 12705
rect 14148 12668 14504 12696
rect 14148 12656 14154 12668
rect 6546 12628 6552 12640
rect 5368 12600 6552 12628
rect 4580 12588 4586 12600
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 7006 12588 7012 12640
rect 7064 12628 7070 12640
rect 10502 12628 10508 12640
rect 7064 12600 10508 12628
rect 7064 12588 7070 12600
rect 10502 12588 10508 12600
rect 10560 12588 10566 12640
rect 10597 12631 10655 12637
rect 10597 12597 10609 12631
rect 10643 12628 10655 12631
rect 10778 12628 10784 12640
rect 10643 12600 10784 12628
rect 10643 12597 10655 12600
rect 10597 12591 10655 12597
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 14182 12588 14188 12640
rect 14240 12628 14246 12640
rect 14369 12631 14427 12637
rect 14369 12628 14381 12631
rect 14240 12600 14381 12628
rect 14240 12588 14246 12600
rect 14369 12597 14381 12600
rect 14415 12597 14427 12631
rect 14476 12628 14504 12668
rect 15105 12665 15117 12699
rect 15151 12696 15163 12699
rect 17218 12696 17224 12708
rect 15151 12668 17224 12696
rect 15151 12665 15163 12668
rect 15105 12659 15163 12665
rect 17218 12656 17224 12668
rect 17276 12656 17282 12708
rect 17678 12656 17684 12708
rect 17736 12656 17742 12708
rect 18248 12628 18276 12736
rect 18690 12656 18696 12708
rect 18748 12696 18754 12708
rect 19076 12696 19104 12795
rect 19242 12792 19248 12795
rect 19300 12792 19306 12844
rect 19518 12792 19524 12844
rect 19576 12792 19582 12844
rect 19705 12835 19763 12841
rect 19705 12801 19717 12835
rect 19751 12801 19763 12835
rect 19705 12795 19763 12801
rect 19720 12764 19748 12795
rect 19886 12792 19892 12844
rect 19944 12792 19950 12844
rect 19306 12736 19748 12764
rect 19996 12764 20024 12940
rect 20070 12928 20076 12980
rect 20128 12928 20134 12980
rect 23014 12928 23020 12980
rect 23072 12928 23078 12980
rect 23198 12928 23204 12980
rect 23256 12968 23262 12980
rect 23569 12971 23627 12977
rect 23256 12940 23520 12968
rect 23256 12928 23262 12940
rect 20714 12860 20720 12912
rect 20772 12900 20778 12912
rect 23492 12900 23520 12940
rect 23569 12937 23581 12971
rect 23615 12968 23627 12971
rect 23750 12968 23756 12980
rect 23615 12940 23756 12968
rect 23615 12937 23627 12940
rect 23569 12931 23627 12937
rect 23750 12928 23756 12940
rect 23808 12928 23814 12980
rect 24486 12928 24492 12980
rect 24544 12968 24550 12980
rect 26053 12971 26111 12977
rect 24544 12940 25912 12968
rect 24544 12928 24550 12940
rect 25884 12900 25912 12940
rect 26053 12937 26065 12971
rect 26099 12968 26111 12971
rect 26142 12968 26148 12980
rect 26099 12940 26148 12968
rect 26099 12937 26111 12940
rect 26053 12931 26111 12937
rect 26142 12928 26148 12940
rect 26200 12928 26206 12980
rect 31478 12928 31484 12980
rect 31536 12928 31542 12980
rect 29454 12900 29460 12912
rect 20772 12872 23336 12900
rect 23492 12872 24072 12900
rect 25884 12872 29460 12900
rect 20772 12860 20778 12872
rect 23198 12792 23204 12844
rect 23256 12792 23262 12844
rect 23308 12841 23336 12872
rect 23293 12835 23351 12841
rect 23293 12801 23305 12835
rect 23339 12801 23351 12835
rect 23293 12795 23351 12801
rect 23474 12792 23480 12844
rect 23532 12792 23538 12844
rect 23842 12792 23848 12844
rect 23900 12792 23906 12844
rect 23934 12792 23940 12844
rect 23992 12792 23998 12844
rect 19996 12736 23244 12764
rect 19306 12708 19334 12736
rect 18748 12668 19104 12696
rect 18748 12656 18754 12668
rect 19242 12656 19248 12708
rect 19300 12668 19334 12708
rect 23216 12696 23244 12736
rect 23492 12696 23520 12792
rect 24044 12764 24072 12872
rect 29454 12860 29460 12872
rect 29512 12860 29518 12912
rect 29730 12860 29736 12912
rect 29788 12900 29794 12912
rect 30282 12900 30288 12912
rect 29788 12872 30288 12900
rect 29788 12860 29794 12872
rect 30282 12860 30288 12872
rect 30340 12900 30346 12912
rect 31021 12903 31079 12909
rect 31021 12900 31033 12903
rect 30340 12872 31033 12900
rect 30340 12860 30346 12872
rect 31021 12869 31033 12872
rect 31067 12900 31079 12903
rect 31110 12900 31116 12912
rect 31067 12872 31116 12900
rect 31067 12869 31079 12872
rect 31021 12863 31079 12869
rect 31110 12860 31116 12872
rect 31168 12860 31174 12912
rect 25406 12792 25412 12844
rect 25464 12832 25470 12844
rect 25682 12832 25688 12844
rect 25464 12804 25688 12832
rect 25464 12792 25470 12804
rect 25682 12792 25688 12804
rect 25740 12792 25746 12844
rect 25869 12835 25927 12841
rect 25869 12801 25881 12835
rect 25915 12801 25927 12835
rect 25869 12795 25927 12801
rect 25774 12764 25780 12776
rect 24044 12736 25780 12764
rect 25774 12724 25780 12736
rect 25832 12764 25838 12776
rect 25884 12764 25912 12795
rect 30926 12792 30932 12844
rect 30984 12832 30990 12844
rect 31297 12835 31355 12841
rect 31297 12832 31309 12835
rect 30984 12804 31309 12832
rect 30984 12792 30990 12804
rect 31297 12801 31309 12804
rect 31343 12801 31355 12835
rect 31297 12795 31355 12801
rect 25832 12736 25912 12764
rect 25832 12724 25838 12736
rect 26050 12724 26056 12776
rect 26108 12764 26114 12776
rect 31113 12767 31171 12773
rect 31113 12764 31125 12767
rect 26108 12736 31125 12764
rect 26108 12724 26114 12736
rect 31113 12733 31125 12736
rect 31159 12764 31171 12767
rect 31662 12764 31668 12776
rect 31159 12736 31668 12764
rect 31159 12733 31171 12736
rect 31113 12727 31171 12733
rect 31662 12724 31668 12736
rect 31720 12724 31726 12776
rect 25498 12696 25504 12708
rect 23216 12668 23520 12696
rect 23860 12668 25504 12696
rect 19300 12656 19306 12668
rect 14476 12600 18276 12628
rect 18601 12631 18659 12637
rect 14369 12591 14427 12597
rect 18601 12597 18613 12631
rect 18647 12628 18659 12631
rect 18874 12628 18880 12640
rect 18647 12600 18880 12628
rect 18647 12597 18659 12600
rect 18601 12591 18659 12597
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 19337 12631 19395 12637
rect 19337 12597 19349 12631
rect 19383 12628 19395 12631
rect 20714 12628 20720 12640
rect 19383 12600 20720 12628
rect 19383 12597 19395 12600
rect 19337 12591 19395 12597
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 23198 12588 23204 12640
rect 23256 12628 23262 12640
rect 23860 12628 23888 12668
rect 25498 12656 25504 12668
rect 25556 12696 25562 12708
rect 25556 12668 25728 12696
rect 25556 12656 25562 12668
rect 23256 12600 23888 12628
rect 23937 12631 23995 12637
rect 23256 12588 23262 12600
rect 23937 12597 23949 12631
rect 23983 12628 23995 12631
rect 24394 12628 24400 12640
rect 23983 12600 24400 12628
rect 23983 12597 23995 12600
rect 23937 12591 23995 12597
rect 24394 12588 24400 12600
rect 24452 12588 24458 12640
rect 25700 12637 25728 12668
rect 25685 12631 25743 12637
rect 25685 12597 25697 12631
rect 25731 12597 25743 12631
rect 25685 12591 25743 12597
rect 31018 12588 31024 12640
rect 31076 12588 31082 12640
rect 1104 12538 44896 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 44896 12538
rect 1104 12464 44896 12486
rect 1578 12384 1584 12436
rect 1636 12384 1642 12436
rect 1857 12427 1915 12433
rect 1857 12393 1869 12427
rect 1903 12424 1915 12427
rect 3050 12424 3056 12436
rect 1903 12396 3056 12424
rect 1903 12393 1915 12396
rect 1857 12387 1915 12393
rect 3050 12384 3056 12396
rect 3108 12384 3114 12436
rect 3970 12384 3976 12436
rect 4028 12424 4034 12436
rect 5537 12427 5595 12433
rect 4028 12396 4844 12424
rect 4028 12384 4034 12396
rect 4816 12368 4844 12396
rect 5537 12393 5549 12427
rect 5583 12424 5595 12427
rect 6270 12424 6276 12436
rect 5583 12396 6276 12424
rect 5583 12393 5595 12396
rect 5537 12387 5595 12393
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 9766 12384 9772 12436
rect 9824 12424 9830 12436
rect 10229 12427 10287 12433
rect 10229 12424 10241 12427
rect 9824 12396 10241 12424
rect 9824 12384 9830 12396
rect 10229 12393 10241 12396
rect 10275 12393 10287 12427
rect 10229 12387 10287 12393
rect 12250 12384 12256 12436
rect 12308 12424 12314 12436
rect 12437 12427 12495 12433
rect 12437 12424 12449 12427
rect 12308 12396 12449 12424
rect 12308 12384 12314 12396
rect 12437 12393 12449 12396
rect 12483 12393 12495 12427
rect 12437 12387 12495 12393
rect 14366 12384 14372 12436
rect 14424 12384 14430 12436
rect 15010 12384 15016 12436
rect 15068 12424 15074 12436
rect 17586 12424 17592 12436
rect 15068 12396 17592 12424
rect 15068 12384 15074 12396
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 17681 12427 17739 12433
rect 17681 12393 17693 12427
rect 17727 12424 17739 12427
rect 30282 12424 30288 12436
rect 17727 12396 30288 12424
rect 17727 12393 17739 12396
rect 17681 12387 17739 12393
rect 30282 12384 30288 12396
rect 30340 12384 30346 12436
rect 4709 12359 4767 12365
rect 4709 12325 4721 12359
rect 4755 12325 4767 12359
rect 4709 12319 4767 12325
rect 4724 12288 4752 12319
rect 4798 12316 4804 12368
rect 4856 12356 4862 12368
rect 5718 12356 5724 12368
rect 4856 12328 5724 12356
rect 4856 12316 4862 12328
rect 5718 12316 5724 12328
rect 5776 12316 5782 12368
rect 6362 12316 6368 12368
rect 6420 12356 6426 12368
rect 6420 12328 8248 12356
rect 6420 12316 6426 12328
rect 6181 12291 6239 12297
rect 6181 12288 6193 12291
rect 4724 12260 6193 12288
rect 6181 12257 6193 12260
rect 6227 12288 6239 12291
rect 6546 12288 6552 12300
rect 6227 12260 6552 12288
rect 6227 12257 6239 12260
rect 6181 12251 6239 12257
rect 6546 12248 6552 12260
rect 6604 12248 6610 12300
rect 7742 12248 7748 12300
rect 7800 12248 7806 12300
rect 1394 12180 1400 12232
rect 1452 12180 1458 12232
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12189 1731 12223
rect 1673 12183 1731 12189
rect 842 12112 848 12164
rect 900 12152 906 12164
rect 1688 12152 1716 12183
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 5169 12223 5227 12229
rect 4120 12192 4844 12220
rect 4120 12180 4126 12192
rect 900 12124 1716 12152
rect 900 12112 906 12124
rect 4706 12112 4712 12164
rect 4764 12112 4770 12164
rect 4816 12152 4844 12192
rect 5169 12189 5181 12223
rect 5215 12220 5227 12223
rect 5442 12220 5448 12232
rect 5215 12192 5448 12220
rect 5215 12189 5227 12192
rect 5169 12183 5227 12189
rect 5442 12180 5448 12192
rect 5500 12220 5506 12232
rect 5813 12223 5871 12229
rect 5813 12220 5825 12223
rect 5500 12192 5825 12220
rect 5500 12180 5506 12192
rect 5813 12189 5825 12192
rect 5859 12189 5871 12223
rect 5813 12183 5871 12189
rect 5902 12180 5908 12232
rect 5960 12180 5966 12232
rect 7282 12180 7288 12232
rect 7340 12220 7346 12232
rect 7653 12223 7711 12229
rect 7653 12220 7665 12223
rect 7340 12192 7665 12220
rect 7340 12180 7346 12192
rect 7653 12189 7665 12192
rect 7699 12189 7711 12223
rect 7653 12183 7711 12189
rect 5718 12161 5724 12164
rect 5261 12155 5319 12161
rect 5261 12152 5273 12155
rect 4816 12124 5273 12152
rect 5261 12121 5273 12124
rect 5307 12152 5319 12155
rect 5696 12155 5724 12161
rect 5307 12124 5580 12152
rect 5307 12121 5319 12124
rect 5261 12115 5319 12121
rect 5442 12044 5448 12096
rect 5500 12044 5506 12096
rect 5552 12084 5580 12124
rect 5696 12121 5708 12155
rect 5696 12115 5724 12121
rect 5718 12112 5724 12115
rect 5776 12112 5782 12164
rect 5920 12084 5948 12180
rect 7668 12152 7696 12183
rect 8018 12180 8024 12232
rect 8076 12180 8082 12232
rect 8220 12229 8248 12328
rect 8754 12316 8760 12368
rect 8812 12356 8818 12368
rect 8812 12328 16574 12356
rect 8812 12316 8818 12328
rect 8662 12248 8668 12300
rect 8720 12248 8726 12300
rect 12158 12248 12164 12300
rect 12216 12288 12222 12300
rect 12216 12260 12940 12288
rect 12216 12248 12222 12260
rect 8205 12223 8263 12229
rect 8205 12189 8217 12223
rect 8251 12220 8263 12223
rect 8251 12192 10088 12220
rect 8251 12189 8263 12192
rect 8205 12183 8263 12189
rect 8294 12152 8300 12164
rect 7668 12124 8300 12152
rect 8294 12112 8300 12124
rect 8352 12112 8358 12164
rect 5552 12056 5948 12084
rect 10060 12084 10088 12192
rect 10594 12180 10600 12232
rect 10652 12220 10658 12232
rect 12345 12223 12403 12229
rect 12345 12220 12357 12223
rect 10652 12192 12357 12220
rect 10652 12180 10658 12192
rect 12345 12189 12357 12192
rect 12391 12189 12403 12223
rect 12345 12183 12403 12189
rect 12912 12164 12940 12260
rect 12986 12248 12992 12300
rect 13044 12288 13050 12300
rect 13044 12260 14320 12288
rect 13044 12248 13050 12260
rect 14185 12223 14243 12229
rect 14185 12220 14197 12223
rect 13004 12192 14197 12220
rect 10502 12112 10508 12164
rect 10560 12112 10566 12164
rect 11054 12112 11060 12164
rect 11112 12152 11118 12164
rect 12713 12155 12771 12161
rect 12713 12152 12725 12155
rect 11112 12124 12725 12152
rect 11112 12112 11118 12124
rect 12713 12121 12725 12124
rect 12759 12121 12771 12155
rect 12713 12115 12771 12121
rect 12894 12112 12900 12164
rect 12952 12112 12958 12164
rect 11238 12084 11244 12096
rect 10060 12056 11244 12084
rect 11238 12044 11244 12056
rect 11296 12084 11302 12096
rect 13004 12084 13032 12192
rect 14185 12189 14197 12192
rect 14231 12189 14243 12223
rect 14292 12220 14320 12260
rect 14734 12248 14740 12300
rect 14792 12248 14798 12300
rect 16546 12288 16574 12328
rect 17034 12316 17040 12368
rect 17092 12356 17098 12368
rect 18230 12356 18236 12368
rect 17092 12328 18236 12356
rect 17092 12316 17098 12328
rect 18230 12316 18236 12328
rect 18288 12316 18294 12368
rect 19794 12316 19800 12368
rect 19852 12316 19858 12368
rect 27706 12288 27712 12300
rect 14844 12260 15424 12288
rect 16546 12260 27712 12288
rect 14844 12220 14872 12260
rect 14292 12192 14872 12220
rect 14185 12183 14243 12189
rect 14918 12180 14924 12232
rect 14976 12220 14982 12232
rect 15105 12223 15163 12229
rect 15105 12220 15117 12223
rect 14976 12192 15117 12220
rect 14976 12180 14982 12192
rect 15105 12189 15117 12192
rect 15151 12189 15163 12223
rect 15105 12183 15163 12189
rect 15194 12180 15200 12232
rect 15252 12220 15258 12232
rect 15289 12223 15347 12229
rect 15289 12220 15301 12223
rect 15252 12192 15301 12220
rect 15252 12180 15258 12192
rect 15289 12189 15301 12192
rect 15335 12189 15347 12223
rect 15396 12220 15424 12260
rect 27706 12248 27712 12260
rect 27764 12248 27770 12300
rect 17129 12223 17187 12229
rect 17129 12220 17141 12223
rect 15396 12192 17141 12220
rect 15289 12183 15347 12189
rect 17129 12189 17141 12192
rect 17175 12189 17187 12223
rect 17129 12183 17187 12189
rect 13078 12112 13084 12164
rect 13136 12152 13142 12164
rect 16942 12152 16948 12164
rect 13136 12124 16948 12152
rect 13136 12112 13142 12124
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 11296 12056 13032 12084
rect 14829 12087 14887 12093
rect 11296 12044 11302 12056
rect 14829 12053 14841 12087
rect 14875 12084 14887 12087
rect 17034 12084 17040 12096
rect 14875 12056 17040 12084
rect 14875 12053 14887 12056
rect 14829 12047 14887 12053
rect 17034 12044 17040 12056
rect 17092 12044 17098 12096
rect 17144 12084 17172 12183
rect 17310 12180 17316 12232
rect 17368 12180 17374 12232
rect 17494 12180 17500 12232
rect 17552 12229 17558 12232
rect 17552 12220 17560 12229
rect 17552 12192 17597 12220
rect 17552 12183 17560 12192
rect 17552 12180 17558 12183
rect 17678 12180 17684 12232
rect 17736 12220 17742 12232
rect 19242 12220 19248 12232
rect 17736 12192 19248 12220
rect 17736 12180 17742 12192
rect 19242 12180 19248 12192
rect 19300 12180 19306 12232
rect 19518 12220 19524 12232
rect 19352 12192 19524 12220
rect 17402 12112 17408 12164
rect 17460 12152 17466 12164
rect 19352 12152 19380 12192
rect 19518 12180 19524 12192
rect 19576 12180 19582 12232
rect 19610 12180 19616 12232
rect 19668 12229 19674 12232
rect 19668 12220 19676 12229
rect 19668 12192 19713 12220
rect 19668 12183 19676 12192
rect 19668 12180 19674 12183
rect 17460 12124 19380 12152
rect 19429 12155 19487 12161
rect 17460 12112 17466 12124
rect 19429 12121 19441 12155
rect 19475 12152 19487 12155
rect 19886 12152 19892 12164
rect 19475 12124 19892 12152
rect 19475 12121 19487 12124
rect 19429 12115 19487 12121
rect 19444 12084 19472 12115
rect 19886 12112 19892 12124
rect 19944 12112 19950 12164
rect 17144 12056 19472 12084
rect 1104 11994 44896 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 44896 11994
rect 1104 11920 44896 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 2774 11880 2780 11892
rect 1627 11852 2780 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 2774 11840 2780 11852
rect 2832 11840 2838 11892
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 15746 11880 15752 11892
rect 8352 11852 15752 11880
rect 8352 11840 8358 11852
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 15838 11840 15844 11892
rect 15896 11880 15902 11892
rect 23842 11880 23848 11892
rect 15896 11852 23848 11880
rect 15896 11840 15902 11852
rect 23842 11840 23848 11852
rect 23900 11840 23906 11892
rect 5442 11772 5448 11824
rect 5500 11812 5506 11824
rect 9950 11812 9956 11824
rect 5500 11784 9956 11812
rect 5500 11772 5506 11784
rect 9950 11772 9956 11784
rect 10008 11772 10014 11824
rect 842 11704 848 11756
rect 900 11744 906 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 900 11716 1409 11744
rect 900 11704 906 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 10502 11704 10508 11756
rect 10560 11744 10566 11756
rect 13170 11744 13176 11756
rect 10560 11716 13176 11744
rect 10560 11704 10566 11716
rect 13170 11704 13176 11716
rect 13228 11744 13234 11756
rect 17402 11744 17408 11756
rect 13228 11716 17408 11744
rect 13228 11704 13234 11716
rect 17402 11704 17408 11716
rect 17460 11704 17466 11756
rect 7926 11636 7932 11688
rect 7984 11676 7990 11688
rect 15838 11676 15844 11688
rect 7984 11648 15844 11676
rect 7984 11636 7990 11648
rect 15838 11636 15844 11648
rect 15896 11636 15902 11688
rect 1104 11450 44896 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 44896 11450
rect 1104 11376 44896 11398
rect 1104 10906 44896 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 44896 10906
rect 1104 10832 44896 10854
rect 1104 10362 44896 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 44896 10362
rect 1104 10288 44896 10310
rect 1104 9818 44896 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 44896 9818
rect 1104 9744 44896 9766
rect 1104 9274 44896 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 44896 9274
rect 1104 9200 44896 9222
rect 1104 8730 44896 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 44896 8730
rect 1104 8656 44896 8678
rect 1104 8186 44896 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 44896 8186
rect 1104 8112 44896 8134
rect 1104 7642 44896 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 44896 7642
rect 1104 7568 44896 7590
rect 1104 7098 44896 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 44896 7098
rect 1104 7024 44896 7046
rect 1104 6554 44896 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 44896 6554
rect 1104 6480 44896 6502
rect 1104 6010 44896 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 44896 6010
rect 1104 5936 44896 5958
rect 1104 5466 44896 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 44896 5466
rect 1104 5392 44896 5414
rect 1104 4922 44896 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 44896 4922
rect 1104 4848 44896 4870
rect 1104 4378 44896 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 44896 4378
rect 1104 4304 44896 4326
rect 1104 3834 44896 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 44896 3834
rect 1104 3760 44896 3782
rect 1104 3290 44896 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 44896 3290
rect 1104 3216 44896 3238
rect 1104 2746 44896 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 44896 2746
rect 1104 2672 44896 2694
rect 1104 2202 44896 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 44896 2202
rect 1104 2128 44896 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 21916 37408 21968 37460
rect 22560 37408 22612 37460
rect 23204 37408 23256 37460
rect 25136 37408 25188 37460
rect 25780 37408 25832 37460
rect 27712 37408 27764 37460
rect 29644 37408 29696 37460
rect 31576 37408 31628 37460
rect 29000 37340 29052 37392
rect 22376 37179 22428 37188
rect 22376 37145 22385 37179
rect 22385 37145 22419 37179
rect 22419 37145 22428 37179
rect 22376 37136 22428 37145
rect 23388 37136 23440 37188
rect 23664 37179 23716 37188
rect 23664 37145 23673 37179
rect 23673 37145 23707 37179
rect 23707 37145 23716 37179
rect 23664 37136 23716 37145
rect 25596 37179 25648 37188
rect 25596 37145 25605 37179
rect 25605 37145 25639 37179
rect 25639 37145 25648 37179
rect 25596 37136 25648 37145
rect 27068 37136 27120 37188
rect 28172 37179 28224 37188
rect 28172 37145 28181 37179
rect 28181 37145 28215 37179
rect 28215 37145 28224 37179
rect 28172 37136 28224 37145
rect 29644 37179 29696 37188
rect 29644 37145 29653 37179
rect 29653 37145 29687 37179
rect 29687 37145 29696 37179
rect 29644 37136 29696 37145
rect 30472 37179 30524 37188
rect 30472 37145 30481 37179
rect 30481 37145 30515 37179
rect 30515 37145 30524 37179
rect 30472 37136 30524 37145
rect 32220 37179 32272 37188
rect 32220 37145 32229 37179
rect 32229 37145 32263 37179
rect 32263 37145 32272 37179
rect 32220 37136 32272 37145
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 22376 35683 22428 35692
rect 22376 35649 22385 35683
rect 22385 35649 22419 35683
rect 22419 35649 22428 35683
rect 22376 35640 22428 35649
rect 22652 35436 22704 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 22284 35232 22336 35284
rect 23664 35096 23716 35148
rect 23204 35071 23256 35080
rect 23204 35037 23213 35071
rect 23213 35037 23247 35071
rect 23247 35037 23256 35071
rect 23204 35028 23256 35037
rect 23296 34960 23348 35012
rect 23572 34960 23624 35012
rect 26976 34960 27028 35012
rect 24124 34892 24176 34944
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 14372 34688 14424 34740
rect 23572 34688 23624 34740
rect 23664 34731 23716 34740
rect 23664 34697 23673 34731
rect 23673 34697 23707 34731
rect 23707 34697 23716 34731
rect 23664 34688 23716 34697
rect 25596 34688 25648 34740
rect 28172 34688 28224 34740
rect 22192 34552 22244 34604
rect 23204 34620 23256 34672
rect 23664 34552 23716 34604
rect 24308 34595 24360 34604
rect 24308 34561 24342 34595
rect 24342 34561 24360 34595
rect 24308 34552 24360 34561
rect 25596 34552 25648 34604
rect 27528 34620 27580 34672
rect 27712 34552 27764 34604
rect 25504 34391 25556 34400
rect 25504 34357 25513 34391
rect 25513 34357 25547 34391
rect 25547 34357 25556 34391
rect 25504 34348 25556 34357
rect 28448 34391 28500 34400
rect 28448 34357 28457 34391
rect 28457 34357 28491 34391
rect 28491 34357 28500 34391
rect 28448 34348 28500 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 16304 34008 16356 34060
rect 22836 34144 22888 34196
rect 23112 34144 23164 34196
rect 23204 34144 23256 34196
rect 23388 34144 23440 34196
rect 23664 34187 23716 34196
rect 23664 34153 23673 34187
rect 23673 34153 23707 34187
rect 23707 34153 23716 34187
rect 23664 34144 23716 34153
rect 24124 34187 24176 34196
rect 24124 34153 24133 34187
rect 24133 34153 24167 34187
rect 24167 34153 24176 34187
rect 24124 34144 24176 34153
rect 24308 34144 24360 34196
rect 27068 34187 27120 34196
rect 27068 34153 27077 34187
rect 27077 34153 27111 34187
rect 27111 34153 27120 34187
rect 27068 34144 27120 34153
rect 22192 34051 22244 34060
rect 22192 34017 22201 34051
rect 22201 34017 22235 34051
rect 22235 34017 22244 34051
rect 22192 34008 22244 34017
rect 21640 33983 21692 33992
rect 21640 33949 21649 33983
rect 21649 33949 21683 33983
rect 21683 33949 21692 33983
rect 21640 33940 21692 33949
rect 21916 33983 21968 33992
rect 21916 33949 21925 33983
rect 21925 33949 21959 33983
rect 21959 33949 21968 33983
rect 21916 33940 21968 33949
rect 23388 33940 23440 33992
rect 29644 34008 29696 34060
rect 23480 33872 23532 33924
rect 22744 33804 22796 33856
rect 24584 33983 24636 33992
rect 24584 33949 24593 33983
rect 24593 33949 24627 33983
rect 24627 33949 24636 33983
rect 24584 33940 24636 33949
rect 24768 33983 24820 33992
rect 24768 33949 24777 33983
rect 24777 33949 24811 33983
rect 24811 33949 24820 33983
rect 24768 33940 24820 33949
rect 25504 33940 25556 33992
rect 27528 33983 27580 33992
rect 27528 33949 27537 33983
rect 27537 33949 27571 33983
rect 27571 33949 27580 33983
rect 27528 33940 27580 33949
rect 26148 33872 26200 33924
rect 27804 33915 27856 33924
rect 27804 33881 27838 33915
rect 27838 33881 27856 33915
rect 27804 33872 27856 33881
rect 26608 33804 26660 33856
rect 29000 33804 29052 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 17776 33600 17828 33652
rect 23112 33600 23164 33652
rect 23296 33643 23348 33652
rect 23296 33609 23305 33643
rect 23305 33609 23339 33643
rect 23339 33609 23348 33643
rect 23296 33600 23348 33609
rect 23388 33643 23440 33652
rect 23388 33609 23397 33643
rect 23397 33609 23431 33643
rect 23431 33609 23440 33643
rect 23388 33600 23440 33609
rect 26148 33643 26200 33652
rect 26148 33609 26157 33643
rect 26157 33609 26191 33643
rect 26191 33609 26200 33643
rect 26148 33600 26200 33609
rect 27712 33643 27764 33652
rect 27712 33609 27721 33643
rect 27721 33609 27755 33643
rect 27755 33609 27764 33643
rect 27712 33600 27764 33609
rect 30472 33600 30524 33652
rect 22652 33507 22704 33516
rect 22652 33473 22661 33507
rect 22661 33473 22695 33507
rect 22695 33473 22704 33507
rect 22652 33464 22704 33473
rect 24584 33532 24636 33584
rect 21640 33396 21692 33448
rect 23204 33464 23256 33516
rect 27068 33464 27120 33516
rect 27896 33507 27948 33516
rect 27896 33473 27905 33507
rect 27905 33473 27939 33507
rect 27939 33473 27948 33507
rect 27896 33464 27948 33473
rect 27988 33507 28040 33516
rect 27988 33473 27997 33507
rect 27997 33473 28031 33507
rect 28031 33473 28040 33507
rect 27988 33464 28040 33473
rect 28264 33507 28316 33516
rect 21916 33328 21968 33380
rect 22744 33328 22796 33380
rect 22928 33439 22980 33448
rect 22928 33405 22937 33439
rect 22937 33405 22971 33439
rect 22971 33405 22980 33439
rect 22928 33396 22980 33405
rect 26516 33439 26568 33448
rect 26516 33405 26525 33439
rect 26525 33405 26559 33439
rect 26559 33405 26568 33439
rect 26516 33396 26568 33405
rect 26608 33439 26660 33448
rect 26608 33405 26617 33439
rect 26617 33405 26651 33439
rect 26651 33405 26660 33439
rect 28264 33473 28273 33507
rect 28273 33473 28307 33507
rect 28307 33473 28316 33507
rect 28264 33464 28316 33473
rect 29552 33464 29604 33516
rect 30472 33464 30524 33516
rect 26608 33396 26660 33405
rect 28448 33396 28500 33448
rect 30656 33396 30708 33448
rect 23572 33328 23624 33380
rect 27436 33328 27488 33380
rect 30196 33260 30248 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 27804 33056 27856 33108
rect 29000 33056 29052 33108
rect 29552 33099 29604 33108
rect 29552 33065 29561 33099
rect 29561 33065 29595 33099
rect 29595 33065 29604 33099
rect 29552 33056 29604 33065
rect 21824 32988 21876 33040
rect 20720 32920 20772 32972
rect 23388 32920 23440 32972
rect 18420 32852 18472 32904
rect 21916 32852 21968 32904
rect 27804 32852 27856 32904
rect 27896 32895 27948 32904
rect 27896 32861 27905 32895
rect 27905 32861 27939 32895
rect 27939 32861 27948 32895
rect 27896 32852 27948 32861
rect 27620 32784 27672 32836
rect 28264 32988 28316 33040
rect 31576 33056 31628 33108
rect 32220 33056 32272 33108
rect 28264 32895 28316 32904
rect 28264 32861 28273 32895
rect 28273 32861 28307 32895
rect 28307 32861 28316 32895
rect 28264 32852 28316 32861
rect 29736 32895 29788 32904
rect 29736 32861 29745 32895
rect 29745 32861 29779 32895
rect 29779 32861 29788 32895
rect 29736 32852 29788 32861
rect 29828 32895 29880 32904
rect 29828 32861 29837 32895
rect 29837 32861 29871 32895
rect 29871 32861 29880 32895
rect 29828 32852 29880 32861
rect 29920 32895 29972 32904
rect 29920 32861 29929 32895
rect 29929 32861 29963 32895
rect 29963 32861 29972 32895
rect 29920 32852 29972 32861
rect 30196 32895 30248 32904
rect 30196 32861 30205 32895
rect 30205 32861 30239 32895
rect 30239 32861 30248 32895
rect 30196 32852 30248 32861
rect 30656 32895 30708 32904
rect 30656 32861 30665 32895
rect 30665 32861 30699 32895
rect 30699 32861 30708 32895
rect 30656 32852 30708 32861
rect 30288 32784 30340 32836
rect 31024 32784 31076 32836
rect 36084 32784 36136 32836
rect 13728 32716 13780 32768
rect 22008 32716 22060 32768
rect 26148 32716 26200 32768
rect 27896 32716 27948 32768
rect 29736 32716 29788 32768
rect 32128 32759 32180 32768
rect 32128 32725 32137 32759
rect 32137 32725 32171 32759
rect 32171 32725 32180 32759
rect 32128 32716 32180 32725
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 14832 32512 14884 32564
rect 12348 32444 12400 32496
rect 19340 32512 19392 32564
rect 23112 32512 23164 32564
rect 23480 32555 23532 32564
rect 23480 32521 23489 32555
rect 23489 32521 23523 32555
rect 23523 32521 23532 32555
rect 23480 32512 23532 32521
rect 23572 32555 23624 32564
rect 23572 32521 23581 32555
rect 23581 32521 23615 32555
rect 23615 32521 23624 32555
rect 23572 32512 23624 32521
rect 29828 32512 29880 32564
rect 31024 32555 31076 32564
rect 31024 32521 31033 32555
rect 31033 32521 31067 32555
rect 31067 32521 31076 32555
rect 31024 32512 31076 32521
rect 11428 32376 11480 32428
rect 15844 32419 15896 32428
rect 15844 32385 15853 32419
rect 15853 32385 15887 32419
rect 15887 32385 15896 32419
rect 15844 32376 15896 32385
rect 19064 32376 19116 32428
rect 19432 32419 19484 32428
rect 19432 32385 19441 32419
rect 19441 32385 19475 32419
rect 19475 32385 19484 32419
rect 19432 32376 19484 32385
rect 13544 32308 13596 32360
rect 16028 32351 16080 32360
rect 16028 32317 16037 32351
rect 16037 32317 16071 32351
rect 16071 32317 16080 32351
rect 16028 32308 16080 32317
rect 16120 32308 16172 32360
rect 20720 32308 20772 32360
rect 21824 32419 21876 32428
rect 21824 32385 21833 32419
rect 21833 32385 21867 32419
rect 21867 32385 21876 32419
rect 21824 32376 21876 32385
rect 13176 32215 13228 32224
rect 13176 32181 13185 32215
rect 13185 32181 13219 32215
rect 13219 32181 13228 32215
rect 13176 32172 13228 32181
rect 13636 32215 13688 32224
rect 13636 32181 13645 32215
rect 13645 32181 13679 32215
rect 13679 32181 13688 32215
rect 13636 32172 13688 32181
rect 15936 32215 15988 32224
rect 15936 32181 15945 32215
rect 15945 32181 15979 32215
rect 15979 32181 15988 32215
rect 15936 32172 15988 32181
rect 19524 32240 19576 32292
rect 23020 32444 23072 32496
rect 23296 32419 23348 32428
rect 23296 32385 23305 32419
rect 23305 32385 23339 32419
rect 23339 32385 23348 32419
rect 23296 32376 23348 32385
rect 31392 32444 31444 32496
rect 37464 32512 37516 32564
rect 23020 32240 23072 32292
rect 23756 32308 23808 32360
rect 24032 32308 24084 32360
rect 26608 32376 26660 32428
rect 28356 32419 28408 32428
rect 28356 32385 28365 32419
rect 28365 32385 28399 32419
rect 28399 32385 28408 32419
rect 28356 32376 28408 32385
rect 28540 32376 28592 32428
rect 26240 32351 26292 32360
rect 26240 32317 26249 32351
rect 26249 32317 26283 32351
rect 26283 32317 26292 32351
rect 26240 32308 26292 32317
rect 27252 32308 27304 32360
rect 29000 32376 29052 32428
rect 29644 32376 29696 32428
rect 25688 32240 25740 32292
rect 29736 32308 29788 32360
rect 32128 32376 32180 32428
rect 30380 32308 30432 32360
rect 31576 32308 31628 32360
rect 37096 32308 37148 32360
rect 22284 32172 22336 32224
rect 23204 32215 23256 32224
rect 23204 32181 23213 32215
rect 23213 32181 23247 32215
rect 23247 32181 23256 32215
rect 23204 32172 23256 32181
rect 23940 32215 23992 32224
rect 23940 32181 23949 32215
rect 23949 32181 23983 32215
rect 23983 32181 23992 32215
rect 23940 32172 23992 32181
rect 26056 32172 26108 32224
rect 27804 32172 27856 32224
rect 29736 32215 29788 32224
rect 29736 32181 29745 32215
rect 29745 32181 29779 32215
rect 29779 32181 29788 32215
rect 29736 32172 29788 32181
rect 32128 32240 32180 32292
rect 36360 32172 36412 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 11060 32011 11112 32020
rect 11060 31977 11069 32011
rect 11069 31977 11103 32011
rect 11103 31977 11112 32011
rect 11060 31968 11112 31977
rect 11428 32011 11480 32020
rect 11428 31977 11437 32011
rect 11437 31977 11471 32011
rect 11471 31977 11480 32011
rect 11428 31968 11480 31977
rect 13544 32011 13596 32020
rect 13544 31977 13553 32011
rect 13553 31977 13587 32011
rect 13587 31977 13596 32011
rect 13544 31968 13596 31977
rect 17224 32011 17276 32020
rect 17224 31977 17233 32011
rect 17233 31977 17267 32011
rect 17267 31977 17276 32011
rect 17224 31968 17276 31977
rect 17684 32011 17736 32020
rect 17684 31977 17693 32011
rect 17693 31977 17727 32011
rect 17727 31977 17736 32011
rect 17684 31968 17736 31977
rect 9128 31900 9180 31952
rect 13636 31832 13688 31884
rect 7932 31764 7984 31816
rect 10968 31807 11020 31816
rect 10968 31773 10977 31807
rect 10977 31773 11011 31807
rect 11011 31773 11020 31807
rect 10968 31764 11020 31773
rect 11152 31764 11204 31816
rect 16120 31764 16172 31816
rect 17040 31900 17092 31952
rect 23020 32011 23072 32020
rect 23020 31977 23029 32011
rect 23029 31977 23063 32011
rect 23063 31977 23072 32011
rect 23020 31968 23072 31977
rect 23204 32011 23256 32020
rect 23204 31977 23213 32011
rect 23213 31977 23247 32011
rect 23247 31977 23256 32011
rect 23204 31968 23256 31977
rect 23756 32011 23808 32020
rect 23756 31977 23765 32011
rect 23765 31977 23799 32011
rect 23799 31977 23808 32011
rect 23756 31968 23808 31977
rect 23940 31968 23992 32020
rect 26056 32011 26108 32020
rect 26056 31977 26065 32011
rect 26065 31977 26099 32011
rect 26099 31977 26108 32011
rect 26056 31968 26108 31977
rect 26516 32011 26568 32020
rect 26516 31977 26525 32011
rect 26525 31977 26559 32011
rect 26559 31977 26568 32011
rect 26516 31968 26568 31977
rect 26608 32011 26660 32020
rect 26608 31977 26617 32011
rect 26617 31977 26651 32011
rect 26651 31977 26660 32011
rect 26608 31968 26660 31977
rect 17868 31764 17920 31816
rect 18972 31764 19024 31816
rect 19340 31807 19392 31816
rect 19340 31773 19349 31807
rect 19349 31773 19383 31807
rect 19383 31773 19392 31807
rect 20812 31832 20864 31884
rect 29736 31900 29788 31952
rect 26424 31832 26476 31884
rect 34428 31968 34480 32020
rect 30932 31832 30984 31884
rect 31392 31832 31444 31884
rect 32772 31832 32824 31884
rect 19340 31764 19392 31773
rect 19984 31807 20036 31816
rect 19984 31773 19993 31807
rect 19993 31773 20027 31807
rect 20027 31773 20036 31807
rect 19984 31764 20036 31773
rect 21916 31807 21968 31816
rect 21916 31773 21925 31807
rect 21925 31773 21959 31807
rect 21959 31773 21968 31807
rect 21916 31764 21968 31773
rect 22008 31764 22060 31816
rect 22744 31764 22796 31816
rect 23020 31807 23072 31816
rect 23020 31773 23029 31807
rect 23029 31773 23063 31807
rect 23063 31773 23072 31807
rect 23020 31764 23072 31773
rect 23940 31807 23992 31816
rect 23940 31773 23949 31807
rect 23949 31773 23983 31807
rect 23983 31773 23992 31807
rect 23940 31764 23992 31773
rect 24124 31764 24176 31816
rect 22468 31696 22520 31748
rect 23480 31696 23532 31748
rect 17500 31628 17552 31680
rect 19616 31671 19668 31680
rect 19616 31637 19625 31671
rect 19625 31637 19659 31671
rect 19659 31637 19668 31671
rect 19616 31628 19668 31637
rect 22376 31628 22428 31680
rect 26148 31696 26200 31748
rect 26976 31807 27028 31816
rect 26976 31773 26985 31807
rect 26985 31773 27019 31807
rect 27019 31773 27028 31807
rect 26976 31764 27028 31773
rect 28816 31764 28868 31816
rect 31024 31764 31076 31816
rect 28356 31696 28408 31748
rect 31484 31807 31536 31816
rect 31484 31773 31493 31807
rect 31493 31773 31527 31807
rect 31527 31773 31536 31807
rect 31484 31764 31536 31773
rect 33324 31696 33376 31748
rect 27528 31628 27580 31680
rect 28080 31671 28132 31680
rect 28080 31637 28089 31671
rect 28089 31637 28123 31671
rect 28123 31637 28132 31671
rect 28080 31628 28132 31637
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 12072 31424 12124 31476
rect 11152 31399 11204 31408
rect 11152 31365 11161 31399
rect 11161 31365 11195 31399
rect 11195 31365 11204 31399
rect 11152 31356 11204 31365
rect 14556 31331 14608 31340
rect 14556 31297 14565 31331
rect 14565 31297 14599 31331
rect 14599 31297 14608 31331
rect 14556 31288 14608 31297
rect 14740 31331 14792 31340
rect 14740 31297 14749 31331
rect 14749 31297 14783 31331
rect 14783 31297 14792 31331
rect 14740 31288 14792 31297
rect 15200 31288 15252 31340
rect 15476 31331 15528 31340
rect 15476 31297 15485 31331
rect 15485 31297 15519 31331
rect 15519 31297 15528 31331
rect 15476 31288 15528 31297
rect 22192 31424 22244 31476
rect 22744 31424 22796 31476
rect 20720 31399 20772 31408
rect 20720 31365 20729 31399
rect 20729 31365 20763 31399
rect 20763 31365 20772 31399
rect 20720 31356 20772 31365
rect 20076 31331 20128 31340
rect 20076 31297 20085 31331
rect 20085 31297 20119 31331
rect 20119 31297 20128 31331
rect 20076 31288 20128 31297
rect 16028 31220 16080 31272
rect 16488 31220 16540 31272
rect 19892 31220 19944 31272
rect 22284 31331 22336 31340
rect 22284 31297 22293 31331
rect 22293 31297 22327 31331
rect 22327 31297 22336 31331
rect 22284 31288 22336 31297
rect 23388 31288 23440 31340
rect 23572 31288 23624 31340
rect 33784 31424 33836 31476
rect 28540 31399 28592 31408
rect 28540 31365 28549 31399
rect 28549 31365 28583 31399
rect 28583 31365 28592 31399
rect 28540 31356 28592 31365
rect 30288 31356 30340 31408
rect 10324 31084 10376 31136
rect 22468 31263 22520 31272
rect 22468 31229 22477 31263
rect 22477 31229 22511 31263
rect 22511 31229 22520 31263
rect 22468 31220 22520 31229
rect 23296 31220 23348 31272
rect 25964 31220 26016 31272
rect 26148 31220 26200 31272
rect 28080 31288 28132 31340
rect 28356 31288 28408 31340
rect 31116 31331 31168 31340
rect 31116 31297 31125 31331
rect 31125 31297 31159 31331
rect 31159 31297 31168 31331
rect 31116 31288 31168 31297
rect 31484 31288 31536 31340
rect 32864 31331 32916 31340
rect 32864 31297 32873 31331
rect 32873 31297 32907 31331
rect 32907 31297 32916 31331
rect 32864 31288 32916 31297
rect 33140 31331 33192 31340
rect 33140 31297 33149 31331
rect 33149 31297 33183 31331
rect 33183 31297 33192 31331
rect 33140 31288 33192 31297
rect 33416 31288 33468 31340
rect 34612 31288 34664 31340
rect 26608 31220 26660 31272
rect 26700 31220 26752 31272
rect 29368 31220 29420 31272
rect 15292 31084 15344 31136
rect 19616 31127 19668 31136
rect 19616 31093 19625 31127
rect 19625 31093 19659 31127
rect 19659 31093 19668 31127
rect 19616 31084 19668 31093
rect 19984 31127 20036 31136
rect 19984 31093 19993 31127
rect 19993 31093 20027 31127
rect 20027 31093 20036 31127
rect 19984 31084 20036 31093
rect 20720 31084 20772 31136
rect 22100 31127 22152 31136
rect 22100 31093 22109 31127
rect 22109 31093 22143 31127
rect 22143 31093 22152 31127
rect 22100 31084 22152 31093
rect 22376 31127 22428 31136
rect 22376 31093 22385 31127
rect 22385 31093 22419 31127
rect 22419 31093 22428 31127
rect 22376 31084 22428 31093
rect 25872 31084 25924 31136
rect 26056 31127 26108 31136
rect 26056 31093 26065 31127
rect 26065 31093 26099 31127
rect 26099 31093 26108 31127
rect 26056 31084 26108 31093
rect 26332 31152 26384 31204
rect 32956 31152 33008 31204
rect 26240 31084 26292 31136
rect 28908 31127 28960 31136
rect 28908 31093 28917 31127
rect 28917 31093 28951 31127
rect 28951 31093 28960 31127
rect 28908 31084 28960 31093
rect 32864 31084 32916 31136
rect 36544 31220 36596 31272
rect 33600 31152 33652 31204
rect 33692 31152 33744 31204
rect 36268 31152 36320 31204
rect 33416 31127 33468 31136
rect 33416 31093 33425 31127
rect 33425 31093 33459 31127
rect 33459 31093 33468 31127
rect 33416 31084 33468 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 11888 30880 11940 30932
rect 12348 30880 12400 30932
rect 14556 30880 14608 30932
rect 12808 30744 12860 30796
rect 19524 30880 19576 30932
rect 22560 30923 22612 30932
rect 22560 30889 22569 30923
rect 22569 30889 22603 30923
rect 22603 30889 22612 30923
rect 22560 30880 22612 30889
rect 23480 30923 23532 30932
rect 23480 30889 23489 30923
rect 23489 30889 23523 30923
rect 23523 30889 23532 30923
rect 23480 30880 23532 30889
rect 23572 30880 23624 30932
rect 24492 30880 24544 30932
rect 26148 30880 26200 30932
rect 27344 30923 27396 30932
rect 27344 30889 27353 30923
rect 27353 30889 27387 30923
rect 27387 30889 27396 30923
rect 27344 30880 27396 30889
rect 27988 30880 28040 30932
rect 28724 30923 28776 30932
rect 28724 30889 28733 30923
rect 28733 30889 28767 30923
rect 28767 30889 28776 30923
rect 28724 30880 28776 30889
rect 32220 30880 32272 30932
rect 33048 30880 33100 30932
rect 33508 30880 33560 30932
rect 34428 30880 34480 30932
rect 38016 30880 38068 30932
rect 17684 30812 17736 30864
rect 18512 30744 18564 30796
rect 13360 30676 13412 30728
rect 15660 30676 15712 30728
rect 23020 30744 23072 30796
rect 22744 30676 22796 30728
rect 23756 30719 23808 30728
rect 23756 30685 23765 30719
rect 23765 30685 23799 30719
rect 23799 30685 23808 30719
rect 23756 30676 23808 30685
rect 24768 30676 24820 30728
rect 12072 30608 12124 30660
rect 14464 30651 14516 30660
rect 14464 30617 14473 30651
rect 14473 30617 14507 30651
rect 14507 30617 14516 30651
rect 14464 30608 14516 30617
rect 12900 30540 12952 30592
rect 13636 30540 13688 30592
rect 14740 30608 14792 30660
rect 19800 30608 19852 30660
rect 18236 30540 18288 30592
rect 19156 30540 19208 30592
rect 20444 30583 20496 30592
rect 20444 30549 20453 30583
rect 20453 30549 20487 30583
rect 20487 30549 20496 30583
rect 23940 30651 23992 30660
rect 23940 30617 23949 30651
rect 23949 30617 23983 30651
rect 23983 30617 23992 30651
rect 23940 30608 23992 30617
rect 25964 30812 26016 30864
rect 28264 30812 28316 30864
rect 26608 30744 26660 30796
rect 31116 30812 31168 30864
rect 33140 30812 33192 30864
rect 20444 30540 20496 30549
rect 21824 30540 21876 30592
rect 25504 30540 25556 30592
rect 26056 30651 26108 30660
rect 26056 30617 26065 30651
rect 26065 30617 26099 30651
rect 26099 30617 26108 30651
rect 26056 30608 26108 30617
rect 26332 30540 26384 30592
rect 27436 30719 27488 30728
rect 27436 30685 27445 30719
rect 27445 30685 27479 30719
rect 27479 30685 27488 30719
rect 27436 30676 27488 30685
rect 27988 30676 28040 30728
rect 26976 30651 27028 30660
rect 26976 30617 26985 30651
rect 26985 30617 27019 30651
rect 27019 30617 27028 30651
rect 26976 30608 27028 30617
rect 27068 30608 27120 30660
rect 33692 30744 33744 30796
rect 33784 30787 33836 30796
rect 33784 30753 33793 30787
rect 33793 30753 33827 30787
rect 33827 30753 33836 30787
rect 33784 30744 33836 30753
rect 28908 30719 28960 30728
rect 28908 30685 28917 30719
rect 28917 30685 28951 30719
rect 28951 30685 28960 30719
rect 28908 30676 28960 30685
rect 33232 30676 33284 30728
rect 33324 30676 33376 30728
rect 34520 30676 34572 30728
rect 35992 30719 36044 30728
rect 35992 30685 36001 30719
rect 36001 30685 36035 30719
rect 36035 30685 36044 30719
rect 35992 30676 36044 30685
rect 36176 30719 36228 30728
rect 36176 30685 36185 30719
rect 36185 30685 36219 30719
rect 36219 30685 36228 30719
rect 36176 30676 36228 30685
rect 33140 30608 33192 30660
rect 28448 30540 28500 30592
rect 29920 30540 29972 30592
rect 31116 30540 31168 30592
rect 32312 30540 32364 30592
rect 32772 30540 32824 30592
rect 33508 30583 33560 30592
rect 33508 30549 33517 30583
rect 33517 30549 33551 30583
rect 33551 30549 33560 30583
rect 33508 30540 33560 30549
rect 33692 30651 33744 30660
rect 33692 30617 33701 30651
rect 33701 30617 33735 30651
rect 33735 30617 33744 30651
rect 33692 30608 33744 30617
rect 33784 30608 33836 30660
rect 34796 30608 34848 30660
rect 35348 30540 35400 30592
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 7840 30268 7892 30320
rect 14464 30336 14516 30388
rect 18512 30379 18564 30388
rect 18512 30345 18521 30379
rect 18521 30345 18555 30379
rect 18555 30345 18564 30379
rect 18512 30336 18564 30345
rect 18788 30336 18840 30388
rect 22468 30336 22520 30388
rect 22560 30336 22612 30388
rect 24308 30336 24360 30388
rect 24492 30379 24544 30388
rect 24492 30345 24501 30379
rect 24501 30345 24535 30379
rect 24535 30345 24544 30379
rect 24492 30336 24544 30345
rect 25964 30336 26016 30388
rect 33692 30336 33744 30388
rect 9772 30243 9824 30252
rect 9772 30209 9781 30243
rect 9781 30209 9815 30243
rect 9815 30209 9824 30243
rect 9772 30200 9824 30209
rect 6552 29996 6604 30048
rect 10876 30268 10928 30320
rect 11060 30132 11112 30184
rect 13452 30132 13504 30184
rect 15752 30243 15804 30252
rect 15752 30209 15761 30243
rect 15761 30209 15795 30243
rect 15795 30209 15804 30243
rect 15752 30200 15804 30209
rect 15844 30200 15896 30252
rect 13820 30132 13872 30184
rect 17408 30200 17460 30252
rect 17592 30200 17644 30252
rect 18052 30243 18104 30252
rect 18052 30209 18061 30243
rect 18061 30209 18095 30243
rect 18095 30209 18104 30243
rect 18052 30200 18104 30209
rect 18236 30200 18288 30252
rect 17316 30175 17368 30184
rect 17316 30141 17325 30175
rect 17325 30141 17359 30175
rect 17359 30141 17368 30175
rect 17316 30132 17368 30141
rect 9772 30064 9824 30116
rect 10876 30064 10928 30116
rect 9680 29996 9732 30048
rect 10048 30039 10100 30048
rect 10048 30005 10057 30039
rect 10057 30005 10091 30039
rect 10091 30005 10100 30039
rect 10048 29996 10100 30005
rect 13728 30064 13780 30116
rect 15752 30064 15804 30116
rect 16856 30064 16908 30116
rect 17684 30107 17736 30116
rect 17684 30073 17693 30107
rect 17693 30073 17727 30107
rect 17727 30073 17736 30107
rect 17684 30064 17736 30073
rect 18696 30268 18748 30320
rect 18788 30243 18840 30252
rect 18788 30209 18797 30243
rect 18797 30209 18831 30243
rect 18831 30209 18840 30243
rect 18788 30200 18840 30209
rect 18972 30311 19024 30320
rect 18972 30277 18981 30311
rect 18981 30277 19015 30311
rect 19015 30277 19024 30311
rect 18972 30268 19024 30277
rect 21640 30268 21692 30320
rect 23848 30268 23900 30320
rect 19432 30200 19484 30252
rect 19524 30200 19576 30252
rect 19892 30200 19944 30252
rect 22652 30243 22704 30252
rect 22652 30209 22661 30243
rect 22661 30209 22695 30243
rect 22695 30209 22704 30243
rect 22652 30200 22704 30209
rect 23020 30200 23072 30252
rect 23480 30200 23532 30252
rect 18880 30132 18932 30184
rect 21916 30132 21968 30184
rect 24032 30243 24084 30252
rect 24032 30209 24041 30243
rect 24041 30209 24075 30243
rect 24075 30209 24084 30243
rect 24032 30200 24084 30209
rect 24216 30268 24268 30320
rect 18604 30064 18656 30116
rect 24216 30175 24268 30184
rect 24216 30141 24225 30175
rect 24225 30141 24259 30175
rect 24259 30141 24268 30175
rect 24216 30132 24268 30141
rect 14556 29996 14608 30048
rect 16028 29996 16080 30048
rect 17224 30039 17276 30048
rect 17224 30005 17233 30039
rect 17233 30005 17267 30039
rect 17267 30005 17276 30039
rect 17224 29996 17276 30005
rect 17868 29996 17920 30048
rect 18144 29996 18196 30048
rect 18788 29996 18840 30048
rect 19156 29996 19208 30048
rect 19524 29996 19576 30048
rect 19616 29996 19668 30048
rect 23480 30064 23532 30116
rect 23940 30064 23992 30116
rect 22376 29996 22428 30048
rect 23388 29996 23440 30048
rect 24492 30064 24544 30116
rect 29092 30243 29144 30252
rect 29092 30209 29101 30243
rect 29101 30209 29135 30243
rect 29135 30209 29144 30243
rect 29092 30200 29144 30209
rect 29368 30243 29420 30252
rect 29368 30209 29377 30243
rect 29377 30209 29411 30243
rect 29411 30209 29420 30243
rect 29368 30200 29420 30209
rect 30196 30243 30248 30252
rect 30196 30209 30205 30243
rect 30205 30209 30239 30243
rect 30239 30209 30248 30243
rect 30196 30200 30248 30209
rect 30380 30200 30432 30252
rect 30748 30243 30800 30252
rect 30748 30209 30757 30243
rect 30757 30209 30791 30243
rect 30791 30209 30800 30243
rect 30748 30200 30800 30209
rect 31668 30268 31720 30320
rect 31852 30268 31904 30320
rect 31484 30243 31536 30252
rect 31484 30209 31493 30243
rect 31493 30209 31527 30243
rect 31527 30209 31536 30243
rect 31484 30200 31536 30209
rect 31760 30200 31812 30252
rect 32404 30200 32456 30252
rect 33416 30268 33468 30320
rect 35992 30268 36044 30320
rect 32680 30200 32732 30252
rect 27712 30132 27764 30184
rect 29276 30175 29328 30184
rect 29276 30141 29285 30175
rect 29285 30141 29319 30175
rect 29319 30141 29328 30175
rect 29276 30132 29328 30141
rect 29828 30132 29880 30184
rect 30104 30175 30156 30184
rect 30104 30141 30113 30175
rect 30113 30141 30147 30175
rect 30147 30141 30156 30175
rect 30104 30132 30156 30141
rect 30564 30175 30616 30184
rect 30564 30141 30573 30175
rect 30573 30141 30607 30175
rect 30607 30141 30616 30175
rect 30564 30132 30616 30141
rect 25872 29996 25924 30048
rect 26240 29996 26292 30048
rect 30288 30064 30340 30116
rect 33784 30132 33836 30184
rect 29460 29996 29512 30048
rect 29552 30039 29604 30048
rect 29552 30005 29561 30039
rect 29561 30005 29595 30039
rect 29595 30005 29604 30039
rect 29552 29996 29604 30005
rect 29920 30039 29972 30048
rect 29920 30005 29929 30039
rect 29929 30005 29963 30039
rect 29963 30005 29972 30039
rect 29920 29996 29972 30005
rect 30472 30039 30524 30048
rect 30472 30005 30481 30039
rect 30481 30005 30515 30039
rect 30515 30005 30524 30039
rect 30472 29996 30524 30005
rect 31116 30064 31168 30116
rect 32128 30107 32180 30116
rect 32128 30073 32137 30107
rect 32137 30073 32171 30107
rect 32171 30073 32180 30107
rect 32128 30064 32180 30073
rect 31944 29996 31996 30048
rect 34796 29996 34848 30048
rect 37004 29996 37056 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 9128 29835 9180 29844
rect 9128 29801 9137 29835
rect 9137 29801 9171 29835
rect 9171 29801 9180 29835
rect 9128 29792 9180 29801
rect 9956 29792 10008 29844
rect 9312 29656 9364 29708
rect 11152 29656 11204 29708
rect 13636 29792 13688 29844
rect 13728 29835 13780 29844
rect 13728 29801 13737 29835
rect 13737 29801 13771 29835
rect 13771 29801 13780 29835
rect 13728 29792 13780 29801
rect 13452 29724 13504 29776
rect 16028 29792 16080 29844
rect 16764 29835 16816 29844
rect 11060 29588 11112 29640
rect 11244 29588 11296 29640
rect 13728 29656 13780 29708
rect 14464 29699 14516 29708
rect 14464 29665 14473 29699
rect 14473 29665 14507 29699
rect 14507 29665 14516 29699
rect 14464 29656 14516 29665
rect 10692 29520 10744 29572
rect 13636 29631 13688 29640
rect 13636 29597 13645 29631
rect 13645 29597 13679 29631
rect 13679 29597 13688 29631
rect 13636 29588 13688 29597
rect 14280 29631 14332 29640
rect 14280 29597 14289 29631
rect 14289 29597 14323 29631
rect 14323 29597 14332 29631
rect 14280 29588 14332 29597
rect 14556 29631 14608 29640
rect 14556 29597 14565 29631
rect 14565 29597 14599 29631
rect 14599 29597 14608 29631
rect 14556 29588 14608 29597
rect 15200 29520 15252 29572
rect 16764 29801 16773 29835
rect 16773 29801 16807 29835
rect 16807 29801 16816 29835
rect 16764 29792 16816 29801
rect 18788 29835 18840 29844
rect 18788 29801 18797 29835
rect 18797 29801 18831 29835
rect 18831 29801 18840 29835
rect 18788 29792 18840 29801
rect 19064 29835 19116 29844
rect 19064 29801 19073 29835
rect 19073 29801 19107 29835
rect 19107 29801 19116 29835
rect 19064 29792 19116 29801
rect 19156 29792 19208 29844
rect 20904 29792 20956 29844
rect 21824 29792 21876 29844
rect 21916 29792 21968 29844
rect 16764 29656 16816 29708
rect 16396 29631 16448 29640
rect 16396 29597 16405 29631
rect 16405 29597 16439 29631
rect 16439 29597 16448 29631
rect 16396 29588 16448 29597
rect 16580 29520 16632 29572
rect 16764 29520 16816 29572
rect 17040 29520 17092 29572
rect 17408 29520 17460 29572
rect 18144 29588 18196 29640
rect 18696 29631 18748 29640
rect 18696 29597 18710 29631
rect 18710 29597 18744 29631
rect 18744 29597 18748 29631
rect 18696 29588 18748 29597
rect 19432 29699 19484 29708
rect 19432 29665 19441 29699
rect 19441 29665 19475 29699
rect 19475 29665 19484 29699
rect 19432 29656 19484 29665
rect 20536 29656 20588 29708
rect 19984 29631 20036 29640
rect 19984 29597 19991 29631
rect 19991 29597 20025 29631
rect 20025 29597 20036 29631
rect 21088 29724 21140 29776
rect 24492 29724 24544 29776
rect 26148 29835 26200 29844
rect 26148 29801 26157 29835
rect 26157 29801 26191 29835
rect 26191 29801 26200 29835
rect 26148 29792 26200 29801
rect 26884 29835 26936 29844
rect 26884 29801 26893 29835
rect 26893 29801 26927 29835
rect 26927 29801 26936 29835
rect 26884 29792 26936 29801
rect 27436 29792 27488 29844
rect 28724 29835 28776 29844
rect 28724 29801 28733 29835
rect 28733 29801 28767 29835
rect 28767 29801 28776 29835
rect 28724 29792 28776 29801
rect 20904 29699 20956 29708
rect 20904 29665 20913 29699
rect 20913 29665 20947 29699
rect 20947 29665 20956 29699
rect 20904 29656 20956 29665
rect 21456 29656 21508 29708
rect 24216 29656 24268 29708
rect 24400 29656 24452 29708
rect 19984 29588 20036 29597
rect 10784 29452 10836 29504
rect 11796 29452 11848 29504
rect 14096 29495 14148 29504
rect 14096 29461 14105 29495
rect 14105 29461 14139 29495
rect 14139 29461 14148 29495
rect 14096 29452 14148 29461
rect 14740 29452 14792 29504
rect 18604 29520 18656 29572
rect 19294 29563 19346 29572
rect 19294 29529 19316 29563
rect 19316 29529 19346 29563
rect 19294 29520 19346 29529
rect 19800 29563 19852 29572
rect 19800 29529 19809 29563
rect 19809 29529 19843 29563
rect 19843 29529 19852 29563
rect 19800 29520 19852 29529
rect 20628 29520 20680 29572
rect 21088 29631 21140 29640
rect 21088 29597 21097 29631
rect 21097 29597 21131 29631
rect 21131 29597 21140 29631
rect 21088 29588 21140 29597
rect 26240 29631 26292 29640
rect 26240 29597 26249 29631
rect 26249 29597 26283 29631
rect 26283 29597 26292 29631
rect 26240 29588 26292 29597
rect 19156 29452 19208 29504
rect 19708 29452 19760 29504
rect 20168 29495 20220 29504
rect 20168 29461 20177 29495
rect 20177 29461 20211 29495
rect 20211 29461 20220 29495
rect 20168 29452 20220 29461
rect 22008 29452 22060 29504
rect 22652 29452 22704 29504
rect 23020 29452 23072 29504
rect 23204 29452 23256 29504
rect 24400 29452 24452 29504
rect 25872 29495 25924 29504
rect 25872 29461 25881 29495
rect 25881 29461 25915 29495
rect 25915 29461 25924 29495
rect 25872 29452 25924 29461
rect 26516 29520 26568 29572
rect 27712 29656 27764 29708
rect 27988 29724 28040 29776
rect 29092 29767 29144 29776
rect 29092 29733 29101 29767
rect 29101 29733 29135 29767
rect 29135 29733 29144 29767
rect 29092 29724 29144 29733
rect 29184 29724 29236 29776
rect 29736 29724 29788 29776
rect 30012 29835 30064 29844
rect 30012 29801 30021 29835
rect 30021 29801 30055 29835
rect 30055 29801 30064 29835
rect 30012 29792 30064 29801
rect 30380 29835 30432 29844
rect 30380 29801 30389 29835
rect 30389 29801 30423 29835
rect 30423 29801 30432 29835
rect 30380 29792 30432 29801
rect 31668 29792 31720 29844
rect 30564 29724 30616 29776
rect 31852 29792 31904 29844
rect 33968 29792 34020 29844
rect 29828 29656 29880 29708
rect 26700 29631 26752 29640
rect 26700 29597 26709 29631
rect 26709 29597 26743 29631
rect 26743 29597 26752 29631
rect 26700 29588 26752 29597
rect 30380 29656 30432 29708
rect 31392 29656 31444 29708
rect 32036 29724 32088 29776
rect 32404 29724 32456 29776
rect 38384 29724 38436 29776
rect 28356 29520 28408 29572
rect 28632 29563 28684 29572
rect 28632 29529 28641 29563
rect 28641 29529 28675 29563
rect 28675 29529 28684 29563
rect 28632 29520 28684 29529
rect 29552 29520 29604 29572
rect 31116 29588 31168 29640
rect 31668 29631 31720 29640
rect 31668 29597 31684 29631
rect 31684 29597 31718 29631
rect 31718 29597 31720 29631
rect 31668 29588 31720 29597
rect 32128 29588 32180 29640
rect 32680 29588 32732 29640
rect 35992 29656 36044 29708
rect 30104 29452 30156 29504
rect 30564 29452 30616 29504
rect 30656 29452 30708 29504
rect 32496 29563 32548 29572
rect 32496 29529 32505 29563
rect 32505 29529 32539 29563
rect 32539 29529 32548 29563
rect 32496 29520 32548 29529
rect 34704 29520 34756 29572
rect 36084 29631 36136 29640
rect 36084 29597 36093 29631
rect 36093 29597 36127 29631
rect 36127 29597 36136 29631
rect 36084 29588 36136 29597
rect 44548 29631 44600 29640
rect 44548 29597 44557 29631
rect 44557 29597 44591 29631
rect 44591 29597 44600 29631
rect 44548 29588 44600 29597
rect 32036 29452 32088 29504
rect 37648 29520 37700 29572
rect 35440 29452 35492 29504
rect 42800 29452 42852 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 7656 29291 7708 29300
rect 7656 29257 7665 29291
rect 7665 29257 7699 29291
rect 7699 29257 7708 29291
rect 7656 29248 7708 29257
rect 9312 29248 9364 29300
rect 8944 29180 8996 29232
rect 10508 29223 10560 29232
rect 10508 29189 10517 29223
rect 10517 29189 10551 29223
rect 10551 29189 10560 29223
rect 10508 29180 10560 29189
rect 11980 29291 12032 29300
rect 11980 29257 11989 29291
rect 11989 29257 12023 29291
rect 12023 29257 12032 29291
rect 11980 29248 12032 29257
rect 12992 29248 13044 29300
rect 17592 29291 17644 29300
rect 17592 29257 17601 29291
rect 17601 29257 17635 29291
rect 17635 29257 17644 29291
rect 17592 29248 17644 29257
rect 19432 29248 19484 29300
rect 19984 29248 20036 29300
rect 17040 29180 17092 29232
rect 17132 29180 17184 29232
rect 17408 29223 17460 29232
rect 17408 29189 17417 29223
rect 17417 29189 17451 29223
rect 17451 29189 17460 29223
rect 17408 29180 17460 29189
rect 18052 29180 18104 29232
rect 21824 29223 21876 29232
rect 21824 29189 21833 29223
rect 21833 29189 21867 29223
rect 21867 29189 21876 29223
rect 21824 29180 21876 29189
rect 23848 29248 23900 29300
rect 22744 29180 22796 29232
rect 25872 29180 25924 29232
rect 6920 29112 6972 29164
rect 10232 29112 10284 29164
rect 11428 29112 11480 29164
rect 11796 29155 11848 29164
rect 11796 29121 11805 29155
rect 11805 29121 11839 29155
rect 11839 29121 11848 29155
rect 11796 29112 11848 29121
rect 12992 29112 13044 29164
rect 13544 29112 13596 29164
rect 13636 29112 13688 29164
rect 7380 29087 7432 29096
rect 7380 29053 7389 29087
rect 7389 29053 7423 29087
rect 7423 29053 7432 29087
rect 7380 29044 7432 29053
rect 10692 29087 10744 29096
rect 10692 29053 10701 29087
rect 10701 29053 10735 29087
rect 10735 29053 10744 29087
rect 10692 29044 10744 29053
rect 11060 29044 11112 29096
rect 13268 29087 13320 29096
rect 13268 29053 13277 29087
rect 13277 29053 13311 29087
rect 13311 29053 13320 29087
rect 13268 29044 13320 29053
rect 13728 29044 13780 29096
rect 16948 29112 17000 29164
rect 18144 29112 18196 29164
rect 19248 29155 19300 29164
rect 19248 29121 19257 29155
rect 19257 29121 19291 29155
rect 19291 29121 19300 29155
rect 19248 29112 19300 29121
rect 19432 29112 19484 29164
rect 22192 29112 22244 29164
rect 23296 29112 23348 29164
rect 23480 29112 23532 29164
rect 7196 28951 7248 28960
rect 7196 28917 7205 28951
rect 7205 28917 7239 28951
rect 7239 28917 7248 28951
rect 7196 28908 7248 28917
rect 9680 28908 9732 28960
rect 10692 28951 10744 28960
rect 10692 28917 10701 28951
rect 10701 28917 10735 28951
rect 10735 28917 10744 28951
rect 10692 28908 10744 28917
rect 11704 28976 11756 29028
rect 16396 28976 16448 29028
rect 21640 29044 21692 29096
rect 21916 29087 21968 29096
rect 21916 29053 21925 29087
rect 21925 29053 21959 29087
rect 21959 29053 21968 29087
rect 21916 29044 21968 29053
rect 19340 28976 19392 29028
rect 24860 29155 24912 29164
rect 24860 29121 24869 29155
rect 24869 29121 24903 29155
rect 24903 29121 24912 29155
rect 24860 29112 24912 29121
rect 27988 29180 28040 29232
rect 28356 29248 28408 29300
rect 29184 29248 29236 29300
rect 29276 29248 29328 29300
rect 29552 29248 29604 29300
rect 31944 29248 31996 29300
rect 34796 29248 34848 29300
rect 28264 29223 28316 29232
rect 28264 29189 28273 29223
rect 28273 29189 28307 29223
rect 28307 29189 28316 29223
rect 28264 29180 28316 29189
rect 29000 29180 29052 29232
rect 29736 29180 29788 29232
rect 26792 29112 26844 29164
rect 28356 29112 28408 29164
rect 29276 29112 29328 29164
rect 29552 29112 29604 29164
rect 30564 29112 30616 29164
rect 30932 29112 30984 29164
rect 31116 29155 31168 29164
rect 31116 29121 31125 29155
rect 31125 29121 31159 29155
rect 31159 29121 31168 29155
rect 31116 29112 31168 29121
rect 31300 29180 31352 29232
rect 35072 29223 35124 29232
rect 35072 29189 35081 29223
rect 35081 29189 35115 29223
rect 35115 29189 35124 29223
rect 35072 29180 35124 29189
rect 28540 29044 28592 29096
rect 29460 29044 29512 29096
rect 23296 28976 23348 29028
rect 23388 28976 23440 29028
rect 28080 28976 28132 29028
rect 28908 28976 28960 29028
rect 31208 29087 31260 29096
rect 31208 29053 31217 29087
rect 31217 29053 31251 29087
rect 31251 29053 31260 29087
rect 31208 29044 31260 29053
rect 29920 28976 29972 29028
rect 31576 29019 31628 29028
rect 31576 28985 31585 29019
rect 31585 28985 31619 29019
rect 31619 28985 31628 29019
rect 31576 28976 31628 28985
rect 33876 29155 33928 29164
rect 33876 29121 33885 29155
rect 33885 29121 33919 29155
rect 33919 29121 33928 29155
rect 33876 29112 33928 29121
rect 34520 29112 34572 29164
rect 34704 29155 34756 29164
rect 34704 29121 34713 29155
rect 34713 29121 34747 29155
rect 34747 29121 34756 29155
rect 34704 29112 34756 29121
rect 35716 29248 35768 29300
rect 35440 29180 35492 29232
rect 35808 29180 35860 29232
rect 37372 29180 37424 29232
rect 38752 29155 38804 29164
rect 38752 29121 38786 29155
rect 38786 29121 38804 29155
rect 38752 29112 38804 29121
rect 34796 29087 34848 29096
rect 34796 29053 34805 29087
rect 34805 29053 34839 29087
rect 34839 29053 34848 29087
rect 34796 29044 34848 29053
rect 35256 29087 35308 29096
rect 35256 29053 35265 29087
rect 35265 29053 35299 29087
rect 35299 29053 35308 29087
rect 35256 29044 35308 29053
rect 35440 29044 35492 29096
rect 34152 28976 34204 29028
rect 35624 28976 35676 29028
rect 36268 29044 36320 29096
rect 37188 29044 37240 29096
rect 36176 28976 36228 29028
rect 37648 29019 37700 29028
rect 37648 28985 37657 29019
rect 37657 28985 37691 29019
rect 37691 28985 37700 29019
rect 37648 28976 37700 28985
rect 38292 28976 38344 29028
rect 44088 28976 44140 29028
rect 13084 28951 13136 28960
rect 13084 28917 13093 28951
rect 13093 28917 13127 28951
rect 13127 28917 13136 28951
rect 13084 28908 13136 28917
rect 17960 28908 18012 28960
rect 20168 28908 20220 28960
rect 21824 28951 21876 28960
rect 21824 28917 21833 28951
rect 21833 28917 21867 28951
rect 21867 28917 21876 28951
rect 21824 28908 21876 28917
rect 22468 28908 22520 28960
rect 23204 28908 23256 28960
rect 24952 28908 25004 28960
rect 25044 28951 25096 28960
rect 25044 28917 25053 28951
rect 25053 28917 25087 28951
rect 25087 28917 25096 28951
rect 25044 28908 25096 28917
rect 26332 28951 26384 28960
rect 26332 28917 26341 28951
rect 26341 28917 26375 28951
rect 26375 28917 26384 28951
rect 26332 28908 26384 28917
rect 26700 28951 26752 28960
rect 26700 28917 26709 28951
rect 26709 28917 26743 28951
rect 26743 28917 26752 28951
rect 26700 28908 26752 28917
rect 26792 28908 26844 28960
rect 28632 28908 28684 28960
rect 29368 28908 29420 28960
rect 29828 28908 29880 28960
rect 33876 28908 33928 28960
rect 34336 28908 34388 28960
rect 34888 28908 34940 28960
rect 36268 28908 36320 28960
rect 39948 28951 40000 28960
rect 39948 28917 39957 28951
rect 39957 28917 39991 28951
rect 39991 28917 40000 28951
rect 39948 28908 40000 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 8944 28747 8996 28756
rect 8944 28713 8953 28747
rect 8953 28713 8987 28747
rect 8987 28713 8996 28747
rect 8944 28704 8996 28713
rect 9312 28747 9364 28756
rect 9312 28713 9321 28747
rect 9321 28713 9355 28747
rect 9355 28713 9364 28747
rect 9312 28704 9364 28713
rect 9680 28704 9732 28756
rect 11060 28704 11112 28756
rect 11336 28747 11388 28756
rect 11336 28713 11345 28747
rect 11345 28713 11379 28747
rect 11379 28713 11388 28747
rect 11336 28704 11388 28713
rect 8024 28636 8076 28688
rect 21824 28704 21876 28756
rect 22836 28704 22888 28756
rect 23296 28747 23348 28756
rect 23296 28713 23305 28747
rect 23305 28713 23339 28747
rect 23339 28713 23348 28747
rect 23296 28704 23348 28713
rect 11520 28636 11572 28688
rect 13176 28636 13228 28688
rect 13728 28636 13780 28688
rect 16120 28636 16172 28688
rect 27436 28704 27488 28756
rect 28816 28747 28868 28756
rect 28816 28713 28825 28747
rect 28825 28713 28859 28747
rect 28859 28713 28868 28747
rect 28816 28704 28868 28713
rect 29736 28704 29788 28756
rect 31116 28704 31168 28756
rect 31668 28704 31720 28756
rect 34336 28704 34388 28756
rect 35348 28704 35400 28756
rect 36084 28704 36136 28756
rect 37188 28704 37240 28756
rect 38384 28704 38436 28756
rect 38752 28704 38804 28756
rect 11428 28568 11480 28620
rect 9128 28543 9180 28552
rect 9128 28509 9137 28543
rect 9137 28509 9171 28543
rect 9171 28509 9180 28543
rect 9128 28500 9180 28509
rect 9588 28500 9640 28552
rect 9956 28500 10008 28552
rect 10692 28500 10744 28552
rect 23204 28568 23256 28620
rect 23388 28568 23440 28620
rect 25504 28568 25556 28620
rect 26148 28568 26200 28620
rect 28908 28636 28960 28688
rect 29000 28636 29052 28688
rect 28816 28568 28868 28620
rect 31300 28636 31352 28688
rect 33140 28636 33192 28688
rect 33324 28636 33376 28688
rect 41144 28636 41196 28688
rect 34060 28568 34112 28620
rect 34612 28568 34664 28620
rect 36728 28568 36780 28620
rect 38016 28611 38068 28620
rect 38016 28577 38025 28611
rect 38025 28577 38059 28611
rect 38059 28577 38068 28611
rect 38016 28568 38068 28577
rect 38568 28568 38620 28620
rect 40040 28568 40092 28620
rect 5724 28432 5776 28484
rect 10600 28475 10652 28484
rect 10600 28441 10609 28475
rect 10609 28441 10643 28475
rect 10643 28441 10652 28475
rect 10600 28432 10652 28441
rect 10784 28475 10836 28484
rect 10784 28441 10793 28475
rect 10793 28441 10827 28475
rect 10827 28441 10836 28475
rect 10784 28432 10836 28441
rect 10876 28475 10928 28484
rect 10876 28441 10885 28475
rect 10885 28441 10919 28475
rect 10919 28441 10928 28475
rect 10876 28432 10928 28441
rect 18052 28432 18104 28484
rect 18236 28475 18288 28484
rect 18236 28441 18245 28475
rect 18245 28441 18279 28475
rect 18279 28441 18288 28475
rect 18236 28432 18288 28441
rect 18420 28475 18472 28484
rect 18420 28441 18429 28475
rect 18429 28441 18463 28475
rect 18463 28441 18472 28475
rect 18420 28432 18472 28441
rect 23112 28543 23164 28552
rect 23112 28509 23121 28543
rect 23121 28509 23155 28543
rect 23155 28509 23164 28543
rect 23112 28500 23164 28509
rect 26700 28500 26752 28552
rect 27252 28543 27304 28552
rect 27252 28509 27261 28543
rect 27261 28509 27295 28543
rect 27295 28509 27304 28543
rect 27252 28500 27304 28509
rect 27896 28500 27948 28552
rect 20260 28432 20312 28484
rect 22192 28432 22244 28484
rect 23388 28475 23440 28484
rect 23388 28441 23397 28475
rect 23397 28441 23431 28475
rect 23431 28441 23440 28475
rect 23388 28432 23440 28441
rect 24952 28432 25004 28484
rect 25596 28432 25648 28484
rect 26148 28432 26200 28484
rect 11520 28364 11572 28416
rect 14924 28364 14976 28416
rect 18512 28364 18564 28416
rect 18604 28407 18656 28416
rect 18604 28373 18613 28407
rect 18613 28373 18647 28407
rect 18647 28373 18656 28407
rect 18604 28364 18656 28373
rect 18788 28364 18840 28416
rect 20076 28364 20128 28416
rect 20168 28364 20220 28416
rect 26792 28364 26844 28416
rect 28264 28432 28316 28484
rect 28448 28432 28500 28484
rect 30288 28500 30340 28552
rect 30748 28500 30800 28552
rect 27712 28364 27764 28416
rect 27988 28407 28040 28416
rect 27988 28373 27997 28407
rect 27997 28373 28031 28407
rect 28031 28373 28040 28407
rect 27988 28364 28040 28373
rect 28724 28407 28776 28416
rect 28724 28373 28733 28407
rect 28733 28373 28767 28407
rect 28767 28373 28776 28407
rect 28724 28364 28776 28373
rect 29000 28364 29052 28416
rect 31392 28475 31444 28484
rect 31392 28441 31401 28475
rect 31401 28441 31435 28475
rect 31435 28441 31444 28475
rect 31392 28432 31444 28441
rect 32864 28475 32916 28484
rect 32864 28441 32873 28475
rect 32873 28441 32907 28475
rect 32907 28441 32916 28475
rect 32864 28432 32916 28441
rect 29368 28364 29420 28416
rect 32680 28407 32732 28416
rect 32680 28373 32689 28407
rect 32689 28373 32723 28407
rect 32723 28373 32732 28407
rect 33508 28432 33560 28484
rect 33876 28432 33928 28484
rect 34612 28432 34664 28484
rect 35716 28500 35768 28552
rect 35808 28543 35860 28552
rect 35808 28509 35817 28543
rect 35817 28509 35851 28543
rect 35851 28509 35860 28543
rect 35808 28500 35860 28509
rect 37004 28500 37056 28552
rect 32680 28364 32732 28373
rect 34336 28364 34388 28416
rect 35624 28475 35676 28484
rect 35624 28441 35633 28475
rect 35633 28441 35667 28475
rect 35667 28441 35676 28475
rect 35624 28432 35676 28441
rect 35992 28432 36044 28484
rect 37464 28432 37516 28484
rect 38752 28432 38804 28484
rect 35348 28407 35400 28416
rect 35348 28373 35357 28407
rect 35357 28373 35391 28407
rect 35391 28373 35400 28407
rect 35348 28364 35400 28373
rect 35532 28364 35584 28416
rect 36452 28364 36504 28416
rect 38200 28364 38252 28416
rect 38660 28364 38712 28416
rect 39948 28500 40000 28552
rect 41236 28543 41288 28552
rect 41236 28509 41245 28543
rect 41245 28509 41279 28543
rect 41279 28509 41288 28543
rect 41236 28500 41288 28509
rect 42064 28432 42116 28484
rect 42984 28364 43036 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 10692 28160 10744 28212
rect 10876 28203 10928 28212
rect 10876 28169 10885 28203
rect 10885 28169 10919 28203
rect 10919 28169 10928 28203
rect 10876 28160 10928 28169
rect 7564 28092 7616 28144
rect 11612 28092 11664 28144
rect 14464 28092 14516 28144
rect 15568 28160 15620 28212
rect 16304 28203 16356 28212
rect 16304 28169 16313 28203
rect 16313 28169 16347 28203
rect 16347 28169 16356 28203
rect 16304 28160 16356 28169
rect 16672 28160 16724 28212
rect 18788 28160 18840 28212
rect 18972 28160 19024 28212
rect 21640 28160 21692 28212
rect 5264 28024 5316 28076
rect 6092 27956 6144 28008
rect 7012 28024 7064 28076
rect 8024 28067 8076 28076
rect 8024 28033 8033 28067
rect 8033 28033 8067 28067
rect 8067 28033 8076 28067
rect 8024 28024 8076 28033
rect 6736 27956 6788 28008
rect 11060 28024 11112 28076
rect 13544 28024 13596 28076
rect 14280 28024 14332 28076
rect 15016 28024 15068 28076
rect 15200 28067 15252 28076
rect 15200 28033 15209 28067
rect 15209 28033 15243 28067
rect 15243 28033 15252 28067
rect 15200 28024 15252 28033
rect 6828 27931 6880 27940
rect 6828 27897 6837 27931
rect 6837 27897 6871 27931
rect 6871 27897 6880 27931
rect 6828 27888 6880 27897
rect 11796 27956 11848 28008
rect 13268 27999 13320 28008
rect 13268 27965 13277 27999
rect 13277 27965 13311 27999
rect 13311 27965 13320 27999
rect 13268 27956 13320 27965
rect 17408 28092 17460 28144
rect 19800 28092 19852 28144
rect 20076 28092 20128 28144
rect 15476 28067 15528 28076
rect 15476 28033 15485 28067
rect 15485 28033 15519 28067
rect 15519 28033 15528 28067
rect 15476 28024 15528 28033
rect 15844 28067 15896 28076
rect 15844 28033 15853 28067
rect 15853 28033 15887 28067
rect 15887 28033 15896 28067
rect 15844 28024 15896 28033
rect 11520 27888 11572 27940
rect 13084 27888 13136 27940
rect 15568 27956 15620 28008
rect 18512 28024 18564 28076
rect 18880 28067 18932 28076
rect 18880 28033 18889 28067
rect 18889 28033 18923 28067
rect 18923 28033 18932 28067
rect 18880 28024 18932 28033
rect 19156 28067 19208 28076
rect 19156 28033 19165 28067
rect 19165 28033 19199 28067
rect 19199 28033 19208 28067
rect 19156 28024 19208 28033
rect 19248 28024 19300 28076
rect 20536 28024 20588 28076
rect 24124 28024 24176 28076
rect 24216 28024 24268 28076
rect 26792 28203 26844 28212
rect 26792 28169 26801 28203
rect 26801 28169 26835 28203
rect 26835 28169 26844 28203
rect 26792 28160 26844 28169
rect 27436 28203 27488 28212
rect 27436 28169 27445 28203
rect 27445 28169 27479 28203
rect 27479 28169 27488 28203
rect 27436 28160 27488 28169
rect 27528 28203 27580 28212
rect 27528 28169 27537 28203
rect 27537 28169 27571 28203
rect 27571 28169 27580 28203
rect 27528 28160 27580 28169
rect 29000 28160 29052 28212
rect 29460 28160 29512 28212
rect 24860 28024 24912 28076
rect 16028 27999 16080 28008
rect 16028 27965 16037 27999
rect 16037 27965 16071 27999
rect 16071 27965 16080 27999
rect 16028 27956 16080 27965
rect 22836 27956 22888 28008
rect 23480 27956 23532 28008
rect 24492 27999 24544 28008
rect 24492 27965 24501 27999
rect 24501 27965 24535 27999
rect 24535 27965 24544 27999
rect 24492 27956 24544 27965
rect 21916 27888 21968 27940
rect 22008 27888 22060 27940
rect 27068 28092 27120 28144
rect 25044 28024 25096 28076
rect 26608 28067 26660 28076
rect 26608 28033 26617 28067
rect 26617 28033 26651 28067
rect 26651 28033 26660 28067
rect 26608 28024 26660 28033
rect 27252 28067 27304 28076
rect 27252 28033 27261 28067
rect 27261 28033 27295 28067
rect 27295 28033 27304 28067
rect 27252 28024 27304 28033
rect 27712 28067 27764 28076
rect 27712 28033 27721 28067
rect 27721 28033 27755 28067
rect 27755 28033 27764 28067
rect 27712 28024 27764 28033
rect 26700 27956 26752 28008
rect 27436 27888 27488 27940
rect 28816 28135 28868 28144
rect 28816 28101 28825 28135
rect 28825 28101 28859 28135
rect 28859 28101 28868 28135
rect 28816 28092 28868 28101
rect 30472 28160 30524 28212
rect 33968 28160 34020 28212
rect 38016 28160 38068 28212
rect 30196 28092 30248 28144
rect 30380 28092 30432 28144
rect 34060 28092 34112 28144
rect 36544 28135 36596 28144
rect 36544 28101 36553 28135
rect 36553 28101 36587 28135
rect 36587 28101 36596 28135
rect 36544 28092 36596 28101
rect 36728 28135 36780 28144
rect 36728 28101 36737 28135
rect 36737 28101 36771 28135
rect 36771 28101 36780 28135
rect 36728 28092 36780 28101
rect 37556 28092 37608 28144
rect 42800 28092 42852 28144
rect 28724 28024 28776 28076
rect 29920 28067 29972 28076
rect 29920 28033 29929 28067
rect 29929 28033 29963 28067
rect 29963 28033 29972 28067
rect 29920 28024 29972 28033
rect 38016 28024 38068 28076
rect 42984 28067 43036 28076
rect 42984 28033 42993 28067
rect 42993 28033 43027 28067
rect 43027 28033 43036 28067
rect 42984 28024 43036 28033
rect 32772 27999 32824 28008
rect 32772 27965 32781 27999
rect 32781 27965 32815 27999
rect 32815 27965 32824 27999
rect 32772 27956 32824 27965
rect 34060 27956 34112 28008
rect 36912 27956 36964 28008
rect 37096 27956 37148 28008
rect 35808 27888 35860 27940
rect 44456 27931 44508 27940
rect 44456 27897 44465 27931
rect 44465 27897 44499 27931
rect 44499 27897 44508 27931
rect 44456 27888 44508 27897
rect 7196 27820 7248 27872
rect 9864 27820 9916 27872
rect 10416 27863 10468 27872
rect 10416 27829 10425 27863
rect 10425 27829 10459 27863
rect 10459 27829 10468 27863
rect 10416 27820 10468 27829
rect 13452 27863 13504 27872
rect 13452 27829 13461 27863
rect 13461 27829 13495 27863
rect 13495 27829 13504 27863
rect 13452 27820 13504 27829
rect 13636 27863 13688 27872
rect 13636 27829 13645 27863
rect 13645 27829 13679 27863
rect 13679 27829 13688 27863
rect 13636 27820 13688 27829
rect 14924 27863 14976 27872
rect 14924 27829 14933 27863
rect 14933 27829 14967 27863
rect 14967 27829 14976 27863
rect 14924 27820 14976 27829
rect 15016 27820 15068 27872
rect 15660 27863 15712 27872
rect 15660 27829 15669 27863
rect 15669 27829 15703 27863
rect 15703 27829 15712 27863
rect 15660 27820 15712 27829
rect 16120 27863 16172 27872
rect 16120 27829 16129 27863
rect 16129 27829 16163 27863
rect 16163 27829 16172 27863
rect 16120 27820 16172 27829
rect 17960 27820 18012 27872
rect 18972 27820 19024 27872
rect 19064 27863 19116 27872
rect 19064 27829 19073 27863
rect 19073 27829 19107 27863
rect 19107 27829 19116 27863
rect 19064 27820 19116 27829
rect 19708 27820 19760 27872
rect 20444 27820 20496 27872
rect 21548 27820 21600 27872
rect 21640 27820 21692 27872
rect 23388 27820 23440 27872
rect 26240 27820 26292 27872
rect 26332 27863 26384 27872
rect 26332 27829 26341 27863
rect 26341 27829 26375 27863
rect 26375 27829 26384 27863
rect 26332 27820 26384 27829
rect 26608 27820 26660 27872
rect 27068 27820 27120 27872
rect 27160 27820 27212 27872
rect 28908 27820 28960 27872
rect 33140 27820 33192 27872
rect 34704 27820 34756 27872
rect 36544 27820 36596 27872
rect 37464 27820 37516 27872
rect 40040 27820 40092 27872
rect 40776 27820 40828 27872
rect 42432 27863 42484 27872
rect 42432 27829 42441 27863
rect 42441 27829 42475 27863
rect 42475 27829 42484 27863
rect 42432 27820 42484 27829
rect 42616 27820 42668 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 5356 27616 5408 27668
rect 6736 27659 6788 27668
rect 6736 27625 6745 27659
rect 6745 27625 6779 27659
rect 6779 27625 6788 27659
rect 6736 27616 6788 27625
rect 7564 27616 7616 27668
rect 7932 27548 7984 27600
rect 10416 27616 10468 27668
rect 6000 27455 6052 27464
rect 6000 27421 6009 27455
rect 6009 27421 6043 27455
rect 6043 27421 6052 27455
rect 6000 27412 6052 27421
rect 6828 27480 6880 27532
rect 9864 27480 9916 27532
rect 11060 27548 11112 27600
rect 18880 27616 18932 27668
rect 19340 27616 19392 27668
rect 19616 27616 19668 27668
rect 21916 27659 21968 27668
rect 21916 27625 21925 27659
rect 21925 27625 21959 27659
rect 21959 27625 21968 27659
rect 21916 27616 21968 27625
rect 22560 27616 22612 27668
rect 26608 27616 26660 27668
rect 26700 27659 26752 27668
rect 26700 27625 26709 27659
rect 26709 27625 26743 27659
rect 26743 27625 26752 27659
rect 26700 27616 26752 27625
rect 26884 27659 26936 27668
rect 26884 27625 26893 27659
rect 26893 27625 26927 27659
rect 26927 27625 26936 27659
rect 26884 27616 26936 27625
rect 13084 27480 13136 27532
rect 13268 27523 13320 27532
rect 13268 27489 13277 27523
rect 13277 27489 13311 27523
rect 13311 27489 13320 27523
rect 13268 27480 13320 27489
rect 5448 27344 5500 27396
rect 8208 27412 8260 27464
rect 8760 27412 8812 27464
rect 12992 27412 13044 27464
rect 19708 27548 19760 27600
rect 14556 27480 14608 27532
rect 15200 27480 15252 27532
rect 17500 27480 17552 27532
rect 19616 27412 19668 27464
rect 19800 27455 19852 27464
rect 19800 27421 19809 27455
rect 19809 27421 19843 27455
rect 19843 27421 19852 27455
rect 19800 27412 19852 27421
rect 9588 27344 9640 27396
rect 13084 27387 13136 27396
rect 13084 27353 13093 27387
rect 13093 27353 13127 27387
rect 13127 27353 13136 27387
rect 13084 27344 13136 27353
rect 15384 27344 15436 27396
rect 15936 27387 15988 27396
rect 15936 27353 15945 27387
rect 15945 27353 15979 27387
rect 15979 27353 15988 27387
rect 15936 27344 15988 27353
rect 16120 27387 16172 27396
rect 16120 27353 16129 27387
rect 16129 27353 16163 27387
rect 16163 27353 16172 27387
rect 16120 27344 16172 27353
rect 16948 27344 17000 27396
rect 17224 27387 17276 27396
rect 17224 27353 17233 27387
rect 17233 27353 17267 27387
rect 17267 27353 17276 27387
rect 17224 27344 17276 27353
rect 17408 27344 17460 27396
rect 19984 27344 20036 27396
rect 6920 27276 6972 27328
rect 11244 27276 11296 27328
rect 15108 27276 15160 27328
rect 16396 27276 16448 27328
rect 20444 27480 20496 27532
rect 22928 27548 22980 27600
rect 26792 27548 26844 27600
rect 27804 27548 27856 27600
rect 25412 27480 25464 27532
rect 26240 27480 26292 27532
rect 22192 27455 22244 27464
rect 22192 27421 22201 27455
rect 22201 27421 22235 27455
rect 22235 27421 22244 27455
rect 22192 27412 22244 27421
rect 25320 27412 25372 27464
rect 26792 27412 26844 27464
rect 27528 27480 27580 27532
rect 30472 27548 30524 27600
rect 31668 27548 31720 27600
rect 32036 27616 32088 27668
rect 32864 27616 32916 27668
rect 34060 27616 34112 27668
rect 34704 27659 34756 27668
rect 34704 27625 34713 27659
rect 34713 27625 34747 27659
rect 34747 27625 34756 27659
rect 34704 27616 34756 27625
rect 35164 27659 35216 27668
rect 35164 27625 35173 27659
rect 35173 27625 35207 27659
rect 35207 27625 35216 27659
rect 35164 27616 35216 27625
rect 35532 27659 35584 27668
rect 35532 27625 35541 27659
rect 35541 27625 35575 27659
rect 35575 27625 35584 27659
rect 35532 27616 35584 27625
rect 37188 27616 37240 27668
rect 29460 27480 29512 27532
rect 29736 27480 29788 27532
rect 27712 27412 27764 27464
rect 28816 27412 28868 27464
rect 21732 27344 21784 27396
rect 21916 27387 21968 27396
rect 21916 27353 21925 27387
rect 21925 27353 21959 27387
rect 21959 27353 21968 27387
rect 21916 27344 21968 27353
rect 23296 27344 23348 27396
rect 26240 27344 26292 27396
rect 26424 27344 26476 27396
rect 29552 27387 29604 27396
rect 29552 27353 29561 27387
rect 29561 27353 29595 27387
rect 29595 27353 29604 27387
rect 29552 27344 29604 27353
rect 20720 27276 20772 27328
rect 21088 27276 21140 27328
rect 22376 27276 22428 27328
rect 24400 27319 24452 27328
rect 24400 27285 24409 27319
rect 24409 27285 24443 27319
rect 24443 27285 24452 27319
rect 24400 27276 24452 27285
rect 24676 27276 24728 27328
rect 29092 27276 29144 27328
rect 29368 27276 29420 27328
rect 30932 27387 30984 27396
rect 30932 27353 30941 27387
rect 30941 27353 30975 27387
rect 30975 27353 30984 27387
rect 30932 27344 30984 27353
rect 31668 27412 31720 27464
rect 32404 27480 32456 27532
rect 32588 27480 32640 27532
rect 33048 27480 33100 27532
rect 33324 27523 33376 27532
rect 33324 27489 33333 27523
rect 33333 27489 33367 27523
rect 33367 27489 33376 27523
rect 33324 27480 33376 27489
rect 32128 27412 32180 27464
rect 33232 27412 33284 27464
rect 37372 27659 37424 27668
rect 37372 27625 37381 27659
rect 37381 27625 37415 27659
rect 37415 27625 37424 27659
rect 37372 27616 37424 27625
rect 34336 27480 34388 27532
rect 35348 27480 35400 27532
rect 40592 27616 40644 27668
rect 41236 27616 41288 27668
rect 42064 27659 42116 27668
rect 42064 27625 42073 27659
rect 42073 27625 42107 27659
rect 42107 27625 42116 27659
rect 42064 27616 42116 27625
rect 42432 27616 42484 27668
rect 34428 27344 34480 27396
rect 36728 27412 36780 27464
rect 37556 27455 37608 27464
rect 37556 27421 37565 27455
rect 37565 27421 37599 27455
rect 37599 27421 37608 27455
rect 37556 27412 37608 27421
rect 40408 27412 40460 27464
rect 36084 27344 36136 27396
rect 39580 27344 39632 27396
rect 42248 27455 42300 27464
rect 42248 27421 42257 27455
rect 42257 27421 42291 27455
rect 42291 27421 42300 27455
rect 42248 27412 42300 27421
rect 42340 27455 42392 27464
rect 42340 27421 42349 27455
rect 42349 27421 42383 27455
rect 42383 27421 42392 27455
rect 42340 27412 42392 27421
rect 42616 27455 42668 27464
rect 42616 27421 42625 27455
rect 42625 27421 42659 27455
rect 42659 27421 42668 27455
rect 42616 27412 42668 27421
rect 31484 27276 31536 27328
rect 32128 27319 32180 27328
rect 32128 27285 32137 27319
rect 32137 27285 32171 27319
rect 32171 27285 32180 27319
rect 32128 27276 32180 27285
rect 32588 27276 32640 27328
rect 32864 27276 32916 27328
rect 33048 27276 33100 27328
rect 34336 27276 34388 27328
rect 35808 27276 35860 27328
rect 41328 27276 41380 27328
rect 44456 27319 44508 27328
rect 44456 27285 44465 27319
rect 44465 27285 44499 27319
rect 44499 27285 44508 27319
rect 44456 27276 44508 27285
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 6000 27072 6052 27124
rect 8760 27072 8812 27124
rect 13268 27072 13320 27124
rect 8484 27004 8536 27056
rect 12992 27004 13044 27056
rect 6828 26936 6880 26988
rect 8208 26979 8260 26988
rect 8208 26945 8217 26979
rect 8217 26945 8251 26979
rect 8251 26945 8260 26979
rect 8208 26936 8260 26945
rect 10876 26936 10928 26988
rect 11428 26936 11480 26988
rect 13268 26979 13320 26988
rect 8392 26911 8444 26920
rect 8392 26877 8401 26911
rect 8401 26877 8435 26911
rect 8435 26877 8444 26911
rect 8392 26868 8444 26877
rect 13268 26945 13294 26979
rect 13294 26945 13320 26979
rect 13268 26936 13320 26945
rect 13636 27004 13688 27056
rect 15108 27072 15160 27124
rect 18052 27072 18104 27124
rect 19708 27115 19760 27124
rect 19708 27081 19717 27115
rect 19717 27081 19751 27115
rect 19751 27081 19760 27115
rect 19708 27072 19760 27081
rect 15476 27004 15528 27056
rect 20904 27047 20956 27056
rect 20904 27013 20913 27047
rect 20913 27013 20947 27047
rect 20947 27013 20956 27047
rect 20904 27004 20956 27013
rect 22192 27072 22244 27124
rect 24676 27072 24728 27124
rect 24400 27004 24452 27056
rect 25596 27072 25648 27124
rect 26056 27072 26108 27124
rect 26700 27115 26752 27124
rect 26700 27081 26709 27115
rect 26709 27081 26743 27115
rect 26743 27081 26752 27115
rect 26700 27072 26752 27081
rect 14740 26936 14792 26988
rect 15016 26936 15068 26988
rect 15200 26936 15252 26988
rect 15660 26936 15712 26988
rect 19524 26979 19576 26988
rect 19524 26945 19533 26979
rect 19533 26945 19567 26979
rect 19567 26945 19576 26979
rect 19524 26936 19576 26945
rect 20628 26979 20680 26988
rect 20628 26945 20637 26979
rect 20637 26945 20671 26979
rect 20671 26945 20680 26979
rect 20628 26936 20680 26945
rect 7196 26800 7248 26852
rect 17224 26868 17276 26920
rect 11428 26800 11480 26852
rect 11704 26800 11756 26852
rect 19432 26868 19484 26920
rect 24676 26936 24728 26988
rect 24768 26979 24820 26988
rect 24768 26945 24777 26979
rect 24777 26945 24811 26979
rect 24811 26945 24820 26979
rect 24768 26936 24820 26945
rect 21180 26868 21232 26920
rect 22376 26911 22428 26920
rect 22376 26877 22385 26911
rect 22385 26877 22419 26911
rect 22419 26877 22428 26911
rect 22376 26868 22428 26877
rect 23204 26868 23256 26920
rect 25964 27004 26016 27056
rect 27436 27115 27488 27124
rect 27436 27081 27445 27115
rect 27445 27081 27479 27115
rect 27479 27081 27488 27115
rect 27436 27072 27488 27081
rect 27804 27072 27856 27124
rect 33416 27072 33468 27124
rect 34520 27072 34572 27124
rect 37372 27072 37424 27124
rect 39580 27115 39632 27124
rect 39580 27081 39589 27115
rect 39589 27081 39623 27115
rect 39623 27081 39632 27115
rect 39580 27072 39632 27081
rect 41052 27072 41104 27124
rect 24952 26911 25004 26920
rect 24952 26877 24961 26911
rect 24961 26877 24995 26911
rect 24995 26877 25004 26911
rect 24952 26868 25004 26877
rect 25504 26911 25556 26920
rect 25504 26877 25513 26911
rect 25513 26877 25547 26911
rect 25547 26877 25556 26911
rect 25504 26868 25556 26877
rect 18604 26800 18656 26852
rect 7748 26732 7800 26784
rect 12256 26732 12308 26784
rect 13728 26732 13780 26784
rect 18512 26732 18564 26784
rect 19064 26732 19116 26784
rect 20444 26775 20496 26784
rect 20444 26741 20453 26775
rect 20453 26741 20487 26775
rect 20487 26741 20496 26775
rect 20444 26732 20496 26741
rect 23296 26800 23348 26852
rect 23940 26800 23992 26852
rect 25136 26800 25188 26852
rect 26424 26936 26476 26988
rect 27068 27004 27120 27056
rect 27620 27004 27672 27056
rect 31484 27004 31536 27056
rect 28448 26936 28500 26988
rect 29368 26936 29420 26988
rect 32128 26979 32180 26988
rect 32128 26945 32137 26979
rect 32137 26945 32171 26979
rect 32171 26945 32180 26979
rect 32128 26936 32180 26945
rect 32496 26936 32548 26988
rect 32588 26936 32640 26988
rect 34244 26936 34296 26988
rect 34336 26936 34388 26988
rect 34796 26936 34848 26988
rect 35256 27004 35308 27056
rect 35164 26979 35216 26988
rect 35164 26945 35173 26979
rect 35173 26945 35207 26979
rect 35207 26945 35216 26979
rect 35164 26936 35216 26945
rect 35440 26936 35492 26988
rect 38752 27004 38804 27056
rect 42432 27047 42484 27056
rect 42432 27013 42441 27047
rect 42441 27013 42475 27047
rect 42475 27013 42484 27047
rect 42432 27004 42484 27013
rect 39764 26979 39816 26988
rect 39764 26945 39773 26979
rect 39773 26945 39807 26979
rect 39807 26945 39816 26979
rect 39764 26936 39816 26945
rect 39856 26979 39908 26988
rect 39856 26945 39865 26979
rect 39865 26945 39899 26979
rect 39899 26945 39908 26979
rect 39856 26936 39908 26945
rect 40040 26979 40092 26988
rect 40040 26945 40049 26979
rect 40049 26945 40083 26979
rect 40083 26945 40092 26979
rect 40040 26936 40092 26945
rect 40408 26936 40460 26988
rect 40500 26979 40552 26988
rect 40500 26945 40509 26979
rect 40509 26945 40543 26979
rect 40543 26945 40552 26979
rect 40500 26936 40552 26945
rect 40776 26979 40828 26988
rect 40776 26945 40785 26979
rect 40785 26945 40819 26979
rect 40819 26945 40828 26979
rect 40776 26936 40828 26945
rect 40960 26979 41012 26988
rect 40960 26945 40969 26979
rect 40969 26945 41003 26979
rect 41003 26945 41012 26979
rect 40960 26936 41012 26945
rect 41052 26979 41104 26988
rect 41052 26945 41059 26979
rect 41059 26945 41093 26979
rect 41093 26945 41104 26979
rect 41052 26936 41104 26945
rect 26608 26800 26660 26852
rect 32036 26868 32088 26920
rect 34520 26911 34572 26920
rect 34520 26877 34529 26911
rect 34529 26877 34563 26911
rect 34563 26877 34572 26911
rect 34520 26868 34572 26877
rect 22560 26732 22612 26784
rect 24216 26732 24268 26784
rect 24584 26732 24636 26784
rect 25228 26732 25280 26784
rect 25596 26775 25648 26784
rect 25596 26741 25605 26775
rect 25605 26741 25639 26775
rect 25639 26741 25648 26775
rect 25596 26732 25648 26741
rect 25780 26775 25832 26784
rect 25780 26741 25789 26775
rect 25789 26741 25823 26775
rect 25823 26741 25832 26775
rect 25780 26732 25832 26741
rect 26240 26732 26292 26784
rect 27528 26800 27580 26852
rect 28356 26843 28408 26852
rect 28356 26809 28365 26843
rect 28365 26809 28399 26843
rect 28399 26809 28408 26843
rect 28356 26800 28408 26809
rect 29000 26843 29052 26852
rect 29000 26809 29009 26843
rect 29009 26809 29043 26843
rect 29043 26809 29052 26843
rect 29000 26800 29052 26809
rect 34888 26843 34940 26852
rect 34888 26809 34897 26843
rect 34897 26809 34931 26843
rect 34931 26809 34940 26843
rect 34888 26800 34940 26809
rect 27252 26775 27304 26784
rect 27252 26741 27261 26775
rect 27261 26741 27295 26775
rect 27295 26741 27304 26775
rect 27252 26732 27304 26741
rect 28264 26732 28316 26784
rect 31024 26732 31076 26784
rect 31392 26732 31444 26784
rect 31760 26732 31812 26784
rect 32588 26775 32640 26784
rect 32588 26741 32597 26775
rect 32597 26741 32631 26775
rect 32631 26741 32640 26775
rect 32588 26732 32640 26741
rect 33140 26732 33192 26784
rect 34520 26732 34572 26784
rect 37188 26868 37240 26920
rect 39948 26911 40000 26920
rect 39948 26877 39957 26911
rect 39957 26877 39991 26911
rect 39991 26877 40000 26911
rect 39948 26868 40000 26877
rect 40132 26868 40184 26920
rect 40684 26911 40736 26920
rect 40684 26877 40693 26911
rect 40693 26877 40727 26911
rect 40727 26877 40736 26911
rect 40684 26868 40736 26877
rect 41236 26911 41288 26920
rect 41236 26877 41245 26911
rect 41245 26877 41279 26911
rect 41279 26877 41288 26911
rect 41236 26868 41288 26877
rect 41328 26911 41380 26920
rect 41328 26877 41337 26911
rect 41337 26877 41371 26911
rect 41371 26877 41380 26911
rect 41328 26868 41380 26877
rect 35072 26800 35124 26852
rect 35440 26732 35492 26784
rect 36912 26732 36964 26784
rect 40316 26775 40368 26784
rect 40316 26741 40325 26775
rect 40325 26741 40359 26775
rect 40359 26741 40368 26775
rect 40316 26732 40368 26741
rect 40500 26732 40552 26784
rect 42248 26936 42300 26988
rect 42064 26868 42116 26920
rect 44272 26800 44324 26852
rect 42248 26732 42300 26784
rect 44456 26775 44508 26784
rect 44456 26741 44465 26775
rect 44465 26741 44499 26775
rect 44499 26741 44508 26775
rect 44456 26732 44508 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 10876 26528 10928 26580
rect 10968 26571 11020 26580
rect 10968 26537 10977 26571
rect 10977 26537 11011 26571
rect 11011 26537 11020 26571
rect 10968 26528 11020 26537
rect 9864 26460 9916 26512
rect 10324 26503 10376 26512
rect 10324 26469 10348 26503
rect 10348 26469 10376 26503
rect 10324 26460 10376 26469
rect 10416 26503 10468 26512
rect 10416 26469 10425 26503
rect 10425 26469 10459 26503
rect 10459 26469 10468 26503
rect 10416 26460 10468 26469
rect 11336 26528 11388 26580
rect 12624 26571 12676 26580
rect 12624 26537 12633 26571
rect 12633 26537 12667 26571
rect 12667 26537 12676 26571
rect 12624 26528 12676 26537
rect 14464 26528 14516 26580
rect 14832 26571 14884 26580
rect 14832 26537 14841 26571
rect 14841 26537 14875 26571
rect 14875 26537 14884 26571
rect 14832 26528 14884 26537
rect 10140 26392 10192 26444
rect 15476 26571 15528 26580
rect 15476 26537 15485 26571
rect 15485 26537 15519 26571
rect 15519 26537 15528 26571
rect 15476 26528 15528 26537
rect 15660 26571 15712 26580
rect 15660 26537 15669 26571
rect 15669 26537 15703 26571
rect 15703 26537 15712 26571
rect 15660 26528 15712 26537
rect 17040 26571 17092 26580
rect 17040 26537 17049 26571
rect 17049 26537 17083 26571
rect 17083 26537 17092 26571
rect 17040 26528 17092 26537
rect 11428 26392 11480 26444
rect 11704 26392 11756 26444
rect 12348 26435 12400 26444
rect 12348 26401 12357 26435
rect 12357 26401 12391 26435
rect 12391 26401 12400 26435
rect 12348 26392 12400 26401
rect 14004 26392 14056 26444
rect 14556 26392 14608 26444
rect 7932 26324 7984 26376
rect 10324 26324 10376 26376
rect 11152 26367 11204 26376
rect 11152 26333 11161 26367
rect 11161 26333 11195 26367
rect 11195 26333 11204 26367
rect 11152 26324 11204 26333
rect 6828 26256 6880 26308
rect 11612 26256 11664 26308
rect 11980 26324 12032 26376
rect 12256 26324 12308 26376
rect 13820 26324 13872 26376
rect 14648 26299 14700 26308
rect 14648 26265 14657 26299
rect 14657 26265 14691 26299
rect 14691 26265 14700 26299
rect 14648 26256 14700 26265
rect 14924 26367 14976 26376
rect 14924 26333 14933 26367
rect 14933 26333 14967 26367
rect 14967 26333 14976 26367
rect 14924 26324 14976 26333
rect 16948 26460 17000 26512
rect 15292 26435 15344 26444
rect 15292 26401 15301 26435
rect 15301 26401 15335 26435
rect 15335 26401 15344 26435
rect 15292 26392 15344 26401
rect 17960 26528 18012 26580
rect 18144 26571 18196 26580
rect 18144 26537 18153 26571
rect 18153 26537 18187 26571
rect 18187 26537 18196 26571
rect 18144 26528 18196 26537
rect 18880 26571 18932 26580
rect 18880 26537 18889 26571
rect 18889 26537 18923 26571
rect 18923 26537 18932 26571
rect 18880 26528 18932 26537
rect 19340 26528 19392 26580
rect 20904 26571 20956 26580
rect 20904 26537 20913 26571
rect 20913 26537 20947 26571
rect 20947 26537 20956 26571
rect 20904 26528 20956 26537
rect 22100 26528 22152 26580
rect 22192 26571 22244 26580
rect 22192 26537 22201 26571
rect 22201 26537 22235 26571
rect 22235 26537 22244 26571
rect 22192 26528 22244 26537
rect 23204 26528 23256 26580
rect 23756 26528 23808 26580
rect 25320 26571 25372 26580
rect 25320 26537 25329 26571
rect 25329 26537 25363 26571
rect 25363 26537 25372 26571
rect 25320 26528 25372 26537
rect 25412 26528 25464 26580
rect 26608 26528 26660 26580
rect 30380 26528 30432 26580
rect 31300 26528 31352 26580
rect 32036 26571 32088 26580
rect 32036 26537 32045 26571
rect 32045 26537 32079 26571
rect 32079 26537 32088 26571
rect 32036 26528 32088 26537
rect 17316 26503 17368 26512
rect 17316 26469 17325 26503
rect 17325 26469 17359 26503
rect 17359 26469 17368 26503
rect 17316 26460 17368 26469
rect 17592 26460 17644 26512
rect 21088 26460 21140 26512
rect 18788 26435 18840 26444
rect 18788 26401 18797 26435
rect 18797 26401 18831 26435
rect 18831 26401 18840 26435
rect 18788 26392 18840 26401
rect 19616 26392 19668 26444
rect 23940 26460 23992 26512
rect 24032 26460 24084 26512
rect 21824 26435 21876 26444
rect 21824 26401 21833 26435
rect 21833 26401 21867 26435
rect 21867 26401 21876 26435
rect 21824 26392 21876 26401
rect 22100 26392 22152 26444
rect 25964 26392 26016 26444
rect 26424 26460 26476 26512
rect 29460 26460 29512 26512
rect 32772 26528 32824 26580
rect 33140 26571 33192 26580
rect 33140 26537 33149 26571
rect 33149 26537 33183 26571
rect 33183 26537 33192 26571
rect 33140 26528 33192 26537
rect 35532 26528 35584 26580
rect 37188 26571 37240 26580
rect 37188 26537 37197 26571
rect 37197 26537 37231 26571
rect 37231 26537 37240 26571
rect 37188 26528 37240 26537
rect 37924 26528 37976 26580
rect 40684 26528 40736 26580
rect 42064 26571 42116 26580
rect 42064 26537 42073 26571
rect 42073 26537 42107 26571
rect 42107 26537 42116 26571
rect 42064 26528 42116 26537
rect 44272 26528 44324 26580
rect 27436 26392 27488 26444
rect 15476 26367 15528 26376
rect 15476 26333 15485 26367
rect 15485 26333 15519 26367
rect 15519 26333 15528 26367
rect 15476 26324 15528 26333
rect 16488 26324 16540 26376
rect 18512 26324 18564 26376
rect 20444 26367 20496 26376
rect 20444 26333 20453 26367
rect 20453 26333 20487 26367
rect 20487 26333 20496 26367
rect 20444 26324 20496 26333
rect 20628 26367 20680 26376
rect 20628 26333 20637 26367
rect 20637 26333 20671 26367
rect 20671 26333 20680 26367
rect 20628 26324 20680 26333
rect 20720 26367 20772 26376
rect 20720 26333 20729 26367
rect 20729 26333 20763 26367
rect 20763 26333 20772 26367
rect 20720 26324 20772 26333
rect 21364 26324 21416 26376
rect 19064 26256 19116 26308
rect 19708 26256 19760 26308
rect 10876 26188 10928 26240
rect 12532 26188 12584 26240
rect 12716 26188 12768 26240
rect 15752 26188 15804 26240
rect 18420 26188 18472 26240
rect 18512 26188 18564 26240
rect 24860 26324 24912 26376
rect 25320 26324 25372 26376
rect 25596 26324 25648 26376
rect 23756 26256 23808 26308
rect 26792 26324 26844 26376
rect 23480 26188 23532 26240
rect 30748 26324 30800 26376
rect 32588 26460 32640 26512
rect 31944 26392 31996 26444
rect 33140 26392 33192 26444
rect 31852 26367 31904 26376
rect 29552 26299 29604 26308
rect 29552 26265 29561 26299
rect 29561 26265 29595 26299
rect 29595 26265 29604 26299
rect 29552 26256 29604 26265
rect 31024 26256 31076 26308
rect 31852 26333 31861 26367
rect 31861 26333 31895 26367
rect 31895 26333 31904 26367
rect 31852 26324 31904 26333
rect 32680 26324 32732 26376
rect 33232 26367 33284 26376
rect 33232 26333 33241 26367
rect 33241 26333 33275 26367
rect 33275 26333 33284 26367
rect 33232 26324 33284 26333
rect 33416 26392 33468 26444
rect 36912 26392 36964 26444
rect 39120 26460 39172 26512
rect 44088 26460 44140 26512
rect 39948 26392 40000 26444
rect 40592 26392 40644 26444
rect 37464 26367 37516 26376
rect 37464 26333 37473 26367
rect 37473 26333 37507 26367
rect 37507 26333 37516 26367
rect 37464 26324 37516 26333
rect 40316 26324 40368 26376
rect 41696 26324 41748 26376
rect 42248 26324 42300 26376
rect 43720 26324 43772 26376
rect 31760 26256 31812 26308
rect 32036 26256 32088 26308
rect 32312 26256 32364 26308
rect 29736 26188 29788 26240
rect 30932 26188 30984 26240
rect 34704 26188 34756 26240
rect 35440 26188 35492 26240
rect 36912 26188 36964 26240
rect 40132 26256 40184 26308
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 5448 25984 5500 26036
rect 5356 25916 5408 25968
rect 10876 25984 10928 26036
rect 12440 26027 12492 26036
rect 12440 25993 12449 26027
rect 12449 25993 12483 26027
rect 12483 25993 12492 26027
rect 12440 25984 12492 25993
rect 13084 25984 13136 26036
rect 16488 26027 16540 26036
rect 16488 25993 16497 26027
rect 16497 25993 16531 26027
rect 16531 25993 16540 26027
rect 16488 25984 16540 25993
rect 17224 25984 17276 26036
rect 18512 25984 18564 26036
rect 21824 26027 21876 26036
rect 21824 25993 21833 26027
rect 21833 25993 21867 26027
rect 21867 25993 21876 26027
rect 21824 25984 21876 25993
rect 10508 25959 10560 25968
rect 10508 25925 10517 25959
rect 10517 25925 10551 25959
rect 10551 25925 10560 25959
rect 10508 25916 10560 25925
rect 5172 25848 5224 25900
rect 5448 25891 5500 25900
rect 5448 25857 5457 25891
rect 5457 25857 5491 25891
rect 5491 25857 5500 25891
rect 5448 25848 5500 25857
rect 7104 25848 7156 25900
rect 7748 25891 7800 25900
rect 7748 25857 7757 25891
rect 7757 25857 7791 25891
rect 7791 25857 7800 25891
rect 7748 25848 7800 25857
rect 7840 25848 7892 25900
rect 9220 25891 9272 25900
rect 9220 25857 9229 25891
rect 9229 25857 9263 25891
rect 9263 25857 9272 25891
rect 9220 25848 9272 25857
rect 9864 25848 9916 25900
rect 10232 25848 10284 25900
rect 10600 25891 10652 25900
rect 10600 25857 10609 25891
rect 10609 25857 10643 25891
rect 10643 25857 10652 25891
rect 10600 25848 10652 25857
rect 10876 25891 10928 25900
rect 10876 25857 10885 25891
rect 10885 25857 10919 25891
rect 10919 25857 10928 25891
rect 10876 25848 10928 25857
rect 11980 25891 12032 25900
rect 11980 25857 11989 25891
rect 11989 25857 12023 25891
rect 12023 25857 12032 25891
rect 11980 25848 12032 25857
rect 12256 25891 12308 25900
rect 12256 25857 12265 25891
rect 12265 25857 12299 25891
rect 12299 25857 12308 25891
rect 12256 25848 12308 25857
rect 7656 25780 7708 25832
rect 7932 25823 7984 25832
rect 7932 25789 7941 25823
rect 7941 25789 7975 25823
rect 7975 25789 7984 25823
rect 7932 25780 7984 25789
rect 9036 25823 9088 25832
rect 9036 25789 9045 25823
rect 9045 25789 9079 25823
rect 9079 25789 9088 25823
rect 9036 25780 9088 25789
rect 10692 25823 10744 25832
rect 10692 25789 10701 25823
rect 10701 25789 10735 25823
rect 10735 25789 10744 25823
rect 10692 25780 10744 25789
rect 12532 25916 12584 25968
rect 19340 25916 19392 25968
rect 23756 25959 23808 25968
rect 23756 25925 23765 25959
rect 23765 25925 23799 25959
rect 23799 25925 23808 25959
rect 23756 25916 23808 25925
rect 25044 25984 25096 26036
rect 25412 25984 25464 26036
rect 25596 25984 25648 26036
rect 24860 25916 24912 25968
rect 12900 25891 12952 25900
rect 12900 25857 12909 25891
rect 12909 25857 12943 25891
rect 12943 25857 12952 25891
rect 12900 25848 12952 25857
rect 13084 25848 13136 25900
rect 13636 25848 13688 25900
rect 14740 25891 14792 25900
rect 14740 25857 14749 25891
rect 14749 25857 14783 25891
rect 14783 25857 14792 25891
rect 14740 25848 14792 25857
rect 14832 25848 14884 25900
rect 15752 25848 15804 25900
rect 16028 25848 16080 25900
rect 12992 25823 13044 25832
rect 12992 25789 13001 25823
rect 13001 25789 13035 25823
rect 13035 25789 13044 25823
rect 12992 25780 13044 25789
rect 20720 25848 20772 25900
rect 22652 25848 22704 25900
rect 23296 25848 23348 25900
rect 23480 25891 23532 25900
rect 23480 25857 23489 25891
rect 23489 25857 23523 25891
rect 23523 25857 23532 25891
rect 23480 25848 23532 25857
rect 18880 25780 18932 25832
rect 22100 25823 22152 25832
rect 22100 25789 22109 25823
rect 22109 25789 22143 25823
rect 22143 25789 22152 25823
rect 22100 25780 22152 25789
rect 23664 25848 23716 25900
rect 10324 25712 10376 25764
rect 10876 25712 10928 25764
rect 15108 25712 15160 25764
rect 19524 25712 19576 25764
rect 8208 25644 8260 25696
rect 10048 25644 10100 25696
rect 10140 25644 10192 25696
rect 11888 25644 11940 25696
rect 13176 25644 13228 25696
rect 13268 25687 13320 25696
rect 13268 25653 13277 25687
rect 13277 25653 13311 25687
rect 13311 25653 13320 25687
rect 13268 25644 13320 25653
rect 15200 25644 15252 25696
rect 22376 25644 22428 25696
rect 22836 25644 22888 25696
rect 23204 25644 23256 25696
rect 23756 25644 23808 25696
rect 24400 25780 24452 25832
rect 24768 25891 24820 25900
rect 24768 25857 24777 25891
rect 24777 25857 24811 25891
rect 24811 25857 24820 25891
rect 24768 25848 24820 25857
rect 24952 25848 25004 25900
rect 26240 25848 26292 25900
rect 26608 25891 26660 25900
rect 26608 25857 26617 25891
rect 26617 25857 26651 25891
rect 26651 25857 26660 25891
rect 26608 25848 26660 25857
rect 26792 25891 26844 25900
rect 26792 25857 26801 25891
rect 26801 25857 26835 25891
rect 26835 25857 26844 25891
rect 26792 25848 26844 25857
rect 32036 25984 32088 26036
rect 32772 25984 32824 26036
rect 31944 25916 31996 25968
rect 34796 26027 34848 26036
rect 34796 25993 34805 26027
rect 34805 25993 34839 26027
rect 34839 25993 34848 26027
rect 34796 25984 34848 25993
rect 36636 25984 36688 26036
rect 36912 25984 36964 26036
rect 37096 25984 37148 26036
rect 37464 25984 37516 26036
rect 29184 25848 29236 25900
rect 32864 25891 32916 25900
rect 32864 25857 32873 25891
rect 32873 25857 32907 25891
rect 32907 25857 32916 25891
rect 32864 25848 32916 25857
rect 25596 25780 25648 25832
rect 26056 25780 26108 25832
rect 31484 25780 31536 25832
rect 32036 25780 32088 25832
rect 33140 25780 33192 25832
rect 31944 25712 31996 25764
rect 34428 25891 34480 25900
rect 34428 25857 34437 25891
rect 34437 25857 34471 25891
rect 34471 25857 34480 25891
rect 34428 25848 34480 25857
rect 36084 25848 36136 25900
rect 37464 25891 37516 25900
rect 37464 25857 37473 25891
rect 37473 25857 37507 25891
rect 37507 25857 37516 25891
rect 37464 25848 37516 25857
rect 35164 25780 35216 25832
rect 24400 25644 24452 25696
rect 24492 25687 24544 25696
rect 24492 25653 24501 25687
rect 24501 25653 24535 25687
rect 24535 25653 24544 25687
rect 24492 25644 24544 25653
rect 25044 25644 25096 25696
rect 27620 25644 27672 25696
rect 28264 25644 28316 25696
rect 28540 25644 28592 25696
rect 29552 25644 29604 25696
rect 32312 25644 32364 25696
rect 33416 25644 33468 25696
rect 33600 25644 33652 25696
rect 34152 25687 34204 25696
rect 34152 25653 34161 25687
rect 34161 25653 34195 25687
rect 34195 25653 34204 25687
rect 34152 25644 34204 25653
rect 34520 25644 34572 25696
rect 36452 25712 36504 25764
rect 37280 25712 37332 25764
rect 38568 25848 38620 25900
rect 37924 25780 37976 25832
rect 35440 25644 35492 25696
rect 37464 25644 37516 25696
rect 38384 25687 38436 25696
rect 38384 25653 38393 25687
rect 38393 25653 38427 25687
rect 38427 25653 38436 25687
rect 38384 25644 38436 25653
rect 39120 25959 39172 25968
rect 39120 25925 39129 25959
rect 39129 25925 39163 25959
rect 39163 25925 39172 25959
rect 39120 25916 39172 25925
rect 39856 25848 39908 25900
rect 41696 25916 41748 25968
rect 40592 25848 40644 25900
rect 41512 25712 41564 25764
rect 40684 25644 40736 25696
rect 44180 25780 44232 25832
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 5264 25483 5316 25492
rect 5264 25449 5273 25483
rect 5273 25449 5307 25483
rect 5307 25449 5316 25483
rect 5264 25440 5316 25449
rect 5724 25483 5776 25492
rect 5724 25449 5733 25483
rect 5733 25449 5767 25483
rect 5767 25449 5776 25483
rect 5724 25440 5776 25449
rect 10048 25440 10100 25492
rect 11704 25372 11756 25424
rect 12256 25372 12308 25424
rect 16028 25372 16080 25424
rect 16304 25440 16356 25492
rect 19524 25483 19576 25492
rect 19524 25449 19533 25483
rect 19533 25449 19567 25483
rect 19567 25449 19576 25483
rect 19524 25440 19576 25449
rect 19708 25483 19760 25492
rect 19708 25449 19717 25483
rect 19717 25449 19751 25483
rect 19751 25449 19760 25483
rect 19708 25440 19760 25449
rect 19800 25440 19852 25492
rect 20628 25440 20680 25492
rect 22376 25440 22428 25492
rect 22560 25440 22612 25492
rect 17684 25372 17736 25424
rect 19616 25372 19668 25424
rect 19984 25372 20036 25424
rect 20536 25372 20588 25424
rect 23756 25483 23808 25492
rect 23756 25449 23765 25483
rect 23765 25449 23799 25483
rect 23799 25449 23808 25483
rect 23756 25440 23808 25449
rect 24860 25440 24912 25492
rect 25044 25483 25096 25492
rect 25044 25449 25053 25483
rect 25053 25449 25087 25483
rect 25087 25449 25096 25483
rect 25044 25440 25096 25449
rect 25504 25483 25556 25492
rect 25504 25449 25513 25483
rect 25513 25449 25547 25483
rect 25547 25449 25556 25483
rect 25504 25440 25556 25449
rect 25596 25440 25648 25492
rect 29828 25483 29880 25492
rect 29828 25449 29837 25483
rect 29837 25449 29871 25483
rect 29871 25449 29880 25483
rect 29828 25440 29880 25449
rect 30104 25440 30156 25492
rect 24768 25372 24820 25424
rect 5632 25347 5684 25356
rect 5632 25313 5641 25347
rect 5641 25313 5675 25347
rect 5675 25313 5684 25347
rect 5632 25304 5684 25313
rect 12992 25304 13044 25356
rect 17316 25304 17368 25356
rect 10232 25236 10284 25288
rect 10416 25279 10468 25288
rect 10416 25245 10425 25279
rect 10425 25245 10459 25279
rect 10459 25245 10468 25279
rect 10416 25236 10468 25245
rect 10508 25236 10560 25288
rect 19432 25304 19484 25356
rect 19800 25304 19852 25356
rect 20352 25304 20404 25356
rect 10324 25168 10376 25220
rect 17684 25236 17736 25288
rect 16120 25211 16172 25220
rect 16120 25177 16129 25211
rect 16129 25177 16163 25211
rect 16163 25177 16172 25211
rect 16120 25168 16172 25177
rect 16304 25211 16356 25220
rect 16304 25177 16313 25211
rect 16313 25177 16347 25211
rect 16347 25177 16356 25211
rect 16304 25168 16356 25177
rect 5908 25100 5960 25152
rect 9220 25100 9272 25152
rect 10048 25100 10100 25152
rect 11612 25100 11664 25152
rect 14280 25100 14332 25152
rect 15660 25100 15712 25152
rect 19524 25279 19576 25288
rect 19524 25245 19533 25279
rect 19533 25245 19567 25279
rect 19567 25245 19576 25279
rect 19524 25236 19576 25245
rect 21088 25304 21140 25356
rect 21456 25304 21508 25356
rect 23388 25347 23440 25356
rect 23388 25313 23397 25347
rect 23397 25313 23431 25347
rect 23431 25313 23440 25347
rect 23388 25304 23440 25313
rect 16488 25143 16540 25152
rect 16488 25109 16497 25143
rect 16497 25109 16531 25143
rect 16531 25109 16540 25143
rect 16488 25100 16540 25109
rect 19616 25100 19668 25152
rect 20536 25168 20588 25220
rect 23572 25279 23624 25288
rect 23572 25245 23581 25279
rect 23581 25245 23615 25279
rect 23615 25245 23624 25279
rect 23572 25236 23624 25245
rect 24952 25236 25004 25288
rect 25320 25279 25372 25288
rect 25320 25245 25329 25279
rect 25329 25245 25363 25279
rect 25363 25245 25372 25279
rect 25320 25236 25372 25245
rect 25780 25236 25832 25288
rect 28632 25415 28684 25424
rect 28632 25381 28641 25415
rect 28641 25381 28675 25415
rect 28675 25381 28684 25415
rect 28632 25372 28684 25381
rect 29920 25372 29972 25424
rect 26516 25304 26568 25356
rect 29552 25279 29604 25288
rect 29552 25245 29561 25279
rect 29561 25245 29595 25279
rect 29595 25245 29604 25279
rect 29552 25236 29604 25245
rect 29736 25279 29788 25288
rect 29736 25245 29745 25279
rect 29745 25245 29779 25279
rect 29779 25245 29788 25279
rect 29736 25236 29788 25245
rect 30104 25304 30156 25356
rect 30288 25304 30340 25356
rect 31116 25440 31168 25492
rect 32036 25483 32088 25492
rect 32036 25449 32045 25483
rect 32045 25449 32079 25483
rect 32079 25449 32088 25483
rect 32036 25440 32088 25449
rect 33416 25440 33468 25492
rect 33692 25440 33744 25492
rect 34152 25440 34204 25492
rect 35164 25483 35216 25492
rect 35164 25449 35173 25483
rect 35173 25449 35207 25483
rect 35207 25449 35216 25483
rect 35164 25440 35216 25449
rect 36452 25440 36504 25492
rect 37556 25440 37608 25492
rect 40592 25440 40644 25492
rect 31392 25372 31444 25424
rect 22284 25168 22336 25220
rect 26148 25168 26200 25220
rect 28448 25211 28500 25220
rect 28448 25177 28457 25211
rect 28457 25177 28491 25211
rect 28491 25177 28500 25211
rect 28448 25168 28500 25177
rect 28908 25211 28960 25220
rect 28908 25177 28917 25211
rect 28917 25177 28951 25211
rect 28951 25177 28960 25211
rect 28908 25168 28960 25177
rect 29092 25211 29144 25220
rect 29092 25177 29101 25211
rect 29101 25177 29135 25211
rect 29135 25177 29144 25211
rect 29092 25168 29144 25177
rect 30932 25236 30984 25288
rect 31760 25347 31812 25356
rect 31760 25313 31769 25347
rect 31769 25313 31803 25347
rect 31803 25313 31812 25347
rect 31760 25304 31812 25313
rect 33692 25304 33744 25356
rect 31484 25236 31536 25288
rect 23204 25100 23256 25152
rect 25228 25100 25280 25152
rect 25320 25100 25372 25152
rect 25412 25100 25464 25152
rect 26056 25100 26108 25152
rect 26240 25100 26292 25152
rect 26976 25100 27028 25152
rect 27436 25100 27488 25152
rect 27528 25100 27580 25152
rect 30012 25143 30064 25152
rect 30012 25109 30021 25143
rect 30021 25109 30055 25143
rect 30055 25109 30064 25143
rect 30012 25100 30064 25109
rect 31392 25168 31444 25220
rect 32220 25236 32272 25288
rect 32772 25168 32824 25220
rect 37740 25372 37792 25424
rect 40684 25415 40736 25424
rect 40684 25381 40693 25415
rect 40693 25381 40727 25415
rect 40727 25381 40736 25415
rect 40684 25372 40736 25381
rect 34520 25304 34572 25356
rect 34888 25236 34940 25288
rect 36176 25236 36228 25288
rect 36912 25304 36964 25356
rect 40868 25347 40920 25356
rect 40868 25313 40877 25347
rect 40877 25313 40911 25347
rect 40911 25313 40920 25347
rect 40868 25304 40920 25313
rect 43720 25347 43772 25356
rect 43720 25313 43729 25347
rect 43729 25313 43763 25347
rect 43763 25313 43772 25347
rect 43720 25304 43772 25313
rect 36636 25279 36688 25288
rect 36636 25245 36645 25279
rect 36645 25245 36679 25279
rect 36679 25245 36688 25279
rect 36636 25236 36688 25245
rect 34060 25100 34112 25152
rect 39304 25236 39356 25288
rect 39764 25236 39816 25288
rect 41512 25236 41564 25288
rect 41696 25236 41748 25288
rect 40868 25100 40920 25152
rect 42800 25236 42852 25288
rect 44272 25279 44324 25288
rect 44272 25245 44281 25279
rect 44281 25245 44315 25279
rect 44315 25245 44324 25279
rect 44272 25236 44324 25245
rect 43168 25168 43220 25220
rect 43812 25211 43864 25220
rect 43812 25177 43821 25211
rect 43821 25177 43855 25211
rect 43855 25177 43864 25211
rect 43812 25168 43864 25177
rect 42984 25143 43036 25152
rect 42984 25109 42993 25143
rect 42993 25109 43027 25143
rect 43027 25109 43036 25143
rect 42984 25100 43036 25109
rect 43076 25143 43128 25152
rect 43076 25109 43085 25143
rect 43085 25109 43119 25143
rect 43119 25109 43128 25143
rect 43076 25100 43128 25109
rect 44456 25143 44508 25152
rect 44456 25109 44465 25143
rect 44465 25109 44499 25143
rect 44499 25109 44508 25143
rect 44456 25100 44508 25109
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 5632 24896 5684 24948
rect 13636 24896 13688 24948
rect 15660 24896 15712 24948
rect 16488 24896 16540 24948
rect 6000 24803 6052 24812
rect 6000 24769 6009 24803
rect 6009 24769 6043 24803
rect 6043 24769 6052 24803
rect 6000 24760 6052 24769
rect 6184 24803 6236 24812
rect 6184 24769 6193 24803
rect 6193 24769 6227 24803
rect 6227 24769 6236 24803
rect 6184 24760 6236 24769
rect 6828 24760 6880 24812
rect 10048 24803 10100 24812
rect 10048 24769 10057 24803
rect 10057 24769 10091 24803
rect 10091 24769 10100 24803
rect 10048 24760 10100 24769
rect 19340 24828 19392 24880
rect 20536 24896 20588 24948
rect 24400 24896 24452 24948
rect 24860 24896 24912 24948
rect 26516 24896 26568 24948
rect 29460 24896 29512 24948
rect 30104 24896 30156 24948
rect 31760 24896 31812 24948
rect 32312 24896 32364 24948
rect 32772 24896 32824 24948
rect 8024 24692 8076 24744
rect 8760 24735 8812 24744
rect 8760 24701 8769 24735
rect 8769 24701 8803 24735
rect 8803 24701 8812 24735
rect 8760 24692 8812 24701
rect 10140 24735 10192 24744
rect 10140 24701 10149 24735
rect 10149 24701 10183 24735
rect 10183 24701 10192 24735
rect 10140 24692 10192 24701
rect 11612 24692 11664 24744
rect 11980 24735 12032 24744
rect 11980 24701 11989 24735
rect 11989 24701 12023 24735
rect 12023 24701 12032 24735
rect 11980 24692 12032 24701
rect 13636 24760 13688 24812
rect 13820 24760 13872 24812
rect 14372 24760 14424 24812
rect 15936 24760 15988 24812
rect 16396 24760 16448 24812
rect 17224 24760 17276 24812
rect 17592 24803 17644 24812
rect 17592 24769 17601 24803
rect 17601 24769 17635 24803
rect 17635 24769 17644 24803
rect 17592 24760 17644 24769
rect 17684 24760 17736 24812
rect 18236 24760 18288 24812
rect 18512 24760 18564 24812
rect 19616 24803 19668 24812
rect 19616 24769 19625 24803
rect 19625 24769 19659 24803
rect 19659 24769 19668 24803
rect 19616 24760 19668 24769
rect 19708 24803 19760 24812
rect 19708 24769 19717 24803
rect 19717 24769 19751 24803
rect 19751 24769 19760 24803
rect 19708 24760 19760 24769
rect 24768 24828 24820 24880
rect 20168 24760 20220 24812
rect 16580 24692 16632 24744
rect 16764 24692 16816 24744
rect 13360 24624 13412 24676
rect 13912 24624 13964 24676
rect 17776 24667 17828 24676
rect 17776 24633 17785 24667
rect 17785 24633 17819 24667
rect 17819 24633 17828 24667
rect 17776 24624 17828 24633
rect 17960 24735 18012 24744
rect 17960 24701 17969 24735
rect 17969 24701 18003 24735
rect 18003 24701 18012 24735
rect 17960 24692 18012 24701
rect 18604 24692 18656 24744
rect 20628 24760 20680 24812
rect 22560 24803 22612 24812
rect 22560 24769 22569 24803
rect 22569 24769 22603 24803
rect 22603 24769 22612 24803
rect 22560 24760 22612 24769
rect 22928 24760 22980 24812
rect 26332 24828 26384 24880
rect 27804 24828 27856 24880
rect 28448 24828 28500 24880
rect 8300 24556 8352 24608
rect 8668 24599 8720 24608
rect 8668 24565 8677 24599
rect 8677 24565 8711 24599
rect 8711 24565 8720 24599
rect 8668 24556 8720 24565
rect 9588 24556 9640 24608
rect 9680 24556 9732 24608
rect 9956 24556 10008 24608
rect 10324 24556 10376 24608
rect 11796 24556 11848 24608
rect 14372 24599 14424 24608
rect 14372 24565 14381 24599
rect 14381 24565 14415 24599
rect 14415 24565 14424 24599
rect 14372 24556 14424 24565
rect 16488 24556 16540 24608
rect 17868 24599 17920 24608
rect 17868 24565 17877 24599
rect 17877 24565 17911 24599
rect 17911 24565 17920 24599
rect 17868 24556 17920 24565
rect 18236 24667 18288 24676
rect 18236 24633 18245 24667
rect 18245 24633 18279 24667
rect 18279 24633 18288 24667
rect 18236 24624 18288 24633
rect 18696 24624 18748 24676
rect 21272 24692 21324 24744
rect 25780 24692 25832 24744
rect 31116 24760 31168 24812
rect 31668 24760 31720 24812
rect 32496 24803 32548 24812
rect 32496 24769 32505 24803
rect 32505 24769 32539 24803
rect 32539 24769 32548 24803
rect 32496 24760 32548 24769
rect 26332 24735 26384 24744
rect 26332 24701 26341 24735
rect 26341 24701 26375 24735
rect 26375 24701 26384 24735
rect 26332 24692 26384 24701
rect 26792 24692 26844 24744
rect 31944 24692 31996 24744
rect 26056 24667 26108 24676
rect 26056 24633 26065 24667
rect 26065 24633 26099 24667
rect 26099 24633 26108 24667
rect 26056 24624 26108 24633
rect 19708 24556 19760 24608
rect 20168 24556 20220 24608
rect 21180 24556 21232 24608
rect 22744 24599 22796 24608
rect 22744 24565 22753 24599
rect 22753 24565 22787 24599
rect 22787 24565 22796 24599
rect 22744 24556 22796 24565
rect 22836 24556 22888 24608
rect 26976 24624 27028 24676
rect 27160 24624 27212 24676
rect 27896 24624 27948 24676
rect 30748 24624 30800 24676
rect 31024 24624 31076 24676
rect 26516 24556 26568 24608
rect 27252 24556 27304 24608
rect 28264 24556 28316 24608
rect 32312 24624 32364 24676
rect 32036 24556 32088 24608
rect 32956 24760 33008 24812
rect 34152 24896 34204 24948
rect 35164 24896 35216 24948
rect 41972 24896 42024 24948
rect 43720 24896 43772 24948
rect 33600 24828 33652 24880
rect 33876 24828 33928 24880
rect 33692 24760 33744 24812
rect 35532 24828 35584 24880
rect 35440 24760 35492 24812
rect 38844 24803 38896 24812
rect 38844 24769 38853 24803
rect 38853 24769 38887 24803
rect 38887 24769 38896 24803
rect 38844 24760 38896 24769
rect 32772 24624 32824 24676
rect 35992 24692 36044 24744
rect 38752 24735 38804 24744
rect 38752 24701 38761 24735
rect 38761 24701 38795 24735
rect 38795 24701 38804 24735
rect 38752 24692 38804 24701
rect 41236 24692 41288 24744
rect 41604 24760 41656 24812
rect 42984 24760 43036 24812
rect 33324 24624 33376 24676
rect 33692 24624 33744 24676
rect 36268 24624 36320 24676
rect 36728 24624 36780 24676
rect 41604 24624 41656 24676
rect 41880 24692 41932 24744
rect 32956 24599 33008 24608
rect 32956 24565 32965 24599
rect 32965 24565 32999 24599
rect 32999 24565 33008 24599
rect 32956 24556 33008 24565
rect 33784 24556 33836 24608
rect 35716 24556 35768 24608
rect 38292 24556 38344 24608
rect 39120 24556 39172 24608
rect 43076 24556 43128 24608
rect 44456 24599 44508 24608
rect 44456 24565 44465 24599
rect 44465 24565 44499 24599
rect 44499 24565 44508 24599
rect 44456 24556 44508 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 9680 24352 9732 24404
rect 9772 24352 9824 24404
rect 9956 24395 10008 24404
rect 9956 24361 9965 24395
rect 9965 24361 9999 24395
rect 9999 24361 10008 24395
rect 9956 24352 10008 24361
rect 11704 24352 11756 24404
rect 12808 24395 12860 24404
rect 12808 24361 12817 24395
rect 12817 24361 12851 24395
rect 12851 24361 12860 24395
rect 12808 24352 12860 24361
rect 13360 24395 13412 24404
rect 13360 24361 13369 24395
rect 13369 24361 13403 24395
rect 13403 24361 13412 24395
rect 13360 24352 13412 24361
rect 13820 24352 13872 24404
rect 14188 24352 14240 24404
rect 14372 24352 14424 24404
rect 5448 24284 5500 24336
rect 7288 24216 7340 24268
rect 10048 24259 10100 24268
rect 10048 24225 10057 24259
rect 10057 24225 10091 24259
rect 10091 24225 10100 24259
rect 10048 24216 10100 24225
rect 7472 24148 7524 24200
rect 10416 24216 10468 24268
rect 10692 24259 10744 24268
rect 10692 24225 10701 24259
rect 10701 24225 10735 24259
rect 10735 24225 10744 24259
rect 10692 24216 10744 24225
rect 7748 24080 7800 24132
rect 10324 24148 10376 24200
rect 10876 24216 10928 24268
rect 2780 24012 2832 24064
rect 9772 24080 9824 24132
rect 11612 24284 11664 24336
rect 11796 24284 11848 24336
rect 14924 24284 14976 24336
rect 15476 24352 15528 24404
rect 16304 24395 16356 24404
rect 16304 24361 16313 24395
rect 16313 24361 16347 24395
rect 16347 24361 16356 24395
rect 16304 24352 16356 24361
rect 16488 24395 16540 24404
rect 16488 24361 16497 24395
rect 16497 24361 16531 24395
rect 16531 24361 16540 24395
rect 16488 24352 16540 24361
rect 16948 24395 17000 24404
rect 16948 24361 16957 24395
rect 16957 24361 16991 24395
rect 16991 24361 17000 24395
rect 16948 24352 17000 24361
rect 17224 24395 17276 24404
rect 17224 24361 17233 24395
rect 17233 24361 17267 24395
rect 17267 24361 17276 24395
rect 17224 24352 17276 24361
rect 14096 24216 14148 24268
rect 14188 24216 14240 24268
rect 14832 24216 14884 24268
rect 12716 24191 12768 24200
rect 12716 24157 12725 24191
rect 12725 24157 12759 24191
rect 12759 24157 12768 24191
rect 12716 24148 12768 24157
rect 12900 24191 12952 24200
rect 12900 24157 12909 24191
rect 12909 24157 12943 24191
rect 12943 24157 12952 24191
rect 12900 24148 12952 24157
rect 15108 24191 15160 24200
rect 15108 24157 15117 24191
rect 15117 24157 15151 24191
rect 15151 24157 15160 24191
rect 15108 24148 15160 24157
rect 15936 24216 15988 24268
rect 16396 24216 16448 24268
rect 16856 24259 16908 24268
rect 16856 24225 16865 24259
rect 16865 24225 16899 24259
rect 16899 24225 16908 24259
rect 16856 24216 16908 24225
rect 8116 24012 8168 24064
rect 9864 24012 9916 24064
rect 10324 24012 10376 24064
rect 10600 24080 10652 24132
rect 10968 24055 11020 24064
rect 10968 24021 10977 24055
rect 10977 24021 11011 24055
rect 11011 24021 11020 24055
rect 10968 24012 11020 24021
rect 14280 24080 14332 24132
rect 14556 24123 14608 24132
rect 14556 24089 14565 24123
rect 14565 24089 14599 24123
rect 14599 24089 14608 24123
rect 14556 24080 14608 24089
rect 16212 24080 16264 24132
rect 16580 24148 16632 24200
rect 17224 24216 17276 24268
rect 17684 24216 17736 24268
rect 17500 24148 17552 24200
rect 17868 24148 17920 24200
rect 18236 24395 18288 24404
rect 18236 24361 18245 24395
rect 18245 24361 18279 24395
rect 18279 24361 18288 24395
rect 18236 24352 18288 24361
rect 18788 24352 18840 24404
rect 19800 24352 19852 24404
rect 20076 24352 20128 24404
rect 20260 24352 20312 24404
rect 22836 24395 22888 24404
rect 22836 24361 22845 24395
rect 22845 24361 22879 24395
rect 22879 24361 22888 24395
rect 22836 24352 22888 24361
rect 23848 24352 23900 24404
rect 24124 24352 24176 24404
rect 27896 24352 27948 24404
rect 19064 24284 19116 24336
rect 18052 24216 18104 24268
rect 18328 24216 18380 24268
rect 19800 24216 19852 24268
rect 21456 24216 21508 24268
rect 21548 24216 21600 24268
rect 22284 24216 22336 24268
rect 23112 24284 23164 24336
rect 24768 24284 24820 24336
rect 25596 24284 25648 24336
rect 27528 24284 27580 24336
rect 27620 24284 27672 24336
rect 28264 24395 28316 24404
rect 28264 24361 28273 24395
rect 28273 24361 28307 24395
rect 28307 24361 28316 24395
rect 28264 24352 28316 24361
rect 29276 24352 29328 24404
rect 29828 24352 29880 24404
rect 30748 24352 30800 24404
rect 28080 24284 28132 24336
rect 31760 24395 31812 24404
rect 31760 24361 31769 24395
rect 31769 24361 31803 24395
rect 31803 24361 31812 24395
rect 31760 24352 31812 24361
rect 31944 24352 31996 24404
rect 33324 24352 33376 24404
rect 33876 24352 33928 24404
rect 34336 24352 34388 24404
rect 34428 24352 34480 24404
rect 23204 24216 23256 24268
rect 16672 24080 16724 24132
rect 17776 24080 17828 24132
rect 18512 24080 18564 24132
rect 18880 24080 18932 24132
rect 21180 24080 21232 24132
rect 22652 24080 22704 24132
rect 22836 24191 22888 24200
rect 22836 24157 22845 24191
rect 22845 24157 22879 24191
rect 22879 24157 22888 24191
rect 22836 24148 22888 24157
rect 23020 24148 23072 24200
rect 23572 24216 23624 24268
rect 24676 24216 24728 24268
rect 25228 24216 25280 24268
rect 30104 24216 30156 24268
rect 24860 24148 24912 24200
rect 27620 24148 27672 24200
rect 27988 24191 28040 24200
rect 27988 24157 27997 24191
rect 27997 24157 28031 24191
rect 28031 24157 28040 24191
rect 27988 24148 28040 24157
rect 23848 24080 23900 24132
rect 25136 24080 25188 24132
rect 26056 24080 26108 24132
rect 13820 24055 13872 24064
rect 13820 24021 13829 24055
rect 13829 24021 13863 24055
rect 13863 24021 13872 24055
rect 13820 24012 13872 24021
rect 14096 24012 14148 24064
rect 16948 24012 17000 24064
rect 17224 24012 17276 24064
rect 19432 24012 19484 24064
rect 19708 24012 19760 24064
rect 23388 24012 23440 24064
rect 24124 24012 24176 24064
rect 24400 24012 24452 24064
rect 24492 24012 24544 24064
rect 24768 24012 24820 24064
rect 24952 24012 25004 24064
rect 26424 24080 26476 24132
rect 26884 24080 26936 24132
rect 27160 24080 27212 24132
rect 27896 24080 27948 24132
rect 28356 24191 28408 24200
rect 28356 24157 28365 24191
rect 28365 24157 28399 24191
rect 28399 24157 28408 24191
rect 28356 24148 28408 24157
rect 28540 24191 28592 24200
rect 28540 24157 28549 24191
rect 28549 24157 28583 24191
rect 28583 24157 28592 24191
rect 28540 24148 28592 24157
rect 29552 24191 29604 24200
rect 29552 24157 29561 24191
rect 29561 24157 29595 24191
rect 29595 24157 29604 24191
rect 29552 24148 29604 24157
rect 30932 24216 30984 24268
rect 32128 24284 32180 24336
rect 32220 24284 32272 24336
rect 35624 24352 35676 24404
rect 31668 24216 31720 24268
rect 31852 24259 31904 24268
rect 31852 24225 31861 24259
rect 31861 24225 31895 24259
rect 31895 24225 31904 24259
rect 31852 24216 31904 24225
rect 32496 24216 32548 24268
rect 33876 24216 33928 24268
rect 33968 24216 34020 24268
rect 34980 24284 35032 24336
rect 29092 24080 29144 24132
rect 26332 24012 26384 24064
rect 32312 24148 32364 24200
rect 30104 24012 30156 24064
rect 34152 24012 34204 24064
rect 34612 24012 34664 24064
rect 34980 24191 35032 24200
rect 34980 24157 34989 24191
rect 34989 24157 35023 24191
rect 35023 24157 35032 24191
rect 34980 24148 35032 24157
rect 35716 24216 35768 24268
rect 42984 24259 43036 24268
rect 42984 24225 42993 24259
rect 42993 24225 43027 24259
rect 43027 24225 43036 24259
rect 42984 24216 43036 24225
rect 35440 24191 35492 24200
rect 35440 24157 35449 24191
rect 35449 24157 35483 24191
rect 35483 24157 35492 24191
rect 35440 24148 35492 24157
rect 35532 24191 35584 24200
rect 35532 24157 35541 24191
rect 35541 24157 35575 24191
rect 35575 24157 35584 24191
rect 35532 24148 35584 24157
rect 35624 24148 35676 24200
rect 36084 24148 36136 24200
rect 36268 24191 36320 24200
rect 36268 24157 36277 24191
rect 36277 24157 36311 24191
rect 36311 24157 36320 24191
rect 36268 24148 36320 24157
rect 36820 24148 36872 24200
rect 37740 24148 37792 24200
rect 40316 24148 40368 24200
rect 41788 24148 41840 24200
rect 37004 24080 37056 24132
rect 41052 24080 41104 24132
rect 36544 24012 36596 24064
rect 41880 24012 41932 24064
rect 42984 24012 43036 24064
rect 43628 24055 43680 24064
rect 43628 24021 43637 24055
rect 43637 24021 43671 24055
rect 43671 24021 43680 24055
rect 43628 24012 43680 24021
rect 44456 24055 44508 24064
rect 44456 24021 44465 24055
rect 44465 24021 44499 24055
rect 44499 24021 44508 24055
rect 44456 24012 44508 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 7196 23808 7248 23860
rect 7380 23851 7432 23860
rect 7380 23817 7389 23851
rect 7389 23817 7423 23851
rect 7423 23817 7432 23851
rect 7380 23808 7432 23817
rect 7472 23851 7524 23860
rect 7472 23817 7481 23851
rect 7481 23817 7515 23851
rect 7515 23817 7524 23851
rect 7472 23808 7524 23817
rect 9772 23808 9824 23860
rect 4620 23740 4672 23792
rect 6276 23740 6328 23792
rect 9680 23740 9732 23792
rect 4252 23672 4304 23724
rect 4436 23715 4488 23724
rect 4436 23681 4445 23715
rect 4445 23681 4479 23715
rect 4479 23681 4488 23715
rect 4436 23672 4488 23681
rect 3424 23604 3476 23656
rect 7288 23604 7340 23656
rect 7748 23647 7800 23656
rect 7748 23613 7757 23647
rect 7757 23613 7791 23647
rect 7791 23613 7800 23647
rect 7748 23604 7800 23613
rect 7932 23715 7984 23724
rect 7932 23681 7941 23715
rect 7941 23681 7975 23715
rect 7975 23681 7984 23715
rect 7932 23672 7984 23681
rect 8576 23604 8628 23656
rect 4436 23536 4488 23588
rect 4804 23536 4856 23588
rect 8024 23536 8076 23588
rect 8116 23536 8168 23588
rect 9772 23672 9824 23724
rect 9956 23672 10008 23724
rect 10324 23808 10376 23860
rect 10784 23808 10836 23860
rect 14280 23808 14332 23860
rect 14556 23808 14608 23860
rect 15660 23851 15712 23860
rect 15660 23817 15669 23851
rect 15669 23817 15703 23851
rect 15703 23817 15712 23851
rect 15660 23808 15712 23817
rect 16948 23808 17000 23860
rect 20076 23808 20128 23860
rect 20996 23808 21048 23860
rect 26976 23808 27028 23860
rect 27436 23808 27488 23860
rect 29000 23808 29052 23860
rect 29552 23808 29604 23860
rect 29920 23808 29972 23860
rect 30104 23808 30156 23860
rect 31852 23808 31904 23860
rect 10876 23740 10928 23792
rect 12716 23740 12768 23792
rect 10324 23672 10376 23724
rect 13544 23672 13596 23724
rect 13636 23715 13688 23724
rect 13636 23681 13645 23715
rect 13645 23681 13679 23715
rect 13679 23681 13688 23715
rect 13636 23672 13688 23681
rect 13912 23672 13964 23724
rect 15016 23672 15068 23724
rect 15384 23672 15436 23724
rect 15476 23715 15528 23724
rect 15476 23681 15485 23715
rect 15485 23681 15519 23715
rect 15519 23681 15528 23715
rect 15476 23672 15528 23681
rect 20168 23672 20220 23724
rect 24124 23740 24176 23792
rect 24492 23672 24544 23724
rect 24952 23740 25004 23792
rect 25136 23740 25188 23792
rect 25596 23672 25648 23724
rect 10140 23536 10192 23588
rect 5356 23468 5408 23520
rect 7196 23511 7248 23520
rect 7196 23477 7205 23511
rect 7205 23477 7239 23511
rect 7239 23477 7248 23511
rect 7196 23468 7248 23477
rect 7472 23468 7524 23520
rect 7656 23468 7708 23520
rect 7840 23511 7892 23520
rect 7840 23477 7849 23511
rect 7849 23477 7883 23511
rect 7883 23477 7892 23511
rect 7840 23468 7892 23477
rect 9496 23468 9548 23520
rect 10968 23604 11020 23656
rect 18604 23604 18656 23656
rect 22652 23604 22704 23656
rect 13084 23536 13136 23588
rect 13636 23536 13688 23588
rect 14556 23536 14608 23588
rect 22284 23536 22336 23588
rect 23572 23604 23624 23656
rect 25872 23672 25924 23724
rect 26148 23740 26200 23792
rect 27528 23740 27580 23792
rect 32312 23808 32364 23860
rect 33324 23808 33376 23860
rect 26700 23672 26752 23724
rect 26976 23672 27028 23724
rect 23756 23536 23808 23588
rect 25228 23579 25280 23588
rect 25228 23545 25237 23579
rect 25237 23545 25271 23579
rect 25271 23545 25280 23579
rect 25228 23536 25280 23545
rect 15200 23511 15252 23520
rect 15200 23477 15209 23511
rect 15209 23477 15243 23511
rect 15243 23477 15252 23511
rect 15200 23468 15252 23477
rect 20168 23468 20220 23520
rect 22100 23468 22152 23520
rect 22928 23468 22980 23520
rect 24400 23468 24452 23520
rect 26424 23604 26476 23656
rect 26608 23604 26660 23656
rect 26884 23604 26936 23656
rect 27436 23715 27488 23724
rect 27436 23681 27445 23715
rect 27445 23681 27479 23715
rect 27479 23681 27488 23715
rect 27436 23672 27488 23681
rect 27804 23672 27856 23724
rect 28816 23672 28868 23724
rect 29552 23672 29604 23724
rect 29920 23672 29972 23724
rect 30288 23672 30340 23724
rect 30748 23672 30800 23724
rect 31484 23715 31536 23724
rect 31484 23681 31493 23715
rect 31493 23681 31527 23715
rect 31527 23681 31536 23715
rect 31484 23672 31536 23681
rect 33232 23740 33284 23792
rect 34428 23783 34480 23792
rect 34428 23749 34437 23783
rect 34437 23749 34471 23783
rect 34471 23749 34480 23783
rect 34428 23740 34480 23749
rect 41604 23808 41656 23860
rect 41788 23851 41840 23860
rect 41788 23817 41797 23851
rect 41797 23817 41831 23851
rect 41831 23817 41840 23851
rect 41788 23808 41840 23817
rect 43168 23851 43220 23860
rect 43168 23817 43177 23851
rect 43177 23817 43211 23851
rect 43211 23817 43220 23851
rect 43168 23808 43220 23817
rect 26516 23536 26568 23588
rect 32220 23604 32272 23656
rect 32588 23715 32640 23724
rect 32588 23681 32597 23715
rect 32597 23681 32631 23715
rect 32631 23681 32640 23715
rect 32588 23672 32640 23681
rect 34336 23672 34388 23724
rect 34520 23715 34572 23724
rect 34520 23681 34529 23715
rect 34529 23681 34563 23715
rect 34563 23681 34572 23715
rect 34520 23672 34572 23681
rect 34612 23672 34664 23724
rect 34796 23715 34848 23724
rect 34796 23681 34805 23715
rect 34805 23681 34839 23715
rect 34839 23681 34848 23715
rect 34796 23672 34848 23681
rect 35992 23740 36044 23792
rect 40316 23783 40368 23792
rect 40316 23749 40325 23783
rect 40325 23749 40359 23783
rect 40359 23749 40368 23783
rect 40316 23740 40368 23749
rect 41880 23740 41932 23792
rect 36728 23715 36780 23724
rect 36728 23681 36737 23715
rect 36737 23681 36771 23715
rect 36771 23681 36780 23715
rect 36728 23672 36780 23681
rect 38936 23715 38988 23724
rect 38936 23681 38945 23715
rect 38945 23681 38979 23715
rect 38979 23681 38988 23715
rect 38936 23672 38988 23681
rect 39396 23715 39448 23724
rect 39396 23681 39405 23715
rect 39405 23681 39439 23715
rect 39439 23681 39448 23715
rect 39396 23672 39448 23681
rect 39672 23672 39724 23724
rect 32404 23647 32456 23656
rect 32404 23613 32413 23647
rect 32413 23613 32447 23647
rect 32447 23613 32456 23647
rect 32404 23604 32456 23613
rect 33600 23604 33652 23656
rect 33968 23604 34020 23656
rect 34152 23604 34204 23656
rect 37556 23604 37608 23656
rect 39212 23647 39264 23656
rect 39212 23613 39221 23647
rect 39221 23613 39255 23647
rect 39255 23613 39264 23647
rect 39212 23604 39264 23613
rect 41236 23604 41288 23656
rect 43812 23672 43864 23724
rect 42984 23647 43036 23656
rect 42984 23613 42993 23647
rect 42993 23613 43027 23647
rect 43027 23613 43036 23647
rect 42984 23604 43036 23613
rect 43628 23647 43680 23656
rect 43628 23613 43637 23647
rect 43637 23613 43671 23647
rect 43671 23613 43680 23647
rect 43628 23604 43680 23613
rect 31852 23536 31904 23588
rect 39856 23536 39908 23588
rect 43536 23536 43588 23588
rect 27160 23468 27212 23520
rect 27436 23468 27488 23520
rect 28264 23468 28316 23520
rect 29184 23468 29236 23520
rect 29644 23468 29696 23520
rect 29828 23511 29880 23520
rect 29828 23477 29837 23511
rect 29837 23477 29871 23511
rect 29871 23477 29880 23511
rect 29828 23468 29880 23477
rect 30932 23511 30984 23520
rect 30932 23477 30941 23511
rect 30941 23477 30975 23511
rect 30975 23477 30984 23511
rect 30932 23468 30984 23477
rect 31576 23511 31628 23520
rect 31576 23477 31585 23511
rect 31585 23477 31619 23511
rect 31619 23477 31628 23511
rect 31576 23468 31628 23477
rect 31944 23511 31996 23520
rect 31944 23477 31953 23511
rect 31953 23477 31987 23511
rect 31987 23477 31996 23511
rect 31944 23468 31996 23477
rect 33048 23468 33100 23520
rect 33784 23468 33836 23520
rect 34520 23511 34572 23520
rect 34520 23477 34529 23511
rect 34529 23477 34563 23511
rect 34563 23477 34572 23511
rect 34520 23468 34572 23477
rect 36452 23511 36504 23520
rect 36452 23477 36461 23511
rect 36461 23477 36495 23511
rect 36495 23477 36504 23511
rect 36452 23468 36504 23477
rect 36728 23468 36780 23520
rect 39120 23511 39172 23520
rect 39120 23477 39129 23511
rect 39129 23477 39163 23511
rect 39163 23477 39172 23511
rect 39120 23468 39172 23477
rect 40684 23468 40736 23520
rect 41696 23468 41748 23520
rect 44088 23468 44140 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 5448 23264 5500 23316
rect 6828 23264 6880 23316
rect 3056 23196 3108 23248
rect 3424 23196 3476 23248
rect 4620 23196 4672 23248
rect 5264 23196 5316 23248
rect 5632 23196 5684 23248
rect 7564 23196 7616 23248
rect 8300 23196 8352 23248
rect 9588 23196 9640 23248
rect 3792 23128 3844 23180
rect 4344 23060 4396 23112
rect 2136 22992 2188 23044
rect 4712 23060 4764 23112
rect 5264 23060 5316 23112
rect 9220 23128 9272 23180
rect 6644 23060 6696 23112
rect 4804 22992 4856 23044
rect 4068 22924 4120 22976
rect 5448 23035 5500 23044
rect 5448 23001 5457 23035
rect 5457 23001 5491 23035
rect 5491 23001 5500 23035
rect 5448 22992 5500 23001
rect 6736 22992 6788 23044
rect 8300 23060 8352 23112
rect 9404 22992 9456 23044
rect 9864 23060 9916 23112
rect 10232 23060 10284 23112
rect 10416 23060 10468 23112
rect 9772 22992 9824 23044
rect 10048 22924 10100 22976
rect 11244 23264 11296 23316
rect 12716 23264 12768 23316
rect 12900 23264 12952 23316
rect 11704 23196 11756 23248
rect 11244 23060 11296 23112
rect 12072 23060 12124 23112
rect 12256 23103 12308 23112
rect 12256 23069 12265 23103
rect 12265 23069 12299 23103
rect 12299 23069 12308 23103
rect 12256 23060 12308 23069
rect 12624 23103 12676 23112
rect 12624 23069 12633 23103
rect 12633 23069 12667 23103
rect 12667 23069 12676 23103
rect 12624 23060 12676 23069
rect 13084 22992 13136 23044
rect 14648 23307 14700 23316
rect 14648 23273 14657 23307
rect 14657 23273 14691 23307
rect 14691 23273 14700 23307
rect 14648 23264 14700 23273
rect 15108 23264 15160 23316
rect 15200 23307 15252 23316
rect 15200 23273 15209 23307
rect 15209 23273 15243 23307
rect 15243 23273 15252 23307
rect 15200 23264 15252 23273
rect 18880 23264 18932 23316
rect 22192 23196 22244 23248
rect 22652 23264 22704 23316
rect 23756 23264 23808 23316
rect 25136 23264 25188 23316
rect 25228 23196 25280 23248
rect 11980 22924 12032 22976
rect 12624 22924 12676 22976
rect 12992 22924 13044 22976
rect 14832 23103 14884 23112
rect 14832 23069 14841 23103
rect 14841 23069 14875 23103
rect 14875 23069 14884 23103
rect 14832 23060 14884 23069
rect 15200 23060 15252 23112
rect 16212 23060 16264 23112
rect 19340 23128 19392 23180
rect 20352 23128 20404 23180
rect 18512 23103 18564 23112
rect 18512 23069 18521 23103
rect 18521 23069 18555 23103
rect 18555 23069 18564 23103
rect 18512 23060 18564 23069
rect 20628 23060 20680 23112
rect 19248 22924 19300 22976
rect 20536 23035 20588 23044
rect 20536 23001 20545 23035
rect 20545 23001 20579 23035
rect 20579 23001 20588 23035
rect 20536 22992 20588 23001
rect 23388 23128 23440 23180
rect 24860 23128 24912 23180
rect 24952 23128 25004 23180
rect 26516 23264 26568 23316
rect 26884 23264 26936 23316
rect 27068 23264 27120 23316
rect 27528 23264 27580 23316
rect 27896 23264 27948 23316
rect 31024 23264 31076 23316
rect 32864 23264 32916 23316
rect 33600 23264 33652 23316
rect 34520 23264 34572 23316
rect 34612 23264 34664 23316
rect 37096 23307 37148 23316
rect 37096 23273 37105 23307
rect 37105 23273 37139 23307
rect 37139 23273 37148 23307
rect 37096 23264 37148 23273
rect 37280 23264 37332 23316
rect 37464 23264 37516 23316
rect 38016 23264 38068 23316
rect 38108 23264 38160 23316
rect 39212 23264 39264 23316
rect 39764 23264 39816 23316
rect 39948 23264 40000 23316
rect 25964 23196 26016 23248
rect 26608 23196 26660 23248
rect 26792 23196 26844 23248
rect 29000 23196 29052 23248
rect 20996 23060 21048 23112
rect 23480 23060 23532 23112
rect 23664 23103 23716 23112
rect 23664 23069 23673 23103
rect 23673 23069 23707 23103
rect 23707 23069 23716 23103
rect 29092 23128 29144 23180
rect 29276 23128 29328 23180
rect 29552 23239 29604 23248
rect 29552 23205 29561 23239
rect 29561 23205 29595 23239
rect 29595 23205 29604 23239
rect 29552 23196 29604 23205
rect 29644 23196 29696 23248
rect 29828 23196 29880 23248
rect 31208 23196 31260 23248
rect 32588 23196 32640 23248
rect 34888 23196 34940 23248
rect 39396 23196 39448 23248
rect 41052 23239 41104 23248
rect 41052 23205 41061 23239
rect 41061 23205 41095 23239
rect 41095 23205 41104 23239
rect 41052 23196 41104 23205
rect 32772 23128 32824 23180
rect 34152 23128 34204 23180
rect 35440 23128 35492 23180
rect 23664 23060 23716 23069
rect 26884 23060 26936 23112
rect 27160 23060 27212 23112
rect 31208 23060 31260 23112
rect 33232 23060 33284 23112
rect 33508 23060 33560 23112
rect 33968 23103 34020 23112
rect 33968 23069 33977 23103
rect 33977 23069 34011 23103
rect 34011 23069 34020 23103
rect 33968 23060 34020 23069
rect 34888 23060 34940 23112
rect 35624 23060 35676 23112
rect 36176 23060 36228 23112
rect 36912 23060 36964 23112
rect 37188 23103 37240 23112
rect 37188 23069 37197 23103
rect 37197 23069 37231 23103
rect 37231 23069 37240 23103
rect 37188 23060 37240 23069
rect 37556 23128 37608 23180
rect 37464 23103 37516 23112
rect 37464 23069 37473 23103
rect 37473 23069 37507 23103
rect 37507 23069 37516 23103
rect 37464 23060 37516 23069
rect 26056 23035 26108 23044
rect 26056 23001 26065 23035
rect 26065 23001 26099 23035
rect 26099 23001 26108 23035
rect 26056 22992 26108 23001
rect 26148 22992 26200 23044
rect 26516 22992 26568 23044
rect 27804 22992 27856 23044
rect 28080 22992 28132 23044
rect 20812 22924 20864 22976
rect 23480 22924 23532 22976
rect 23664 22924 23716 22976
rect 23848 22924 23900 22976
rect 26884 22924 26936 22976
rect 29000 22992 29052 23044
rect 31024 22992 31076 23044
rect 31392 22992 31444 23044
rect 32956 23035 33008 23044
rect 32956 23001 32965 23035
rect 32965 23001 32999 23035
rect 32999 23001 33008 23035
rect 32956 22992 33008 23001
rect 33784 22992 33836 23044
rect 35440 22992 35492 23044
rect 38568 23060 38620 23112
rect 40684 23171 40736 23180
rect 40684 23137 40693 23171
rect 40693 23137 40727 23171
rect 40727 23137 40736 23171
rect 40684 23128 40736 23137
rect 40776 23171 40828 23180
rect 40776 23137 40785 23171
rect 40785 23137 40819 23171
rect 40819 23137 40828 23171
rect 40776 23128 40828 23137
rect 39856 23103 39908 23112
rect 39856 23069 39865 23103
rect 39865 23069 39899 23103
rect 39899 23069 39908 23103
rect 39856 23060 39908 23069
rect 40868 23060 40920 23112
rect 41144 23128 41196 23180
rect 41512 23171 41564 23180
rect 41512 23137 41521 23171
rect 41521 23137 41555 23171
rect 41555 23137 41564 23171
rect 41512 23128 41564 23137
rect 31852 22924 31904 22976
rect 32128 22924 32180 22976
rect 34612 22924 34664 22976
rect 35624 22924 35676 22976
rect 38476 22924 38528 22976
rect 40408 22924 40460 22976
rect 41236 23103 41288 23112
rect 41236 23069 41245 23103
rect 41245 23069 41279 23103
rect 41279 23069 41288 23103
rect 41236 23060 41288 23069
rect 41696 23103 41748 23112
rect 41696 23069 41705 23103
rect 41705 23069 41739 23103
rect 41739 23069 41748 23103
rect 41696 23060 41748 23069
rect 42432 23103 42484 23112
rect 42432 23069 42441 23103
rect 42441 23069 42475 23103
rect 42475 23069 42484 23103
rect 42432 23060 42484 23069
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 5264 22720 5316 22772
rect 5632 22695 5684 22704
rect 5632 22661 5641 22695
rect 5641 22661 5675 22695
rect 5675 22661 5684 22695
rect 5632 22652 5684 22661
rect 9036 22720 9088 22772
rect 9128 22720 9180 22772
rect 8116 22652 8168 22704
rect 9404 22695 9456 22704
rect 9404 22661 9413 22695
rect 9413 22661 9447 22695
rect 9447 22661 9456 22695
rect 9404 22652 9456 22661
rect 11888 22652 11940 22704
rect 13360 22763 13412 22772
rect 13360 22729 13369 22763
rect 13369 22729 13403 22763
rect 13403 22729 13412 22763
rect 13360 22720 13412 22729
rect 14832 22720 14884 22772
rect 15016 22720 15068 22772
rect 4804 22584 4856 22636
rect 3792 22516 3844 22568
rect 5172 22584 5224 22636
rect 5448 22627 5500 22636
rect 5448 22593 5457 22627
rect 5457 22593 5491 22627
rect 5491 22593 5500 22627
rect 5448 22584 5500 22593
rect 5816 22627 5868 22636
rect 5816 22593 5825 22627
rect 5825 22593 5859 22627
rect 5859 22593 5868 22627
rect 5816 22584 5868 22593
rect 8392 22584 8444 22636
rect 8208 22516 8260 22568
rect 8852 22516 8904 22568
rect 9036 22584 9088 22636
rect 9220 22627 9272 22636
rect 9220 22593 9229 22627
rect 9229 22593 9263 22627
rect 9263 22593 9272 22627
rect 9220 22584 9272 22593
rect 9588 22627 9640 22636
rect 9588 22593 9602 22627
rect 9602 22593 9636 22627
rect 9636 22593 9640 22627
rect 9588 22584 9640 22593
rect 9772 22584 9824 22636
rect 9956 22584 10008 22636
rect 10048 22627 10100 22636
rect 10048 22593 10057 22627
rect 10057 22593 10091 22627
rect 10091 22593 10100 22627
rect 10048 22584 10100 22593
rect 10140 22584 10192 22636
rect 9128 22516 9180 22568
rect 10692 22584 10744 22636
rect 9404 22516 9456 22568
rect 10324 22516 10376 22568
rect 11704 22516 11756 22568
rect 12440 22584 12492 22636
rect 12808 22584 12860 22636
rect 19340 22652 19392 22704
rect 12164 22516 12216 22568
rect 14372 22584 14424 22636
rect 14556 22584 14608 22636
rect 18512 22584 18564 22636
rect 13820 22516 13872 22568
rect 5632 22448 5684 22500
rect 6000 22491 6052 22500
rect 6000 22457 6009 22491
rect 6009 22457 6043 22491
rect 6043 22457 6052 22491
rect 6000 22448 6052 22457
rect 13544 22448 13596 22500
rect 5080 22380 5132 22432
rect 8668 22423 8720 22432
rect 8668 22389 8677 22423
rect 8677 22389 8711 22423
rect 8711 22389 8720 22423
rect 8668 22380 8720 22389
rect 10508 22380 10560 22432
rect 10784 22380 10836 22432
rect 12716 22380 12768 22432
rect 13176 22380 13228 22432
rect 14188 22559 14240 22568
rect 14188 22525 14197 22559
rect 14197 22525 14231 22559
rect 14231 22525 14240 22559
rect 14188 22516 14240 22525
rect 14372 22448 14424 22500
rect 16948 22448 17000 22500
rect 20352 22652 20404 22704
rect 19800 22584 19852 22636
rect 20812 22627 20864 22636
rect 20812 22593 20821 22627
rect 20821 22593 20855 22627
rect 20855 22593 20864 22627
rect 20812 22584 20864 22593
rect 21548 22652 21600 22704
rect 21456 22627 21508 22636
rect 21456 22593 21465 22627
rect 21465 22593 21499 22627
rect 21499 22593 21508 22627
rect 23664 22720 23716 22772
rect 22100 22652 22152 22704
rect 24492 22695 24544 22704
rect 24492 22661 24501 22695
rect 24501 22661 24535 22695
rect 24535 22661 24544 22695
rect 24492 22652 24544 22661
rect 27344 22652 27396 22704
rect 29092 22652 29144 22704
rect 29368 22652 29420 22704
rect 29552 22652 29604 22704
rect 29828 22652 29880 22704
rect 31484 22652 31536 22704
rect 31852 22720 31904 22772
rect 32956 22720 33008 22772
rect 33416 22720 33468 22772
rect 33968 22720 34020 22772
rect 36544 22720 36596 22772
rect 38476 22720 38528 22772
rect 42432 22720 42484 22772
rect 33324 22652 33376 22704
rect 36360 22652 36412 22704
rect 38108 22652 38160 22704
rect 40868 22652 40920 22704
rect 41788 22652 41840 22704
rect 21456 22584 21508 22593
rect 22192 22627 22244 22636
rect 22192 22593 22201 22627
rect 22201 22593 22235 22627
rect 22235 22593 22244 22627
rect 22192 22584 22244 22593
rect 22836 22584 22888 22636
rect 24400 22584 24452 22636
rect 25228 22584 25280 22636
rect 26148 22584 26200 22636
rect 26240 22627 26292 22636
rect 26240 22593 26249 22627
rect 26249 22593 26283 22627
rect 26283 22593 26292 22627
rect 26240 22584 26292 22593
rect 26516 22627 26568 22636
rect 26516 22593 26525 22627
rect 26525 22593 26559 22627
rect 26559 22593 26568 22627
rect 26516 22584 26568 22593
rect 26884 22584 26936 22636
rect 20996 22516 21048 22568
rect 16304 22380 16356 22432
rect 20536 22380 20588 22432
rect 20812 22423 20864 22432
rect 20812 22389 20821 22423
rect 20821 22389 20855 22423
rect 20855 22389 20864 22423
rect 20812 22380 20864 22389
rect 24860 22516 24912 22568
rect 26056 22516 26108 22568
rect 26332 22559 26384 22568
rect 21824 22380 21876 22432
rect 22284 22380 22336 22432
rect 22376 22423 22428 22432
rect 22376 22389 22385 22423
rect 22385 22389 22419 22423
rect 22419 22389 22428 22423
rect 22376 22380 22428 22389
rect 23940 22380 23992 22432
rect 25596 22380 25648 22432
rect 26332 22525 26341 22559
rect 26341 22525 26375 22559
rect 26375 22525 26384 22559
rect 26332 22516 26384 22525
rect 27344 22516 27396 22568
rect 29000 22516 29052 22568
rect 29276 22627 29328 22636
rect 29276 22593 29285 22627
rect 29285 22593 29319 22627
rect 29319 22593 29328 22627
rect 29276 22584 29328 22593
rect 31024 22627 31076 22636
rect 31024 22593 31033 22627
rect 31033 22593 31067 22627
rect 31067 22593 31076 22627
rect 31024 22584 31076 22593
rect 31208 22627 31260 22636
rect 31208 22593 31217 22627
rect 31217 22593 31251 22627
rect 31251 22593 31260 22627
rect 31208 22584 31260 22593
rect 31300 22584 31352 22636
rect 35624 22584 35676 22636
rect 38016 22584 38068 22636
rect 38384 22584 38436 22636
rect 40316 22627 40368 22636
rect 40316 22593 40325 22627
rect 40325 22593 40359 22627
rect 40359 22593 40368 22627
rect 40316 22584 40368 22593
rect 40408 22584 40460 22636
rect 42432 22584 42484 22636
rect 26332 22380 26384 22432
rect 27436 22380 27488 22432
rect 29000 22380 29052 22432
rect 30932 22516 30984 22568
rect 29276 22448 29328 22500
rect 29736 22448 29788 22500
rect 32956 22516 33008 22568
rect 37924 22516 37976 22568
rect 29184 22423 29236 22432
rect 29184 22389 29193 22423
rect 29193 22389 29227 22423
rect 29227 22389 29236 22423
rect 29184 22380 29236 22389
rect 30932 22380 30984 22432
rect 31300 22380 31352 22432
rect 31392 22423 31444 22432
rect 31392 22389 31401 22423
rect 31401 22389 31435 22423
rect 31435 22389 31444 22423
rect 31392 22380 31444 22389
rect 31484 22380 31536 22432
rect 33416 22448 33468 22500
rect 35532 22448 35584 22500
rect 44456 22491 44508 22500
rect 44456 22457 44465 22491
rect 44465 22457 44499 22491
rect 44499 22457 44508 22491
rect 44456 22448 44508 22457
rect 32036 22380 32088 22432
rect 36820 22380 36872 22432
rect 39764 22380 39816 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 5724 22176 5776 22228
rect 7380 22176 7432 22228
rect 5816 22108 5868 22160
rect 7748 22176 7800 22228
rect 10692 22176 10744 22228
rect 13544 22176 13596 22228
rect 14556 22176 14608 22228
rect 14924 22219 14976 22228
rect 14924 22185 14933 22219
rect 14933 22185 14967 22219
rect 14967 22185 14976 22219
rect 14924 22176 14976 22185
rect 15568 22176 15620 22228
rect 15844 22219 15896 22228
rect 15844 22185 15853 22219
rect 15853 22185 15887 22219
rect 15887 22185 15896 22219
rect 15844 22176 15896 22185
rect 16304 22176 16356 22228
rect 10140 22108 10192 22160
rect 10416 22108 10468 22160
rect 12164 22151 12216 22160
rect 12164 22117 12173 22151
rect 12173 22117 12207 22151
rect 12207 22117 12216 22151
rect 12164 22108 12216 22117
rect 6460 22040 6512 22092
rect 5080 22015 5132 22024
rect 5080 21981 5089 22015
rect 5089 21981 5123 22015
rect 5123 21981 5132 22015
rect 5080 21972 5132 21981
rect 5264 22015 5316 22024
rect 5264 21981 5273 22015
rect 5273 21981 5307 22015
rect 5307 21981 5316 22015
rect 5264 21972 5316 21981
rect 5908 21972 5960 22024
rect 7932 22083 7984 22092
rect 7932 22049 7941 22083
rect 7941 22049 7975 22083
rect 7975 22049 7984 22083
rect 7932 22040 7984 22049
rect 11060 22040 11112 22092
rect 11336 22040 11388 22092
rect 13912 22108 13964 22160
rect 14004 22108 14056 22160
rect 14280 22108 14332 22160
rect 5540 21879 5592 21888
rect 5540 21845 5549 21879
rect 5549 21845 5583 21879
rect 5583 21845 5592 21879
rect 5540 21836 5592 21845
rect 6920 21904 6972 21956
rect 7012 21947 7064 21956
rect 7012 21913 7021 21947
rect 7021 21913 7055 21947
rect 7055 21913 7064 21947
rect 7012 21904 7064 21913
rect 10048 21972 10100 22024
rect 10416 21972 10468 22024
rect 15844 22083 15896 22092
rect 15844 22049 15853 22083
rect 15853 22049 15887 22083
rect 15887 22049 15896 22083
rect 15844 22040 15896 22049
rect 16488 22040 16540 22092
rect 11980 22015 12032 22024
rect 11980 21981 11989 22015
rect 11989 21981 12023 22015
rect 12023 21981 12032 22015
rect 11980 21972 12032 21981
rect 12072 21972 12124 22024
rect 12440 22015 12492 22024
rect 12440 21981 12449 22015
rect 12449 21981 12483 22015
rect 12483 21981 12492 22015
rect 12440 21972 12492 21981
rect 7380 21904 7432 21956
rect 8208 21904 8260 21956
rect 9680 21904 9732 21956
rect 10876 21904 10928 21956
rect 11336 21904 11388 21956
rect 11704 21904 11756 21956
rect 11888 21947 11940 21956
rect 11888 21913 11897 21947
rect 11897 21913 11931 21947
rect 11931 21913 11940 21947
rect 11888 21904 11940 21913
rect 12532 21947 12584 21956
rect 12532 21913 12541 21947
rect 12541 21913 12575 21947
rect 12575 21913 12584 21947
rect 12532 21904 12584 21913
rect 7288 21836 7340 21888
rect 8484 21836 8536 21888
rect 14924 22015 14976 22024
rect 14924 21981 14933 22015
rect 14933 21981 14967 22015
rect 14967 21981 14976 22015
rect 14924 21972 14976 21981
rect 15016 22015 15068 22024
rect 15016 21981 15025 22015
rect 15025 21981 15059 22015
rect 15059 21981 15068 22015
rect 15016 21972 15068 21981
rect 15752 21972 15804 22024
rect 17132 22176 17184 22228
rect 16948 22108 17000 22160
rect 20812 22176 20864 22228
rect 21180 22176 21232 22228
rect 21548 22176 21600 22228
rect 25136 22219 25188 22228
rect 25136 22185 25145 22219
rect 25145 22185 25179 22219
rect 25179 22185 25188 22219
rect 25136 22176 25188 22185
rect 25228 22176 25280 22228
rect 19616 22108 19668 22160
rect 20444 22108 20496 22160
rect 18052 22040 18104 22092
rect 21272 22040 21324 22092
rect 21640 22040 21692 22092
rect 24676 22108 24728 22160
rect 26056 22219 26108 22228
rect 26056 22185 26065 22219
rect 26065 22185 26099 22219
rect 26099 22185 26108 22219
rect 26056 22176 26108 22185
rect 26332 22108 26384 22160
rect 26424 22108 26476 22160
rect 26608 22108 26660 22160
rect 26792 22219 26844 22228
rect 26792 22185 26801 22219
rect 26801 22185 26835 22219
rect 26835 22185 26844 22219
rect 26792 22176 26844 22185
rect 27252 22176 27304 22228
rect 27804 22219 27856 22228
rect 27804 22185 27813 22219
rect 27813 22185 27847 22219
rect 27847 22185 27856 22219
rect 27804 22176 27856 22185
rect 27988 22176 28040 22228
rect 28172 22176 28224 22228
rect 28448 22176 28500 22228
rect 33048 22176 33100 22228
rect 33232 22219 33284 22228
rect 33232 22185 33241 22219
rect 33241 22185 33275 22219
rect 33275 22185 33284 22219
rect 33232 22176 33284 22185
rect 33508 22176 33560 22228
rect 24584 22040 24636 22092
rect 16856 21972 16908 22024
rect 18236 21972 18288 22024
rect 19156 21972 19208 22024
rect 19248 22015 19300 22024
rect 19248 21981 19257 22015
rect 19257 21981 19291 22015
rect 19291 21981 19300 22015
rect 19248 21972 19300 21981
rect 19524 22015 19576 22024
rect 19524 21981 19533 22015
rect 19533 21981 19567 22015
rect 19567 21981 19576 22015
rect 19524 21972 19576 21981
rect 21180 21972 21232 22024
rect 24216 21972 24268 22024
rect 14556 21904 14608 21956
rect 14832 21904 14884 21956
rect 16488 21904 16540 21956
rect 16948 21947 17000 21956
rect 16948 21913 16957 21947
rect 16957 21913 16991 21947
rect 16991 21913 17000 21947
rect 16948 21904 17000 21913
rect 12716 21836 12768 21888
rect 12808 21836 12860 21888
rect 13544 21836 13596 21888
rect 18144 21879 18196 21888
rect 18144 21845 18153 21879
rect 18153 21845 18187 21879
rect 18187 21845 18196 21879
rect 18144 21836 18196 21845
rect 18328 21947 18380 21956
rect 18328 21913 18337 21947
rect 18337 21913 18371 21947
rect 18371 21913 18380 21947
rect 18328 21904 18380 21913
rect 18512 21947 18564 21956
rect 18512 21913 18521 21947
rect 18521 21913 18555 21947
rect 18555 21913 18564 21947
rect 18512 21904 18564 21913
rect 18880 21904 18932 21956
rect 24400 21947 24452 21956
rect 24400 21913 24409 21947
rect 24409 21913 24443 21947
rect 24443 21913 24452 21947
rect 24400 21904 24452 21913
rect 20628 21836 20680 21888
rect 21824 21836 21876 21888
rect 24492 21836 24544 21888
rect 24860 21947 24912 21956
rect 24860 21913 24869 21947
rect 24869 21913 24903 21947
rect 24903 21913 24912 21947
rect 24860 21904 24912 21913
rect 25136 22015 25188 22024
rect 25136 21981 25145 22015
rect 25145 21981 25179 22015
rect 25179 21981 25188 22015
rect 25136 21972 25188 21981
rect 25228 21904 25280 21956
rect 25044 21836 25096 21888
rect 25964 22040 26016 22092
rect 26148 22083 26200 22092
rect 26148 22049 26157 22083
rect 26157 22049 26191 22083
rect 26191 22049 26200 22083
rect 26148 22040 26200 22049
rect 27160 22040 27212 22092
rect 25964 21904 26016 21956
rect 25688 21836 25740 21888
rect 26792 22015 26844 22024
rect 26792 21981 26801 22015
rect 26801 21981 26835 22015
rect 26835 21981 26844 22015
rect 26792 21972 26844 21981
rect 27988 22083 28040 22092
rect 27988 22049 27997 22083
rect 27997 22049 28031 22083
rect 28031 22049 28040 22083
rect 27988 22040 28040 22049
rect 30564 22108 30616 22160
rect 31116 22108 31168 22160
rect 31208 22108 31260 22160
rect 31484 22108 31536 22160
rect 31024 22040 31076 22092
rect 34152 22108 34204 22160
rect 34520 22176 34572 22228
rect 35164 22176 35216 22228
rect 35440 22176 35492 22228
rect 36360 22176 36412 22228
rect 35256 22108 35308 22160
rect 36084 22108 36136 22160
rect 28080 22015 28132 22024
rect 28080 21981 28089 22015
rect 28089 21981 28123 22015
rect 28123 21981 28132 22015
rect 28080 21972 28132 21981
rect 29000 21972 29052 22024
rect 26976 21879 27028 21888
rect 26976 21845 26985 21879
rect 26985 21845 27019 21879
rect 27019 21845 27028 21879
rect 26976 21836 27028 21845
rect 32496 21904 32548 21956
rect 32036 21836 32088 21888
rect 33048 21904 33100 21956
rect 33692 21972 33744 22024
rect 35532 22040 35584 22092
rect 38384 22040 38436 22092
rect 34060 21904 34112 21956
rect 34520 21904 34572 21956
rect 34704 21947 34756 21956
rect 34704 21913 34713 21947
rect 34713 21913 34747 21947
rect 34747 21913 34756 21947
rect 34704 21904 34756 21913
rect 35440 21972 35492 22024
rect 40040 21972 40092 22024
rect 41236 22176 41288 22228
rect 40316 22108 40368 22160
rect 40408 22015 40460 22024
rect 40408 21981 40417 22015
rect 40417 21981 40451 22015
rect 40451 21981 40460 22015
rect 40408 21972 40460 21981
rect 35532 21947 35584 21956
rect 35532 21913 35541 21947
rect 35541 21913 35575 21947
rect 35575 21913 35584 21947
rect 35532 21904 35584 21913
rect 38660 21904 38712 21956
rect 38936 21904 38988 21956
rect 40684 21972 40736 22024
rect 43536 22015 43588 22024
rect 43536 21981 43545 22015
rect 43545 21981 43579 22015
rect 43579 21981 43588 22015
rect 43536 21972 43588 21981
rect 43352 21904 43404 21956
rect 35992 21879 36044 21888
rect 35992 21845 36001 21879
rect 36001 21845 36035 21879
rect 36035 21845 36044 21879
rect 35992 21836 36044 21845
rect 36452 21836 36504 21888
rect 39948 21836 40000 21888
rect 40132 21879 40184 21888
rect 40132 21845 40141 21879
rect 40141 21845 40175 21879
rect 40175 21845 40184 21879
rect 40132 21836 40184 21845
rect 43076 21836 43128 21888
rect 44456 21879 44508 21888
rect 44456 21845 44465 21879
rect 44465 21845 44499 21879
rect 44499 21845 44508 21879
rect 44456 21836 44508 21845
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 6920 21632 6972 21684
rect 7380 21632 7432 21684
rect 7840 21632 7892 21684
rect 8484 21632 8536 21684
rect 9036 21632 9088 21684
rect 9864 21675 9916 21684
rect 9864 21641 9873 21675
rect 9873 21641 9907 21675
rect 9907 21641 9916 21675
rect 9864 21632 9916 21641
rect 3976 21564 4028 21616
rect 11060 21632 11112 21684
rect 2688 21539 2740 21548
rect 2688 21505 2697 21539
rect 2697 21505 2731 21539
rect 2731 21505 2740 21539
rect 2688 21496 2740 21505
rect 2504 21428 2556 21480
rect 5632 21539 5684 21548
rect 5632 21505 5641 21539
rect 5641 21505 5675 21539
rect 5675 21505 5684 21539
rect 5632 21496 5684 21505
rect 5816 21539 5868 21548
rect 5816 21505 5825 21539
rect 5825 21505 5859 21539
rect 5859 21505 5868 21539
rect 5816 21496 5868 21505
rect 5908 21539 5960 21548
rect 5908 21505 5917 21539
rect 5917 21505 5951 21539
rect 5951 21505 5960 21539
rect 5908 21496 5960 21505
rect 4896 21428 4948 21480
rect 6368 21496 6420 21548
rect 10048 21564 10100 21616
rect 11612 21564 11664 21616
rect 11888 21564 11940 21616
rect 12808 21632 12860 21684
rect 14372 21632 14424 21684
rect 20812 21675 20864 21684
rect 20812 21641 20821 21675
rect 20821 21641 20855 21675
rect 20855 21641 20864 21675
rect 20812 21632 20864 21641
rect 13728 21564 13780 21616
rect 14556 21564 14608 21616
rect 8760 21496 8812 21548
rect 9956 21539 10008 21548
rect 9956 21505 9965 21539
rect 9965 21505 9999 21539
rect 9999 21505 10008 21539
rect 9956 21496 10008 21505
rect 9496 21428 9548 21480
rect 10692 21496 10744 21548
rect 12164 21496 12216 21548
rect 12440 21496 12492 21548
rect 12716 21539 12768 21548
rect 12716 21505 12725 21539
rect 12725 21505 12759 21539
rect 12759 21505 12768 21539
rect 12716 21496 12768 21505
rect 13268 21496 13320 21548
rect 17684 21496 17736 21548
rect 18144 21564 18196 21616
rect 31024 21632 31076 21684
rect 32036 21632 32088 21684
rect 32312 21632 32364 21684
rect 23940 21607 23992 21616
rect 23940 21573 23949 21607
rect 23949 21573 23983 21607
rect 23983 21573 23992 21607
rect 23940 21564 23992 21573
rect 24584 21564 24636 21616
rect 10968 21428 11020 21480
rect 14832 21428 14884 21480
rect 14924 21428 14976 21480
rect 17500 21428 17552 21480
rect 20628 21539 20680 21548
rect 20628 21505 20637 21539
rect 20637 21505 20671 21539
rect 20671 21505 20680 21539
rect 20628 21496 20680 21505
rect 21272 21496 21324 21548
rect 20720 21428 20772 21480
rect 23848 21496 23900 21548
rect 24400 21496 24452 21548
rect 23112 21428 23164 21480
rect 9680 21360 9732 21412
rect 11980 21360 12032 21412
rect 15476 21360 15528 21412
rect 17224 21360 17276 21412
rect 23848 21360 23900 21412
rect 24400 21403 24452 21412
rect 24400 21369 24409 21403
rect 24409 21369 24443 21403
rect 24443 21369 24452 21403
rect 24400 21360 24452 21369
rect 24676 21496 24728 21548
rect 24584 21471 24636 21480
rect 24584 21437 24593 21471
rect 24593 21437 24627 21471
rect 24627 21437 24636 21471
rect 24584 21428 24636 21437
rect 24860 21496 24912 21548
rect 26976 21496 27028 21548
rect 30564 21496 30616 21548
rect 30748 21539 30800 21548
rect 30748 21505 30757 21539
rect 30757 21505 30791 21539
rect 30791 21505 30800 21539
rect 30748 21496 30800 21505
rect 30840 21496 30892 21548
rect 25964 21428 26016 21480
rect 27804 21428 27856 21480
rect 5632 21292 5684 21344
rect 6368 21292 6420 21344
rect 8576 21292 8628 21344
rect 8852 21292 8904 21344
rect 10232 21292 10284 21344
rect 11428 21292 11480 21344
rect 14924 21292 14976 21344
rect 15016 21292 15068 21344
rect 19524 21292 19576 21344
rect 19616 21292 19668 21344
rect 20076 21292 20128 21344
rect 20812 21292 20864 21344
rect 20996 21292 21048 21344
rect 21548 21335 21600 21344
rect 21548 21301 21557 21335
rect 21557 21301 21591 21335
rect 21591 21301 21600 21335
rect 21548 21292 21600 21301
rect 23480 21292 23532 21344
rect 24032 21292 24084 21344
rect 24216 21292 24268 21344
rect 24768 21360 24820 21412
rect 24860 21360 24912 21412
rect 27068 21360 27120 21412
rect 29736 21360 29788 21412
rect 27344 21292 27396 21344
rect 30012 21335 30064 21344
rect 30012 21301 30021 21335
rect 30021 21301 30055 21335
rect 30055 21301 30064 21335
rect 30012 21292 30064 21301
rect 30196 21335 30248 21344
rect 30196 21301 30205 21335
rect 30205 21301 30239 21335
rect 30239 21301 30248 21335
rect 30196 21292 30248 21301
rect 30932 21428 30984 21480
rect 31208 21539 31260 21548
rect 31208 21505 31217 21539
rect 31217 21505 31251 21539
rect 31251 21505 31260 21539
rect 31208 21496 31260 21505
rect 31576 21496 31628 21548
rect 32312 21496 32364 21548
rect 33048 21632 33100 21684
rect 33232 21675 33284 21684
rect 33232 21641 33241 21675
rect 33241 21641 33275 21675
rect 33275 21641 33284 21675
rect 33232 21632 33284 21641
rect 32404 21471 32456 21480
rect 32404 21437 32413 21471
rect 32413 21437 32447 21471
rect 32447 21437 32456 21471
rect 33508 21539 33560 21548
rect 33508 21505 33517 21539
rect 33517 21505 33551 21539
rect 33551 21505 33560 21539
rect 33508 21496 33560 21505
rect 35348 21632 35400 21684
rect 35072 21564 35124 21616
rect 37280 21607 37332 21616
rect 37280 21573 37289 21607
rect 37289 21573 37323 21607
rect 37323 21573 37332 21607
rect 37280 21564 37332 21573
rect 37372 21564 37424 21616
rect 38936 21675 38988 21684
rect 38936 21641 38945 21675
rect 38945 21641 38979 21675
rect 38979 21641 38988 21675
rect 38936 21632 38988 21641
rect 43536 21632 43588 21684
rect 32404 21428 32456 21437
rect 33048 21428 33100 21480
rect 35256 21496 35308 21548
rect 37464 21496 37516 21548
rect 38108 21564 38160 21616
rect 40132 21564 40184 21616
rect 35164 21428 35216 21480
rect 35532 21428 35584 21480
rect 37740 21428 37792 21480
rect 38016 21471 38068 21480
rect 38016 21437 38025 21471
rect 38025 21437 38059 21471
rect 38059 21437 38068 21471
rect 38016 21428 38068 21437
rect 38292 21496 38344 21548
rect 38752 21539 38804 21548
rect 38752 21505 38761 21539
rect 38761 21505 38795 21539
rect 38795 21505 38804 21539
rect 38752 21496 38804 21505
rect 38844 21496 38896 21548
rect 39120 21471 39172 21480
rect 39120 21437 39129 21471
rect 39129 21437 39163 21471
rect 39163 21437 39172 21471
rect 39120 21428 39172 21437
rect 30472 21335 30524 21344
rect 30472 21301 30481 21335
rect 30481 21301 30515 21335
rect 30515 21301 30524 21335
rect 30472 21292 30524 21301
rect 31024 21292 31076 21344
rect 40408 21496 40460 21548
rect 42800 21539 42852 21548
rect 42800 21505 42809 21539
rect 42809 21505 42843 21539
rect 42843 21505 42852 21539
rect 42800 21496 42852 21505
rect 43076 21539 43128 21548
rect 43076 21505 43085 21539
rect 43085 21505 43119 21539
rect 43119 21505 43128 21539
rect 43076 21496 43128 21505
rect 44180 21496 44232 21548
rect 40316 21471 40368 21480
rect 40316 21437 40325 21471
rect 40325 21437 40359 21471
rect 40359 21437 40368 21471
rect 40316 21428 40368 21437
rect 41328 21360 41380 21412
rect 43904 21360 43956 21412
rect 32312 21335 32364 21344
rect 32312 21301 32321 21335
rect 32321 21301 32355 21335
rect 32355 21301 32364 21335
rect 32312 21292 32364 21301
rect 33048 21292 33100 21344
rect 33692 21292 33744 21344
rect 37372 21292 37424 21344
rect 37556 21335 37608 21344
rect 37556 21301 37565 21335
rect 37565 21301 37599 21335
rect 37599 21301 37608 21335
rect 37556 21292 37608 21301
rect 38108 21292 38160 21344
rect 38292 21292 38344 21344
rect 38384 21335 38436 21344
rect 38384 21301 38393 21335
rect 38393 21301 38427 21335
rect 38427 21301 38436 21335
rect 38384 21292 38436 21301
rect 39028 21335 39080 21344
rect 39028 21301 39037 21335
rect 39037 21301 39071 21335
rect 39071 21301 39080 21335
rect 39028 21292 39080 21301
rect 39396 21335 39448 21344
rect 39396 21301 39405 21335
rect 39405 21301 39439 21335
rect 39439 21301 39448 21335
rect 39396 21292 39448 21301
rect 43812 21292 43864 21344
rect 44456 21335 44508 21344
rect 44456 21301 44465 21335
rect 44465 21301 44499 21335
rect 44499 21301 44508 21335
rect 44456 21292 44508 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 3976 21088 4028 21140
rect 4620 21088 4672 21140
rect 5816 21088 5868 21140
rect 7196 21088 7248 21140
rect 2136 20927 2188 20936
rect 2136 20893 2145 20927
rect 2145 20893 2179 20927
rect 2179 20893 2188 20927
rect 2136 20884 2188 20893
rect 3056 20952 3108 21004
rect 7840 21088 7892 21140
rect 8852 21088 8904 21140
rect 9772 21131 9824 21140
rect 9772 21097 9781 21131
rect 9781 21097 9815 21131
rect 9815 21097 9824 21131
rect 9772 21088 9824 21097
rect 11520 21088 11572 21140
rect 13084 21131 13136 21140
rect 13084 21097 13093 21131
rect 13093 21097 13127 21131
rect 13127 21097 13136 21131
rect 13084 21088 13136 21097
rect 13268 21088 13320 21140
rect 2596 20884 2648 20936
rect 3240 20884 3292 20936
rect 3884 20884 3936 20936
rect 3976 20859 4028 20868
rect 3976 20825 3985 20859
rect 3985 20825 4019 20859
rect 4019 20825 4028 20859
rect 3976 20816 4028 20825
rect 4160 20884 4212 20936
rect 4896 20884 4948 20936
rect 5264 20884 5316 20936
rect 5632 20884 5684 20936
rect 6460 20884 6512 20936
rect 8208 20927 8260 20936
rect 8208 20893 8217 20927
rect 8217 20893 8251 20927
rect 8251 20893 8260 20927
rect 8208 20884 8260 20893
rect 9496 21020 9548 21072
rect 9128 20952 9180 21004
rect 10876 21020 10928 21072
rect 10324 20952 10376 21004
rect 7288 20816 7340 20868
rect 8852 20816 8904 20868
rect 8208 20748 8260 20800
rect 8944 20748 8996 20800
rect 9496 20927 9548 20936
rect 9496 20893 9505 20927
rect 9505 20893 9539 20927
rect 9539 20893 9548 20927
rect 9496 20884 9548 20893
rect 9680 20927 9732 20936
rect 9680 20893 9683 20927
rect 9683 20893 9732 20927
rect 9680 20884 9732 20893
rect 9772 20884 9824 20936
rect 10968 20884 11020 20936
rect 12072 21020 12124 21072
rect 12256 21020 12308 21072
rect 12808 21020 12860 21072
rect 13452 21088 13504 21140
rect 14648 21088 14700 21140
rect 17132 21088 17184 21140
rect 18144 21131 18196 21140
rect 18144 21097 18153 21131
rect 18153 21097 18187 21131
rect 18187 21097 18196 21131
rect 18144 21088 18196 21097
rect 19248 21131 19300 21140
rect 19248 21097 19257 21131
rect 19257 21097 19291 21131
rect 19291 21097 19300 21131
rect 19248 21088 19300 21097
rect 19708 21131 19760 21140
rect 19708 21097 19717 21131
rect 19717 21097 19751 21131
rect 19751 21097 19760 21131
rect 19708 21088 19760 21097
rect 20812 21088 20864 21140
rect 14096 21020 14148 21072
rect 15016 21020 15068 21072
rect 15476 21020 15528 21072
rect 12440 20952 12492 21004
rect 12256 20927 12308 20936
rect 12256 20893 12259 20927
rect 12259 20893 12308 20927
rect 9404 20859 9456 20868
rect 9404 20825 9413 20859
rect 9413 20825 9447 20859
rect 9447 20825 9456 20859
rect 9404 20816 9456 20825
rect 10416 20816 10468 20868
rect 10692 20816 10744 20868
rect 12256 20884 12308 20893
rect 14004 20952 14056 21004
rect 12808 20927 12860 20936
rect 12808 20893 12817 20927
rect 12817 20893 12851 20927
rect 12851 20893 12860 20927
rect 12808 20884 12860 20893
rect 13360 20884 13412 20936
rect 13544 20884 13596 20936
rect 13820 20884 13872 20936
rect 14464 20884 14516 20936
rect 18420 20952 18472 21004
rect 20904 20952 20956 21004
rect 24584 21088 24636 21140
rect 24860 21088 24912 21140
rect 26976 21131 27028 21140
rect 26976 21097 26985 21131
rect 26985 21097 27019 21131
rect 27019 21097 27028 21131
rect 26976 21088 27028 21097
rect 30564 21088 30616 21140
rect 34060 21088 34112 21140
rect 34888 21088 34940 21140
rect 35532 21088 35584 21140
rect 35992 21131 36044 21140
rect 35992 21097 36001 21131
rect 36001 21097 36035 21131
rect 36035 21097 36044 21131
rect 35992 21088 36044 21097
rect 36268 21088 36320 21140
rect 38384 21131 38436 21140
rect 38384 21097 38393 21131
rect 38393 21097 38427 21131
rect 38427 21097 38436 21131
rect 38384 21088 38436 21097
rect 38844 21088 38896 21140
rect 39396 21088 39448 21140
rect 21548 21020 21600 21072
rect 33416 21020 33468 21072
rect 33968 21020 34020 21072
rect 36360 21020 36412 21072
rect 37096 21020 37148 21072
rect 14740 20884 14792 20936
rect 11888 20816 11940 20868
rect 12440 20816 12492 20868
rect 13176 20816 13228 20868
rect 13452 20859 13504 20868
rect 13452 20825 13461 20859
rect 13461 20825 13495 20859
rect 13495 20825 13504 20859
rect 13452 20816 13504 20825
rect 15292 20884 15344 20936
rect 17224 20884 17276 20936
rect 17592 20927 17644 20936
rect 17592 20893 17601 20927
rect 17601 20893 17635 20927
rect 17635 20893 17644 20927
rect 17592 20884 17644 20893
rect 17684 20927 17736 20936
rect 17684 20893 17693 20927
rect 17693 20893 17727 20927
rect 17727 20893 17736 20927
rect 17684 20884 17736 20893
rect 10968 20748 11020 20800
rect 11428 20748 11480 20800
rect 11980 20748 12032 20800
rect 12624 20748 12676 20800
rect 13544 20748 13596 20800
rect 14096 20748 14148 20800
rect 14832 20748 14884 20800
rect 15108 20859 15160 20868
rect 15108 20825 15117 20859
rect 15117 20825 15151 20859
rect 15151 20825 15160 20859
rect 15108 20816 15160 20825
rect 18328 20927 18380 20936
rect 18328 20893 18337 20927
rect 18337 20893 18371 20927
rect 18371 20893 18380 20927
rect 18328 20884 18380 20893
rect 19432 20884 19484 20936
rect 21180 20927 21232 20936
rect 21180 20893 21189 20927
rect 21189 20893 21223 20927
rect 21223 20893 21232 20927
rect 21180 20884 21232 20893
rect 18696 20816 18748 20868
rect 18328 20748 18380 20800
rect 20628 20816 20680 20868
rect 21548 20927 21600 20936
rect 21548 20893 21557 20927
rect 21557 20893 21591 20927
rect 21591 20893 21600 20927
rect 21548 20884 21600 20893
rect 21732 20952 21784 21004
rect 23112 20995 23164 21004
rect 23112 20961 23121 20995
rect 23121 20961 23155 20995
rect 23155 20961 23164 20995
rect 23112 20952 23164 20961
rect 24584 20995 24636 21004
rect 24584 20961 24593 20995
rect 24593 20961 24627 20995
rect 24627 20961 24636 20995
rect 24584 20952 24636 20961
rect 23296 20927 23348 20936
rect 23296 20893 23305 20927
rect 23305 20893 23339 20927
rect 23339 20893 23348 20927
rect 23296 20884 23348 20893
rect 24400 20884 24452 20936
rect 19524 20748 19576 20800
rect 19892 20748 19944 20800
rect 20812 20748 20864 20800
rect 21364 20791 21416 20800
rect 21364 20757 21373 20791
rect 21373 20757 21407 20791
rect 21407 20757 21416 20791
rect 21364 20748 21416 20757
rect 21824 20748 21876 20800
rect 23664 20816 23716 20868
rect 24860 20884 24912 20936
rect 25320 20952 25372 21004
rect 25320 20816 25372 20868
rect 25780 20816 25832 20868
rect 25136 20748 25188 20800
rect 26332 20927 26384 20936
rect 26332 20893 26341 20927
rect 26341 20893 26375 20927
rect 26375 20893 26384 20927
rect 26332 20884 26384 20893
rect 30196 20952 30248 21004
rect 33692 20952 33744 21004
rect 35348 20952 35400 21004
rect 40316 20952 40368 21004
rect 27068 20884 27120 20936
rect 27804 20884 27856 20936
rect 30840 20884 30892 20936
rect 34612 20884 34664 20936
rect 36176 20927 36228 20936
rect 36176 20893 36185 20927
rect 36185 20893 36219 20927
rect 36219 20893 36228 20927
rect 36176 20884 36228 20893
rect 36268 20927 36320 20936
rect 36268 20893 36277 20927
rect 36277 20893 36311 20927
rect 36311 20893 36320 20927
rect 36268 20884 36320 20893
rect 38200 20927 38252 20936
rect 38200 20893 38209 20927
rect 38209 20893 38243 20927
rect 38243 20893 38252 20927
rect 38200 20884 38252 20893
rect 38292 20927 38344 20936
rect 38292 20893 38301 20927
rect 38301 20893 38335 20927
rect 38335 20893 38344 20927
rect 38292 20884 38344 20893
rect 43352 21063 43404 21072
rect 43352 21029 43361 21063
rect 43361 21029 43395 21063
rect 43395 21029 43404 21063
rect 43352 21020 43404 21029
rect 43260 20927 43312 20936
rect 43260 20893 43269 20927
rect 43269 20893 43303 20927
rect 43303 20893 43312 20927
rect 43260 20884 43312 20893
rect 43812 21131 43864 21140
rect 43812 21097 43821 21131
rect 43821 21097 43855 21131
rect 43855 21097 43864 21131
rect 43812 21088 43864 21097
rect 26516 20859 26568 20868
rect 26516 20825 26525 20859
rect 26525 20825 26559 20859
rect 26559 20825 26568 20859
rect 26516 20816 26568 20825
rect 27068 20748 27120 20800
rect 27620 20748 27672 20800
rect 29736 20816 29788 20868
rect 34888 20816 34940 20868
rect 35348 20816 35400 20868
rect 31024 20748 31076 20800
rect 41604 20816 41656 20868
rect 41788 20816 41840 20868
rect 43904 20927 43956 20936
rect 43904 20893 43913 20927
rect 43913 20893 43947 20927
rect 43947 20893 43956 20927
rect 43904 20884 43956 20893
rect 44272 20927 44324 20936
rect 44272 20893 44281 20927
rect 44281 20893 44315 20927
rect 44315 20893 44324 20927
rect 44272 20884 44324 20893
rect 42616 20791 42668 20800
rect 42616 20757 42625 20791
rect 42625 20757 42659 20791
rect 42659 20757 42668 20791
rect 42616 20748 42668 20757
rect 44088 20748 44140 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 6092 20587 6144 20596
rect 6092 20553 6101 20587
rect 6101 20553 6135 20587
rect 6135 20553 6144 20587
rect 6092 20544 6144 20553
rect 8576 20544 8628 20596
rect 2688 20476 2740 20528
rect 8484 20476 8536 20528
rect 9036 20476 9088 20528
rect 9864 20476 9916 20528
rect 11336 20544 11388 20596
rect 12440 20544 12492 20596
rect 13268 20544 13320 20596
rect 13360 20544 13412 20596
rect 14556 20544 14608 20596
rect 16028 20544 16080 20596
rect 19524 20544 19576 20596
rect 3332 20408 3384 20460
rect 4160 20408 4212 20460
rect 5724 20451 5776 20460
rect 5724 20417 5733 20451
rect 5733 20417 5767 20451
rect 5767 20417 5776 20451
rect 5724 20408 5776 20417
rect 5908 20451 5960 20460
rect 5908 20417 5917 20451
rect 5917 20417 5951 20451
rect 5951 20417 5960 20451
rect 5908 20408 5960 20417
rect 7564 20408 7616 20460
rect 3424 20383 3476 20392
rect 3424 20349 3433 20383
rect 3433 20349 3467 20383
rect 3467 20349 3476 20383
rect 3424 20340 3476 20349
rect 6000 20340 6052 20392
rect 8116 20340 8168 20392
rect 9588 20451 9640 20460
rect 9588 20417 9597 20451
rect 9597 20417 9631 20451
rect 9631 20417 9640 20451
rect 9588 20408 9640 20417
rect 9772 20408 9824 20460
rect 10048 20408 10100 20460
rect 10232 20451 10284 20460
rect 10232 20417 10241 20451
rect 10241 20417 10275 20451
rect 10275 20417 10284 20451
rect 10232 20408 10284 20417
rect 10324 20451 10376 20460
rect 10324 20417 10338 20451
rect 10338 20417 10372 20451
rect 10372 20417 10376 20451
rect 10324 20408 10376 20417
rect 10968 20476 11020 20528
rect 13176 20476 13228 20528
rect 11888 20408 11940 20460
rect 9956 20272 10008 20324
rect 10232 20272 10284 20324
rect 10508 20315 10560 20324
rect 10508 20281 10517 20315
rect 10517 20281 10551 20315
rect 10551 20281 10560 20315
rect 10508 20272 10560 20281
rect 10692 20340 10744 20392
rect 13084 20408 13136 20460
rect 15568 20476 15620 20528
rect 13728 20408 13780 20460
rect 13912 20408 13964 20460
rect 14740 20451 14792 20460
rect 14740 20417 14749 20451
rect 14749 20417 14783 20451
rect 14783 20417 14792 20451
rect 14740 20408 14792 20417
rect 15660 20451 15712 20460
rect 15660 20417 15669 20451
rect 15669 20417 15703 20451
rect 15703 20417 15712 20451
rect 15660 20408 15712 20417
rect 15844 20408 15896 20460
rect 18236 20476 18288 20528
rect 19340 20476 19392 20528
rect 20536 20544 20588 20596
rect 23112 20544 23164 20596
rect 23664 20544 23716 20596
rect 24216 20587 24268 20596
rect 24216 20553 24225 20587
rect 24225 20553 24259 20587
rect 24259 20553 24268 20587
rect 24216 20544 24268 20553
rect 24860 20544 24912 20596
rect 26516 20544 26568 20596
rect 26608 20544 26660 20596
rect 18420 20451 18472 20460
rect 18420 20417 18429 20451
rect 18429 20417 18463 20451
rect 18463 20417 18472 20451
rect 18420 20408 18472 20417
rect 19708 20408 19760 20460
rect 19892 20408 19944 20460
rect 19984 20408 20036 20460
rect 20904 20408 20956 20460
rect 21180 20451 21232 20460
rect 21180 20417 21189 20451
rect 21189 20417 21223 20451
rect 21223 20417 21232 20451
rect 21180 20408 21232 20417
rect 21548 20408 21600 20460
rect 22100 20408 22152 20460
rect 22652 20408 22704 20460
rect 23388 20408 23440 20460
rect 23756 20451 23808 20460
rect 23756 20417 23765 20451
rect 23765 20417 23799 20451
rect 23799 20417 23808 20451
rect 23756 20408 23808 20417
rect 24032 20451 24084 20460
rect 24032 20417 24041 20451
rect 24041 20417 24075 20451
rect 24075 20417 24084 20451
rect 24032 20408 24084 20417
rect 25596 20408 25648 20460
rect 13636 20340 13688 20392
rect 15476 20383 15528 20392
rect 15476 20349 15485 20383
rect 15485 20349 15519 20383
rect 15519 20349 15528 20383
rect 15476 20340 15528 20349
rect 6000 20204 6052 20256
rect 6552 20204 6604 20256
rect 9772 20204 9824 20256
rect 10784 20204 10836 20256
rect 14648 20247 14700 20256
rect 14648 20213 14657 20247
rect 14657 20213 14691 20247
rect 14691 20213 14700 20247
rect 14648 20204 14700 20213
rect 14924 20247 14976 20256
rect 14924 20213 14933 20247
rect 14933 20213 14967 20247
rect 14967 20213 14976 20247
rect 14924 20204 14976 20213
rect 16304 20247 16356 20256
rect 16304 20213 16313 20247
rect 16313 20213 16347 20247
rect 16347 20213 16356 20247
rect 16304 20204 16356 20213
rect 16856 20272 16908 20324
rect 17500 20340 17552 20392
rect 18696 20340 18748 20392
rect 18972 20340 19024 20392
rect 20352 20340 20404 20392
rect 21364 20340 21416 20392
rect 22008 20340 22060 20392
rect 23020 20340 23072 20392
rect 24124 20340 24176 20392
rect 25136 20340 25188 20392
rect 26056 20451 26108 20460
rect 26056 20417 26065 20451
rect 26065 20417 26099 20451
rect 26099 20417 26108 20451
rect 26056 20408 26108 20417
rect 26332 20451 26384 20460
rect 26332 20417 26341 20451
rect 26341 20417 26375 20451
rect 26375 20417 26384 20451
rect 26332 20408 26384 20417
rect 26792 20408 26844 20460
rect 27988 20587 28040 20596
rect 27988 20553 27997 20587
rect 27997 20553 28031 20587
rect 28031 20553 28040 20587
rect 27988 20544 28040 20553
rect 29092 20544 29144 20596
rect 26148 20340 26200 20392
rect 26424 20383 26476 20392
rect 26424 20349 26433 20383
rect 26433 20349 26467 20383
rect 26467 20349 26476 20383
rect 26424 20340 26476 20349
rect 17776 20204 17828 20256
rect 19984 20272 20036 20324
rect 18512 20204 18564 20256
rect 19616 20204 19668 20256
rect 21456 20272 21508 20324
rect 20996 20247 21048 20256
rect 20996 20213 21005 20247
rect 21005 20213 21039 20247
rect 21039 20213 21048 20247
rect 20996 20204 21048 20213
rect 22652 20204 22704 20256
rect 23112 20272 23164 20324
rect 23664 20204 23716 20256
rect 24860 20272 24912 20324
rect 25044 20272 25096 20324
rect 28724 20476 28776 20528
rect 29736 20476 29788 20528
rect 33600 20544 33652 20596
rect 33876 20544 33928 20596
rect 36176 20544 36228 20596
rect 28080 20451 28132 20460
rect 28080 20417 28089 20451
rect 28089 20417 28123 20451
rect 28123 20417 28132 20451
rect 28080 20408 28132 20417
rect 28264 20451 28316 20460
rect 28264 20417 28273 20451
rect 28273 20417 28307 20451
rect 28307 20417 28316 20451
rect 28264 20408 28316 20417
rect 29000 20451 29052 20460
rect 29000 20417 29009 20451
rect 29009 20417 29043 20451
rect 29043 20417 29052 20451
rect 29000 20408 29052 20417
rect 29276 20408 29328 20460
rect 29092 20383 29144 20392
rect 29092 20349 29101 20383
rect 29101 20349 29135 20383
rect 29135 20349 29144 20383
rect 29092 20340 29144 20349
rect 29736 20272 29788 20324
rect 30196 20476 30248 20528
rect 32404 20476 32456 20528
rect 32680 20476 32732 20528
rect 38292 20544 38344 20596
rect 39120 20544 39172 20596
rect 41604 20587 41656 20596
rect 41604 20553 41613 20587
rect 41613 20553 41647 20587
rect 41647 20553 41656 20587
rect 41604 20544 41656 20553
rect 30012 20272 30064 20324
rect 23848 20204 23900 20256
rect 25964 20204 26016 20256
rect 26056 20204 26108 20256
rect 26976 20247 27028 20256
rect 26976 20213 26985 20247
rect 26985 20213 27019 20247
rect 27019 20213 27028 20247
rect 26976 20204 27028 20213
rect 27620 20247 27672 20256
rect 27620 20213 27629 20247
rect 27629 20213 27663 20247
rect 27663 20213 27672 20247
rect 27620 20204 27672 20213
rect 29000 20247 29052 20256
rect 29000 20213 29009 20247
rect 29009 20213 29043 20247
rect 29043 20213 29052 20247
rect 29000 20204 29052 20213
rect 29276 20204 29328 20256
rect 29368 20204 29420 20256
rect 34428 20408 34480 20460
rect 36820 20476 36872 20528
rect 38476 20476 38528 20528
rect 40776 20476 40828 20528
rect 34612 20340 34664 20392
rect 36176 20340 36228 20392
rect 37096 20408 37148 20460
rect 41788 20451 41840 20460
rect 41788 20417 41797 20451
rect 41797 20417 41831 20451
rect 41831 20417 41840 20451
rect 41788 20408 41840 20417
rect 41972 20408 42024 20460
rect 36912 20383 36964 20392
rect 36912 20349 36921 20383
rect 36921 20349 36955 20383
rect 36955 20349 36964 20383
rect 36912 20340 36964 20349
rect 37188 20340 37240 20392
rect 37924 20340 37976 20392
rect 31852 20272 31904 20324
rect 42616 20340 42668 20392
rect 30288 20247 30340 20256
rect 30288 20213 30297 20247
rect 30297 20213 30331 20247
rect 30331 20213 30340 20247
rect 30288 20204 30340 20213
rect 30840 20204 30892 20256
rect 31668 20204 31720 20256
rect 33876 20204 33928 20256
rect 34796 20204 34848 20256
rect 36360 20204 36412 20256
rect 38660 20272 38712 20324
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 5908 20000 5960 20052
rect 9220 20000 9272 20052
rect 9404 20000 9456 20052
rect 10232 20000 10284 20052
rect 12716 20000 12768 20052
rect 5724 19932 5776 19984
rect 3884 19864 3936 19916
rect 6644 19864 6696 19916
rect 6736 19907 6788 19916
rect 6736 19873 6745 19907
rect 6745 19873 6779 19907
rect 6779 19873 6788 19907
rect 6736 19864 6788 19873
rect 3332 19839 3384 19848
rect 3332 19805 3341 19839
rect 3341 19805 3375 19839
rect 3375 19805 3384 19839
rect 3332 19796 3384 19805
rect 4804 19839 4856 19848
rect 4804 19805 4813 19839
rect 4813 19805 4847 19839
rect 4847 19805 4856 19839
rect 4804 19796 4856 19805
rect 5264 19839 5316 19848
rect 5264 19805 5267 19839
rect 5267 19805 5316 19839
rect 5264 19796 5316 19805
rect 6368 19796 6420 19848
rect 7472 19907 7524 19916
rect 7472 19873 7481 19907
rect 7481 19873 7515 19907
rect 7515 19873 7524 19907
rect 7472 19864 7524 19873
rect 8300 19864 8352 19916
rect 8852 19864 8904 19916
rect 2412 19660 2464 19712
rect 3240 19771 3292 19780
rect 3240 19737 3249 19771
rect 3249 19737 3283 19771
rect 3283 19737 3292 19771
rect 3240 19728 3292 19737
rect 4068 19728 4120 19780
rect 4620 19728 4672 19780
rect 5356 19728 5408 19780
rect 6552 19728 6604 19780
rect 8484 19796 8536 19848
rect 7472 19728 7524 19780
rect 8944 19839 8996 19848
rect 8944 19805 8953 19839
rect 8953 19805 8987 19839
rect 8987 19805 8996 19839
rect 8944 19796 8996 19805
rect 9036 19796 9088 19848
rect 10876 19932 10928 19984
rect 13360 20000 13412 20052
rect 13636 20000 13688 20052
rect 14740 20000 14792 20052
rect 15384 20000 15436 20052
rect 16028 20043 16080 20052
rect 16028 20009 16037 20043
rect 16037 20009 16071 20043
rect 16071 20009 16080 20043
rect 16028 20000 16080 20009
rect 16488 20000 16540 20052
rect 18972 20000 19024 20052
rect 23848 20000 23900 20052
rect 24308 20000 24360 20052
rect 25504 20043 25556 20052
rect 25504 20009 25513 20043
rect 25513 20009 25547 20043
rect 25547 20009 25556 20043
rect 25504 20000 25556 20009
rect 25596 20000 25648 20052
rect 25872 20000 25924 20052
rect 26332 20000 26384 20052
rect 26516 20043 26568 20052
rect 26516 20009 26525 20043
rect 26525 20009 26559 20043
rect 26559 20009 26568 20043
rect 26516 20000 26568 20009
rect 28816 20000 28868 20052
rect 13084 19932 13136 19984
rect 13728 19932 13780 19984
rect 13820 19932 13872 19984
rect 18512 19932 18564 19984
rect 9772 19864 9824 19916
rect 11520 19864 11572 19916
rect 9496 19796 9548 19848
rect 10416 19796 10468 19848
rect 10968 19796 11020 19848
rect 12164 19796 12216 19848
rect 14464 19864 14516 19916
rect 14556 19864 14608 19916
rect 15108 19864 15160 19916
rect 15568 19864 15620 19916
rect 13084 19839 13136 19848
rect 13084 19805 13093 19839
rect 13093 19805 13127 19839
rect 13127 19805 13136 19839
rect 13084 19796 13136 19805
rect 15200 19796 15252 19848
rect 15936 19839 15988 19848
rect 15936 19805 15945 19839
rect 15945 19805 15979 19839
rect 15979 19805 15988 19839
rect 15936 19796 15988 19805
rect 16488 19796 16540 19848
rect 18052 19839 18104 19848
rect 18052 19805 18061 19839
rect 18061 19805 18095 19839
rect 18095 19805 18104 19839
rect 18052 19796 18104 19805
rect 18236 19839 18288 19848
rect 18236 19805 18245 19839
rect 18245 19805 18279 19839
rect 18279 19805 18288 19839
rect 18236 19796 18288 19805
rect 9404 19728 9456 19780
rect 13820 19728 13872 19780
rect 15016 19728 15068 19780
rect 15844 19728 15896 19780
rect 16396 19728 16448 19780
rect 8208 19660 8260 19712
rect 8300 19703 8352 19712
rect 8300 19669 8309 19703
rect 8309 19669 8343 19703
rect 8343 19669 8352 19703
rect 8300 19660 8352 19669
rect 8392 19660 8444 19712
rect 15660 19660 15712 19712
rect 17868 19660 17920 19712
rect 18512 19796 18564 19848
rect 19616 19864 19668 19916
rect 19800 19864 19852 19916
rect 20076 19864 20128 19916
rect 24124 19864 24176 19916
rect 23480 19796 23532 19848
rect 23572 19839 23624 19848
rect 23572 19805 23581 19839
rect 23581 19805 23615 19839
rect 23615 19805 23624 19839
rect 23572 19796 23624 19805
rect 23756 19796 23808 19848
rect 25412 19932 25464 19984
rect 24584 19864 24636 19916
rect 25688 19907 25740 19916
rect 25688 19873 25697 19907
rect 25697 19873 25731 19907
rect 25731 19873 25740 19907
rect 25688 19864 25740 19873
rect 26424 19864 26476 19916
rect 25596 19796 25648 19848
rect 25780 19839 25832 19848
rect 25780 19805 25789 19839
rect 25789 19805 25823 19839
rect 25823 19805 25832 19839
rect 25780 19796 25832 19805
rect 27252 19864 27304 19916
rect 29368 19907 29420 19916
rect 29368 19873 29377 19907
rect 29377 19873 29411 19907
rect 29411 19873 29420 19907
rect 29368 19864 29420 19873
rect 29828 19907 29880 19916
rect 29828 19873 29837 19907
rect 29837 19873 29871 19907
rect 29871 19873 29880 19907
rect 29828 19864 29880 19873
rect 30564 20000 30616 20052
rect 31392 20000 31444 20052
rect 33600 20043 33652 20052
rect 33600 20009 33609 20043
rect 33609 20009 33643 20043
rect 33643 20009 33652 20043
rect 33600 20000 33652 20009
rect 33876 20000 33928 20052
rect 35440 20000 35492 20052
rect 35532 20043 35584 20052
rect 35532 20009 35541 20043
rect 35541 20009 35575 20043
rect 35575 20009 35584 20043
rect 35532 20000 35584 20009
rect 37004 20000 37056 20052
rect 37188 20000 37240 20052
rect 30288 19932 30340 19984
rect 26792 19839 26844 19848
rect 26792 19805 26801 19839
rect 26801 19805 26835 19839
rect 26835 19805 26844 19839
rect 26792 19796 26844 19805
rect 28908 19796 28960 19848
rect 31576 19864 31628 19916
rect 32220 19864 32272 19916
rect 22100 19728 22152 19780
rect 22192 19728 22244 19780
rect 19156 19660 19208 19712
rect 20996 19660 21048 19712
rect 22008 19660 22060 19712
rect 23112 19728 23164 19780
rect 23388 19728 23440 19780
rect 24584 19771 24636 19780
rect 24584 19737 24593 19771
rect 24593 19737 24627 19771
rect 24627 19737 24636 19771
rect 24584 19728 24636 19737
rect 29000 19771 29052 19780
rect 29000 19737 29009 19771
rect 29009 19737 29043 19771
rect 29043 19737 29052 19771
rect 29000 19728 29052 19737
rect 29092 19728 29144 19780
rect 30012 19771 30064 19780
rect 30012 19737 30021 19771
rect 30021 19737 30055 19771
rect 30055 19737 30064 19771
rect 30012 19728 30064 19737
rect 30472 19728 30524 19780
rect 26332 19703 26384 19712
rect 26332 19669 26341 19703
rect 26341 19669 26375 19703
rect 26375 19669 26384 19703
rect 26332 19660 26384 19669
rect 26516 19660 26568 19712
rect 30196 19660 30248 19712
rect 32680 19864 32732 19916
rect 34060 19907 34112 19916
rect 34060 19873 34069 19907
rect 34069 19873 34103 19907
rect 34103 19873 34112 19907
rect 34060 19864 34112 19873
rect 33140 19796 33192 19848
rect 33416 19796 33468 19848
rect 33508 19839 33560 19848
rect 33508 19805 33517 19839
rect 33517 19805 33551 19839
rect 33551 19805 33560 19839
rect 33508 19796 33560 19805
rect 34520 19864 34572 19916
rect 34612 19864 34664 19916
rect 34428 19796 34480 19848
rect 35440 19839 35492 19848
rect 35440 19805 35449 19839
rect 35449 19805 35483 19839
rect 35483 19805 35492 19839
rect 35440 19796 35492 19805
rect 32220 19728 32272 19780
rect 32772 19703 32824 19712
rect 32772 19669 32781 19703
rect 32781 19669 32815 19703
rect 32815 19669 32824 19703
rect 32772 19660 32824 19669
rect 32956 19728 33008 19780
rect 33968 19771 34020 19780
rect 33968 19737 33977 19771
rect 33977 19737 34011 19771
rect 34011 19737 34020 19771
rect 33968 19728 34020 19737
rect 35532 19728 35584 19780
rect 33048 19660 33100 19712
rect 34060 19660 34112 19712
rect 34244 19660 34296 19712
rect 38752 19864 38804 19916
rect 39672 19839 39724 19848
rect 39672 19805 39681 19839
rect 39681 19805 39715 19839
rect 39715 19805 39724 19839
rect 39672 19796 39724 19805
rect 40776 19839 40828 19848
rect 40776 19805 40785 19839
rect 40785 19805 40819 19839
rect 40819 19805 40828 19839
rect 44180 19864 44232 19916
rect 40776 19796 40828 19805
rect 43260 19796 43312 19848
rect 37464 19703 37516 19712
rect 37464 19669 37473 19703
rect 37473 19669 37507 19703
rect 37507 19669 37516 19703
rect 37464 19660 37516 19669
rect 38568 19660 38620 19712
rect 40408 19660 40460 19712
rect 44456 19703 44508 19712
rect 44456 19669 44465 19703
rect 44465 19669 44499 19703
rect 44499 19669 44508 19703
rect 44456 19660 44508 19669
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 2688 19456 2740 19508
rect 2412 19431 2464 19440
rect 2412 19397 2421 19431
rect 2421 19397 2455 19431
rect 2455 19397 2464 19431
rect 2412 19388 2464 19397
rect 8392 19456 8444 19508
rect 8944 19456 8996 19508
rect 9772 19456 9824 19508
rect 10692 19456 10744 19508
rect 12164 19456 12216 19508
rect 12440 19456 12492 19508
rect 12808 19456 12860 19508
rect 6184 19388 6236 19440
rect 8024 19388 8076 19440
rect 2596 19363 2648 19372
rect 2596 19329 2610 19363
rect 2610 19329 2644 19363
rect 2644 19329 2648 19363
rect 2596 19320 2648 19329
rect 2780 19363 2832 19372
rect 2780 19329 2806 19363
rect 2806 19329 2832 19363
rect 2780 19320 2832 19329
rect 3148 19320 3200 19372
rect 6460 19320 6512 19372
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 6736 19363 6788 19372
rect 6736 19329 6745 19363
rect 6745 19329 6779 19363
rect 6779 19329 6788 19363
rect 6736 19320 6788 19329
rect 8576 19363 8628 19372
rect 8576 19329 8585 19363
rect 8585 19329 8619 19363
rect 8619 19329 8628 19363
rect 8576 19320 8628 19329
rect 10140 19320 10192 19372
rect 10416 19363 10468 19372
rect 10416 19329 10425 19363
rect 10425 19329 10459 19363
rect 10459 19329 10468 19363
rect 10416 19320 10468 19329
rect 10692 19363 10744 19372
rect 10692 19329 10695 19363
rect 10695 19329 10744 19363
rect 2504 19252 2556 19304
rect 8484 19252 8536 19304
rect 9312 19252 9364 19304
rect 9680 19252 9732 19304
rect 10692 19320 10744 19329
rect 3608 19184 3660 19236
rect 6000 19184 6052 19236
rect 6092 19184 6144 19236
rect 6644 19184 6696 19236
rect 10876 19320 10928 19372
rect 12072 19320 12124 19372
rect 14372 19388 14424 19440
rect 14648 19388 14700 19440
rect 18420 19456 18472 19508
rect 12716 19320 12768 19372
rect 12164 19184 12216 19236
rect 12624 19184 12676 19236
rect 13544 19363 13596 19372
rect 13544 19329 13547 19363
rect 13547 19329 13596 19363
rect 13268 19252 13320 19304
rect 13544 19320 13596 19329
rect 13820 19320 13872 19372
rect 14832 19320 14884 19372
rect 15200 19363 15252 19372
rect 15200 19329 15203 19363
rect 15203 19329 15252 19363
rect 14556 19252 14608 19304
rect 13728 19184 13780 19236
rect 15200 19320 15252 19329
rect 15476 19363 15528 19372
rect 15476 19329 15485 19363
rect 15485 19329 15519 19363
rect 15519 19329 15528 19363
rect 15476 19320 15528 19329
rect 15292 19252 15344 19304
rect 16672 19388 16724 19440
rect 19248 19456 19300 19508
rect 20168 19499 20220 19508
rect 20168 19465 20177 19499
rect 20177 19465 20211 19499
rect 20211 19465 20220 19499
rect 20168 19456 20220 19465
rect 20720 19456 20772 19508
rect 15936 19320 15988 19372
rect 18788 19363 18840 19372
rect 18788 19329 18797 19363
rect 18797 19329 18831 19363
rect 18831 19329 18840 19363
rect 18788 19320 18840 19329
rect 18880 19363 18932 19372
rect 18880 19329 18889 19363
rect 18889 19329 18923 19363
rect 18923 19329 18932 19363
rect 18880 19320 18932 19329
rect 19524 19320 19576 19372
rect 19616 19363 19668 19372
rect 19616 19329 19625 19363
rect 19625 19329 19659 19363
rect 19659 19329 19668 19363
rect 19616 19320 19668 19329
rect 21548 19388 21600 19440
rect 23664 19456 23716 19508
rect 24584 19456 24636 19508
rect 29920 19456 29972 19508
rect 32128 19456 32180 19508
rect 32404 19456 32456 19508
rect 34704 19456 34756 19508
rect 40776 19456 40828 19508
rect 44088 19456 44140 19508
rect 19984 19363 20036 19372
rect 19984 19329 19993 19363
rect 19993 19329 20027 19363
rect 20027 19329 20036 19363
rect 19984 19320 20036 19329
rect 20720 19320 20772 19372
rect 15936 19184 15988 19236
rect 4620 19116 4672 19168
rect 8300 19116 8352 19168
rect 11704 19116 11756 19168
rect 16856 19184 16908 19236
rect 17408 19184 17460 19236
rect 18144 19184 18196 19236
rect 19524 19184 19576 19236
rect 16580 19116 16632 19168
rect 18512 19116 18564 19168
rect 18604 19159 18656 19168
rect 18604 19125 18613 19159
rect 18613 19125 18647 19159
rect 18647 19125 18656 19159
rect 18604 19116 18656 19125
rect 19248 19116 19300 19168
rect 20168 19252 20220 19304
rect 20628 19252 20680 19304
rect 22008 19363 22060 19372
rect 22008 19329 22017 19363
rect 22017 19329 22051 19363
rect 22051 19329 22060 19363
rect 22008 19320 22060 19329
rect 23112 19388 23164 19440
rect 23388 19388 23440 19440
rect 33508 19388 33560 19440
rect 34060 19431 34112 19440
rect 34060 19397 34069 19431
rect 34069 19397 34103 19431
rect 34103 19397 34112 19431
rect 34060 19388 34112 19397
rect 34152 19388 34204 19440
rect 22192 19320 22244 19372
rect 25964 19320 26016 19372
rect 26976 19320 27028 19372
rect 27804 19320 27856 19372
rect 27988 19320 28040 19372
rect 31300 19320 31352 19372
rect 34244 19363 34296 19372
rect 34244 19329 34253 19363
rect 34253 19329 34287 19363
rect 34287 19329 34296 19363
rect 34244 19320 34296 19329
rect 41052 19388 41104 19440
rect 38568 19363 38620 19372
rect 38568 19329 38577 19363
rect 38577 19329 38611 19363
rect 38611 19329 38620 19363
rect 38568 19320 38620 19329
rect 38660 19320 38712 19372
rect 40316 19320 40368 19372
rect 40408 19363 40460 19372
rect 40408 19329 40417 19363
rect 40417 19329 40451 19363
rect 40451 19329 40460 19363
rect 40408 19320 40460 19329
rect 42432 19363 42484 19372
rect 42432 19329 42441 19363
rect 42441 19329 42475 19363
rect 42475 19329 42484 19363
rect 42432 19320 42484 19329
rect 42708 19363 42760 19372
rect 42708 19329 42742 19363
rect 42742 19329 42760 19363
rect 42708 19320 42760 19329
rect 22928 19252 22980 19304
rect 24032 19252 24084 19304
rect 26240 19252 26292 19304
rect 27896 19252 27948 19304
rect 28080 19252 28132 19304
rect 29000 19252 29052 19304
rect 21456 19184 21508 19236
rect 21272 19159 21324 19168
rect 21272 19125 21281 19159
rect 21281 19125 21315 19159
rect 21315 19125 21324 19159
rect 21272 19116 21324 19125
rect 21732 19116 21784 19168
rect 21916 19116 21968 19168
rect 22100 19159 22152 19168
rect 22100 19125 22109 19159
rect 22109 19125 22143 19159
rect 22143 19125 22152 19159
rect 22100 19116 22152 19125
rect 22284 19184 22336 19236
rect 31668 19184 31720 19236
rect 31852 19184 31904 19236
rect 32220 19295 32272 19304
rect 32220 19261 32229 19295
rect 32229 19261 32263 19295
rect 32263 19261 32272 19295
rect 32220 19252 32272 19261
rect 36544 19252 36596 19304
rect 38292 19252 38344 19304
rect 38476 19184 38528 19236
rect 25136 19116 25188 19168
rect 25688 19116 25740 19168
rect 27068 19116 27120 19168
rect 31392 19116 31444 19168
rect 31484 19159 31536 19168
rect 31484 19125 31493 19159
rect 31493 19125 31527 19159
rect 31527 19125 31536 19159
rect 31484 19116 31536 19125
rect 32128 19159 32180 19168
rect 32128 19125 32137 19159
rect 32137 19125 32171 19159
rect 32171 19125 32180 19159
rect 32128 19116 32180 19125
rect 33508 19116 33560 19168
rect 43812 19227 43864 19236
rect 43812 19193 43821 19227
rect 43821 19193 43855 19227
rect 43855 19193 43864 19227
rect 43812 19184 43864 19193
rect 38844 19116 38896 19168
rect 40040 19159 40092 19168
rect 40040 19125 40049 19159
rect 40049 19125 40083 19159
rect 40083 19125 40092 19159
rect 40040 19116 40092 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 2504 18955 2556 18964
rect 2504 18921 2513 18955
rect 2513 18921 2547 18955
rect 2547 18921 2556 18955
rect 2504 18912 2556 18921
rect 3424 18955 3476 18964
rect 3424 18921 3433 18955
rect 3433 18921 3467 18955
rect 3467 18921 3476 18955
rect 3424 18912 3476 18921
rect 4620 18912 4672 18964
rect 6276 18912 6328 18964
rect 7196 18912 7248 18964
rect 2872 18844 2924 18896
rect 4068 18844 4120 18896
rect 6368 18844 6420 18896
rect 6552 18844 6604 18896
rect 6184 18819 6236 18828
rect 3240 18751 3292 18760
rect 3240 18717 3249 18751
rect 3249 18717 3283 18751
rect 3283 18717 3292 18751
rect 3240 18708 3292 18717
rect 3424 18708 3476 18760
rect 3884 18751 3936 18760
rect 3884 18717 3893 18751
rect 3893 18717 3927 18751
rect 3927 18717 3936 18751
rect 3884 18708 3936 18717
rect 3976 18708 4028 18760
rect 4804 18708 4856 18760
rect 5264 18708 5316 18760
rect 6184 18785 6193 18819
rect 6193 18785 6227 18819
rect 6227 18785 6236 18819
rect 6184 18776 6236 18785
rect 7104 18819 7156 18828
rect 7104 18785 7113 18819
rect 7113 18785 7147 18819
rect 7147 18785 7156 18819
rect 7104 18776 7156 18785
rect 6276 18708 6328 18760
rect 6460 18751 6512 18760
rect 6460 18717 6469 18751
rect 6469 18717 6503 18751
rect 6503 18717 6512 18751
rect 6460 18708 6512 18717
rect 2412 18683 2464 18692
rect 2412 18649 2421 18683
rect 2421 18649 2455 18683
rect 2455 18649 2464 18683
rect 2412 18640 2464 18649
rect 3332 18640 3384 18692
rect 4712 18640 4764 18692
rect 5080 18640 5132 18692
rect 5816 18640 5868 18692
rect 5908 18572 5960 18624
rect 6092 18572 6144 18624
rect 7564 18708 7616 18760
rect 8208 18844 8260 18896
rect 9220 18844 9272 18896
rect 7932 18776 7984 18828
rect 8024 18751 8076 18760
rect 8024 18717 8033 18751
rect 8033 18717 8067 18751
rect 8067 18717 8076 18751
rect 8024 18708 8076 18717
rect 8300 18751 8352 18760
rect 8300 18717 8309 18751
rect 8309 18717 8343 18751
rect 8343 18717 8352 18751
rect 8300 18708 8352 18717
rect 8208 18572 8260 18624
rect 8484 18708 8536 18760
rect 8944 18708 8996 18760
rect 9864 18912 9916 18964
rect 10508 18955 10560 18964
rect 10508 18921 10517 18955
rect 10517 18921 10551 18955
rect 10551 18921 10560 18955
rect 10508 18912 10560 18921
rect 9956 18844 10008 18896
rect 9680 18751 9732 18760
rect 9680 18717 9683 18751
rect 9683 18717 9732 18751
rect 9680 18708 9732 18717
rect 9864 18708 9916 18760
rect 9036 18572 9088 18624
rect 10140 18683 10192 18692
rect 10140 18649 10149 18683
rect 10149 18649 10183 18683
rect 10183 18649 10192 18683
rect 10140 18640 10192 18649
rect 10232 18683 10284 18692
rect 10232 18649 10241 18683
rect 10241 18649 10275 18683
rect 10275 18649 10284 18683
rect 10232 18640 10284 18649
rect 10692 18751 10744 18760
rect 10692 18717 10701 18751
rect 10701 18717 10735 18751
rect 10735 18717 10744 18751
rect 10692 18708 10744 18717
rect 11980 18844 12032 18896
rect 12440 18776 12492 18828
rect 12164 18708 12216 18760
rect 10968 18683 11020 18692
rect 10968 18649 10977 18683
rect 10977 18649 11011 18683
rect 11011 18649 11020 18683
rect 10968 18640 11020 18649
rect 12348 18640 12400 18692
rect 12808 18887 12860 18896
rect 12808 18853 12817 18887
rect 12817 18853 12851 18887
rect 12851 18853 12860 18887
rect 12808 18844 12860 18853
rect 12716 18776 12768 18828
rect 13360 18844 13412 18896
rect 13452 18844 13504 18896
rect 15476 18844 15528 18896
rect 17040 18955 17092 18964
rect 17040 18921 17049 18955
rect 17049 18921 17083 18955
rect 17083 18921 17092 18955
rect 17040 18912 17092 18921
rect 20628 18912 20680 18964
rect 21732 18955 21784 18964
rect 21732 18921 21741 18955
rect 21741 18921 21775 18955
rect 21775 18921 21784 18955
rect 21732 18912 21784 18921
rect 23480 18912 23532 18964
rect 27528 18912 27580 18964
rect 27896 18912 27948 18964
rect 28908 18955 28960 18964
rect 19248 18844 19300 18896
rect 21180 18844 21232 18896
rect 13268 18776 13320 18828
rect 14924 18776 14976 18828
rect 22100 18844 22152 18896
rect 12716 18640 12768 18692
rect 13636 18708 13688 18760
rect 14464 18751 14516 18760
rect 14464 18717 14473 18751
rect 14473 18717 14507 18751
rect 14507 18717 14516 18751
rect 14464 18708 14516 18717
rect 14648 18751 14700 18760
rect 14648 18717 14657 18751
rect 14657 18717 14691 18751
rect 14691 18717 14700 18751
rect 14648 18708 14700 18717
rect 14832 18751 14884 18760
rect 14832 18717 14841 18751
rect 14841 18717 14875 18751
rect 14875 18717 14884 18751
rect 14832 18708 14884 18717
rect 13176 18683 13228 18692
rect 13176 18649 13185 18683
rect 13185 18649 13219 18683
rect 13219 18649 13228 18683
rect 13176 18640 13228 18649
rect 11888 18572 11940 18624
rect 12164 18572 12216 18624
rect 14372 18640 14424 18692
rect 13452 18572 13504 18624
rect 16948 18708 17000 18760
rect 17224 18708 17276 18760
rect 19156 18708 19208 18760
rect 19984 18708 20036 18760
rect 21548 18751 21600 18760
rect 21548 18717 21557 18751
rect 21557 18717 21591 18751
rect 21591 18717 21600 18751
rect 21548 18708 21600 18717
rect 21916 18776 21968 18828
rect 23480 18776 23532 18828
rect 24860 18776 24912 18828
rect 28908 18921 28917 18955
rect 28917 18921 28951 18955
rect 28951 18921 28960 18955
rect 28908 18912 28960 18921
rect 30104 18912 30156 18964
rect 31852 18912 31904 18964
rect 37464 18955 37516 18964
rect 37464 18921 37473 18955
rect 37473 18921 37507 18955
rect 37507 18921 37516 18955
rect 37464 18912 37516 18921
rect 36544 18844 36596 18896
rect 38660 18912 38712 18964
rect 40040 18844 40092 18896
rect 41788 18912 41840 18964
rect 21824 18751 21876 18760
rect 21824 18717 21833 18751
rect 21833 18717 21867 18751
rect 21867 18717 21876 18751
rect 21824 18708 21876 18717
rect 24032 18708 24084 18760
rect 28264 18751 28316 18760
rect 28264 18717 28273 18751
rect 28273 18717 28307 18751
rect 28307 18717 28316 18751
rect 28264 18708 28316 18717
rect 28540 18708 28592 18760
rect 28816 18708 28868 18760
rect 28908 18708 28960 18760
rect 29552 18776 29604 18828
rect 31024 18776 31076 18828
rect 31760 18776 31812 18828
rect 37280 18776 37332 18828
rect 29092 18751 29144 18760
rect 29092 18717 29101 18751
rect 29101 18717 29135 18751
rect 29135 18717 29144 18751
rect 29092 18708 29144 18717
rect 29184 18751 29236 18760
rect 29184 18717 29193 18751
rect 29193 18717 29227 18751
rect 29227 18717 29236 18751
rect 29184 18708 29236 18717
rect 30748 18708 30800 18760
rect 20720 18640 20772 18692
rect 20904 18640 20956 18692
rect 32588 18708 32640 18760
rect 37004 18708 37056 18760
rect 37096 18708 37148 18760
rect 41052 18819 41104 18828
rect 41052 18785 41061 18819
rect 41061 18785 41095 18819
rect 41095 18785 41104 18819
rect 41052 18776 41104 18785
rect 43812 18819 43864 18828
rect 43812 18785 43821 18819
rect 43821 18785 43855 18819
rect 43855 18785 43864 18819
rect 43812 18776 43864 18785
rect 38108 18751 38160 18760
rect 38108 18717 38117 18751
rect 38117 18717 38151 18751
rect 38151 18717 38160 18751
rect 38108 18708 38160 18717
rect 38292 18751 38344 18760
rect 38292 18717 38301 18751
rect 38301 18717 38335 18751
rect 38335 18717 38344 18751
rect 38292 18708 38344 18717
rect 38936 18708 38988 18760
rect 22100 18640 22152 18692
rect 16580 18615 16632 18624
rect 16580 18581 16589 18615
rect 16589 18581 16623 18615
rect 16623 18581 16632 18615
rect 16580 18572 16632 18581
rect 17224 18572 17276 18624
rect 17500 18572 17552 18624
rect 17776 18572 17828 18624
rect 19524 18572 19576 18624
rect 21548 18572 21600 18624
rect 22376 18572 22428 18624
rect 28540 18572 28592 18624
rect 28724 18615 28776 18624
rect 28724 18581 28733 18615
rect 28733 18581 28767 18615
rect 28767 18581 28776 18615
rect 28724 18572 28776 18581
rect 29368 18683 29420 18692
rect 29368 18649 29377 18683
rect 29377 18649 29411 18683
rect 29411 18649 29420 18683
rect 29368 18640 29420 18649
rect 30656 18640 30708 18692
rect 31484 18640 31536 18692
rect 34980 18640 35032 18692
rect 38752 18640 38804 18692
rect 40316 18751 40368 18760
rect 40316 18717 40325 18751
rect 40325 18717 40359 18751
rect 40359 18717 40368 18751
rect 40316 18708 40368 18717
rect 40868 18708 40920 18760
rect 43168 18751 43220 18760
rect 43168 18717 43177 18751
rect 43177 18717 43211 18751
rect 43211 18717 43220 18751
rect 43168 18708 43220 18717
rect 41144 18640 41196 18692
rect 41604 18640 41656 18692
rect 41696 18640 41748 18692
rect 32312 18572 32364 18624
rect 34060 18572 34112 18624
rect 37188 18572 37240 18624
rect 39580 18572 39632 18624
rect 40132 18572 40184 18624
rect 42524 18615 42576 18624
rect 42524 18581 42533 18615
rect 42533 18581 42567 18615
rect 42567 18581 42576 18615
rect 42524 18572 42576 18581
rect 43260 18615 43312 18624
rect 43260 18581 43269 18615
rect 43269 18581 43303 18615
rect 43303 18581 43312 18615
rect 43260 18572 43312 18581
rect 44456 18615 44508 18624
rect 44456 18581 44465 18615
rect 44465 18581 44499 18615
rect 44499 18581 44508 18615
rect 44456 18572 44508 18581
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 3608 18368 3660 18420
rect 4804 18368 4856 18420
rect 2136 18232 2188 18284
rect 2504 18275 2556 18284
rect 2504 18241 2513 18275
rect 2513 18241 2547 18275
rect 2547 18241 2556 18275
rect 2504 18232 2556 18241
rect 2872 18275 2924 18284
rect 2872 18241 2881 18275
rect 2881 18241 2915 18275
rect 2915 18241 2924 18275
rect 2872 18232 2924 18241
rect 3424 18232 3476 18284
rect 2596 18207 2648 18216
rect 2596 18173 2605 18207
rect 2605 18173 2639 18207
rect 2639 18173 2648 18207
rect 2596 18164 2648 18173
rect 3056 18207 3108 18216
rect 3056 18173 3065 18207
rect 3065 18173 3099 18207
rect 3099 18173 3108 18207
rect 3056 18164 3108 18173
rect 4620 18232 4672 18284
rect 5908 18300 5960 18352
rect 6828 18368 6880 18420
rect 10140 18368 10192 18420
rect 10232 18368 10284 18420
rect 11888 18368 11940 18420
rect 12348 18368 12400 18420
rect 13268 18368 13320 18420
rect 13360 18368 13412 18420
rect 8208 18300 8260 18352
rect 8300 18343 8352 18352
rect 8300 18309 8309 18343
rect 8309 18309 8343 18343
rect 8343 18309 8352 18343
rect 8300 18300 8352 18309
rect 8392 18343 8444 18352
rect 8392 18309 8401 18343
rect 8401 18309 8435 18343
rect 8435 18309 8444 18343
rect 8392 18300 8444 18309
rect 9680 18300 9732 18352
rect 10692 18300 10744 18352
rect 13452 18300 13504 18352
rect 13912 18343 13964 18352
rect 13912 18309 13921 18343
rect 13921 18309 13955 18343
rect 13955 18309 13964 18343
rect 13912 18300 13964 18309
rect 16028 18368 16080 18420
rect 16948 18368 17000 18420
rect 18144 18411 18196 18420
rect 18144 18377 18153 18411
rect 18153 18377 18187 18411
rect 18187 18377 18196 18411
rect 18144 18368 18196 18377
rect 19616 18368 19668 18420
rect 20904 18368 20956 18420
rect 15384 18300 15436 18352
rect 5172 18275 5224 18284
rect 5172 18241 5176 18275
rect 5176 18241 5210 18275
rect 5210 18241 5224 18275
rect 5172 18232 5224 18241
rect 5724 18275 5776 18284
rect 5724 18241 5733 18275
rect 5733 18241 5767 18275
rect 5767 18241 5776 18275
rect 5724 18232 5776 18241
rect 5816 18164 5868 18216
rect 6368 18232 6420 18284
rect 6828 18275 6880 18284
rect 6828 18241 6842 18275
rect 6842 18241 6876 18275
rect 6876 18241 6880 18275
rect 6828 18232 6880 18241
rect 7564 18232 7616 18284
rect 7932 18232 7984 18284
rect 8484 18275 8536 18284
rect 8484 18241 8498 18275
rect 8498 18241 8532 18275
rect 8532 18241 8536 18275
rect 8484 18232 8536 18241
rect 7840 18164 7892 18216
rect 9036 18275 9088 18284
rect 9036 18241 9045 18275
rect 9045 18241 9079 18275
rect 9079 18241 9088 18275
rect 9036 18232 9088 18241
rect 9220 18275 9272 18284
rect 9220 18241 9234 18275
rect 9234 18241 9268 18275
rect 9268 18241 9272 18275
rect 9220 18232 9272 18241
rect 8944 18164 8996 18216
rect 10324 18232 10376 18284
rect 9956 18164 10008 18216
rect 10140 18164 10192 18216
rect 11980 18232 12032 18284
rect 12164 18275 12216 18284
rect 12164 18241 12173 18275
rect 12173 18241 12207 18275
rect 12207 18241 12216 18275
rect 12164 18232 12216 18241
rect 12624 18232 12676 18284
rect 13176 18232 13228 18284
rect 13360 18232 13412 18284
rect 12808 18207 12860 18216
rect 12808 18173 12817 18207
rect 12817 18173 12851 18207
rect 12851 18173 12860 18207
rect 12808 18164 12860 18173
rect 12992 18164 13044 18216
rect 5448 18096 5500 18148
rect 3976 18028 4028 18080
rect 6828 18096 6880 18148
rect 7012 18139 7064 18148
rect 7012 18105 7021 18139
rect 7021 18105 7055 18139
rect 7055 18105 7064 18139
rect 7012 18096 7064 18105
rect 8484 18096 8536 18148
rect 10416 18096 10468 18148
rect 14096 18275 14148 18284
rect 14096 18241 14105 18275
rect 14105 18241 14139 18275
rect 14139 18241 14148 18275
rect 14096 18232 14148 18241
rect 14740 18275 14792 18284
rect 14740 18241 14749 18275
rect 14749 18241 14783 18275
rect 14783 18241 14792 18275
rect 14740 18232 14792 18241
rect 14924 18275 14976 18284
rect 14924 18241 14933 18275
rect 14933 18241 14967 18275
rect 14967 18241 14976 18275
rect 14924 18232 14976 18241
rect 15108 18275 15160 18284
rect 15108 18241 15117 18275
rect 15117 18241 15151 18275
rect 15151 18241 15160 18275
rect 15108 18232 15160 18241
rect 17868 18300 17920 18352
rect 18512 18300 18564 18352
rect 21456 18300 21508 18352
rect 16672 18164 16724 18216
rect 17316 18275 17368 18284
rect 17316 18241 17325 18275
rect 17325 18241 17359 18275
rect 17359 18241 17368 18275
rect 17316 18232 17368 18241
rect 17592 18232 17644 18284
rect 17684 18275 17736 18284
rect 17684 18241 17693 18275
rect 17693 18241 17727 18275
rect 17727 18241 17736 18275
rect 17684 18232 17736 18241
rect 18236 18232 18288 18284
rect 19248 18232 19300 18284
rect 19616 18275 19668 18284
rect 19616 18241 19625 18275
rect 19625 18241 19659 18275
rect 19659 18241 19668 18275
rect 19616 18232 19668 18241
rect 19800 18232 19852 18284
rect 17132 18164 17184 18216
rect 17776 18207 17828 18216
rect 17776 18173 17785 18207
rect 17785 18173 17819 18207
rect 17819 18173 17828 18207
rect 17776 18164 17828 18173
rect 19984 18164 20036 18216
rect 20168 18164 20220 18216
rect 21548 18164 21600 18216
rect 22928 18300 22980 18352
rect 23296 18411 23348 18420
rect 23296 18377 23305 18411
rect 23305 18377 23339 18411
rect 23339 18377 23348 18411
rect 23296 18368 23348 18377
rect 24032 18411 24084 18420
rect 24032 18377 24041 18411
rect 24041 18377 24075 18411
rect 24075 18377 24084 18411
rect 24032 18368 24084 18377
rect 24860 18368 24912 18420
rect 25596 18368 25648 18420
rect 22192 18275 22244 18284
rect 22192 18241 22201 18275
rect 22201 18241 22235 18275
rect 22235 18241 22244 18275
rect 22192 18232 22244 18241
rect 22376 18275 22428 18284
rect 22376 18241 22385 18275
rect 22385 18241 22419 18275
rect 22419 18241 22428 18275
rect 22376 18232 22428 18241
rect 22468 18275 22520 18284
rect 22468 18241 22477 18275
rect 22477 18241 22511 18275
rect 22511 18241 22520 18275
rect 22468 18232 22520 18241
rect 22836 18275 22888 18284
rect 22836 18241 22845 18275
rect 22845 18241 22879 18275
rect 22879 18241 22888 18275
rect 22836 18232 22888 18241
rect 23572 18275 23624 18284
rect 23572 18241 23581 18275
rect 23581 18241 23615 18275
rect 23615 18241 23624 18275
rect 23572 18232 23624 18241
rect 24032 18232 24084 18284
rect 26240 18300 26292 18352
rect 25412 18275 25464 18284
rect 25412 18241 25421 18275
rect 25421 18241 25455 18275
rect 25455 18241 25464 18275
rect 25412 18232 25464 18241
rect 26148 18232 26200 18284
rect 26516 18232 26568 18284
rect 26976 18343 27028 18352
rect 26976 18309 26985 18343
rect 26985 18309 27019 18343
rect 27019 18309 27028 18343
rect 26976 18300 27028 18309
rect 27896 18368 27948 18420
rect 29000 18368 29052 18420
rect 28264 18232 28316 18284
rect 28540 18300 28592 18352
rect 29276 18343 29328 18352
rect 29276 18309 29292 18343
rect 29292 18309 29326 18343
rect 29326 18309 29328 18343
rect 29276 18300 29328 18309
rect 30748 18368 30800 18420
rect 32588 18411 32640 18420
rect 32588 18377 32597 18411
rect 32597 18377 32631 18411
rect 32631 18377 32640 18411
rect 32588 18368 32640 18377
rect 22928 18207 22980 18216
rect 22928 18173 22937 18207
rect 22937 18173 22971 18207
rect 22971 18173 22980 18207
rect 22928 18164 22980 18173
rect 23388 18164 23440 18216
rect 27068 18207 27120 18216
rect 27068 18173 27077 18207
rect 27077 18173 27111 18207
rect 27111 18173 27120 18207
rect 27068 18164 27120 18173
rect 28448 18164 28500 18216
rect 29368 18207 29420 18216
rect 29368 18173 29377 18207
rect 29377 18173 29411 18207
rect 29411 18173 29420 18207
rect 29368 18164 29420 18173
rect 29552 18275 29604 18284
rect 29552 18241 29561 18275
rect 29561 18241 29595 18275
rect 29595 18241 29604 18275
rect 29552 18232 29604 18241
rect 31208 18275 31260 18284
rect 31208 18241 31217 18275
rect 31217 18241 31251 18275
rect 31251 18241 31260 18275
rect 31208 18232 31260 18241
rect 31392 18232 31444 18284
rect 32956 18300 33008 18352
rect 37096 18411 37148 18420
rect 37096 18377 37105 18411
rect 37105 18377 37139 18411
rect 37139 18377 37148 18411
rect 37096 18368 37148 18377
rect 40868 18411 40920 18420
rect 40868 18377 40877 18411
rect 40877 18377 40911 18411
rect 40911 18377 40920 18411
rect 40868 18368 40920 18377
rect 41604 18411 41656 18420
rect 41604 18377 41613 18411
rect 41613 18377 41647 18411
rect 41647 18377 41656 18411
rect 41604 18368 41656 18377
rect 36636 18343 36688 18352
rect 36636 18309 36645 18343
rect 36645 18309 36679 18343
rect 36679 18309 36688 18343
rect 36636 18300 36688 18309
rect 41328 18300 41380 18352
rect 31668 18232 31720 18284
rect 32312 18275 32364 18284
rect 32312 18241 32321 18275
rect 32321 18241 32355 18275
rect 32355 18241 32364 18275
rect 32312 18232 32364 18241
rect 32772 18232 32824 18284
rect 6368 18028 6420 18080
rect 12164 18028 12216 18080
rect 12992 18028 13044 18080
rect 14096 18028 14148 18080
rect 16856 18028 16908 18080
rect 17224 18028 17276 18080
rect 17592 18028 17644 18080
rect 19340 18071 19392 18080
rect 19340 18037 19349 18071
rect 19349 18037 19383 18071
rect 19383 18037 19392 18071
rect 19340 18028 19392 18037
rect 19892 18028 19944 18080
rect 22376 18071 22428 18080
rect 22376 18037 22385 18071
rect 22385 18037 22419 18071
rect 22419 18037 22428 18071
rect 22376 18028 22428 18037
rect 22652 18139 22704 18148
rect 22652 18105 22661 18139
rect 22661 18105 22695 18139
rect 22695 18105 22704 18139
rect 22652 18096 22704 18105
rect 27252 18096 27304 18148
rect 27620 18096 27672 18148
rect 28724 18096 28776 18148
rect 33140 18164 33192 18216
rect 33324 18164 33376 18216
rect 34060 18232 34112 18284
rect 34244 18275 34296 18284
rect 34244 18241 34253 18275
rect 34253 18241 34287 18275
rect 34287 18241 34296 18275
rect 34244 18232 34296 18241
rect 23020 18028 23072 18080
rect 23480 18028 23532 18080
rect 23756 18071 23808 18080
rect 23756 18037 23765 18071
rect 23765 18037 23799 18071
rect 23799 18037 23808 18071
rect 23756 18028 23808 18037
rect 25412 18071 25464 18080
rect 25412 18037 25421 18071
rect 25421 18037 25455 18071
rect 25455 18037 25464 18071
rect 25412 18028 25464 18037
rect 25688 18071 25740 18080
rect 25688 18037 25697 18071
rect 25697 18037 25731 18071
rect 25731 18037 25740 18071
rect 25688 18028 25740 18037
rect 26884 18028 26936 18080
rect 27712 18028 27764 18080
rect 29184 18028 29236 18080
rect 33048 18096 33100 18148
rect 34060 18096 34112 18148
rect 34704 18275 34756 18284
rect 34704 18241 34713 18275
rect 34713 18241 34747 18275
rect 34747 18241 34756 18275
rect 34704 18232 34756 18241
rect 36912 18275 36964 18284
rect 36912 18241 36921 18275
rect 36921 18241 36955 18275
rect 36955 18241 36964 18275
rect 36912 18232 36964 18241
rect 37372 18275 37424 18284
rect 37372 18241 37381 18275
rect 37381 18241 37415 18275
rect 37415 18241 37424 18275
rect 37372 18232 37424 18241
rect 37464 18232 37516 18284
rect 41696 18232 41748 18284
rect 41788 18275 41840 18284
rect 41788 18241 41797 18275
rect 41797 18241 41831 18275
rect 41831 18241 41840 18275
rect 41788 18232 41840 18241
rect 41880 18275 41932 18284
rect 41880 18241 41889 18275
rect 41889 18241 41923 18275
rect 41923 18241 41932 18275
rect 41880 18232 41932 18241
rect 43168 18232 43220 18284
rect 34888 18164 34940 18216
rect 37280 18164 37332 18216
rect 40316 18207 40368 18216
rect 40316 18173 40325 18207
rect 40325 18173 40359 18207
rect 40359 18173 40368 18207
rect 40316 18164 40368 18173
rect 42524 18164 42576 18216
rect 35348 18096 35400 18148
rect 38200 18096 38252 18148
rect 31668 18028 31720 18080
rect 32312 18028 32364 18080
rect 33784 18028 33836 18080
rect 33968 18071 34020 18080
rect 33968 18037 33977 18071
rect 33977 18037 34011 18071
rect 34011 18037 34020 18071
rect 33968 18028 34020 18037
rect 34152 18071 34204 18080
rect 34152 18037 34161 18071
rect 34161 18037 34195 18071
rect 34195 18037 34204 18071
rect 34152 18028 34204 18037
rect 34520 18071 34572 18080
rect 34520 18037 34529 18071
rect 34529 18037 34563 18071
rect 34563 18037 34572 18071
rect 34520 18028 34572 18037
rect 34704 18028 34756 18080
rect 34888 18071 34940 18080
rect 34888 18037 34897 18071
rect 34897 18037 34931 18071
rect 34931 18037 34940 18071
rect 34888 18028 34940 18037
rect 34980 18028 35032 18080
rect 37464 18028 37516 18080
rect 38108 18028 38160 18080
rect 38660 18028 38712 18080
rect 41788 18028 41840 18080
rect 42524 18028 42576 18080
rect 44088 18028 44140 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 2412 17867 2464 17876
rect 2412 17833 2421 17867
rect 2421 17833 2455 17867
rect 2455 17833 2464 17867
rect 2412 17824 2464 17833
rect 2504 17824 2556 17876
rect 2596 17663 2648 17672
rect 2596 17629 2605 17663
rect 2605 17629 2639 17663
rect 2639 17629 2648 17663
rect 2596 17620 2648 17629
rect 3056 17824 3108 17876
rect 4804 17824 4856 17876
rect 6276 17824 6328 17876
rect 6552 17756 6604 17808
rect 6920 17756 6972 17808
rect 7288 17824 7340 17876
rect 7748 17824 7800 17876
rect 8024 17824 8076 17876
rect 8208 17824 8260 17876
rect 9680 17824 9732 17876
rect 9956 17867 10008 17876
rect 9956 17833 9965 17867
rect 9965 17833 9999 17867
rect 9999 17833 10008 17867
rect 9956 17824 10008 17833
rect 10324 17824 10376 17876
rect 10968 17824 11020 17876
rect 11704 17824 11756 17876
rect 12624 17824 12676 17876
rect 13544 17824 13596 17876
rect 15200 17867 15252 17876
rect 15200 17833 15209 17867
rect 15209 17833 15243 17867
rect 15243 17833 15252 17867
rect 15200 17824 15252 17833
rect 16304 17824 16356 17876
rect 22836 17824 22888 17876
rect 8392 17756 8444 17808
rect 13728 17756 13780 17808
rect 17776 17756 17828 17808
rect 23572 17824 23624 17876
rect 24032 17824 24084 17876
rect 24952 17756 25004 17808
rect 25964 17867 26016 17876
rect 25964 17833 25973 17867
rect 25973 17833 26007 17867
rect 26007 17833 26016 17867
rect 25964 17824 26016 17833
rect 26240 17867 26292 17876
rect 26240 17833 26249 17867
rect 26249 17833 26283 17867
rect 26283 17833 26292 17867
rect 26240 17824 26292 17833
rect 26976 17867 27028 17876
rect 26976 17833 26985 17867
rect 26985 17833 27019 17867
rect 27019 17833 27028 17867
rect 26976 17824 27028 17833
rect 27528 17824 27580 17876
rect 2872 17620 2924 17672
rect 3332 17663 3384 17672
rect 3332 17629 3341 17663
rect 3341 17629 3375 17663
rect 3375 17629 3384 17663
rect 3332 17620 3384 17629
rect 4620 17620 4672 17672
rect 4712 17620 4764 17672
rect 4896 17620 4948 17672
rect 6000 17620 6052 17672
rect 6184 17663 6236 17672
rect 6184 17629 6193 17663
rect 6193 17629 6227 17663
rect 6227 17629 6236 17663
rect 6184 17620 6236 17629
rect 6460 17663 6512 17672
rect 3240 17552 3292 17604
rect 5908 17595 5960 17604
rect 5908 17561 5917 17595
rect 5917 17561 5951 17595
rect 5951 17561 5960 17595
rect 6460 17629 6469 17663
rect 6469 17629 6503 17663
rect 6503 17629 6512 17663
rect 6460 17620 6512 17629
rect 6736 17620 6788 17672
rect 7656 17620 7708 17672
rect 8208 17620 8260 17672
rect 5908 17552 5960 17561
rect 6368 17595 6420 17604
rect 6368 17561 6377 17595
rect 6377 17561 6411 17595
rect 6411 17561 6420 17595
rect 6368 17552 6420 17561
rect 7840 17595 7892 17604
rect 7840 17561 7849 17595
rect 7849 17561 7883 17595
rect 7883 17561 7892 17595
rect 7840 17552 7892 17561
rect 8300 17552 8352 17604
rect 7196 17484 7248 17536
rect 7288 17484 7340 17536
rect 9772 17663 9824 17672
rect 9772 17629 9786 17663
rect 9786 17629 9820 17663
rect 9820 17629 9824 17663
rect 9772 17620 9824 17629
rect 9220 17552 9272 17604
rect 9496 17552 9548 17604
rect 11336 17552 11388 17604
rect 11520 17552 11572 17604
rect 9956 17484 10008 17536
rect 11704 17663 11756 17672
rect 11704 17629 11713 17663
rect 11713 17629 11747 17663
rect 11747 17629 11756 17663
rect 11704 17620 11756 17629
rect 11980 17663 12032 17672
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 11888 17595 11940 17604
rect 11888 17561 11897 17595
rect 11897 17561 11931 17595
rect 11931 17561 11940 17595
rect 11888 17552 11940 17561
rect 12164 17484 12216 17536
rect 12900 17688 12952 17740
rect 17040 17688 17092 17740
rect 12992 17620 13044 17672
rect 13360 17552 13412 17604
rect 14924 17595 14976 17604
rect 14924 17561 14933 17595
rect 14933 17561 14967 17595
rect 14967 17561 14976 17595
rect 14924 17552 14976 17561
rect 15108 17595 15160 17604
rect 15108 17561 15117 17595
rect 15117 17561 15151 17595
rect 15151 17561 15160 17595
rect 15108 17552 15160 17561
rect 15292 17620 15344 17672
rect 16120 17620 16172 17672
rect 16580 17620 16632 17672
rect 16856 17620 16908 17672
rect 19616 17663 19668 17672
rect 19616 17629 19625 17663
rect 19625 17629 19659 17663
rect 19659 17629 19668 17663
rect 19616 17620 19668 17629
rect 19800 17731 19852 17740
rect 19800 17697 19809 17731
rect 19809 17697 19843 17731
rect 19843 17697 19852 17731
rect 19800 17688 19852 17697
rect 23020 17731 23072 17740
rect 23020 17697 23029 17731
rect 23029 17697 23063 17731
rect 23063 17697 23072 17731
rect 23020 17688 23072 17697
rect 20260 17620 20312 17672
rect 22192 17620 22244 17672
rect 22376 17620 22428 17672
rect 22560 17620 22612 17672
rect 26148 17688 26200 17740
rect 23204 17663 23256 17672
rect 23204 17629 23213 17663
rect 23213 17629 23247 17663
rect 23247 17629 23256 17663
rect 23204 17620 23256 17629
rect 25228 17620 25280 17672
rect 25688 17620 25740 17672
rect 26332 17620 26384 17672
rect 27252 17756 27304 17808
rect 27620 17688 27672 17740
rect 28172 17824 28224 17876
rect 29736 17824 29788 17876
rect 29828 17867 29880 17876
rect 29828 17833 29837 17867
rect 29837 17833 29871 17867
rect 29871 17833 29880 17867
rect 29828 17824 29880 17833
rect 31392 17867 31444 17876
rect 31392 17833 31401 17867
rect 31401 17833 31435 17867
rect 31435 17833 31444 17867
rect 31392 17824 31444 17833
rect 32312 17824 32364 17876
rect 32956 17824 33008 17876
rect 27988 17756 28040 17808
rect 33416 17824 33468 17876
rect 33876 17867 33928 17876
rect 33876 17833 33885 17867
rect 33885 17833 33919 17867
rect 33919 17833 33928 17867
rect 33876 17824 33928 17833
rect 34060 17867 34112 17876
rect 34060 17833 34069 17867
rect 34069 17833 34103 17867
rect 34103 17833 34112 17867
rect 34060 17824 34112 17833
rect 34244 17824 34296 17876
rect 36268 17824 36320 17876
rect 37188 17824 37240 17876
rect 38752 17824 38804 17876
rect 28172 17688 28224 17740
rect 28632 17688 28684 17740
rect 31208 17731 31260 17740
rect 31208 17697 31217 17731
rect 31217 17697 31251 17731
rect 31251 17697 31260 17731
rect 31208 17688 31260 17697
rect 31760 17731 31812 17740
rect 31760 17697 31769 17731
rect 31769 17697 31803 17731
rect 31803 17697 31812 17731
rect 31760 17688 31812 17697
rect 32404 17731 32456 17740
rect 32404 17697 32413 17731
rect 32413 17697 32447 17731
rect 32447 17697 32456 17731
rect 32404 17688 32456 17697
rect 19340 17552 19392 17604
rect 23020 17552 23072 17604
rect 13176 17484 13228 17536
rect 14464 17484 14516 17536
rect 17132 17484 17184 17536
rect 17776 17484 17828 17536
rect 17868 17484 17920 17536
rect 22100 17484 22152 17536
rect 22192 17484 22244 17536
rect 24584 17484 24636 17536
rect 26792 17552 26844 17604
rect 27528 17620 27580 17672
rect 27988 17663 28040 17672
rect 27988 17629 27997 17663
rect 27997 17629 28031 17663
rect 28031 17629 28040 17663
rect 27988 17620 28040 17629
rect 28080 17620 28132 17672
rect 29368 17620 29420 17672
rect 29736 17663 29788 17672
rect 29736 17629 29745 17663
rect 29745 17629 29779 17663
rect 29779 17629 29788 17663
rect 29736 17620 29788 17629
rect 30288 17620 30340 17672
rect 31116 17663 31168 17672
rect 31116 17629 31125 17663
rect 31125 17629 31159 17663
rect 31159 17629 31168 17663
rect 31116 17620 31168 17629
rect 31392 17663 31444 17672
rect 31392 17629 31401 17663
rect 31401 17629 31435 17663
rect 31435 17629 31444 17663
rect 31392 17620 31444 17629
rect 31944 17663 31996 17672
rect 31944 17629 31953 17663
rect 31953 17629 31987 17663
rect 31987 17629 31996 17663
rect 31944 17620 31996 17629
rect 32588 17620 32640 17672
rect 26424 17484 26476 17536
rect 26700 17527 26752 17536
rect 26700 17493 26709 17527
rect 26709 17493 26743 17527
rect 26743 17493 26752 17527
rect 26700 17484 26752 17493
rect 27252 17484 27304 17536
rect 29552 17595 29604 17604
rect 29552 17561 29567 17595
rect 29567 17561 29601 17595
rect 29601 17561 29604 17595
rect 29552 17552 29604 17561
rect 31668 17595 31720 17604
rect 31668 17561 31677 17595
rect 31677 17561 31711 17595
rect 31711 17561 31720 17595
rect 31668 17552 31720 17561
rect 28448 17484 28500 17536
rect 28816 17484 28868 17536
rect 31024 17484 31076 17536
rect 36544 17756 36596 17808
rect 33140 17731 33192 17740
rect 33140 17697 33149 17731
rect 33149 17697 33183 17731
rect 33183 17697 33192 17731
rect 33140 17688 33192 17697
rect 33232 17663 33284 17672
rect 33232 17629 33241 17663
rect 33241 17629 33275 17663
rect 33275 17629 33284 17663
rect 33232 17620 33284 17629
rect 35164 17688 35216 17740
rect 33784 17620 33836 17672
rect 33968 17663 34020 17672
rect 33968 17629 33977 17663
rect 33977 17629 34011 17663
rect 34011 17629 34020 17663
rect 33968 17620 34020 17629
rect 32128 17527 32180 17536
rect 32128 17493 32137 17527
rect 32137 17493 32171 17527
rect 32171 17493 32180 17527
rect 32128 17484 32180 17493
rect 33600 17552 33652 17604
rect 33876 17552 33928 17604
rect 34428 17620 34480 17672
rect 36728 17688 36780 17740
rect 37832 17756 37884 17808
rect 38476 17756 38528 17808
rect 40040 17824 40092 17876
rect 43260 17824 43312 17876
rect 41696 17756 41748 17808
rect 42708 17756 42760 17808
rect 38936 17688 38988 17740
rect 35348 17663 35400 17672
rect 35348 17629 35357 17663
rect 35357 17629 35391 17663
rect 35391 17629 35400 17663
rect 35348 17620 35400 17629
rect 36452 17663 36504 17672
rect 36452 17629 36461 17663
rect 36461 17629 36495 17663
rect 36495 17629 36504 17663
rect 36452 17620 36504 17629
rect 34152 17484 34204 17536
rect 35072 17595 35124 17604
rect 35072 17561 35081 17595
rect 35081 17561 35115 17595
rect 35115 17561 35124 17595
rect 35072 17552 35124 17561
rect 35164 17552 35216 17604
rect 35348 17484 35400 17536
rect 36084 17552 36136 17604
rect 37556 17663 37608 17672
rect 37556 17629 37565 17663
rect 37565 17629 37599 17663
rect 37599 17629 37608 17663
rect 37556 17620 37608 17629
rect 38200 17663 38252 17672
rect 38200 17629 38209 17663
rect 38209 17629 38243 17663
rect 38243 17629 38252 17663
rect 38200 17620 38252 17629
rect 38844 17663 38896 17672
rect 38844 17629 38853 17663
rect 38853 17629 38887 17663
rect 38887 17629 38896 17663
rect 38844 17620 38896 17629
rect 39856 17663 39908 17672
rect 39856 17629 39865 17663
rect 39865 17629 39899 17663
rect 39899 17629 39908 17663
rect 39856 17620 39908 17629
rect 40132 17663 40184 17672
rect 40132 17629 40166 17663
rect 40166 17629 40184 17663
rect 40132 17620 40184 17629
rect 41328 17620 41380 17672
rect 38752 17552 38804 17604
rect 39028 17595 39080 17604
rect 39028 17561 39037 17595
rect 39037 17561 39071 17595
rect 39071 17561 39080 17595
rect 39028 17552 39080 17561
rect 39580 17552 39632 17604
rect 41788 17663 41840 17672
rect 41788 17629 41797 17663
rect 41797 17629 41831 17663
rect 41831 17629 41840 17663
rect 41788 17620 41840 17629
rect 37004 17484 37056 17536
rect 42524 17620 42576 17672
rect 43812 17620 43864 17672
rect 42708 17484 42760 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 3792 17323 3844 17332
rect 3792 17289 3801 17323
rect 3801 17289 3835 17323
rect 3835 17289 3844 17323
rect 3792 17280 3844 17289
rect 3976 17280 4028 17332
rect 5172 17280 5224 17332
rect 5448 17280 5500 17332
rect 8576 17280 8628 17332
rect 9036 17280 9088 17332
rect 9312 17323 9364 17332
rect 9312 17289 9321 17323
rect 9321 17289 9355 17323
rect 9355 17289 9364 17323
rect 9312 17280 9364 17289
rect 4712 17212 4764 17264
rect 4988 17212 5040 17264
rect 7840 17212 7892 17264
rect 8208 17212 8260 17264
rect 11704 17323 11756 17332
rect 11704 17289 11713 17323
rect 11713 17289 11747 17323
rect 11747 17289 11756 17323
rect 11704 17280 11756 17289
rect 2228 17187 2280 17196
rect 2228 17153 2237 17187
rect 2237 17153 2271 17187
rect 2271 17153 2280 17187
rect 2228 17144 2280 17153
rect 3608 17187 3660 17196
rect 3608 17153 3617 17187
rect 3617 17153 3651 17187
rect 3651 17153 3660 17187
rect 3608 17144 3660 17153
rect 5448 17144 5500 17196
rect 6828 17144 6880 17196
rect 4712 17076 4764 17128
rect 5080 17076 5132 17128
rect 7932 17144 7984 17196
rect 8760 17187 8812 17196
rect 8760 17153 8769 17187
rect 8769 17153 8803 17187
rect 8803 17153 8812 17187
rect 8760 17144 8812 17153
rect 9128 17187 9180 17196
rect 9128 17153 9137 17187
rect 9137 17153 9171 17187
rect 9171 17153 9180 17187
rect 9128 17144 9180 17153
rect 9496 17187 9548 17196
rect 9496 17153 9505 17187
rect 9505 17153 9539 17187
rect 9539 17153 9548 17187
rect 9496 17144 9548 17153
rect 7564 17076 7616 17128
rect 7748 17076 7800 17128
rect 9772 17187 9824 17196
rect 9772 17153 9781 17187
rect 9781 17153 9815 17187
rect 9815 17153 9824 17187
rect 9772 17144 9824 17153
rect 9864 17187 9916 17196
rect 9864 17153 9878 17187
rect 9878 17153 9912 17187
rect 9912 17153 9916 17187
rect 9864 17144 9916 17153
rect 10140 17144 10192 17196
rect 10508 17144 10560 17196
rect 10692 17144 10744 17196
rect 11428 17144 11480 17196
rect 12624 17212 12676 17264
rect 10232 17076 10284 17128
rect 11060 17076 11112 17128
rect 11888 17076 11940 17128
rect 3700 17008 3752 17060
rect 5540 17008 5592 17060
rect 6276 17008 6328 17060
rect 8300 17008 8352 17060
rect 10968 17008 11020 17060
rect 2320 16983 2372 16992
rect 2320 16949 2329 16983
rect 2329 16949 2363 16983
rect 2363 16949 2372 16983
rect 2320 16940 2372 16949
rect 3884 16940 3936 16992
rect 4896 16940 4948 16992
rect 5356 16940 5408 16992
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 13176 17187 13228 17196
rect 13176 17153 13185 17187
rect 13185 17153 13219 17187
rect 13219 17153 13228 17187
rect 13176 17144 13228 17153
rect 13268 17187 13320 17196
rect 13268 17153 13277 17187
rect 13277 17153 13311 17187
rect 13311 17153 13320 17187
rect 13268 17144 13320 17153
rect 14464 17212 14516 17264
rect 13728 17187 13780 17196
rect 13728 17153 13737 17187
rect 13737 17153 13771 17187
rect 13771 17153 13780 17187
rect 13728 17144 13780 17153
rect 13912 17187 13964 17196
rect 13912 17153 13921 17187
rect 13921 17153 13955 17187
rect 13955 17153 13964 17187
rect 13912 17144 13964 17153
rect 14096 17187 14148 17196
rect 14096 17153 14110 17187
rect 14110 17153 14144 17187
rect 14144 17153 14148 17187
rect 14096 17144 14148 17153
rect 13544 17051 13596 17060
rect 13544 17017 13553 17051
rect 13553 17017 13587 17051
rect 13587 17017 13596 17051
rect 13544 17008 13596 17017
rect 14188 17008 14240 17060
rect 19616 17280 19668 17332
rect 22100 17280 22152 17332
rect 23112 17280 23164 17332
rect 16856 17212 16908 17264
rect 23204 17255 23256 17264
rect 23204 17221 23213 17255
rect 23213 17221 23247 17255
rect 23247 17221 23256 17255
rect 23204 17212 23256 17221
rect 24400 17280 24452 17332
rect 24768 17280 24820 17332
rect 26792 17280 26844 17332
rect 27160 17280 27212 17332
rect 31668 17280 31720 17332
rect 31944 17280 31996 17332
rect 34060 17280 34112 17332
rect 26240 17212 26292 17264
rect 15016 17187 15068 17196
rect 15016 17153 15025 17187
rect 15025 17153 15059 17187
rect 15059 17153 15068 17187
rect 15016 17144 15068 17153
rect 17776 17144 17828 17196
rect 18696 17187 18748 17196
rect 18696 17153 18705 17187
rect 18705 17153 18739 17187
rect 18739 17153 18748 17187
rect 18696 17144 18748 17153
rect 18788 17187 18840 17196
rect 18788 17153 18797 17187
rect 18797 17153 18831 17187
rect 18831 17153 18840 17187
rect 18788 17144 18840 17153
rect 15844 17076 15896 17128
rect 17960 17076 18012 17128
rect 19156 17144 19208 17196
rect 20260 17144 20312 17196
rect 22744 17144 22796 17196
rect 24768 17187 24820 17196
rect 24768 17153 24777 17187
rect 24777 17153 24811 17187
rect 24811 17153 24820 17187
rect 24768 17144 24820 17153
rect 26332 17144 26384 17196
rect 19064 17076 19116 17128
rect 24308 17076 24360 17128
rect 24860 17119 24912 17128
rect 24860 17085 24869 17119
rect 24869 17085 24903 17119
rect 24903 17085 24912 17119
rect 24860 17076 24912 17085
rect 24032 17008 24084 17060
rect 12900 16940 12952 16992
rect 14096 16940 14148 16992
rect 14372 16940 14424 16992
rect 18788 16940 18840 16992
rect 19156 16940 19208 16992
rect 19340 16983 19392 16992
rect 19340 16949 19349 16983
rect 19349 16949 19383 16983
rect 19383 16949 19392 16983
rect 19340 16940 19392 16949
rect 19432 16940 19484 16992
rect 19800 16940 19852 16992
rect 24584 16940 24636 16992
rect 25320 17076 25372 17128
rect 26700 17212 26752 17264
rect 26516 17144 26568 17196
rect 27712 17255 27764 17264
rect 27712 17221 27721 17255
rect 27721 17221 27755 17255
rect 27755 17221 27764 17255
rect 27712 17212 27764 17221
rect 28080 17144 28132 17196
rect 27160 17076 27212 17128
rect 29644 17144 29696 17196
rect 32128 17255 32180 17264
rect 32128 17221 32137 17255
rect 32137 17221 32171 17255
rect 32171 17221 32180 17255
rect 32128 17212 32180 17221
rect 32312 17255 32364 17264
rect 32312 17221 32321 17255
rect 32321 17221 32355 17255
rect 32355 17221 32364 17255
rect 32312 17212 32364 17221
rect 36084 17323 36136 17332
rect 36084 17289 36093 17323
rect 36093 17289 36127 17323
rect 36127 17289 36136 17323
rect 36084 17280 36136 17289
rect 37280 17280 37332 17332
rect 35716 17212 35768 17264
rect 36360 17255 36412 17264
rect 36360 17221 36369 17255
rect 36369 17221 36403 17255
rect 36403 17221 36412 17255
rect 36360 17212 36412 17221
rect 36912 17212 36964 17264
rect 38476 17280 38528 17332
rect 31392 17144 31444 17196
rect 29552 17119 29604 17128
rect 29552 17085 29561 17119
rect 29561 17085 29595 17119
rect 29595 17085 29604 17119
rect 29552 17076 29604 17085
rect 30288 17076 30340 17128
rect 25044 16940 25096 16992
rect 26884 16940 26936 16992
rect 27160 16983 27212 16992
rect 27160 16949 27169 16983
rect 27169 16949 27203 16983
rect 27203 16949 27212 16983
rect 27160 16940 27212 16949
rect 27988 16940 28040 16992
rect 30196 17008 30248 17060
rect 31484 17008 31536 17060
rect 35532 17144 35584 17196
rect 35900 17187 35952 17196
rect 35900 17153 35909 17187
rect 35909 17153 35943 17187
rect 35943 17153 35952 17187
rect 35900 17144 35952 17153
rect 36636 17187 36688 17196
rect 36636 17153 36645 17187
rect 36645 17153 36679 17187
rect 36679 17153 36688 17187
rect 36636 17144 36688 17153
rect 37648 17187 37700 17196
rect 37648 17153 37657 17187
rect 37657 17153 37691 17187
rect 37691 17153 37700 17187
rect 37648 17144 37700 17153
rect 38384 17187 38436 17196
rect 38384 17153 38393 17187
rect 38393 17153 38427 17187
rect 38427 17153 38436 17187
rect 38384 17144 38436 17153
rect 38660 17144 38712 17196
rect 40224 17280 40276 17332
rect 40316 17280 40368 17332
rect 41236 17280 41288 17332
rect 41788 17280 41840 17332
rect 43812 17323 43864 17332
rect 43812 17289 43821 17323
rect 43821 17289 43855 17323
rect 43855 17289 43864 17323
rect 43812 17280 43864 17289
rect 38844 17212 38896 17264
rect 38936 17144 38988 17196
rect 39856 17212 39908 17264
rect 35440 17076 35492 17128
rect 35716 17119 35768 17128
rect 35716 17085 35725 17119
rect 35725 17085 35759 17119
rect 35759 17085 35768 17119
rect 35716 17076 35768 17085
rect 36452 17119 36504 17128
rect 36452 17085 36461 17119
rect 36461 17085 36495 17119
rect 36495 17085 36504 17119
rect 36452 17076 36504 17085
rect 36544 17076 36596 17128
rect 42432 17187 42484 17196
rect 42432 17153 42441 17187
rect 42441 17153 42475 17187
rect 42475 17153 42484 17187
rect 42432 17144 42484 17153
rect 42708 17187 42760 17196
rect 42708 17153 42742 17187
rect 42742 17153 42760 17187
rect 42708 17144 42760 17153
rect 36728 17008 36780 17060
rect 37740 17008 37792 17060
rect 29368 16940 29420 16992
rect 29460 16983 29512 16992
rect 29460 16949 29469 16983
rect 29469 16949 29503 16983
rect 29503 16949 29512 16983
rect 29460 16940 29512 16949
rect 29736 16940 29788 16992
rect 31668 16983 31720 16992
rect 31668 16949 31677 16983
rect 31677 16949 31711 16983
rect 31711 16949 31720 16983
rect 31668 16940 31720 16949
rect 33140 16940 33192 16992
rect 35716 16940 35768 16992
rect 37188 16940 37240 16992
rect 37648 16940 37700 16992
rect 38292 16940 38344 16992
rect 38476 16940 38528 16992
rect 44456 17051 44508 17060
rect 44456 17017 44465 17051
rect 44465 17017 44499 17051
rect 44499 17017 44508 17051
rect 44456 17008 44508 17017
rect 41236 16940 41288 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3240 16736 3292 16788
rect 3700 16736 3752 16788
rect 4620 16736 4672 16788
rect 2136 16668 2188 16720
rect 3976 16668 4028 16720
rect 2320 16643 2372 16652
rect 2320 16609 2329 16643
rect 2329 16609 2363 16643
rect 2363 16609 2372 16643
rect 4160 16668 4212 16720
rect 5080 16668 5132 16720
rect 5264 16668 5316 16720
rect 5448 16668 5500 16720
rect 2320 16600 2372 16609
rect 848 16532 900 16584
rect 6000 16668 6052 16720
rect 6184 16668 6236 16720
rect 7472 16668 7524 16720
rect 8300 16668 8352 16720
rect 8576 16668 8628 16720
rect 8760 16779 8812 16788
rect 8760 16745 8769 16779
rect 8769 16745 8803 16779
rect 8803 16745 8812 16779
rect 8760 16736 8812 16745
rect 10140 16736 10192 16788
rect 19800 16736 19852 16788
rect 21088 16779 21140 16788
rect 21088 16745 21097 16779
rect 21097 16745 21131 16779
rect 21131 16745 21140 16779
rect 21088 16736 21140 16745
rect 22284 16736 22336 16788
rect 22560 16736 22612 16788
rect 23112 16736 23164 16788
rect 24308 16736 24360 16788
rect 3516 16532 3568 16584
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 1768 16507 1820 16516
rect 1768 16473 1777 16507
rect 1777 16473 1811 16507
rect 1811 16473 1820 16507
rect 1768 16464 1820 16473
rect 2964 16464 3016 16516
rect 3056 16464 3108 16516
rect 4988 16532 5040 16584
rect 5356 16532 5408 16584
rect 5540 16532 5592 16584
rect 5908 16532 5960 16584
rect 6460 16575 6512 16584
rect 6460 16541 6469 16575
rect 6469 16541 6503 16575
rect 6503 16541 6512 16575
rect 6460 16532 6512 16541
rect 7380 16532 7432 16584
rect 7472 16532 7524 16584
rect 7840 16532 7892 16584
rect 8944 16532 8996 16584
rect 9864 16668 9916 16720
rect 9312 16600 9364 16652
rect 10600 16643 10652 16652
rect 10600 16609 10609 16643
rect 10609 16609 10643 16643
rect 10643 16609 10652 16643
rect 10600 16600 10652 16609
rect 10968 16643 11020 16652
rect 10968 16609 10977 16643
rect 10977 16609 11011 16643
rect 11011 16609 11020 16643
rect 10968 16600 11020 16609
rect 11612 16668 11664 16720
rect 11704 16668 11756 16720
rect 17040 16668 17092 16720
rect 17408 16711 17460 16720
rect 17408 16677 17417 16711
rect 17417 16677 17451 16711
rect 17451 16677 17460 16711
rect 17408 16668 17460 16677
rect 17868 16711 17920 16720
rect 17868 16677 17877 16711
rect 17877 16677 17911 16711
rect 17911 16677 17920 16711
rect 17868 16668 17920 16677
rect 25504 16779 25556 16788
rect 25504 16745 25513 16779
rect 25513 16745 25547 16779
rect 25547 16745 25556 16779
rect 25504 16736 25556 16745
rect 26792 16736 26844 16788
rect 28172 16736 28224 16788
rect 28448 16779 28500 16788
rect 28448 16745 28457 16779
rect 28457 16745 28491 16779
rect 28491 16745 28500 16779
rect 28448 16736 28500 16745
rect 31668 16779 31720 16788
rect 25136 16668 25188 16720
rect 25872 16711 25924 16720
rect 25872 16677 25881 16711
rect 25881 16677 25915 16711
rect 25915 16677 25924 16711
rect 25872 16668 25924 16677
rect 26884 16668 26936 16720
rect 27344 16668 27396 16720
rect 31668 16745 31677 16779
rect 31677 16745 31711 16779
rect 31711 16745 31720 16779
rect 31668 16736 31720 16745
rect 31944 16736 31996 16788
rect 32496 16779 32548 16788
rect 32496 16745 32505 16779
rect 32505 16745 32539 16779
rect 32539 16745 32548 16779
rect 32496 16736 32548 16745
rect 33416 16736 33468 16788
rect 34060 16736 34112 16788
rect 35900 16736 35952 16788
rect 37188 16736 37240 16788
rect 37464 16736 37516 16788
rect 3240 16396 3292 16448
rect 3516 16396 3568 16448
rect 4068 16396 4120 16448
rect 5540 16396 5592 16448
rect 5908 16396 5960 16448
rect 7564 16464 7616 16516
rect 7748 16464 7800 16516
rect 9036 16464 9088 16516
rect 10140 16532 10192 16584
rect 11244 16575 11296 16584
rect 11244 16541 11253 16575
rect 11253 16541 11287 16575
rect 11287 16541 11296 16575
rect 11244 16532 11296 16541
rect 12716 16600 12768 16652
rect 10600 16464 10652 16516
rect 11428 16507 11480 16516
rect 11428 16473 11437 16507
rect 11437 16473 11471 16507
rect 11471 16473 11480 16507
rect 11428 16464 11480 16473
rect 15292 16600 15344 16652
rect 15844 16600 15896 16652
rect 12992 16464 13044 16516
rect 16120 16575 16172 16584
rect 16120 16541 16129 16575
rect 16129 16541 16163 16575
rect 16163 16541 16172 16575
rect 16120 16532 16172 16541
rect 19524 16600 19576 16652
rect 22284 16600 22336 16652
rect 15936 16507 15988 16516
rect 15936 16473 15945 16507
rect 15945 16473 15979 16507
rect 15979 16473 15988 16507
rect 15936 16464 15988 16473
rect 16028 16507 16080 16516
rect 16028 16473 16037 16507
rect 16037 16473 16071 16507
rect 16071 16473 16080 16507
rect 16028 16464 16080 16473
rect 6460 16396 6512 16448
rect 7380 16439 7432 16448
rect 7380 16405 7389 16439
rect 7389 16405 7423 16439
rect 7423 16405 7432 16439
rect 7380 16396 7432 16405
rect 8208 16396 8260 16448
rect 9496 16396 9548 16448
rect 10968 16396 11020 16448
rect 11152 16396 11204 16448
rect 15108 16396 15160 16448
rect 17224 16507 17276 16516
rect 17224 16473 17233 16507
rect 17233 16473 17267 16507
rect 17267 16473 17276 16507
rect 17224 16464 17276 16473
rect 17592 16464 17644 16516
rect 20536 16464 20588 16516
rect 21180 16575 21232 16584
rect 21180 16541 21189 16575
rect 21189 16541 21223 16575
rect 21223 16541 21232 16575
rect 21180 16532 21232 16541
rect 22192 16532 22244 16584
rect 22652 16575 22704 16584
rect 22652 16541 22661 16575
rect 22661 16541 22695 16575
rect 22695 16541 22704 16575
rect 22652 16532 22704 16541
rect 24308 16600 24360 16652
rect 25044 16643 25096 16652
rect 25044 16609 25053 16643
rect 25053 16609 25087 16643
rect 25087 16609 25096 16643
rect 25044 16600 25096 16609
rect 25412 16600 25464 16652
rect 26332 16643 26384 16652
rect 26332 16609 26341 16643
rect 26341 16609 26375 16643
rect 26375 16609 26384 16643
rect 29368 16668 29420 16720
rect 31392 16668 31444 16720
rect 32036 16711 32088 16720
rect 32036 16677 32045 16711
rect 32045 16677 32079 16711
rect 32079 16677 32088 16711
rect 32036 16668 32088 16677
rect 26332 16600 26384 16609
rect 28540 16643 28592 16652
rect 28540 16609 28549 16643
rect 28549 16609 28583 16643
rect 28583 16609 28592 16643
rect 28540 16600 28592 16609
rect 30840 16600 30892 16652
rect 25136 16575 25188 16584
rect 25136 16541 25145 16575
rect 25145 16541 25179 16575
rect 25179 16541 25188 16575
rect 25136 16532 25188 16541
rect 25780 16532 25832 16584
rect 29000 16532 29052 16584
rect 22284 16464 22336 16516
rect 24124 16464 24176 16516
rect 24952 16464 25004 16516
rect 25964 16507 26016 16516
rect 25964 16473 25973 16507
rect 25973 16473 26007 16507
rect 26007 16473 26016 16507
rect 25964 16464 26016 16473
rect 26148 16507 26200 16516
rect 26148 16473 26157 16507
rect 26157 16473 26191 16507
rect 26191 16473 26200 16507
rect 26148 16464 26200 16473
rect 26884 16464 26936 16516
rect 28264 16464 28316 16516
rect 31300 16532 31352 16584
rect 31760 16643 31812 16652
rect 31760 16609 31769 16643
rect 31769 16609 31803 16643
rect 31803 16609 31812 16643
rect 32404 16668 32456 16720
rect 38476 16736 38528 16788
rect 38384 16711 38436 16720
rect 38384 16677 38393 16711
rect 38393 16677 38427 16711
rect 38427 16677 38436 16711
rect 38384 16668 38436 16677
rect 39304 16668 39356 16720
rect 31760 16600 31812 16609
rect 32312 16600 32364 16652
rect 37740 16643 37792 16652
rect 37740 16609 37749 16643
rect 37749 16609 37783 16643
rect 37783 16609 37792 16643
rect 37740 16600 37792 16609
rect 38752 16600 38804 16652
rect 32036 16532 32088 16584
rect 33232 16532 33284 16584
rect 33416 16532 33468 16584
rect 40224 16532 40276 16584
rect 40316 16532 40368 16584
rect 22192 16396 22244 16448
rect 22744 16396 22796 16448
rect 29368 16464 29420 16516
rect 29920 16464 29972 16516
rect 28908 16439 28960 16448
rect 28908 16405 28917 16439
rect 28917 16405 28951 16439
rect 28951 16405 28960 16439
rect 28908 16396 28960 16405
rect 29184 16396 29236 16448
rect 36820 16464 36872 16516
rect 37832 16464 37884 16516
rect 38568 16464 38620 16516
rect 42432 16464 42484 16516
rect 35992 16396 36044 16448
rect 36912 16396 36964 16448
rect 37372 16439 37424 16448
rect 37372 16405 37381 16439
rect 37381 16405 37415 16439
rect 37415 16405 37424 16439
rect 37372 16396 37424 16405
rect 44456 16439 44508 16448
rect 44456 16405 44465 16439
rect 44465 16405 44499 16439
rect 44499 16405 44508 16439
rect 44456 16396 44508 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 2228 16192 2280 16244
rect 848 16056 900 16108
rect 1768 16056 1820 16108
rect 2964 16124 3016 16176
rect 2320 16056 2372 16108
rect 2780 16099 2832 16108
rect 2780 16065 2789 16099
rect 2789 16065 2823 16099
rect 2823 16065 2832 16099
rect 2780 16056 2832 16065
rect 2228 16031 2280 16040
rect 2228 15997 2237 16031
rect 2237 15997 2271 16031
rect 2271 15997 2280 16031
rect 2228 15988 2280 15997
rect 3424 15988 3476 16040
rect 3056 15852 3108 15904
rect 3424 15852 3476 15904
rect 3884 16099 3936 16108
rect 3884 16065 3893 16099
rect 3893 16065 3927 16099
rect 3927 16065 3936 16099
rect 5264 16124 5316 16176
rect 3884 16056 3936 16065
rect 4620 16099 4672 16108
rect 4620 16065 4629 16099
rect 4629 16065 4663 16099
rect 4663 16065 4672 16099
rect 4620 16056 4672 16065
rect 6368 16192 6420 16244
rect 6644 16235 6696 16244
rect 6644 16201 6653 16235
rect 6653 16201 6687 16235
rect 6687 16201 6696 16235
rect 6644 16192 6696 16201
rect 6920 16192 6972 16244
rect 6000 16124 6052 16176
rect 6736 16124 6788 16176
rect 9128 16192 9180 16244
rect 9496 16192 9548 16244
rect 3700 15988 3752 16040
rect 3792 15988 3844 16040
rect 5816 16099 5868 16108
rect 5816 16065 5825 16099
rect 5825 16065 5859 16099
rect 5859 16065 5868 16099
rect 5816 16056 5868 16065
rect 6368 16056 6420 16108
rect 6920 16031 6972 16040
rect 6920 15997 6929 16031
rect 6929 15997 6963 16031
rect 6963 15997 6972 16031
rect 6920 15988 6972 15997
rect 7288 16056 7340 16108
rect 7840 16056 7892 16108
rect 8852 16124 8904 16176
rect 7288 15920 7340 15972
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 6368 15852 6420 15904
rect 8024 15988 8076 16040
rect 8208 16031 8260 16040
rect 8208 15997 8217 16031
rect 8217 15997 8251 16031
rect 8251 15997 8260 16031
rect 8208 15988 8260 15997
rect 7748 15920 7800 15972
rect 8392 16031 8444 16040
rect 8392 15997 8426 16031
rect 8426 15997 8444 16031
rect 8760 16099 8812 16108
rect 8760 16065 8769 16099
rect 8769 16065 8803 16099
rect 8803 16065 8812 16099
rect 8760 16056 8812 16065
rect 9036 16056 9088 16108
rect 8392 15988 8444 15997
rect 9128 15988 9180 16040
rect 9404 16124 9456 16176
rect 10508 16167 10560 16176
rect 10508 16133 10517 16167
rect 10517 16133 10551 16167
rect 10551 16133 10560 16167
rect 10508 16124 10560 16133
rect 9036 15920 9088 15972
rect 9404 15920 9456 15972
rect 10324 16099 10376 16108
rect 10324 16065 10333 16099
rect 10333 16065 10367 16099
rect 10367 16065 10376 16099
rect 10324 16056 10376 16065
rect 10600 16099 10652 16108
rect 10600 16065 10609 16099
rect 10609 16065 10643 16099
rect 10643 16065 10652 16099
rect 10600 16056 10652 16065
rect 10784 16192 10836 16244
rect 11152 16192 11204 16244
rect 11428 16192 11480 16244
rect 11612 16192 11664 16244
rect 11060 16124 11112 16176
rect 12164 16124 12216 16176
rect 15384 16192 15436 16244
rect 15844 16192 15896 16244
rect 16764 16192 16816 16244
rect 17776 16192 17828 16244
rect 20076 16192 20128 16244
rect 20536 16235 20588 16244
rect 20536 16201 20545 16235
rect 20545 16201 20579 16235
rect 20579 16201 20588 16235
rect 20536 16192 20588 16201
rect 22008 16192 22060 16244
rect 22744 16192 22796 16244
rect 15200 16167 15252 16176
rect 15200 16133 15209 16167
rect 15209 16133 15243 16167
rect 15243 16133 15252 16167
rect 15200 16124 15252 16133
rect 11612 16099 11664 16108
rect 11612 16065 11621 16099
rect 11621 16065 11655 16099
rect 11655 16065 11664 16099
rect 11612 16056 11664 16065
rect 11888 16099 11940 16108
rect 11888 16065 11897 16099
rect 11897 16065 11931 16099
rect 11931 16065 11940 16099
rect 11888 16056 11940 16065
rect 12072 16099 12124 16108
rect 12072 16065 12075 16099
rect 12075 16065 12124 16099
rect 12072 16056 12124 16065
rect 12348 16099 12400 16108
rect 12348 16065 12357 16099
rect 12357 16065 12391 16099
rect 12391 16065 12400 16099
rect 12348 16056 12400 16065
rect 12624 16056 12676 16108
rect 12992 16099 13044 16108
rect 12992 16065 13001 16099
rect 13001 16065 13035 16099
rect 13035 16065 13044 16099
rect 12992 16056 13044 16065
rect 10784 15988 10836 16040
rect 15108 15988 15160 16040
rect 9220 15852 9272 15904
rect 10232 15920 10284 15972
rect 11336 15920 11388 15972
rect 12992 15920 13044 15972
rect 17592 16124 17644 16176
rect 15844 16099 15896 16108
rect 15844 16065 15853 16099
rect 15853 16065 15887 16099
rect 15887 16065 15896 16099
rect 15844 16056 15896 16065
rect 15936 16099 15988 16108
rect 15936 16065 15945 16099
rect 15945 16065 15979 16099
rect 15979 16065 15988 16099
rect 15936 16056 15988 16065
rect 16396 16056 16448 16108
rect 16672 16056 16724 16108
rect 16948 15988 17000 16040
rect 17316 16099 17368 16108
rect 17316 16065 17325 16099
rect 17325 16065 17359 16099
rect 17359 16065 17368 16099
rect 17316 16056 17368 16065
rect 22284 16124 22336 16176
rect 22468 16124 22520 16176
rect 18880 16099 18932 16108
rect 18880 16065 18889 16099
rect 18889 16065 18923 16099
rect 18923 16065 18932 16099
rect 18880 16056 18932 16065
rect 20076 16099 20128 16108
rect 20076 16065 20085 16099
rect 20085 16065 20119 16099
rect 20119 16065 20128 16099
rect 20076 16056 20128 16065
rect 20352 16099 20404 16108
rect 20352 16065 20361 16099
rect 20361 16065 20395 16099
rect 20395 16065 20404 16099
rect 20352 16056 20404 16065
rect 22376 16099 22428 16108
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 22652 16099 22704 16108
rect 22652 16065 22661 16099
rect 22661 16065 22695 16099
rect 22695 16065 22704 16099
rect 22652 16056 22704 16065
rect 18604 15988 18656 16040
rect 9956 15895 10008 15904
rect 9956 15861 9965 15895
rect 9965 15861 9999 15895
rect 9999 15861 10008 15895
rect 9956 15852 10008 15861
rect 10324 15852 10376 15904
rect 10876 15852 10928 15904
rect 11152 15852 11204 15904
rect 15752 15920 15804 15972
rect 16120 15920 16172 15972
rect 16212 15963 16264 15972
rect 16212 15929 16221 15963
rect 16221 15929 16255 15963
rect 16255 15929 16264 15963
rect 16212 15920 16264 15929
rect 18328 15920 18380 15972
rect 13268 15852 13320 15904
rect 13728 15852 13780 15904
rect 17040 15852 17092 15904
rect 17224 15895 17276 15904
rect 17224 15861 17233 15895
rect 17233 15861 17267 15895
rect 17267 15861 17276 15895
rect 17224 15852 17276 15861
rect 18788 15895 18840 15904
rect 18788 15861 18797 15895
rect 18797 15861 18831 15895
rect 18831 15861 18840 15895
rect 18788 15852 18840 15861
rect 19064 15895 19116 15904
rect 19064 15861 19073 15895
rect 19073 15861 19107 15895
rect 19107 15861 19116 15895
rect 19064 15852 19116 15861
rect 21640 15988 21692 16040
rect 22560 15988 22612 16040
rect 23388 16056 23440 16108
rect 25136 16192 25188 16244
rect 24952 16124 25004 16176
rect 26608 16192 26660 16244
rect 28080 16192 28132 16244
rect 29000 16235 29052 16244
rect 29000 16201 29009 16235
rect 29009 16201 29043 16235
rect 29043 16201 29052 16235
rect 29000 16192 29052 16201
rect 26332 16124 26384 16176
rect 30840 16192 30892 16244
rect 32404 16235 32456 16244
rect 32404 16201 32413 16235
rect 32413 16201 32447 16235
rect 32447 16201 32456 16235
rect 32404 16192 32456 16201
rect 32588 16192 32640 16244
rect 30748 16124 30800 16176
rect 25504 16056 25556 16108
rect 25596 16056 25648 16108
rect 27528 16056 27580 16108
rect 29368 16031 29420 16040
rect 29368 15997 29377 16031
rect 29377 15997 29411 16031
rect 29411 15997 29420 16031
rect 29368 15988 29420 15997
rect 29644 16056 29696 16108
rect 29828 16056 29880 16108
rect 32588 16099 32640 16108
rect 32588 16065 32597 16099
rect 32597 16065 32631 16099
rect 32631 16065 32640 16099
rect 32588 16056 32640 16065
rect 30104 15988 30156 16040
rect 32404 15988 32456 16040
rect 32956 16235 33008 16244
rect 32956 16201 32965 16235
rect 32965 16201 32999 16235
rect 32999 16201 33008 16235
rect 32956 16192 33008 16201
rect 36544 16192 36596 16244
rect 33692 16124 33744 16176
rect 34888 16056 34940 16108
rect 35348 16099 35400 16108
rect 35348 16065 35357 16099
rect 35357 16065 35391 16099
rect 35391 16065 35400 16099
rect 35348 16056 35400 16065
rect 35808 16099 35860 16108
rect 35808 16065 35817 16099
rect 35817 16065 35851 16099
rect 35851 16065 35860 16099
rect 35808 16056 35860 16065
rect 38752 16235 38804 16244
rect 38752 16201 38761 16235
rect 38761 16201 38795 16235
rect 38795 16201 38804 16235
rect 38752 16192 38804 16201
rect 42800 16124 42852 16176
rect 34336 15988 34388 16040
rect 34796 15988 34848 16040
rect 36544 16031 36596 16040
rect 36544 15997 36553 16031
rect 36553 15997 36587 16031
rect 36587 15997 36596 16031
rect 36544 15988 36596 15997
rect 36636 16031 36688 16040
rect 36636 15997 36645 16031
rect 36645 15997 36679 16031
rect 36679 15997 36688 16031
rect 36636 15988 36688 15997
rect 36912 16056 36964 16108
rect 39028 16056 39080 16108
rect 20168 15852 20220 15904
rect 22652 15920 22704 15972
rect 22744 15920 22796 15972
rect 25228 15920 25280 15972
rect 25872 15920 25924 15972
rect 22100 15852 22152 15904
rect 23020 15895 23072 15904
rect 23020 15861 23029 15895
rect 23029 15861 23063 15895
rect 23063 15861 23072 15895
rect 23020 15852 23072 15861
rect 23204 15895 23256 15904
rect 23204 15861 23213 15895
rect 23213 15861 23247 15895
rect 23247 15861 23256 15895
rect 23204 15852 23256 15861
rect 24124 15852 24176 15904
rect 26332 15852 26384 15904
rect 26516 15852 26568 15904
rect 29736 15895 29788 15904
rect 29736 15861 29745 15895
rect 29745 15861 29779 15895
rect 29779 15861 29788 15895
rect 29736 15852 29788 15861
rect 30104 15852 30156 15904
rect 32312 15852 32364 15904
rect 32588 15895 32640 15904
rect 32588 15861 32597 15895
rect 32597 15861 32631 15895
rect 32631 15861 32640 15895
rect 32588 15852 32640 15861
rect 32772 15852 32824 15904
rect 33600 15852 33652 15904
rect 35440 15920 35492 15972
rect 36728 15963 36780 15972
rect 36728 15929 36737 15963
rect 36737 15929 36771 15963
rect 36771 15929 36780 15963
rect 36728 15920 36780 15929
rect 37004 15988 37056 16040
rect 38660 16031 38712 16040
rect 38660 15997 38669 16031
rect 38669 15997 38703 16031
rect 38703 15997 38712 16031
rect 38660 15988 38712 15997
rect 44272 15920 44324 15972
rect 35808 15852 35860 15904
rect 37188 15852 37240 15904
rect 44456 15895 44508 15904
rect 44456 15861 44465 15895
rect 44465 15861 44499 15895
rect 44499 15861 44508 15895
rect 44456 15852 44508 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2780 15648 2832 15700
rect 5724 15648 5776 15700
rect 5908 15691 5960 15700
rect 5908 15657 5917 15691
rect 5917 15657 5951 15691
rect 5951 15657 5960 15691
rect 5908 15648 5960 15657
rect 6644 15691 6696 15700
rect 6644 15657 6653 15691
rect 6653 15657 6687 15691
rect 6687 15657 6696 15691
rect 6644 15648 6696 15657
rect 2964 15580 3016 15632
rect 3976 15580 4028 15632
rect 5448 15580 5500 15632
rect 6276 15512 6328 15564
rect 6644 15512 6696 15564
rect 7196 15648 7248 15700
rect 7564 15648 7616 15700
rect 8760 15648 8812 15700
rect 8852 15648 8904 15700
rect 7104 15580 7156 15632
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 2412 15487 2464 15496
rect 2412 15453 2421 15487
rect 2421 15453 2455 15487
rect 2455 15453 2464 15487
rect 2412 15444 2464 15453
rect 2688 15444 2740 15496
rect 4068 15444 4120 15496
rect 2228 15308 2280 15360
rect 2780 15308 2832 15360
rect 5632 15376 5684 15428
rect 3240 15308 3292 15360
rect 3516 15308 3568 15360
rect 5908 15444 5960 15496
rect 6736 15444 6788 15496
rect 6920 15444 6972 15496
rect 7380 15444 7432 15496
rect 7656 15512 7708 15564
rect 6276 15419 6328 15428
rect 6276 15385 6285 15419
rect 6285 15385 6319 15419
rect 6319 15385 6328 15419
rect 6276 15376 6328 15385
rect 7012 15419 7064 15428
rect 7012 15385 7021 15419
rect 7021 15385 7055 15419
rect 7055 15385 7064 15419
rect 7012 15376 7064 15385
rect 7104 15419 7156 15428
rect 7104 15385 7113 15419
rect 7113 15385 7147 15419
rect 7147 15385 7156 15419
rect 7104 15376 7156 15385
rect 5908 15308 5960 15360
rect 6736 15308 6788 15360
rect 7932 15444 7984 15496
rect 8116 15487 8168 15496
rect 8116 15453 8125 15487
rect 8125 15453 8159 15487
rect 8159 15453 8168 15487
rect 8116 15444 8168 15453
rect 8576 15444 8628 15496
rect 9680 15580 9732 15632
rect 10600 15648 10652 15700
rect 10876 15580 10928 15632
rect 9496 15555 9548 15564
rect 9496 15521 9505 15555
rect 9505 15521 9539 15555
rect 9539 15521 9548 15555
rect 9496 15512 9548 15521
rect 10324 15512 10376 15564
rect 10416 15555 10468 15564
rect 10416 15521 10425 15555
rect 10425 15521 10459 15555
rect 10459 15521 10468 15555
rect 10416 15512 10468 15521
rect 11612 15580 11664 15632
rect 12624 15648 12676 15700
rect 12716 15580 12768 15632
rect 12900 15580 12952 15632
rect 12992 15580 13044 15632
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 12808 15512 12860 15564
rect 14924 15648 14976 15700
rect 14372 15580 14424 15632
rect 15936 15580 15988 15632
rect 16120 15580 16172 15632
rect 20168 15648 20220 15700
rect 22284 15691 22336 15700
rect 22284 15657 22293 15691
rect 22293 15657 22327 15691
rect 22327 15657 22336 15691
rect 22284 15648 22336 15657
rect 22560 15648 22612 15700
rect 23848 15691 23900 15700
rect 23848 15657 23857 15691
rect 23857 15657 23891 15691
rect 23891 15657 23900 15691
rect 23848 15648 23900 15657
rect 25596 15691 25648 15700
rect 25596 15657 25605 15691
rect 25605 15657 25639 15691
rect 25639 15657 25648 15691
rect 25596 15648 25648 15657
rect 17776 15580 17828 15632
rect 17960 15580 18012 15632
rect 9772 15444 9824 15453
rect 11152 15487 11204 15496
rect 11152 15453 11161 15487
rect 11161 15453 11195 15487
rect 11195 15453 11204 15487
rect 11152 15444 11204 15453
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 12716 15487 12768 15496
rect 12716 15453 12725 15487
rect 12725 15453 12759 15487
rect 12759 15453 12768 15487
rect 12716 15444 12768 15453
rect 12900 15487 12952 15496
rect 12900 15453 12914 15487
rect 12914 15453 12948 15487
rect 12948 15453 12952 15487
rect 15108 15555 15160 15564
rect 15108 15521 15117 15555
rect 15117 15521 15151 15555
rect 15151 15521 15160 15555
rect 15108 15512 15160 15521
rect 16028 15512 16080 15564
rect 14096 15487 14148 15496
rect 12900 15444 12952 15453
rect 14096 15453 14105 15487
rect 14105 15453 14139 15487
rect 14139 15453 14148 15487
rect 14096 15444 14148 15453
rect 14188 15444 14240 15496
rect 14740 15444 14792 15496
rect 15936 15487 15988 15496
rect 15936 15453 15945 15487
rect 15945 15453 15979 15487
rect 15979 15453 15988 15487
rect 15936 15444 15988 15453
rect 16396 15487 16448 15496
rect 16396 15453 16399 15487
rect 16399 15453 16448 15487
rect 16396 15444 16448 15453
rect 16764 15444 16816 15496
rect 17960 15487 18012 15496
rect 17960 15453 17969 15487
rect 17969 15453 18003 15487
rect 18003 15453 18012 15487
rect 17960 15444 18012 15453
rect 18052 15487 18104 15496
rect 19064 15580 19116 15632
rect 28080 15691 28132 15700
rect 28080 15657 28089 15691
rect 28089 15657 28123 15691
rect 28123 15657 28132 15691
rect 28080 15648 28132 15657
rect 28264 15691 28316 15700
rect 28264 15657 28273 15691
rect 28273 15657 28307 15691
rect 28307 15657 28316 15691
rect 28264 15648 28316 15657
rect 29092 15648 29144 15700
rect 29920 15691 29972 15700
rect 29920 15657 29929 15691
rect 29929 15657 29963 15691
rect 29963 15657 29972 15691
rect 29920 15648 29972 15657
rect 31852 15648 31904 15700
rect 22468 15555 22520 15564
rect 22468 15521 22477 15555
rect 22477 15521 22511 15555
rect 22511 15521 22520 15555
rect 31760 15580 31812 15632
rect 22468 15512 22520 15521
rect 18052 15453 18066 15487
rect 18066 15453 18100 15487
rect 18100 15453 18104 15487
rect 18052 15444 18104 15453
rect 8484 15308 8536 15360
rect 9036 15308 9088 15360
rect 10048 15308 10100 15360
rect 10784 15351 10836 15360
rect 10784 15317 10793 15351
rect 10793 15317 10827 15351
rect 10827 15317 10836 15351
rect 10784 15308 10836 15317
rect 10876 15308 10928 15360
rect 12348 15376 12400 15428
rect 12808 15419 12860 15428
rect 12808 15385 12817 15419
rect 12817 15385 12851 15419
rect 12851 15385 12860 15419
rect 12808 15376 12860 15385
rect 13728 15419 13780 15428
rect 13728 15385 13737 15419
rect 13737 15385 13771 15419
rect 13771 15385 13780 15419
rect 13728 15376 13780 15385
rect 13912 15376 13964 15428
rect 14372 15419 14424 15428
rect 14372 15385 14381 15419
rect 14381 15385 14415 15419
rect 14415 15385 14424 15419
rect 14372 15376 14424 15385
rect 11980 15308 12032 15360
rect 14740 15308 14792 15360
rect 15844 15308 15896 15360
rect 16212 15419 16264 15428
rect 16212 15385 16221 15419
rect 16221 15385 16255 15419
rect 16255 15385 16264 15419
rect 16212 15376 16264 15385
rect 16304 15308 16356 15360
rect 16488 15308 16540 15360
rect 17500 15308 17552 15360
rect 18144 15376 18196 15428
rect 18512 15444 18564 15496
rect 18696 15487 18748 15496
rect 18696 15453 18705 15487
rect 18705 15453 18739 15487
rect 18739 15453 18748 15487
rect 18696 15444 18748 15453
rect 18880 15487 18932 15496
rect 18880 15453 18883 15487
rect 18883 15453 18932 15487
rect 18880 15444 18932 15453
rect 22376 15444 22428 15496
rect 23204 15444 23256 15496
rect 19432 15376 19484 15428
rect 22284 15419 22336 15428
rect 22284 15385 22293 15419
rect 22293 15385 22327 15419
rect 22327 15385 22336 15419
rect 22284 15376 22336 15385
rect 23296 15376 23348 15428
rect 26332 15444 26384 15496
rect 26700 15487 26752 15496
rect 26700 15453 26709 15487
rect 26709 15453 26743 15487
rect 26743 15453 26752 15487
rect 29184 15512 29236 15564
rect 32588 15691 32640 15700
rect 32588 15657 32597 15691
rect 32597 15657 32631 15691
rect 32631 15657 32640 15691
rect 32588 15648 32640 15657
rect 32864 15691 32916 15700
rect 32864 15657 32873 15691
rect 32873 15657 32907 15691
rect 32907 15657 32916 15691
rect 32864 15648 32916 15657
rect 33324 15691 33376 15700
rect 33324 15657 33333 15691
rect 33333 15657 33367 15691
rect 33367 15657 33376 15691
rect 33324 15648 33376 15657
rect 33508 15691 33560 15700
rect 33508 15657 33517 15691
rect 33517 15657 33551 15691
rect 33551 15657 33560 15691
rect 33508 15648 33560 15657
rect 34336 15648 34388 15700
rect 34796 15691 34848 15700
rect 34796 15657 34805 15691
rect 34805 15657 34839 15691
rect 34839 15657 34848 15691
rect 34796 15648 34848 15657
rect 32680 15580 32732 15632
rect 33048 15580 33100 15632
rect 33232 15580 33284 15632
rect 37004 15691 37056 15700
rect 37004 15657 37013 15691
rect 37013 15657 37047 15691
rect 37047 15657 37056 15691
rect 37004 15648 37056 15657
rect 37280 15648 37332 15700
rect 34704 15512 34756 15564
rect 34796 15555 34848 15564
rect 34796 15521 34805 15555
rect 34805 15521 34839 15555
rect 34839 15521 34848 15555
rect 34796 15512 34848 15521
rect 41420 15512 41472 15564
rect 26700 15444 26752 15453
rect 23756 15308 23808 15360
rect 26240 15376 26292 15428
rect 26976 15376 27028 15428
rect 27804 15419 27856 15428
rect 27804 15385 27813 15419
rect 27813 15385 27847 15419
rect 27847 15385 27856 15419
rect 27804 15376 27856 15385
rect 29552 15487 29604 15496
rect 29552 15453 29561 15487
rect 29561 15453 29595 15487
rect 29595 15453 29604 15487
rect 29552 15444 29604 15453
rect 29644 15487 29696 15496
rect 29644 15453 29653 15487
rect 29653 15453 29687 15487
rect 29687 15453 29696 15487
rect 29644 15444 29696 15453
rect 32772 15444 32824 15496
rect 32956 15487 33008 15496
rect 32956 15453 32965 15487
rect 32965 15453 32999 15487
rect 32999 15453 33008 15487
rect 32956 15444 33008 15453
rect 33048 15487 33100 15496
rect 33048 15453 33057 15487
rect 33057 15453 33091 15487
rect 33091 15453 33100 15487
rect 33048 15444 33100 15453
rect 33324 15487 33376 15496
rect 33324 15453 33333 15487
rect 33333 15453 33367 15487
rect 33367 15453 33376 15487
rect 33324 15444 33376 15453
rect 33600 15487 33652 15496
rect 33600 15453 33609 15487
rect 33609 15453 33643 15487
rect 33643 15453 33652 15487
rect 33600 15444 33652 15453
rect 32220 15376 32272 15428
rect 32864 15376 32916 15428
rect 33784 15419 33836 15428
rect 33784 15385 33793 15419
rect 33793 15385 33827 15419
rect 33827 15385 33836 15419
rect 33784 15376 33836 15385
rect 24216 15351 24268 15360
rect 24216 15317 24225 15351
rect 24225 15317 24259 15351
rect 24259 15317 24268 15351
rect 24216 15308 24268 15317
rect 25228 15351 25280 15360
rect 25228 15317 25237 15351
rect 25237 15317 25271 15351
rect 25271 15317 25280 15351
rect 25228 15308 25280 15317
rect 25688 15308 25740 15360
rect 26148 15308 26200 15360
rect 27068 15351 27120 15360
rect 27068 15317 27077 15351
rect 27077 15317 27111 15351
rect 27111 15317 27120 15351
rect 27068 15308 27120 15317
rect 27528 15308 27580 15360
rect 30748 15308 30800 15360
rect 31208 15308 31260 15360
rect 34244 15487 34296 15496
rect 34244 15453 34253 15487
rect 34253 15453 34287 15487
rect 34287 15453 34296 15487
rect 34244 15444 34296 15453
rect 35808 15376 35860 15428
rect 37648 15444 37700 15496
rect 38568 15444 38620 15496
rect 40224 15444 40276 15496
rect 37188 15376 37240 15428
rect 41236 15487 41288 15496
rect 41236 15453 41245 15487
rect 41245 15453 41279 15487
rect 41279 15453 41288 15487
rect 41236 15444 41288 15453
rect 42340 15444 42392 15496
rect 37096 15308 37148 15360
rect 38660 15308 38712 15360
rect 43076 15308 43128 15360
rect 44088 15308 44140 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 2596 15104 2648 15156
rect 3240 15104 3292 15156
rect 3608 15036 3660 15088
rect 8116 15104 8168 15156
rect 8392 15104 8444 15156
rect 8852 15147 8904 15156
rect 8852 15113 8861 15147
rect 8861 15113 8895 15147
rect 8895 15113 8904 15147
rect 8852 15104 8904 15113
rect 10692 15104 10744 15156
rect 11060 15147 11112 15156
rect 11060 15113 11069 15147
rect 11069 15113 11103 15147
rect 11103 15113 11112 15147
rect 11060 15104 11112 15113
rect 11612 15104 11664 15156
rect 11980 15104 12032 15156
rect 12164 15147 12216 15156
rect 12164 15113 12173 15147
rect 12173 15113 12207 15147
rect 12207 15113 12216 15147
rect 12164 15104 12216 15113
rect 6920 15036 6972 15088
rect 2504 14968 2556 15020
rect 3516 14968 3568 15020
rect 2688 14943 2740 14952
rect 2688 14909 2697 14943
rect 2697 14909 2731 14943
rect 2731 14909 2740 14943
rect 2688 14900 2740 14909
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 7104 15011 7156 15020
rect 7104 14977 7113 15011
rect 7113 14977 7147 15011
rect 7147 14977 7156 15011
rect 7104 14968 7156 14977
rect 7748 15036 7800 15088
rect 7932 14968 7984 15020
rect 8024 14968 8076 15020
rect 9220 15036 9272 15088
rect 10048 15036 10100 15088
rect 13728 15104 13780 15156
rect 8852 14968 8904 15020
rect 9312 14968 9364 15020
rect 9864 14968 9916 15020
rect 10508 14968 10560 15020
rect 8484 14900 8536 14952
rect 6920 14832 6972 14884
rect 7840 14832 7892 14884
rect 9496 14900 9548 14952
rect 9956 14900 10008 14952
rect 10600 14943 10652 14952
rect 10600 14909 10609 14943
rect 10609 14909 10643 14943
rect 10643 14909 10652 14943
rect 10600 14900 10652 14909
rect 10876 14968 10928 15020
rect 11888 14968 11940 15020
rect 11980 14968 12032 15020
rect 13084 15036 13136 15088
rect 14004 15036 14056 15088
rect 15108 15104 15160 15156
rect 15200 15104 15252 15156
rect 18420 15104 18472 15156
rect 18696 15104 18748 15156
rect 14556 14968 14608 15020
rect 18512 15036 18564 15088
rect 21180 15104 21232 15156
rect 23756 15104 23808 15156
rect 23848 15147 23900 15156
rect 23848 15113 23857 15147
rect 23857 15113 23891 15147
rect 23891 15113 23900 15147
rect 23848 15104 23900 15113
rect 14924 15011 14976 15020
rect 14924 14977 14933 15011
rect 14933 14977 14967 15011
rect 14967 14977 14976 15011
rect 14924 14968 14976 14977
rect 15384 14968 15436 15020
rect 15844 14968 15896 15020
rect 11612 14900 11664 14952
rect 16764 14900 16816 14952
rect 3976 14764 4028 14816
rect 6092 14807 6144 14816
rect 6092 14773 6101 14807
rect 6101 14773 6135 14807
rect 6135 14773 6144 14807
rect 6092 14764 6144 14773
rect 6276 14764 6328 14816
rect 7012 14807 7064 14816
rect 7012 14773 7021 14807
rect 7021 14773 7055 14807
rect 7055 14773 7064 14807
rect 7012 14764 7064 14773
rect 7196 14764 7248 14816
rect 11152 14832 11204 14884
rect 11704 14832 11756 14884
rect 9772 14807 9824 14816
rect 9772 14773 9781 14807
rect 9781 14773 9815 14807
rect 9815 14773 9824 14807
rect 9772 14764 9824 14773
rect 10508 14764 10560 14816
rect 11520 14764 11572 14816
rect 12072 14764 12124 14816
rect 14832 14832 14884 14884
rect 15108 14832 15160 14884
rect 16672 14832 16724 14884
rect 19892 15036 19944 15088
rect 26240 15104 26292 15156
rect 19248 14968 19300 15020
rect 19524 14900 19576 14952
rect 23020 14968 23072 15020
rect 23572 14968 23624 15020
rect 23664 14968 23716 15020
rect 24308 15011 24360 15020
rect 24308 14977 24317 15011
rect 24317 14977 24351 15011
rect 24351 14977 24360 15011
rect 24308 14968 24360 14977
rect 26148 15011 26200 15020
rect 26148 14977 26157 15011
rect 26157 14977 26191 15011
rect 26191 14977 26200 15011
rect 26148 14968 26200 14977
rect 26424 15011 26476 15020
rect 26424 14977 26433 15011
rect 26433 14977 26467 15011
rect 26467 14977 26476 15011
rect 26424 14968 26476 14977
rect 15752 14764 15804 14816
rect 19432 14832 19484 14884
rect 23756 14900 23808 14952
rect 25228 14900 25280 14952
rect 27344 15147 27396 15156
rect 27344 15113 27353 15147
rect 27353 15113 27387 15147
rect 27387 15113 27396 15147
rect 27344 15104 27396 15113
rect 27804 15104 27856 15156
rect 26884 15036 26936 15088
rect 29460 15036 29512 15088
rect 29552 15036 29604 15088
rect 31300 15104 31352 15156
rect 27712 14968 27764 15020
rect 28724 14968 28776 15020
rect 30840 15011 30892 15020
rect 30840 14977 30849 15011
rect 30849 14977 30883 15011
rect 30883 14977 30892 15011
rect 30840 14968 30892 14977
rect 31116 14968 31168 15020
rect 31208 15011 31260 15020
rect 31208 14977 31217 15011
rect 31217 14977 31251 15011
rect 31251 14977 31260 15011
rect 31208 14968 31260 14977
rect 31576 15104 31628 15156
rect 32956 15104 33008 15156
rect 33784 15104 33836 15156
rect 36176 15104 36228 15156
rect 39028 15147 39080 15156
rect 39028 15113 39037 15147
rect 39037 15113 39071 15147
rect 39071 15113 39080 15147
rect 39028 15104 39080 15113
rect 41420 15104 41472 15156
rect 33508 15079 33560 15088
rect 33508 15045 33517 15079
rect 33517 15045 33551 15079
rect 33551 15045 33560 15079
rect 33508 15036 33560 15045
rect 37372 15036 37424 15088
rect 31576 14968 31628 15020
rect 31760 15011 31812 15020
rect 31760 14977 31769 15011
rect 31769 14977 31803 15011
rect 31803 14977 31812 15011
rect 31760 14968 31812 14977
rect 33140 14968 33192 15020
rect 33692 15011 33744 15020
rect 33692 14977 33701 15011
rect 33701 14977 33735 15011
rect 33735 14977 33744 15011
rect 33692 14968 33744 14977
rect 27344 14900 27396 14952
rect 27804 14900 27856 14952
rect 30656 14900 30708 14952
rect 31024 14943 31076 14952
rect 31024 14909 31033 14943
rect 31033 14909 31067 14943
rect 31067 14909 31076 14943
rect 31024 14900 31076 14909
rect 31392 14900 31444 14952
rect 37648 15011 37700 15020
rect 37648 14977 37657 15011
rect 37657 14977 37691 15011
rect 37691 14977 37700 15011
rect 37648 14968 37700 14977
rect 37740 14968 37792 15020
rect 43076 14943 43128 14952
rect 43076 14909 43085 14943
rect 43085 14909 43119 14943
rect 43119 14909 43128 14943
rect 43076 14900 43128 14909
rect 19984 14832 20036 14884
rect 20720 14832 20772 14884
rect 21640 14832 21692 14884
rect 20812 14764 20864 14816
rect 23572 14764 23624 14816
rect 23664 14764 23716 14816
rect 24124 14764 24176 14816
rect 31208 14832 31260 14884
rect 31300 14832 31352 14884
rect 26332 14807 26384 14816
rect 26332 14773 26341 14807
rect 26341 14773 26375 14807
rect 26375 14773 26384 14807
rect 26332 14764 26384 14773
rect 26884 14764 26936 14816
rect 27068 14807 27120 14816
rect 27068 14773 27077 14807
rect 27077 14773 27111 14807
rect 27111 14773 27120 14807
rect 27068 14764 27120 14773
rect 27804 14764 27856 14816
rect 30932 14807 30984 14816
rect 30932 14773 30941 14807
rect 30941 14773 30975 14807
rect 30975 14773 30984 14807
rect 30932 14764 30984 14773
rect 31576 14764 31628 14816
rect 31852 14764 31904 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2412 14560 2464 14612
rect 7104 14560 7156 14612
rect 7840 14560 7892 14612
rect 7656 14492 7708 14544
rect 6092 14424 6144 14476
rect 7748 14424 7800 14476
rect 8208 14492 8260 14544
rect 9128 14492 9180 14544
rect 8024 14467 8076 14476
rect 8024 14433 8033 14467
rect 8033 14433 8067 14467
rect 8067 14433 8076 14467
rect 8024 14424 8076 14433
rect 848 14356 900 14408
rect 2320 14331 2372 14340
rect 2320 14297 2329 14331
rect 2329 14297 2363 14331
rect 2363 14297 2372 14331
rect 2320 14288 2372 14297
rect 3976 14288 4028 14340
rect 6920 14356 6972 14408
rect 8392 14356 8444 14408
rect 2780 14220 2832 14272
rect 4804 14220 4856 14272
rect 7748 14288 7800 14340
rect 8760 14356 8812 14408
rect 9220 14424 9272 14476
rect 9772 14560 9824 14612
rect 12624 14560 12676 14612
rect 16580 14560 16632 14612
rect 9588 14535 9640 14544
rect 9588 14501 9597 14535
rect 9597 14501 9631 14535
rect 9631 14501 9640 14535
rect 9588 14492 9640 14501
rect 11704 14424 11756 14476
rect 13360 14424 13412 14476
rect 13912 14424 13964 14476
rect 9312 14399 9364 14408
rect 9312 14365 9321 14399
rect 9321 14365 9355 14399
rect 9355 14365 9364 14399
rect 9312 14356 9364 14365
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 14188 14356 14240 14408
rect 15016 14424 15068 14476
rect 16672 14492 16724 14544
rect 18604 14492 18656 14544
rect 19248 14492 19300 14544
rect 19984 14560 20036 14612
rect 20260 14492 20312 14544
rect 22100 14492 22152 14544
rect 15752 14424 15804 14476
rect 16028 14356 16080 14408
rect 16120 14399 16172 14408
rect 16120 14365 16129 14399
rect 16129 14365 16163 14399
rect 16163 14365 16172 14399
rect 16120 14356 16172 14365
rect 20352 14424 20404 14476
rect 16764 14356 16816 14408
rect 19616 14356 19668 14408
rect 19800 14356 19852 14408
rect 20076 14399 20128 14408
rect 20076 14365 20085 14399
rect 20085 14365 20119 14399
rect 20119 14365 20128 14399
rect 20076 14356 20128 14365
rect 20168 14399 20220 14408
rect 20168 14365 20177 14399
rect 20177 14365 20211 14399
rect 20211 14365 20220 14399
rect 20168 14356 20220 14365
rect 20536 14356 20588 14408
rect 21732 14399 21784 14408
rect 21732 14365 21741 14399
rect 21741 14365 21775 14399
rect 21775 14365 21784 14399
rect 21732 14356 21784 14365
rect 6736 14220 6788 14272
rect 7012 14263 7064 14272
rect 7012 14229 7021 14263
rect 7021 14229 7055 14263
rect 7055 14229 7064 14263
rect 7012 14220 7064 14229
rect 7472 14220 7524 14272
rect 7932 14220 7984 14272
rect 9496 14288 9548 14340
rect 16856 14288 16908 14340
rect 14832 14220 14884 14272
rect 15108 14220 15160 14272
rect 15660 14263 15712 14272
rect 15660 14229 15669 14263
rect 15669 14229 15703 14263
rect 15703 14229 15712 14263
rect 15660 14220 15712 14229
rect 17040 14220 17092 14272
rect 19248 14220 19300 14272
rect 20352 14331 20404 14340
rect 20352 14297 20361 14331
rect 20361 14297 20395 14331
rect 20395 14297 20404 14331
rect 20352 14288 20404 14297
rect 21916 14220 21968 14272
rect 22008 14263 22060 14272
rect 22008 14229 22017 14263
rect 22017 14229 22051 14263
rect 22051 14229 22060 14263
rect 22008 14220 22060 14229
rect 22560 14467 22612 14476
rect 22560 14433 22569 14467
rect 22569 14433 22603 14467
rect 22603 14433 22612 14467
rect 22560 14424 22612 14433
rect 22928 14603 22980 14612
rect 22928 14569 22937 14603
rect 22937 14569 22971 14603
rect 22971 14569 22980 14603
rect 22928 14560 22980 14569
rect 23572 14603 23624 14612
rect 23572 14569 23581 14603
rect 23581 14569 23615 14603
rect 23615 14569 23624 14603
rect 23572 14560 23624 14569
rect 24308 14560 24360 14612
rect 30932 14603 30984 14612
rect 25596 14492 25648 14544
rect 30932 14569 30941 14603
rect 30941 14569 30975 14603
rect 30975 14569 30984 14603
rect 30932 14560 30984 14569
rect 31116 14603 31168 14612
rect 31116 14569 31125 14603
rect 31125 14569 31159 14603
rect 31159 14569 31168 14603
rect 31116 14560 31168 14569
rect 23020 14356 23072 14408
rect 22468 14331 22520 14340
rect 22468 14297 22477 14331
rect 22477 14297 22511 14331
rect 22511 14297 22520 14331
rect 22468 14288 22520 14297
rect 24032 14424 24084 14476
rect 24124 14424 24176 14476
rect 27344 14424 27396 14476
rect 31760 14492 31812 14544
rect 31576 14424 31628 14476
rect 33692 14424 33744 14476
rect 24676 14356 24728 14408
rect 26424 14356 26476 14408
rect 27436 14356 27488 14408
rect 30840 14399 30892 14408
rect 30840 14365 30849 14399
rect 30849 14365 30883 14399
rect 30883 14365 30892 14399
rect 30840 14356 30892 14365
rect 44272 14399 44324 14408
rect 44272 14365 44281 14399
rect 44281 14365 44315 14399
rect 44315 14365 44324 14399
rect 44272 14356 44324 14365
rect 28816 14288 28868 14340
rect 30288 14288 30340 14340
rect 31852 14288 31904 14340
rect 30472 14220 30524 14272
rect 44456 14263 44508 14272
rect 44456 14229 44465 14263
rect 44465 14229 44499 14263
rect 44499 14229 44508 14263
rect 44456 14220 44508 14229
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 2320 14016 2372 14068
rect 2504 14059 2556 14068
rect 2504 14025 2513 14059
rect 2513 14025 2547 14059
rect 2547 14025 2556 14059
rect 2504 14016 2556 14025
rect 2780 14016 2832 14068
rect 2688 13948 2740 14000
rect 4620 14016 4672 14068
rect 4804 14016 4856 14068
rect 5724 14059 5776 14068
rect 5724 14025 5733 14059
rect 5733 14025 5767 14059
rect 5767 14025 5776 14059
rect 5724 14016 5776 14025
rect 5816 14016 5868 14068
rect 10876 14016 10928 14068
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 3240 13880 3292 13932
rect 1584 13676 1636 13728
rect 2044 13855 2096 13864
rect 2044 13821 2053 13855
rect 2053 13821 2087 13855
rect 2087 13821 2096 13855
rect 2044 13812 2096 13821
rect 2136 13855 2188 13864
rect 2136 13821 2145 13855
rect 2145 13821 2179 13855
rect 2179 13821 2188 13855
rect 2136 13812 2188 13821
rect 2780 13744 2832 13796
rect 2964 13812 3016 13864
rect 5264 13948 5316 14000
rect 7840 13948 7892 14000
rect 11980 14016 12032 14068
rect 12072 14059 12124 14068
rect 12072 14025 12089 14059
rect 12089 14025 12123 14059
rect 12123 14025 12124 14059
rect 12072 14016 12124 14025
rect 15844 14016 15896 14068
rect 16856 14016 16908 14068
rect 17132 14059 17184 14068
rect 17132 14025 17141 14059
rect 17141 14025 17175 14059
rect 17175 14025 17184 14059
rect 17132 14016 17184 14025
rect 5908 13880 5960 13932
rect 8208 13923 8260 13932
rect 8208 13889 8217 13923
rect 8217 13889 8251 13923
rect 8251 13889 8260 13923
rect 8208 13880 8260 13889
rect 4804 13855 4856 13864
rect 4804 13821 4813 13855
rect 4813 13821 4847 13855
rect 4847 13821 4856 13855
rect 4804 13812 4856 13821
rect 4896 13855 4948 13864
rect 4896 13821 4905 13855
rect 4905 13821 4939 13855
rect 4939 13821 4948 13855
rect 4896 13812 4948 13821
rect 5448 13812 5500 13864
rect 5816 13812 5868 13864
rect 6092 13812 6144 13864
rect 5356 13744 5408 13796
rect 6644 13744 6696 13796
rect 8116 13812 8168 13864
rect 8576 13923 8628 13932
rect 8576 13889 8585 13923
rect 8585 13889 8619 13923
rect 8619 13889 8628 13923
rect 8576 13880 8628 13889
rect 8760 13855 8812 13864
rect 8760 13821 8769 13855
rect 8769 13821 8803 13855
rect 8803 13821 8812 13855
rect 8760 13812 8812 13821
rect 9588 13880 9640 13932
rect 10416 13923 10468 13932
rect 10416 13889 10425 13923
rect 10425 13889 10459 13923
rect 10459 13889 10468 13923
rect 10416 13880 10468 13889
rect 12716 13948 12768 14000
rect 9220 13812 9272 13864
rect 11980 13923 12032 13932
rect 11980 13889 11983 13923
rect 11983 13889 12032 13923
rect 10968 13812 11020 13864
rect 11980 13880 12032 13889
rect 12900 13880 12952 13932
rect 14556 13923 14608 13932
rect 14556 13889 14565 13923
rect 14565 13889 14599 13923
rect 14599 13889 14608 13923
rect 14556 13880 14608 13889
rect 14924 13880 14976 13932
rect 15200 13948 15252 14000
rect 15660 13880 15712 13932
rect 8576 13744 8628 13796
rect 12164 13812 12216 13864
rect 15108 13855 15160 13864
rect 15108 13821 15117 13855
rect 15117 13821 15151 13855
rect 15151 13821 15160 13855
rect 15108 13812 15160 13821
rect 15936 13923 15988 13932
rect 15936 13889 15945 13923
rect 15945 13889 15979 13923
rect 15979 13889 15988 13923
rect 15936 13880 15988 13889
rect 16028 13923 16080 13932
rect 16028 13889 16037 13923
rect 16037 13889 16071 13923
rect 16071 13889 16080 13923
rect 16028 13880 16080 13889
rect 16212 13880 16264 13932
rect 17408 13923 17460 13932
rect 17408 13889 17417 13923
rect 17417 13889 17451 13923
rect 17451 13889 17460 13923
rect 17408 13880 17460 13889
rect 17592 13923 17644 13932
rect 17592 13889 17601 13923
rect 17601 13889 17635 13923
rect 17635 13889 17644 13923
rect 17592 13880 17644 13889
rect 17684 13923 17736 13932
rect 17684 13889 17693 13923
rect 17693 13889 17727 13923
rect 17727 13889 17736 13923
rect 17684 13880 17736 13889
rect 17960 13880 18012 13932
rect 18696 13923 18748 13932
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 19616 13948 19668 14000
rect 23112 14016 23164 14068
rect 28080 14059 28132 14068
rect 28080 14025 28089 14059
rect 28089 14025 28123 14059
rect 28123 14025 28132 14059
rect 28080 14016 28132 14025
rect 22008 13991 22060 14000
rect 22008 13957 22017 13991
rect 22017 13957 22051 13991
rect 22051 13957 22060 13991
rect 22008 13948 22060 13957
rect 22192 13991 22244 14000
rect 22192 13957 22201 13991
rect 22201 13957 22235 13991
rect 22235 13957 22244 13991
rect 22192 13948 22244 13957
rect 19156 13923 19208 13932
rect 19156 13889 19159 13923
rect 19159 13889 19208 13923
rect 12348 13744 12400 13796
rect 13820 13744 13872 13796
rect 14188 13744 14240 13796
rect 17868 13812 17920 13864
rect 16948 13744 17000 13796
rect 18604 13812 18656 13864
rect 18788 13812 18840 13864
rect 19156 13880 19208 13889
rect 19708 13880 19760 13932
rect 22468 13880 22520 13932
rect 22836 13991 22888 14000
rect 22836 13957 22845 13991
rect 22845 13957 22879 13991
rect 22879 13957 22888 13991
rect 22836 13948 22888 13957
rect 26148 13948 26200 14000
rect 25596 13880 25648 13932
rect 25872 13923 25924 13932
rect 25872 13889 25881 13923
rect 25881 13889 25915 13923
rect 25915 13889 25924 13923
rect 25872 13880 25924 13889
rect 26240 13880 26292 13932
rect 26516 13880 26568 13932
rect 26608 13923 26660 13932
rect 26608 13889 26617 13923
rect 26617 13889 26651 13923
rect 26651 13889 26660 13923
rect 26608 13880 26660 13889
rect 26792 13923 26844 13932
rect 26792 13889 26801 13923
rect 26801 13889 26835 13923
rect 26835 13889 26844 13923
rect 26792 13880 26844 13889
rect 21732 13812 21784 13864
rect 25320 13812 25372 13864
rect 26332 13812 26384 13864
rect 4620 13676 4672 13728
rect 6000 13676 6052 13728
rect 9588 13676 9640 13728
rect 10600 13719 10652 13728
rect 10600 13685 10609 13719
rect 10609 13685 10643 13719
rect 10643 13685 10652 13719
rect 10600 13676 10652 13685
rect 10876 13676 10928 13728
rect 17408 13676 17460 13728
rect 22284 13744 22336 13796
rect 27160 13923 27212 13932
rect 27160 13889 27169 13923
rect 27169 13889 27203 13923
rect 27203 13889 27212 13923
rect 27160 13880 27212 13889
rect 27528 13923 27580 13932
rect 27528 13889 27537 13923
rect 27537 13889 27571 13923
rect 27571 13889 27580 13923
rect 27528 13880 27580 13889
rect 29000 14059 29052 14068
rect 29000 14025 29009 14059
rect 29009 14025 29043 14059
rect 29043 14025 29052 14059
rect 29000 14016 29052 14025
rect 34612 14016 34664 14068
rect 44088 14016 44140 14068
rect 28908 13948 28960 14000
rect 31668 13948 31720 14000
rect 32312 13991 32364 14000
rect 32312 13957 32321 13991
rect 32321 13957 32355 13991
rect 32355 13957 32364 13991
rect 32312 13948 32364 13957
rect 33324 13948 33376 14000
rect 27712 13855 27764 13864
rect 27712 13821 27721 13855
rect 27721 13821 27755 13855
rect 27755 13821 27764 13855
rect 27712 13812 27764 13821
rect 28540 13880 28592 13932
rect 33232 13880 33284 13932
rect 43076 13880 43128 13932
rect 34060 13812 34112 13864
rect 28816 13744 28868 13796
rect 28908 13744 28960 13796
rect 30288 13744 30340 13796
rect 25688 13676 25740 13728
rect 26424 13676 26476 13728
rect 26700 13676 26752 13728
rect 32312 13744 32364 13796
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2872 13472 2924 13524
rect 4712 13472 4764 13524
rect 4896 13515 4948 13524
rect 4896 13481 4905 13515
rect 4905 13481 4939 13515
rect 4939 13481 4948 13515
rect 4896 13472 4948 13481
rect 5356 13472 5408 13524
rect 5724 13472 5776 13524
rect 6552 13472 6604 13524
rect 1584 13379 1636 13388
rect 1584 13345 1593 13379
rect 1593 13345 1627 13379
rect 1627 13345 1636 13379
rect 1584 13336 1636 13345
rect 2044 13379 2096 13388
rect 2044 13345 2078 13379
rect 2078 13345 2096 13379
rect 2780 13404 2832 13456
rect 4068 13404 4120 13456
rect 5080 13404 5132 13456
rect 2044 13336 2096 13345
rect 2688 13336 2740 13388
rect 4528 13336 4580 13388
rect 5816 13404 5868 13456
rect 5908 13404 5960 13456
rect 6920 13472 6972 13524
rect 10416 13472 10468 13524
rect 11796 13472 11848 13524
rect 11888 13515 11940 13524
rect 11888 13481 11897 13515
rect 11897 13481 11931 13515
rect 11931 13481 11940 13515
rect 11888 13472 11940 13481
rect 12624 13472 12676 13524
rect 13084 13515 13136 13524
rect 13084 13481 13093 13515
rect 13093 13481 13127 13515
rect 13127 13481 13136 13515
rect 13084 13472 13136 13481
rect 13912 13472 13964 13524
rect 2872 13268 2924 13320
rect 2780 13200 2832 13252
rect 2136 13132 2188 13184
rect 2596 13132 2648 13184
rect 3148 13175 3200 13184
rect 3148 13141 3157 13175
rect 3157 13141 3191 13175
rect 3191 13141 3200 13175
rect 3148 13132 3200 13141
rect 3976 13200 4028 13252
rect 4804 13268 4856 13320
rect 6000 13379 6052 13388
rect 6000 13345 6009 13379
rect 6009 13345 6043 13379
rect 6043 13345 6052 13379
rect 6000 13336 6052 13345
rect 6644 13336 6696 13388
rect 4344 13243 4396 13252
rect 4344 13209 4353 13243
rect 4353 13209 4387 13243
rect 4387 13209 4396 13243
rect 4344 13200 4396 13209
rect 4528 13132 4580 13184
rect 5264 13243 5316 13252
rect 5264 13209 5273 13243
rect 5273 13209 5307 13243
rect 5307 13209 5316 13243
rect 5264 13200 5316 13209
rect 5908 13200 5960 13252
rect 6552 13268 6604 13320
rect 8852 13404 8904 13456
rect 9128 13447 9180 13456
rect 9128 13413 9137 13447
rect 9137 13413 9171 13447
rect 9171 13413 9180 13447
rect 9128 13404 9180 13413
rect 9312 13404 9364 13456
rect 9496 13404 9548 13456
rect 10968 13404 11020 13456
rect 11520 13447 11572 13456
rect 11520 13413 11529 13447
rect 11529 13413 11563 13447
rect 11563 13413 11572 13447
rect 11520 13404 11572 13413
rect 11980 13404 12032 13456
rect 8024 13336 8076 13388
rect 7472 13311 7524 13320
rect 7472 13277 7481 13311
rect 7481 13277 7515 13311
rect 7515 13277 7524 13311
rect 7472 13268 7524 13277
rect 7564 13268 7616 13320
rect 8576 13268 8628 13320
rect 9404 13311 9456 13320
rect 9404 13277 9434 13311
rect 9434 13277 9456 13311
rect 9404 13268 9456 13277
rect 9588 13336 9640 13388
rect 13820 13404 13872 13456
rect 14188 13404 14240 13456
rect 15476 13404 15528 13456
rect 17408 13515 17460 13524
rect 17408 13481 17417 13515
rect 17417 13481 17451 13515
rect 17451 13481 17460 13515
rect 17408 13472 17460 13481
rect 22284 13515 22336 13524
rect 22284 13481 22293 13515
rect 22293 13481 22327 13515
rect 22327 13481 22336 13515
rect 22284 13472 22336 13481
rect 22468 13515 22520 13524
rect 22468 13481 22477 13515
rect 22477 13481 22511 13515
rect 22511 13481 22520 13515
rect 22468 13472 22520 13481
rect 26056 13472 26108 13524
rect 26608 13472 26660 13524
rect 17776 13404 17828 13456
rect 22100 13404 22152 13456
rect 27160 13472 27212 13524
rect 29000 13472 29052 13524
rect 30012 13472 30064 13524
rect 36084 13472 36136 13524
rect 9956 13311 10008 13320
rect 9956 13277 9965 13311
rect 9965 13277 9999 13311
rect 9999 13277 10008 13311
rect 9956 13268 10008 13277
rect 10048 13268 10100 13320
rect 10968 13311 11020 13320
rect 10968 13277 10977 13311
rect 10977 13277 11011 13311
rect 11011 13277 11020 13311
rect 10968 13268 11020 13277
rect 11520 13268 11572 13320
rect 11704 13311 11756 13320
rect 11704 13277 11713 13311
rect 11713 13277 11747 13311
rect 11747 13277 11756 13311
rect 11704 13268 11756 13277
rect 11980 13311 12032 13320
rect 11980 13277 12029 13311
rect 12029 13277 12032 13311
rect 11980 13268 12032 13277
rect 12164 13311 12216 13320
rect 12164 13277 12176 13311
rect 12176 13277 12210 13311
rect 12210 13277 12216 13311
rect 12164 13268 12216 13277
rect 12348 13268 12400 13320
rect 12624 13336 12676 13388
rect 6920 13200 6972 13252
rect 10876 13243 10928 13252
rect 10876 13209 10885 13243
rect 10885 13209 10919 13243
rect 10919 13209 10928 13243
rect 10876 13200 10928 13209
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 12900 13311 12952 13320
rect 12900 13277 12914 13311
rect 12914 13277 12948 13311
rect 12948 13277 12952 13311
rect 12900 13268 12952 13277
rect 13636 13311 13688 13320
rect 13636 13277 13645 13311
rect 13645 13277 13679 13311
rect 13679 13277 13688 13311
rect 13636 13268 13688 13277
rect 5356 13132 5408 13184
rect 6092 13175 6144 13184
rect 6092 13141 6101 13175
rect 6101 13141 6135 13175
rect 6135 13141 6144 13175
rect 6092 13132 6144 13141
rect 6552 13132 6604 13184
rect 8116 13175 8168 13184
rect 8116 13141 8125 13175
rect 8125 13141 8159 13175
rect 8159 13141 8168 13175
rect 8116 13132 8168 13141
rect 9864 13132 9916 13184
rect 10416 13132 10468 13184
rect 11152 13132 11204 13184
rect 13452 13243 13504 13252
rect 13452 13209 13461 13243
rect 13461 13209 13495 13243
rect 13495 13209 13504 13243
rect 13452 13200 13504 13209
rect 14648 13311 14700 13320
rect 14648 13277 14657 13311
rect 14657 13277 14691 13311
rect 14691 13277 14700 13311
rect 14648 13268 14700 13277
rect 15016 13311 15068 13320
rect 15016 13277 15025 13311
rect 15025 13277 15059 13311
rect 15059 13277 15068 13311
rect 15016 13268 15068 13277
rect 15660 13268 15712 13320
rect 16028 13200 16080 13252
rect 13912 13132 13964 13184
rect 14280 13132 14332 13184
rect 16948 13268 17000 13320
rect 17500 13268 17552 13320
rect 17960 13268 18012 13320
rect 26608 13336 26660 13388
rect 28908 13379 28960 13388
rect 17040 13243 17092 13252
rect 17040 13209 17049 13243
rect 17049 13209 17083 13243
rect 17083 13209 17092 13243
rect 17040 13200 17092 13209
rect 17132 13243 17184 13252
rect 17132 13209 17141 13243
rect 17141 13209 17175 13243
rect 17175 13209 17184 13243
rect 17132 13200 17184 13209
rect 19156 13200 19208 13252
rect 20076 13200 20128 13252
rect 23480 13200 23532 13252
rect 18328 13132 18380 13184
rect 22100 13132 22152 13184
rect 25872 13200 25924 13252
rect 26332 13268 26384 13320
rect 28908 13345 28917 13379
rect 28917 13345 28951 13379
rect 28951 13345 28960 13379
rect 28908 13336 28960 13345
rect 28540 13311 28592 13320
rect 28540 13277 28549 13311
rect 28549 13277 28583 13311
rect 28583 13277 28592 13311
rect 28540 13268 28592 13277
rect 29644 13336 29696 13388
rect 31024 13336 31076 13388
rect 31392 13268 31444 13320
rect 28356 13243 28408 13252
rect 28356 13209 28365 13243
rect 28365 13209 28399 13243
rect 28399 13209 28408 13243
rect 28356 13200 28408 13209
rect 28816 13243 28868 13252
rect 28816 13209 28825 13243
rect 28825 13209 28859 13243
rect 28859 13209 28868 13243
rect 28816 13200 28868 13209
rect 29460 13200 29512 13252
rect 30932 13243 30984 13252
rect 30932 13209 30941 13243
rect 30941 13209 30975 13243
rect 30975 13209 30984 13243
rect 30932 13200 30984 13209
rect 31116 13243 31168 13252
rect 31116 13209 31125 13243
rect 31125 13209 31159 13243
rect 31159 13209 31168 13243
rect 31116 13200 31168 13209
rect 31576 13336 31628 13388
rect 37924 13336 37976 13388
rect 31668 13243 31720 13252
rect 31668 13209 31677 13243
rect 31677 13209 31711 13243
rect 31711 13209 31720 13243
rect 31668 13200 31720 13209
rect 37556 13132 37608 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 1584 12928 1636 12980
rect 2688 12928 2740 12980
rect 3332 12928 3384 12980
rect 4804 12928 4856 12980
rect 5540 12928 5592 12980
rect 10048 12928 10100 12980
rect 10508 12928 10560 12980
rect 2504 12860 2556 12912
rect 1584 12792 1636 12844
rect 2964 12835 3016 12844
rect 2964 12801 2973 12835
rect 2973 12801 3007 12835
rect 3007 12801 3016 12835
rect 2964 12792 3016 12801
rect 3240 12835 3292 12844
rect 3240 12801 3249 12835
rect 3249 12801 3283 12835
rect 3283 12801 3292 12835
rect 3240 12792 3292 12801
rect 5356 12903 5408 12912
rect 5356 12869 5365 12903
rect 5365 12869 5399 12903
rect 5399 12869 5408 12903
rect 5356 12860 5408 12869
rect 1676 12724 1728 12776
rect 2504 12767 2556 12776
rect 2504 12733 2513 12767
rect 2513 12733 2547 12767
rect 2547 12733 2556 12767
rect 2504 12724 2556 12733
rect 2596 12724 2648 12776
rect 4344 12724 4396 12776
rect 2872 12656 2924 12708
rect 5264 12792 5316 12844
rect 5724 12792 5776 12844
rect 5448 12724 5500 12776
rect 5908 12767 5960 12776
rect 5908 12733 5917 12767
rect 5917 12733 5951 12767
rect 5951 12733 5960 12767
rect 5908 12724 5960 12733
rect 6552 12767 6604 12776
rect 6552 12733 6561 12767
rect 6561 12733 6595 12767
rect 6595 12733 6604 12767
rect 6552 12724 6604 12733
rect 7196 12792 7248 12844
rect 8024 12792 8076 12844
rect 9588 12860 9640 12912
rect 10324 12903 10376 12912
rect 10324 12869 10333 12903
rect 10333 12869 10367 12903
rect 10367 12869 10376 12903
rect 11612 12971 11664 12980
rect 11612 12937 11621 12971
rect 11621 12937 11655 12971
rect 11655 12937 11664 12971
rect 11612 12928 11664 12937
rect 12440 12928 12492 12980
rect 14372 12928 14424 12980
rect 14556 12928 14608 12980
rect 17592 12928 17644 12980
rect 10324 12860 10376 12869
rect 8852 12792 8904 12844
rect 7932 12767 7984 12776
rect 7932 12733 7941 12767
rect 7941 12733 7975 12767
rect 7975 12733 7984 12767
rect 7932 12724 7984 12733
rect 8116 12724 8168 12776
rect 9680 12835 9732 12844
rect 9680 12801 9689 12835
rect 9689 12801 9723 12835
rect 9723 12801 9732 12835
rect 9680 12792 9732 12801
rect 9772 12792 9824 12844
rect 10692 12792 10744 12844
rect 13268 12903 13320 12912
rect 13268 12869 13277 12903
rect 13277 12869 13311 12903
rect 13311 12869 13320 12903
rect 13268 12860 13320 12869
rect 14004 12903 14056 12912
rect 14004 12869 14013 12903
rect 14013 12869 14047 12903
rect 14047 12869 14056 12903
rect 14004 12860 14056 12869
rect 15016 12860 15068 12912
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 12164 12835 12216 12844
rect 12164 12801 12173 12835
rect 12173 12801 12207 12835
rect 12207 12801 12216 12835
rect 12164 12792 12216 12801
rect 12440 12792 12492 12844
rect 4620 12699 4672 12708
rect 4620 12665 4629 12699
rect 4629 12665 4663 12699
rect 4663 12665 4672 12699
rect 4620 12656 4672 12665
rect 4712 12699 4764 12708
rect 4712 12665 4721 12699
rect 4721 12665 4755 12699
rect 4755 12665 4764 12699
rect 4712 12656 4764 12665
rect 2504 12588 2556 12640
rect 3976 12588 4028 12640
rect 4528 12588 4580 12640
rect 5632 12656 5684 12708
rect 7380 12656 7432 12708
rect 7748 12656 7800 12708
rect 9496 12699 9548 12708
rect 9496 12665 9505 12699
rect 9505 12665 9539 12699
rect 9539 12665 9548 12699
rect 9496 12656 9548 12665
rect 9588 12656 9640 12708
rect 12256 12767 12308 12776
rect 12256 12733 12265 12767
rect 12265 12733 12299 12767
rect 12299 12733 12308 12767
rect 12256 12724 12308 12733
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 14740 12835 14792 12844
rect 14740 12801 14749 12835
rect 14749 12801 14783 12835
rect 14783 12801 14792 12835
rect 14740 12792 14792 12801
rect 14832 12835 14884 12844
rect 14832 12801 14841 12835
rect 14841 12801 14875 12835
rect 14875 12801 14884 12835
rect 14832 12792 14884 12801
rect 15292 12835 15344 12844
rect 15292 12801 15301 12835
rect 15301 12801 15335 12835
rect 15335 12801 15344 12835
rect 15292 12792 15344 12801
rect 15752 12792 15804 12844
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 17316 12903 17368 12912
rect 17316 12869 17325 12903
rect 17325 12869 17359 12903
rect 17359 12869 17368 12903
rect 17316 12860 17368 12869
rect 17408 12903 17460 12912
rect 17408 12869 17417 12903
rect 17417 12869 17451 12903
rect 17451 12869 17460 12903
rect 17408 12860 17460 12869
rect 17500 12835 17552 12844
rect 18788 12928 18840 12980
rect 18880 12928 18932 12980
rect 18328 12903 18380 12912
rect 18328 12869 18337 12903
rect 18337 12869 18371 12903
rect 18371 12869 18380 12903
rect 18328 12860 18380 12869
rect 19616 12860 19668 12912
rect 17500 12801 17514 12835
rect 17514 12801 17548 12835
rect 17548 12801 17552 12835
rect 17500 12792 17552 12801
rect 16028 12724 16080 12776
rect 17960 12724 18012 12776
rect 18512 12835 18564 12844
rect 18512 12801 18515 12835
rect 18515 12801 18564 12835
rect 18512 12792 18564 12801
rect 18788 12835 18840 12844
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 19248 12835 19300 12844
rect 19248 12801 19251 12835
rect 19251 12801 19300 12835
rect 13452 12656 13504 12708
rect 14096 12656 14148 12708
rect 6552 12588 6604 12640
rect 7012 12588 7064 12640
rect 10508 12588 10560 12640
rect 10784 12588 10836 12640
rect 14188 12588 14240 12640
rect 17224 12656 17276 12708
rect 17684 12699 17736 12708
rect 17684 12665 17693 12699
rect 17693 12665 17727 12699
rect 17727 12665 17736 12699
rect 17684 12656 17736 12665
rect 18696 12656 18748 12708
rect 19248 12792 19300 12801
rect 19524 12835 19576 12844
rect 19524 12801 19533 12835
rect 19533 12801 19567 12835
rect 19567 12801 19576 12835
rect 19524 12792 19576 12801
rect 19892 12835 19944 12844
rect 19892 12801 19901 12835
rect 19901 12801 19935 12835
rect 19935 12801 19944 12835
rect 19892 12792 19944 12801
rect 20076 12971 20128 12980
rect 20076 12937 20085 12971
rect 20085 12937 20119 12971
rect 20119 12937 20128 12971
rect 20076 12928 20128 12937
rect 23020 12971 23072 12980
rect 23020 12937 23029 12971
rect 23029 12937 23063 12971
rect 23063 12937 23072 12971
rect 23020 12928 23072 12937
rect 23204 12928 23256 12980
rect 20720 12860 20772 12912
rect 23756 12928 23808 12980
rect 24492 12928 24544 12980
rect 26148 12928 26200 12980
rect 31484 12971 31536 12980
rect 31484 12937 31493 12971
rect 31493 12937 31527 12971
rect 31527 12937 31536 12971
rect 31484 12928 31536 12937
rect 23204 12835 23256 12844
rect 23204 12801 23213 12835
rect 23213 12801 23247 12835
rect 23247 12801 23256 12835
rect 23204 12792 23256 12801
rect 23480 12835 23532 12844
rect 23480 12801 23489 12835
rect 23489 12801 23523 12835
rect 23523 12801 23532 12835
rect 23480 12792 23532 12801
rect 23848 12835 23900 12844
rect 23848 12801 23857 12835
rect 23857 12801 23891 12835
rect 23891 12801 23900 12835
rect 23848 12792 23900 12801
rect 23940 12835 23992 12844
rect 23940 12801 23949 12835
rect 23949 12801 23983 12835
rect 23983 12801 23992 12835
rect 23940 12792 23992 12801
rect 19248 12656 19300 12708
rect 29460 12860 29512 12912
rect 29736 12860 29788 12912
rect 30288 12860 30340 12912
rect 31116 12860 31168 12912
rect 25412 12792 25464 12844
rect 25688 12835 25740 12844
rect 25688 12801 25697 12835
rect 25697 12801 25731 12835
rect 25731 12801 25740 12835
rect 25688 12792 25740 12801
rect 25780 12724 25832 12776
rect 30932 12792 30984 12844
rect 26056 12724 26108 12776
rect 31668 12724 31720 12776
rect 18880 12588 18932 12640
rect 20720 12588 20772 12640
rect 23204 12631 23256 12640
rect 23204 12597 23213 12631
rect 23213 12597 23247 12631
rect 23247 12597 23256 12631
rect 25504 12656 25556 12708
rect 23204 12588 23256 12597
rect 24400 12588 24452 12640
rect 31024 12631 31076 12640
rect 31024 12597 31033 12631
rect 31033 12597 31067 12631
rect 31067 12597 31076 12631
rect 31024 12588 31076 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 1584 12427 1636 12436
rect 1584 12393 1593 12427
rect 1593 12393 1627 12427
rect 1627 12393 1636 12427
rect 1584 12384 1636 12393
rect 3056 12384 3108 12436
rect 3976 12384 4028 12436
rect 6276 12384 6328 12436
rect 9772 12384 9824 12436
rect 12256 12384 12308 12436
rect 14372 12427 14424 12436
rect 14372 12393 14381 12427
rect 14381 12393 14415 12427
rect 14415 12393 14424 12427
rect 14372 12384 14424 12393
rect 15016 12384 15068 12436
rect 17592 12384 17644 12436
rect 30288 12384 30340 12436
rect 4804 12316 4856 12368
rect 5724 12316 5776 12368
rect 6368 12316 6420 12368
rect 6552 12248 6604 12300
rect 7748 12291 7800 12300
rect 7748 12257 7757 12291
rect 7757 12257 7791 12291
rect 7791 12257 7800 12291
rect 7748 12248 7800 12257
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 848 12112 900 12164
rect 4068 12180 4120 12232
rect 4712 12155 4764 12164
rect 4712 12121 4721 12155
rect 4721 12121 4755 12155
rect 4755 12121 4764 12155
rect 4712 12112 4764 12121
rect 5448 12180 5500 12232
rect 5908 12223 5960 12232
rect 5908 12189 5917 12223
rect 5917 12189 5951 12223
rect 5951 12189 5960 12223
rect 5908 12180 5960 12189
rect 7288 12180 7340 12232
rect 5724 12155 5776 12164
rect 5448 12087 5500 12096
rect 5448 12053 5457 12087
rect 5457 12053 5491 12087
rect 5491 12053 5500 12087
rect 5448 12044 5500 12053
rect 5724 12121 5742 12155
rect 5742 12121 5776 12155
rect 5724 12112 5776 12121
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 8760 12316 8812 12368
rect 8668 12291 8720 12300
rect 8668 12257 8677 12291
rect 8677 12257 8711 12291
rect 8711 12257 8720 12291
rect 8668 12248 8720 12257
rect 12164 12248 12216 12300
rect 8300 12112 8352 12164
rect 10600 12180 10652 12232
rect 12992 12248 13044 12300
rect 10508 12155 10560 12164
rect 10508 12121 10517 12155
rect 10517 12121 10551 12155
rect 10551 12121 10560 12155
rect 10508 12112 10560 12121
rect 11060 12112 11112 12164
rect 12900 12155 12952 12164
rect 12900 12121 12909 12155
rect 12909 12121 12943 12155
rect 12943 12121 12952 12155
rect 12900 12112 12952 12121
rect 11244 12044 11296 12096
rect 14740 12291 14792 12300
rect 14740 12257 14749 12291
rect 14749 12257 14783 12291
rect 14783 12257 14792 12291
rect 14740 12248 14792 12257
rect 17040 12316 17092 12368
rect 18236 12316 18288 12368
rect 19800 12359 19852 12368
rect 19800 12325 19809 12359
rect 19809 12325 19843 12359
rect 19843 12325 19852 12359
rect 19800 12316 19852 12325
rect 14924 12180 14976 12232
rect 15200 12180 15252 12232
rect 27712 12248 27764 12300
rect 13084 12112 13136 12164
rect 16948 12112 17000 12164
rect 17040 12044 17092 12096
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 17500 12223 17552 12232
rect 17500 12189 17514 12223
rect 17514 12189 17548 12223
rect 17548 12189 17552 12223
rect 17500 12180 17552 12189
rect 17684 12180 17736 12232
rect 19248 12223 19300 12232
rect 19248 12189 19257 12223
rect 19257 12189 19291 12223
rect 19291 12189 19300 12223
rect 19248 12180 19300 12189
rect 19524 12223 19576 12232
rect 17408 12155 17460 12164
rect 17408 12121 17417 12155
rect 17417 12121 17451 12155
rect 17451 12121 17460 12155
rect 19524 12189 19533 12223
rect 19533 12189 19567 12223
rect 19567 12189 19576 12223
rect 19524 12180 19576 12189
rect 19616 12223 19668 12232
rect 19616 12189 19630 12223
rect 19630 12189 19664 12223
rect 19664 12189 19668 12223
rect 19616 12180 19668 12189
rect 17408 12112 17460 12121
rect 19892 12112 19944 12164
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 2780 11840 2832 11892
rect 8300 11840 8352 11892
rect 15752 11840 15804 11892
rect 15844 11840 15896 11892
rect 23848 11840 23900 11892
rect 5448 11772 5500 11824
rect 9956 11772 10008 11824
rect 848 11704 900 11756
rect 10508 11704 10560 11756
rect 13176 11704 13228 11756
rect 17408 11704 17460 11756
rect 7932 11636 7984 11688
rect 15844 11636 15896 11688
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
<< metal2 >>
rect 21914 39200 21970 40000
rect 22558 39200 22614 40000
rect 23202 39200 23258 40000
rect 25134 39200 25190 40000
rect 25778 39200 25834 40000
rect 27710 39200 27766 40000
rect 28998 39200 29054 40000
rect 29642 39200 29698 40000
rect 31574 39200 31630 40000
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 21928 37466 21956 39200
rect 22572 37466 22600 39200
rect 23216 37466 23244 39200
rect 25148 37466 25176 39200
rect 25792 37466 25820 39200
rect 27724 37466 27752 39200
rect 21916 37460 21968 37466
rect 21916 37402 21968 37408
rect 22560 37460 22612 37466
rect 22560 37402 22612 37408
rect 23204 37460 23256 37466
rect 23204 37402 23256 37408
rect 25136 37460 25188 37466
rect 25136 37402 25188 37408
rect 25780 37460 25832 37466
rect 25780 37402 25832 37408
rect 27712 37460 27764 37466
rect 27712 37402 27764 37408
rect 29012 37398 29040 39200
rect 29656 37466 29684 39200
rect 31588 37466 31616 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 29644 37460 29696 37466
rect 29644 37402 29696 37408
rect 31576 37460 31628 37466
rect 31576 37402 31628 37408
rect 29000 37392 29052 37398
rect 29000 37334 29052 37340
rect 22376 37188 22428 37194
rect 22376 37130 22428 37136
rect 23388 37188 23440 37194
rect 23388 37130 23440 37136
rect 23664 37188 23716 37194
rect 23664 37130 23716 37136
rect 25596 37188 25648 37194
rect 25596 37130 25648 37136
rect 27068 37188 27120 37194
rect 27068 37130 27120 37136
rect 28172 37188 28224 37194
rect 28172 37130 28224 37136
rect 29644 37188 29696 37194
rect 29644 37130 29696 37136
rect 30472 37188 30524 37194
rect 30472 37130 30524 37136
rect 32220 37188 32272 37194
rect 32220 37130 32272 37136
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 22388 35698 22416 37130
rect 22376 35692 22428 35698
rect 22376 35634 22428 35640
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 22388 35306 22416 35634
rect 22652 35488 22704 35494
rect 22652 35430 22704 35436
rect 22296 35290 22416 35306
rect 22284 35284 22416 35290
rect 22336 35278 22416 35284
rect 22284 35226 22336 35232
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 14372 34740 14424 34746
rect 14372 34682 14424 34688
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 13728 32768 13780 32774
rect 13728 32710 13780 32716
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 12348 32496 12400 32502
rect 12348 32438 12400 32444
rect 11428 32428 11480 32434
rect 11428 32370 11480 32376
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 11440 32026 11468 32370
rect 11060 32020 11112 32026
rect 11060 31962 11112 31968
rect 11428 32020 11480 32026
rect 11428 31962 11480 31968
rect 9128 31952 9180 31958
rect 9128 31894 9180 31900
rect 7932 31816 7984 31822
rect 7932 31758 7984 31764
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 7840 30320 7892 30326
rect 7840 30262 7892 30268
rect 6552 30048 6604 30054
rect 6552 29990 6604 29996
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 5724 28484 5776 28490
rect 5724 28426 5776 28432
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 5264 28076 5316 28082
rect 5264 28018 5316 28024
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 5172 25900 5224 25906
rect 5172 25842 5224 25848
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 5184 25242 5212 25842
rect 5276 25498 5304 28018
rect 5356 27668 5408 27674
rect 5356 27610 5408 27616
rect 5368 25974 5396 27610
rect 5448 27396 5500 27402
rect 5448 27338 5500 27344
rect 5460 26042 5488 27338
rect 5448 26036 5500 26042
rect 5448 25978 5500 25984
rect 5356 25968 5408 25974
rect 5356 25910 5408 25916
rect 5446 25936 5502 25945
rect 5264 25492 5316 25498
rect 5264 25434 5316 25440
rect 5184 25214 5304 25242
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 2780 24064 2832 24070
rect 2780 24006 2832 24012
rect 2136 23044 2188 23050
rect 2136 22986 2188 22992
rect 2148 20942 2176 22986
rect 2688 21548 2740 21554
rect 2688 21490 2740 21496
rect 2504 21480 2556 21486
rect 2504 21422 2556 21428
rect 2136 20936 2188 20942
rect 2136 20878 2188 20884
rect 2148 18290 2176 20878
rect 2412 19712 2464 19718
rect 2412 19654 2464 19660
rect 2424 19446 2452 19654
rect 2412 19440 2464 19446
rect 2516 19417 2544 21422
rect 2596 20936 2648 20942
rect 2596 20878 2648 20884
rect 2412 19382 2464 19388
rect 2502 19408 2558 19417
rect 2608 19378 2636 20878
rect 2700 20534 2728 21490
rect 2688 20528 2740 20534
rect 2688 20470 2740 20476
rect 2700 19514 2728 20470
rect 2688 19508 2740 19514
rect 2688 19450 2740 19456
rect 2792 19378 2820 24006
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4620 23792 4672 23798
rect 4620 23734 4672 23740
rect 4252 23724 4304 23730
rect 4252 23666 4304 23672
rect 4436 23724 4488 23730
rect 4436 23666 4488 23672
rect 3424 23656 3476 23662
rect 4264 23610 4292 23666
rect 3424 23598 3476 23604
rect 3436 23254 3464 23598
rect 4080 23582 4292 23610
rect 4448 23594 4476 23666
rect 4436 23588 4488 23594
rect 3056 23248 3108 23254
rect 3056 23190 3108 23196
rect 3424 23248 3476 23254
rect 3424 23190 3476 23196
rect 3068 21010 3096 23190
rect 3792 23180 3844 23186
rect 3792 23122 3844 23128
rect 3804 22574 3832 23122
rect 4080 22982 4108 23582
rect 4436 23530 4488 23536
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23254 4660 23734
rect 4804 23588 4856 23594
rect 4804 23530 4856 23536
rect 4620 23248 4672 23254
rect 4620 23190 4672 23196
rect 4344 23112 4396 23118
rect 4344 23054 4396 23060
rect 4712 23112 4764 23118
rect 4712 23054 4764 23060
rect 4068 22976 4120 22982
rect 4068 22918 4120 22924
rect 4356 22681 4384 23054
rect 4342 22672 4398 22681
rect 4342 22607 4398 22616
rect 3792 22568 3844 22574
rect 3792 22510 3844 22516
rect 3056 21004 3108 21010
rect 3056 20946 3108 20952
rect 2502 19343 2558 19352
rect 2596 19372 2648 19378
rect 2516 19310 2544 19343
rect 2596 19314 2648 19320
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2504 19304 2556 19310
rect 2504 19246 2556 19252
rect 2516 18970 2544 19246
rect 2504 18964 2556 18970
rect 2504 18906 2556 18912
rect 2412 18692 2464 18698
rect 2412 18634 2464 18640
rect 2136 18284 2188 18290
rect 2136 18226 2188 18232
rect 2424 17882 2452 18634
rect 2504 18284 2556 18290
rect 2504 18226 2556 18232
rect 2516 17882 2544 18226
rect 2608 18222 2636 19314
rect 2872 18896 2924 18902
rect 2872 18838 2924 18844
rect 2884 18290 2912 18838
rect 2872 18284 2924 18290
rect 2872 18226 2924 18232
rect 3068 18222 3096 20946
rect 3240 20936 3292 20942
rect 3240 20878 3292 20884
rect 3252 19786 3280 20878
rect 3332 20460 3384 20466
rect 3332 20402 3384 20408
rect 3344 19854 3372 20402
rect 3424 20392 3476 20398
rect 3424 20334 3476 20340
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 3240 19780 3292 19786
rect 3240 19722 3292 19728
rect 3148 19372 3200 19378
rect 3252 19360 3280 19722
rect 3252 19332 3372 19360
rect 3148 19314 3200 19320
rect 2596 18216 2648 18222
rect 2596 18158 2648 18164
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 3068 17882 3096 18158
rect 2412 17876 2464 17882
rect 2412 17818 2464 17824
rect 2504 17876 2556 17882
rect 2504 17818 2556 17824
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2228 17196 2280 17202
rect 2228 17138 2280 17144
rect 2136 16720 2188 16726
rect 2136 16662 2188 16668
rect 848 16584 900 16590
rect 846 16552 848 16561
rect 900 16552 902 16561
rect 846 16487 902 16496
rect 1768 16516 1820 16522
rect 1768 16458 1820 16464
rect 1780 16114 1808 16458
rect 848 16108 900 16114
rect 848 16050 900 16056
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 860 15881 888 16050
rect 2148 16028 2176 16662
rect 2240 16250 2268 17138
rect 2320 16992 2372 16998
rect 2320 16934 2372 16940
rect 2332 16658 2360 16934
rect 2320 16652 2372 16658
rect 2320 16594 2372 16600
rect 2228 16244 2280 16250
rect 2228 16186 2280 16192
rect 2332 16114 2360 16594
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2228 16040 2280 16046
rect 2148 16000 2228 16028
rect 2228 15982 2280 15988
rect 846 15872 902 15881
rect 846 15807 902 15816
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15065 1440 15438
rect 2240 15366 2268 15982
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2228 15360 2280 15366
rect 2228 15302 2280 15308
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 2424 14618 2452 15438
rect 2608 15162 2636 17614
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2792 15706 2820 16050
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2596 15156 2648 15162
rect 2596 15098 2648 15104
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 846 14512 902 14521
rect 846 14447 902 14456
rect 860 14414 888 14447
rect 848 14408 900 14414
rect 848 14350 900 14356
rect 2320 14340 2372 14346
rect 2320 14282 2372 14288
rect 2332 14074 2360 14282
rect 2516 14074 2544 14962
rect 2700 14958 2728 15438
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2792 14958 2820 15302
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2792 14074 2820 14214
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 2504 14068 2556 14074
rect 2504 14010 2556 14016
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2688 14000 2740 14006
rect 2688 13942 2740 13948
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 1584 13728 1636 13734
rect 1398 13696 1454 13705
rect 1584 13670 1636 13676
rect 1398 13631 1454 13640
rect 1596 13394 1624 13670
rect 2056 13394 2084 13806
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 1398 13016 1454 13025
rect 1596 13002 1624 13330
rect 2148 13190 2176 13806
rect 2700 13394 2728 13942
rect 2792 13802 2820 14010
rect 2780 13796 2832 13802
rect 2780 13738 2832 13744
rect 2792 13462 2820 13738
rect 2884 13530 2912 17614
rect 2964 16516 3016 16522
rect 2964 16458 3016 16464
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 2976 16182 3004 16458
rect 2964 16176 3016 16182
rect 2964 16118 3016 16124
rect 2976 15638 3004 16118
rect 3068 15910 3096 16458
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 2964 15632 3016 15638
rect 2964 15574 3016 15580
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2780 13456 2832 13462
rect 2832 13404 2912 13410
rect 2780 13398 2912 13404
rect 2688 13388 2740 13394
rect 2792 13382 2912 13398
rect 2688 13330 2740 13336
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2596 13184 2648 13190
rect 2596 13126 2648 13132
rect 1596 12986 1716 13002
rect 1398 12951 1454 12960
rect 1584 12980 1716 12986
rect 1412 12238 1440 12951
rect 1636 12974 1716 12980
rect 1584 12922 1636 12928
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1596 12442 1624 12786
rect 1688 12782 1716 12974
rect 2504 12912 2556 12918
rect 2608 12866 2636 13126
rect 2700 12986 2728 13330
rect 2884 13326 2912 13382
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2556 12860 2636 12866
rect 2504 12854 2636 12860
rect 2516 12838 2636 12854
rect 2608 12782 2636 12838
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 2504 12776 2556 12782
rect 2504 12718 2556 12724
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2516 12646 2544 12718
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1400 12232 1452 12238
rect 846 12200 902 12209
rect 1400 12174 1452 12180
rect 846 12135 848 12144
rect 900 12135 902 12144
rect 848 12106 900 12112
rect 2792 11898 2820 13194
rect 2884 12714 2912 13262
rect 2976 12850 3004 13806
rect 3160 13297 3188 19314
rect 3240 18760 3292 18766
rect 3240 18702 3292 18708
rect 3252 17610 3280 18702
rect 3344 18698 3372 19332
rect 3436 18970 3464 20334
rect 3608 19236 3660 19242
rect 3608 19178 3660 19184
rect 3424 18964 3476 18970
rect 3424 18906 3476 18912
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3332 18692 3384 18698
rect 3332 18634 3384 18640
rect 3436 18290 3464 18702
rect 3620 18426 3648 19178
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3240 17604 3292 17610
rect 3240 17546 3292 17552
rect 3252 16794 3280 17546
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 3240 16448 3292 16454
rect 3240 16390 3292 16396
rect 3252 15366 3280 16390
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3252 15162 3280 15302
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 3240 13932 3292 13938
rect 3240 13874 3292 13880
rect 3146 13288 3202 13297
rect 3146 13223 3202 13232
rect 3160 13190 3188 13223
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3252 12850 3280 13874
rect 3344 12986 3372 17614
rect 3436 16046 3464 18226
rect 3804 17338 3832 22510
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3976 21616 4028 21622
rect 3976 21558 4028 21564
rect 3988 21146 4016 21558
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 3976 21140 4028 21146
rect 3976 21082 4028 21088
rect 4620 21140 4672 21146
rect 4620 21082 4672 21088
rect 3884 20936 3936 20942
rect 3884 20878 3936 20884
rect 3896 19922 3924 20878
rect 3988 20874 4016 21082
rect 4160 20936 4212 20942
rect 4160 20878 4212 20884
rect 3976 20868 4028 20874
rect 3976 20810 4028 20816
rect 4172 20466 4200 20878
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3884 19916 3936 19922
rect 3884 19858 3936 19864
rect 3896 18766 3924 19858
rect 4632 19786 4660 21082
rect 4068 19780 4120 19786
rect 4068 19722 4120 19728
rect 4620 19780 4672 19786
rect 4620 19722 4672 19728
rect 4080 18902 4108 19722
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4632 18970 4660 19110
rect 4620 18964 4672 18970
rect 4620 18906 4672 18912
rect 4068 18896 4120 18902
rect 4724 18850 4752 23054
rect 4816 23050 4844 23530
rect 5276 23254 5304 25214
rect 5368 23526 5396 25910
rect 5446 25871 5448 25880
rect 5500 25871 5502 25880
rect 5448 25842 5500 25848
rect 5736 25498 5764 28426
rect 6092 28008 6144 28014
rect 6092 27950 6144 27956
rect 6000 27464 6052 27470
rect 6000 27406 6052 27412
rect 6012 27130 6040 27406
rect 6000 27124 6052 27130
rect 6000 27066 6052 27072
rect 5724 25492 5776 25498
rect 5724 25434 5776 25440
rect 6104 25401 6132 27950
rect 6090 25392 6146 25401
rect 5632 25356 5684 25362
rect 6090 25327 6146 25336
rect 5632 25298 5684 25304
rect 5644 24954 5672 25298
rect 5908 25152 5960 25158
rect 5908 25094 5960 25100
rect 5632 24948 5684 24954
rect 5632 24890 5684 24896
rect 5448 24336 5500 24342
rect 5448 24278 5500 24284
rect 5356 23520 5408 23526
rect 5356 23462 5408 23468
rect 5460 23322 5488 24278
rect 5538 23760 5594 23769
rect 5538 23695 5594 23704
rect 5448 23316 5500 23322
rect 5448 23258 5500 23264
rect 5264 23248 5316 23254
rect 5264 23190 5316 23196
rect 5264 23112 5316 23118
rect 5264 23054 5316 23060
rect 4804 23044 4856 23050
rect 4804 22986 4856 22992
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5276 22778 5304 23054
rect 5448 23044 5500 23050
rect 5448 22986 5500 22992
rect 5264 22772 5316 22778
rect 5264 22714 5316 22720
rect 5170 22672 5226 22681
rect 4804 22636 4856 22642
rect 5460 22642 5488 22986
rect 5448 22636 5500 22642
rect 5170 22607 5172 22616
rect 4804 22578 4856 22584
rect 5224 22607 5226 22616
rect 5172 22578 5224 22584
rect 5368 22596 5448 22624
rect 4816 19854 4844 22578
rect 5080 22432 5132 22438
rect 5078 22400 5080 22409
rect 5132 22400 5134 22409
rect 5078 22335 5134 22344
rect 5092 22030 5120 22335
rect 5080 22024 5132 22030
rect 5080 21966 5132 21972
rect 5264 22024 5316 22030
rect 5264 21966 5316 21972
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5276 21593 5304 21966
rect 5262 21584 5318 21593
rect 5262 21519 5318 21528
rect 4896 21480 4948 21486
rect 4896 21422 4948 21428
rect 4908 20942 4936 21422
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 5264 20936 5316 20942
rect 5264 20878 5316 20884
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 5276 19854 5304 20878
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5368 19786 5396 22596
rect 5448 22578 5500 22584
rect 5552 21894 5580 23695
rect 5632 23248 5684 23254
rect 5632 23190 5684 23196
rect 5644 22710 5672 23190
rect 5632 22704 5684 22710
rect 5632 22646 5684 22652
rect 5814 22672 5870 22681
rect 5644 22506 5672 22646
rect 5814 22607 5816 22616
rect 5868 22607 5870 22616
rect 5816 22578 5868 22584
rect 5632 22500 5684 22506
rect 5632 22442 5684 22448
rect 5724 22228 5776 22234
rect 5724 22170 5776 22176
rect 5540 21888 5592 21894
rect 5540 21830 5592 21836
rect 5446 21584 5502 21593
rect 5446 21519 5502 21528
rect 5632 21548 5684 21554
rect 5356 19780 5408 19786
rect 5356 19722 5408 19728
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5460 19224 5488 21519
rect 5632 21490 5684 21496
rect 5644 21350 5672 21490
rect 5632 21344 5684 21350
rect 5632 21286 5684 21292
rect 5632 20936 5684 20942
rect 5632 20878 5684 20884
rect 5460 19196 5580 19224
rect 5446 19136 5502 19145
rect 5446 19071 5502 19080
rect 4068 18838 4120 18844
rect 3884 18760 3936 18766
rect 3884 18702 3936 18708
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 3608 17196 3660 17202
rect 3608 17138 3660 17144
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3528 16454 3556 16526
rect 3516 16448 3568 16454
rect 3516 16390 3568 16396
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 3424 15904 3476 15910
rect 3476 15864 3556 15892
rect 3424 15846 3476 15852
rect 3528 15366 3556 15864
rect 3516 15360 3568 15366
rect 3516 15302 3568 15308
rect 3528 15026 3556 15302
rect 3620 15094 3648 17138
rect 3700 17060 3752 17066
rect 3700 17002 3752 17008
rect 3712 16794 3740 17002
rect 3896 16998 3924 18702
rect 3988 18086 4016 18702
rect 3976 18080 4028 18086
rect 3976 18022 4028 18028
rect 3976 17332 4028 17338
rect 3976 17274 4028 17280
rect 3884 16992 3936 16998
rect 3804 16952 3884 16980
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3698 16688 3754 16697
rect 3698 16623 3754 16632
rect 3712 16046 3740 16623
rect 3804 16046 3832 16952
rect 3884 16934 3936 16940
rect 3988 16810 4016 17274
rect 3896 16782 4016 16810
rect 3896 16114 3924 16782
rect 3976 16720 4028 16726
rect 3976 16662 4028 16668
rect 3988 16590 4016 16662
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 3700 16040 3752 16046
rect 3700 15982 3752 15988
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3988 15638 4016 16526
rect 4080 16454 4108 18838
rect 4632 18822 4752 18850
rect 5184 18822 5396 18850
rect 4632 18465 4660 18822
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4712 18692 4764 18698
rect 4712 18634 4764 18640
rect 4618 18456 4674 18465
rect 4618 18391 4674 18400
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17678 4660 18226
rect 4724 17762 4752 18634
rect 4816 18426 4844 18702
rect 5080 18692 5132 18698
rect 5184 18680 5212 18822
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 5132 18652 5212 18680
rect 5080 18634 5132 18640
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4816 17882 4844 18362
rect 4894 18320 4950 18329
rect 4894 18255 4950 18264
rect 5172 18284 5224 18290
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4724 17734 4844 17762
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16794 4660 17614
rect 4724 17270 4752 17614
rect 4712 17264 4764 17270
rect 4712 17206 4764 17212
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4160 16720 4212 16726
rect 4160 16662 4212 16668
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4172 15892 4200 16662
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4080 15864 4200 15892
rect 3976 15632 4028 15638
rect 3976 15574 4028 15580
rect 3608 15088 3660 15094
rect 3608 15030 3660 15036
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3988 14822 4016 15574
rect 4080 15502 4108 15864
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3988 14346 4016 14758
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3976 14340 4028 14346
rect 3976 14282 4028 14288
rect 4632 14074 4660 16050
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2976 12434 3004 12786
rect 3988 12646 4016 13194
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3988 12442 4016 12582
rect 3056 12436 3108 12442
rect 2976 12406 3056 12434
rect 3056 12378 3108 12384
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 4080 12238 4108 13398
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 4356 12782 4384 13194
rect 4540 13190 4568 13330
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4540 12646 4568 13126
rect 4632 12714 4660 13670
rect 4724 13530 4752 17070
rect 4816 15910 4844 17734
rect 4908 17678 4936 18255
rect 5276 18272 5304 18702
rect 5224 18244 5304 18272
rect 5172 18226 5224 18232
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 4988 17264 5040 17270
rect 4986 17232 4988 17241
rect 5040 17232 5042 17241
rect 4986 17167 5042 17176
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4908 16697 4936 16934
rect 4894 16688 4950 16697
rect 4894 16623 4950 16632
rect 5000 16590 5028 17167
rect 5080 17128 5132 17134
rect 5080 17070 5132 17076
rect 5092 16726 5120 17070
rect 5080 16720 5132 16726
rect 5080 16662 5132 16668
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 5184 16538 5212 17274
rect 5276 16726 5304 18244
rect 5368 16998 5396 18822
rect 5460 18154 5488 19071
rect 5448 18148 5500 18154
rect 5448 18090 5500 18096
rect 5552 18034 5580 19196
rect 5460 18006 5580 18034
rect 5460 17338 5488 18006
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5460 16726 5488 17138
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 5264 16720 5316 16726
rect 5264 16662 5316 16668
rect 5448 16720 5500 16726
rect 5448 16662 5500 16668
rect 5356 16584 5408 16590
rect 5184 16510 5304 16538
rect 5356 16526 5408 16532
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5276 16182 5304 16510
rect 5264 16176 5316 16182
rect 5264 16118 5316 16124
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4816 14074 4844 14214
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4816 13870 4844 14010
rect 5264 14000 5316 14006
rect 5264 13942 5316 13948
rect 5368 13954 5396 16526
rect 5460 15638 5488 16662
rect 5552 16590 5580 17002
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5540 16448 5592 16454
rect 5644 16402 5672 20878
rect 5736 20466 5764 22170
rect 5828 22166 5856 22578
rect 5816 22160 5868 22166
rect 5816 22102 5868 22108
rect 5920 22030 5948 25094
rect 6000 24812 6052 24818
rect 6000 24754 6052 24760
rect 6012 22506 6040 24754
rect 6000 22500 6052 22506
rect 6000 22442 6052 22448
rect 5908 22024 5960 22030
rect 5908 21966 5960 21972
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 5908 21548 5960 21554
rect 5960 21508 6040 21536
rect 5908 21490 5960 21496
rect 5828 21146 5856 21490
rect 5816 21140 5868 21146
rect 5816 21082 5868 21088
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5908 20460 5960 20466
rect 5908 20402 5960 20408
rect 5736 19990 5764 20402
rect 5920 20058 5948 20402
rect 6012 20398 6040 21508
rect 6104 20602 6132 25327
rect 6184 24812 6236 24818
rect 6184 24754 6236 24760
rect 6092 20596 6144 20602
rect 6092 20538 6144 20544
rect 6000 20392 6052 20398
rect 6000 20334 6052 20340
rect 6000 20256 6052 20262
rect 5998 20224 6000 20233
rect 6052 20224 6054 20233
rect 5998 20159 6054 20168
rect 5908 20052 5960 20058
rect 5908 19994 5960 20000
rect 5724 19984 5776 19990
rect 5724 19926 5776 19932
rect 5736 19689 5764 19926
rect 5722 19680 5778 19689
rect 5722 19615 5778 19624
rect 6012 19242 6040 20159
rect 6196 19530 6224 24754
rect 6276 23792 6328 23798
rect 6276 23734 6328 23740
rect 6104 19502 6224 19530
rect 6104 19242 6132 19502
rect 6184 19440 6236 19446
rect 6184 19382 6236 19388
rect 6000 19236 6052 19242
rect 6000 19178 6052 19184
rect 6092 19236 6144 19242
rect 6092 19178 6144 19184
rect 6196 18834 6224 19382
rect 6288 18970 6316 23734
rect 6460 22092 6512 22098
rect 6460 22034 6512 22040
rect 6368 21548 6420 21554
rect 6368 21490 6420 21496
rect 6380 21350 6408 21490
rect 6368 21344 6420 21350
rect 6368 21286 6420 21292
rect 6472 20942 6500 22034
rect 6460 20936 6512 20942
rect 6460 20878 6512 20884
rect 6564 20262 6592 29990
rect 7654 29472 7710 29481
rect 7654 29407 7710 29416
rect 7668 29306 7696 29407
rect 7656 29300 7708 29306
rect 7656 29242 7708 29248
rect 6920 29164 6972 29170
rect 6920 29106 6972 29112
rect 6736 28008 6788 28014
rect 6736 27950 6788 27956
rect 6826 27976 6882 27985
rect 6748 27713 6776 27950
rect 6826 27911 6828 27920
rect 6880 27911 6882 27920
rect 6828 27882 6880 27888
rect 6734 27704 6790 27713
rect 6734 27639 6736 27648
rect 6788 27639 6790 27648
rect 6736 27610 6788 27616
rect 6828 27532 6880 27538
rect 6828 27474 6880 27480
rect 6840 26994 6868 27474
rect 6932 27334 6960 29106
rect 7380 29096 7432 29102
rect 7380 29038 7432 29044
rect 7196 28960 7248 28966
rect 7196 28902 7248 28908
rect 7012 28076 7064 28082
rect 7012 28018 7064 28024
rect 6920 27328 6972 27334
rect 6920 27270 6972 27276
rect 6828 26988 6880 26994
rect 6828 26930 6880 26936
rect 6840 26314 6868 26930
rect 6932 26489 6960 27270
rect 6918 26480 6974 26489
rect 6918 26415 6974 26424
rect 6828 26308 6880 26314
rect 6828 26250 6880 26256
rect 6840 24818 6868 26250
rect 6828 24812 6880 24818
rect 6828 24754 6880 24760
rect 6840 23322 6868 24754
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6644 23112 6696 23118
rect 6644 23054 6696 23060
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 6656 20040 6684 23054
rect 6736 23044 6788 23050
rect 6736 22986 6788 22992
rect 6380 20012 6684 20040
rect 6380 19854 6408 20012
rect 6748 19922 6776 22986
rect 7024 22094 7052 28018
rect 7208 27878 7236 28902
rect 7196 27872 7248 27878
rect 7196 27814 7248 27820
rect 7196 26852 7248 26858
rect 7196 26794 7248 26800
rect 7104 25900 7156 25906
rect 7104 25842 7156 25848
rect 6840 22066 7052 22094
rect 6840 21026 6868 22066
rect 6920 21956 6972 21962
rect 6920 21898 6972 21904
rect 7012 21956 7064 21962
rect 7012 21898 7064 21904
rect 6932 21690 6960 21898
rect 6920 21684 6972 21690
rect 6920 21626 6972 21632
rect 7024 21185 7052 21898
rect 7010 21176 7066 21185
rect 7010 21111 7066 21120
rect 6840 20998 7052 21026
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 6736 19916 6788 19922
rect 6736 19858 6788 19864
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6276 18964 6328 18970
rect 6276 18906 6328 18912
rect 6380 18902 6408 19790
rect 6552 19780 6604 19786
rect 6552 19722 6604 19728
rect 6564 19378 6592 19722
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 6552 19372 6604 19378
rect 6656 19360 6684 19858
rect 6748 19496 6776 19858
rect 6748 19468 6868 19496
rect 6736 19372 6788 19378
rect 6656 19332 6736 19360
rect 6552 19314 6604 19320
rect 6736 19314 6788 19320
rect 6368 18896 6420 18902
rect 6368 18838 6420 18844
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 5816 18692 5868 18698
rect 5816 18634 5868 18640
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5592 16396 5672 16402
rect 5540 16390 5672 16396
rect 5552 16374 5672 16390
rect 5448 15632 5500 15638
rect 5552 15609 5580 16374
rect 5736 15706 5764 18226
rect 5828 18222 5856 18634
rect 5908 18624 5960 18630
rect 5908 18566 5960 18572
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 5920 18358 5948 18566
rect 5908 18352 5960 18358
rect 5908 18294 5960 18300
rect 5816 18216 5868 18222
rect 5816 18158 5868 18164
rect 5920 17610 5948 18294
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 5908 17604 5960 17610
rect 5908 17546 5960 17552
rect 5920 16590 5948 17546
rect 6012 16726 6040 17614
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 5908 16584 5960 16590
rect 5908 16526 5960 16532
rect 5908 16448 5960 16454
rect 6104 16402 6132 18566
rect 6196 17678 6224 18770
rect 6276 18760 6328 18766
rect 6276 18702 6328 18708
rect 6288 17882 6316 18702
rect 6380 18290 6408 18838
rect 6472 18766 6500 19314
rect 6644 19236 6696 19242
rect 6644 19178 6696 19184
rect 6552 18896 6604 18902
rect 6552 18838 6604 18844
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6380 18086 6408 18226
rect 6368 18080 6420 18086
rect 6368 18022 6420 18028
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6288 17066 6316 17818
rect 6472 17678 6500 18702
rect 6564 17814 6592 18838
rect 6552 17808 6604 17814
rect 6552 17750 6604 17756
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6368 17604 6420 17610
rect 6368 17546 6420 17552
rect 6276 17060 6328 17066
rect 6276 17002 6328 17008
rect 6184 16720 6236 16726
rect 6184 16662 6236 16668
rect 5960 16396 6132 16402
rect 5908 16390 6132 16396
rect 5920 16374 6132 16390
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5448 15574 5500 15580
rect 5538 15600 5594 15609
rect 5538 15535 5594 15544
rect 5632 15428 5684 15434
rect 5632 15370 5684 15376
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4816 13410 4844 13806
rect 4908 13530 4936 13806
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 5080 13456 5132 13462
rect 4724 13382 4844 13410
rect 5078 13424 5080 13433
rect 5132 13424 5134 13433
rect 4724 12714 4752 13382
rect 5078 13359 5134 13368
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4816 12986 4844 13262
rect 5276 13258 5304 13942
rect 5368 13926 5580 13954
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5356 13796 5408 13802
rect 5356 13738 5408 13744
rect 5368 13530 5396 13738
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 5276 12850 5304 13194
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5368 12918 5396 13126
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4528 12640 4580 12646
rect 4528 12582 4580 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 5368 12434 5396 12854
rect 5460 12782 5488 13806
rect 5552 12986 5580 13926
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5644 12714 5672 15370
rect 5828 14074 5856 16050
rect 5920 15706 5948 16374
rect 6000 16176 6052 16182
rect 6000 16118 6052 16124
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 5920 15502 5948 15642
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5908 15360 5960 15366
rect 5908 15302 5960 15308
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5736 13530 5764 14010
rect 5920 13938 5948 15302
rect 6012 14362 6040 16118
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 6104 14482 6132 14758
rect 6196 14657 6224 16662
rect 6288 15570 6316 17002
rect 6380 16250 6408 17546
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 6472 16454 6500 16526
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6380 16114 6408 16186
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 6276 15428 6328 15434
rect 6276 15370 6328 15376
rect 6288 14822 6316 15370
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 6182 14648 6238 14657
rect 6182 14583 6238 14592
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 6012 14334 6132 14362
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 6104 13870 6132 14334
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5828 13462 5856 13806
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5908 13456 5960 13462
rect 5908 13398 5960 13404
rect 5920 13258 5948 13398
rect 6012 13394 6040 13670
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 5908 13252 5960 13258
rect 5908 13194 5960 13200
rect 6104 13190 6132 13806
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5368 12406 5488 12434
rect 4804 12368 4856 12374
rect 4724 12316 4804 12322
rect 4724 12310 4856 12316
rect 4724 12294 4844 12310
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4724 12170 4752 12294
rect 5460 12238 5488 12406
rect 5736 12374 5764 12786
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5736 12170 5764 12310
rect 5920 12238 5948 12718
rect 6196 12434 6224 14583
rect 6276 12436 6328 12442
rect 6196 12406 6276 12434
rect 6276 12378 6328 12384
rect 6380 12374 6408 15846
rect 6564 15552 6592 17750
rect 6656 17513 6684 19178
rect 6748 17678 6776 19314
rect 6840 18426 6868 19468
rect 7024 18601 7052 20998
rect 7116 18834 7144 25842
rect 7208 23866 7236 26794
rect 7288 24268 7340 24274
rect 7288 24210 7340 24216
rect 7196 23860 7248 23866
rect 7196 23802 7248 23808
rect 7300 23662 7328 24210
rect 7392 23866 7420 29038
rect 7564 28144 7616 28150
rect 7564 28086 7616 28092
rect 7576 27674 7604 28086
rect 7564 27668 7616 27674
rect 7564 27610 7616 27616
rect 7472 24200 7524 24206
rect 7472 24142 7524 24148
rect 7484 23866 7512 24142
rect 7380 23860 7432 23866
rect 7380 23802 7432 23808
rect 7472 23860 7524 23866
rect 7472 23802 7524 23808
rect 7288 23656 7340 23662
rect 7288 23598 7340 23604
rect 7196 23520 7248 23526
rect 7196 23462 7248 23468
rect 7208 21146 7236 23462
rect 7300 21894 7328 23598
rect 7472 23520 7524 23526
rect 7472 23462 7524 23468
rect 7380 22228 7432 22234
rect 7380 22170 7432 22176
rect 7392 21962 7420 22170
rect 7484 22094 7512 23462
rect 7576 23254 7604 27610
rect 7748 26784 7800 26790
rect 7748 26726 7800 26732
rect 7760 25906 7788 26726
rect 7852 25906 7880 30262
rect 7944 27606 7972 31758
rect 9140 29850 9168 31894
rect 10968 31816 11020 31822
rect 10968 31758 11020 31764
rect 10324 31136 10376 31142
rect 10324 31078 10376 31084
rect 9772 30252 9824 30258
rect 9772 30194 9824 30200
rect 9784 30122 9812 30194
rect 10046 30152 10102 30161
rect 9772 30116 9824 30122
rect 10046 30087 10102 30096
rect 9772 30058 9824 30064
rect 9680 30048 9732 30054
rect 9680 29990 9732 29996
rect 9128 29844 9180 29850
rect 9128 29786 9180 29792
rect 8944 29232 8996 29238
rect 8944 29174 8996 29180
rect 8956 28762 8984 29174
rect 8944 28756 8996 28762
rect 8944 28698 8996 28704
rect 8024 28688 8076 28694
rect 8024 28630 8076 28636
rect 8036 28082 8064 28630
rect 9140 28558 9168 29786
rect 9312 29708 9364 29714
rect 9312 29650 9364 29656
rect 9324 29306 9352 29650
rect 9312 29300 9364 29306
rect 9312 29242 9364 29248
rect 9324 28762 9352 29242
rect 9692 28966 9720 29990
rect 9680 28960 9732 28966
rect 9680 28902 9732 28908
rect 9692 28762 9720 28902
rect 9312 28756 9364 28762
rect 9312 28698 9364 28704
rect 9680 28756 9732 28762
rect 9680 28698 9732 28704
rect 9128 28552 9180 28558
rect 9128 28494 9180 28500
rect 8024 28076 8076 28082
rect 8024 28018 8076 28024
rect 7932 27600 7984 27606
rect 7932 27542 7984 27548
rect 7944 26382 7972 27542
rect 8208 27464 8260 27470
rect 8114 27432 8170 27441
rect 8208 27406 8260 27412
rect 8760 27464 8812 27470
rect 8760 27406 8812 27412
rect 8114 27367 8170 27376
rect 7932 26376 7984 26382
rect 7932 26318 7984 26324
rect 7944 25922 7972 26318
rect 7748 25900 7800 25906
rect 7748 25842 7800 25848
rect 7840 25900 7892 25906
rect 7944 25894 8064 25922
rect 7840 25842 7892 25848
rect 7656 25832 7708 25838
rect 7656 25774 7708 25780
rect 7932 25832 7984 25838
rect 7932 25774 7984 25780
rect 7668 23526 7696 25774
rect 7944 24993 7972 25774
rect 7930 24984 7986 24993
rect 7930 24919 7986 24928
rect 8036 24750 8064 25894
rect 8024 24744 8076 24750
rect 8024 24686 8076 24692
rect 7748 24132 7800 24138
rect 7748 24074 7800 24080
rect 7760 23662 7788 24074
rect 8128 24070 8156 27367
rect 8220 26994 8248 27406
rect 8772 27130 8800 27406
rect 8760 27124 8812 27130
rect 8760 27066 8812 27072
rect 8484 27056 8536 27062
rect 8484 26998 8536 27004
rect 8208 26988 8260 26994
rect 8208 26930 8260 26936
rect 8220 26874 8248 26930
rect 8392 26920 8444 26926
rect 8390 26888 8392 26897
rect 8444 26888 8446 26897
rect 8220 26846 8340 26874
rect 8208 25696 8260 25702
rect 8206 25664 8208 25673
rect 8260 25664 8262 25673
rect 8206 25599 8262 25608
rect 8312 24614 8340 26846
rect 8390 26823 8446 26832
rect 8300 24608 8352 24614
rect 8300 24550 8352 24556
rect 8116 24064 8168 24070
rect 8116 24006 8168 24012
rect 8022 23896 8078 23905
rect 8022 23831 8078 23840
rect 7932 23724 7984 23730
rect 7932 23666 7984 23672
rect 7748 23656 7800 23662
rect 7944 23633 7972 23666
rect 7748 23598 7800 23604
rect 7930 23624 7986 23633
rect 7656 23520 7708 23526
rect 7656 23462 7708 23468
rect 7760 23338 7788 23598
rect 8036 23594 8064 23831
rect 7930 23559 7986 23568
rect 8024 23588 8076 23594
rect 8024 23530 8076 23536
rect 8116 23588 8168 23594
rect 8116 23530 8168 23536
rect 7840 23520 7892 23526
rect 7838 23488 7840 23497
rect 7892 23488 7894 23497
rect 7838 23423 7894 23432
rect 7668 23310 7788 23338
rect 7564 23248 7616 23254
rect 7564 23190 7616 23196
rect 7484 22066 7604 22094
rect 7470 21992 7526 22001
rect 7380 21956 7432 21962
rect 7470 21927 7526 21936
rect 7380 21898 7432 21904
rect 7288 21888 7340 21894
rect 7288 21830 7340 21836
rect 7196 21140 7248 21146
rect 7196 21082 7248 21088
rect 7300 20874 7328 21830
rect 7392 21690 7420 21898
rect 7380 21684 7432 21690
rect 7380 21626 7432 21632
rect 7484 21570 7512 21927
rect 7392 21542 7512 21570
rect 7288 20868 7340 20874
rect 7288 20810 7340 20816
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 7104 18828 7156 18834
rect 7104 18770 7156 18776
rect 7102 18728 7158 18737
rect 7102 18663 7158 18672
rect 7010 18592 7066 18601
rect 7010 18527 7066 18536
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 6840 18290 6868 18362
rect 6828 18284 6880 18290
rect 6828 18226 6880 18232
rect 6840 18154 6868 18226
rect 7024 18154 7052 18527
rect 6828 18148 6880 18154
rect 6828 18090 6880 18096
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 6920 17808 6972 17814
rect 6918 17776 6920 17785
rect 6972 17776 6974 17785
rect 6918 17711 6974 17720
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 6642 17504 6698 17513
rect 6642 17439 6698 17448
rect 6656 16250 6684 17439
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6748 16182 6776 17614
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6736 16176 6788 16182
rect 6736 16118 6788 16124
rect 6642 16008 6698 16017
rect 6642 15943 6698 15952
rect 6656 15706 6684 15943
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6644 15564 6696 15570
rect 6564 15524 6644 15552
rect 6644 15506 6696 15512
rect 6736 15496 6788 15502
rect 6734 15464 6736 15473
rect 6788 15464 6790 15473
rect 6734 15399 6790 15408
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 6748 14278 6776 15302
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 6564 13326 6592 13466
rect 6656 13394 6684 13738
rect 6840 13546 6868 17138
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6932 16046 6960 16186
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 7116 15638 7144 18663
rect 7208 17542 7236 18906
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7300 17542 7328 17818
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7288 17536 7340 17542
rect 7288 17478 7340 17484
rect 7208 15706 7236 17478
rect 7300 16697 7328 17478
rect 7286 16688 7342 16697
rect 7286 16623 7342 16632
rect 7300 16114 7328 16623
rect 7392 16590 7420 21542
rect 7470 21448 7526 21457
rect 7470 21383 7526 21392
rect 7484 19922 7512 21383
rect 7576 20466 7604 22066
rect 7564 20460 7616 20466
rect 7564 20402 7616 20408
rect 7472 19916 7524 19922
rect 7472 19858 7524 19864
rect 7472 19780 7524 19786
rect 7472 19722 7524 19728
rect 7484 16726 7512 19722
rect 7564 18760 7616 18766
rect 7668 18737 7696 23310
rect 7930 23080 7986 23089
rect 7930 23015 7986 23024
rect 7748 22228 7800 22234
rect 7748 22170 7800 22176
rect 7564 18702 7616 18708
rect 7654 18728 7710 18737
rect 7576 18290 7604 18702
rect 7654 18663 7710 18672
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7760 17882 7788 22170
rect 7944 22098 7972 23015
rect 8128 22710 8156 23530
rect 8300 23248 8352 23254
rect 8300 23190 8352 23196
rect 8312 23118 8340 23190
rect 8300 23112 8352 23118
rect 8300 23054 8352 23060
rect 8116 22704 8168 22710
rect 8116 22646 8168 22652
rect 8208 22568 8260 22574
rect 8208 22510 8260 22516
rect 7932 22092 7984 22098
rect 7932 22034 7984 22040
rect 8220 21962 8248 22510
rect 8208 21956 8260 21962
rect 8208 21898 8260 21904
rect 7840 21684 7892 21690
rect 7840 21626 7892 21632
rect 7852 21146 7880 21626
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 8220 20942 8248 21898
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 8208 20800 8260 20806
rect 8206 20768 8208 20777
rect 8260 20768 8262 20777
rect 8206 20703 8262 20712
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 8024 19440 8076 19446
rect 8024 19382 8076 19388
rect 7932 18828 7984 18834
rect 7932 18770 7984 18776
rect 7944 18465 7972 18770
rect 8036 18766 8064 19382
rect 8024 18760 8076 18766
rect 8024 18702 8076 18708
rect 7930 18456 7986 18465
rect 7852 18414 7930 18442
rect 7852 18222 7880 18414
rect 7930 18391 7986 18400
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 7840 18216 7892 18222
rect 7840 18158 7892 18164
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7944 17785 7972 18226
rect 8036 17882 8064 18702
rect 8024 17876 8076 17882
rect 8024 17818 8076 17824
rect 7930 17776 7986 17785
rect 7930 17711 7986 17720
rect 7656 17672 7708 17678
rect 7708 17632 7788 17660
rect 7656 17614 7708 17620
rect 7760 17134 7788 17632
rect 7840 17604 7892 17610
rect 7840 17546 7892 17552
rect 7852 17270 7880 17546
rect 8128 17377 8156 20334
rect 8312 19922 8340 23054
rect 8392 22636 8444 22642
rect 8392 22578 8444 22584
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 8298 19816 8354 19825
rect 8404 19802 8432 22578
rect 8496 21894 8524 26998
rect 8772 24750 8800 27066
rect 9220 25900 9272 25906
rect 9220 25842 9272 25848
rect 9036 25832 9088 25838
rect 9036 25774 9088 25780
rect 8760 24744 8812 24750
rect 8758 24712 8760 24721
rect 8812 24712 8814 24721
rect 8758 24647 8814 24656
rect 8668 24608 8720 24614
rect 8668 24550 8720 24556
rect 8576 23656 8628 23662
rect 8576 23598 8628 23604
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8484 21684 8536 21690
rect 8484 21626 8536 21632
rect 8496 20534 8524 21626
rect 8588 21350 8616 23598
rect 8680 22438 8708 24550
rect 9048 22778 9076 25774
rect 9232 25158 9260 25842
rect 9220 25152 9272 25158
rect 9220 25094 9272 25100
rect 9220 23180 9272 23186
rect 9220 23122 9272 23128
rect 9036 22772 9088 22778
rect 9036 22714 9088 22720
rect 9128 22772 9180 22778
rect 9128 22714 9180 22720
rect 9036 22636 9088 22642
rect 9036 22578 9088 22584
rect 8852 22568 8904 22574
rect 8852 22510 8904 22516
rect 8668 22432 8720 22438
rect 8668 22374 8720 22380
rect 8760 21548 8812 21554
rect 8760 21490 8812 21496
rect 8576 21344 8628 21350
rect 8576 21286 8628 21292
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 8484 20528 8536 20534
rect 8484 20470 8536 20476
rect 8354 19774 8432 19802
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 8298 19751 8354 19760
rect 8312 19718 8340 19751
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8220 18902 8248 19654
rect 8404 19514 8432 19654
rect 8392 19508 8444 19514
rect 8392 19450 8444 19456
rect 8496 19310 8524 19790
rect 8588 19378 8616 20538
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8484 19304 8536 19310
rect 8298 19272 8354 19281
rect 8484 19246 8536 19252
rect 8298 19207 8354 19216
rect 8312 19174 8340 19207
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8208 18896 8260 18902
rect 8208 18838 8260 18844
rect 8220 18748 8248 18838
rect 8300 18760 8352 18766
rect 8220 18720 8300 18748
rect 8300 18702 8352 18708
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8220 18358 8248 18566
rect 8312 18358 8340 18702
rect 8208 18352 8260 18358
rect 8208 18294 8260 18300
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 8392 18352 8444 18358
rect 8392 18294 8444 18300
rect 8220 17882 8248 18294
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 8404 17814 8432 18294
rect 8496 18290 8524 18702
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8482 18184 8538 18193
rect 8482 18119 8484 18128
rect 8536 18119 8538 18128
rect 8484 18090 8536 18096
rect 8392 17808 8444 17814
rect 8392 17750 8444 17756
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8114 17368 8170 17377
rect 8114 17303 8170 17312
rect 8220 17270 8248 17614
rect 8300 17604 8352 17610
rect 8300 17546 8352 17552
rect 7840 17264 7892 17270
rect 7840 17206 7892 17212
rect 8208 17264 8260 17270
rect 8208 17206 8260 17212
rect 7564 17128 7616 17134
rect 7748 17128 7800 17134
rect 7616 17088 7696 17116
rect 7564 17070 7616 17076
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7562 16552 7618 16561
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 7288 15972 7340 15978
rect 7288 15914 7340 15920
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7104 15632 7156 15638
rect 7104 15574 7156 15580
rect 6920 15496 6972 15502
rect 7208 15450 7236 15642
rect 6920 15438 6972 15444
rect 6932 15094 6960 15438
rect 7116 15434 7236 15450
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 7104 15428 7236 15434
rect 7156 15422 7236 15428
rect 7104 15370 7156 15376
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6932 14414 6960 14826
rect 7024 14822 7052 15370
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7116 14618 7144 14962
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6840 13530 6960 13546
rect 6840 13524 6972 13530
rect 6840 13518 6920 13524
rect 6920 13466 6972 13472
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6564 13190 6592 13262
rect 6656 13240 6684 13330
rect 6920 13252 6972 13258
rect 6656 13212 6920 13240
rect 6920 13194 6972 13200
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6564 12646 6592 12718
rect 7024 12646 7052 14214
rect 7208 12850 7236 14758
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 6368 12368 6420 12374
rect 6368 12310 6420 12316
rect 6564 12306 6592 12582
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 7300 12238 7328 15914
rect 7392 15502 7420 16390
rect 7380 15496 7432 15502
rect 7378 15464 7380 15473
rect 7432 15464 7434 15473
rect 7378 15399 7434 15408
rect 7392 12714 7420 15399
rect 7484 14278 7512 16526
rect 7562 16487 7564 16496
rect 7616 16487 7618 16496
rect 7564 16458 7616 16464
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7470 13424 7526 13433
rect 7470 13359 7526 13368
rect 7484 13326 7512 13359
rect 7576 13326 7604 15642
rect 7668 15570 7696 17088
rect 7748 17070 7800 17076
rect 7760 16522 7788 17070
rect 7852 16590 7880 17206
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7840 16584 7892 16590
rect 7840 16526 7892 16532
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 7760 15978 7788 16458
rect 7852 16114 7880 16526
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7748 15972 7800 15978
rect 7748 15914 7800 15920
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7668 14550 7696 15506
rect 7760 15094 7788 15914
rect 7748 15088 7800 15094
rect 7748 15030 7800 15036
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 7760 14482 7788 15030
rect 7852 14890 7880 16050
rect 7944 15502 7972 17138
rect 8220 16454 8248 17206
rect 8312 17066 8340 17546
rect 8588 17338 8616 19314
rect 8666 18864 8722 18873
rect 8666 18799 8722 18808
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8312 16726 8340 17002
rect 8680 16810 8708 18799
rect 8772 17202 8800 21490
rect 8864 21457 8892 22510
rect 9048 21690 9076 22578
rect 9140 22574 9168 22714
rect 9232 22642 9260 23122
rect 9220 22636 9272 22642
rect 9220 22578 9272 22584
rect 9128 22568 9180 22574
rect 9126 22536 9128 22545
rect 9180 22536 9182 22545
rect 9324 22522 9352 28698
rect 9588 28552 9640 28558
rect 9588 28494 9640 28500
rect 9600 27402 9628 28494
rect 9588 27396 9640 27402
rect 9588 27338 9640 27344
rect 9600 27169 9628 27338
rect 9586 27160 9642 27169
rect 9586 27095 9642 27104
rect 9784 26738 9812 30058
rect 10060 30054 10088 30087
rect 10048 30048 10100 30054
rect 10048 29990 10100 29996
rect 9956 29844 10008 29850
rect 9956 29786 10008 29792
rect 9968 28558 9996 29786
rect 10232 29164 10284 29170
rect 10232 29106 10284 29112
rect 9956 28552 10008 28558
rect 9956 28494 10008 28500
rect 10046 28112 10102 28121
rect 10046 28047 10102 28056
rect 9864 27872 9916 27878
rect 9864 27814 9916 27820
rect 9876 27538 9904 27814
rect 9864 27532 9916 27538
rect 9864 27474 9916 27480
rect 9692 26710 9812 26738
rect 9692 24614 9720 26710
rect 9876 26602 9904 27474
rect 9784 26574 9904 26602
rect 9588 24608 9640 24614
rect 9588 24550 9640 24556
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9600 24449 9628 24550
rect 9586 24440 9642 24449
rect 9784 24410 9812 26574
rect 9864 26512 9916 26518
rect 9864 26454 9916 26460
rect 9876 25906 9904 26454
rect 9864 25900 9916 25906
rect 9864 25842 9916 25848
rect 9586 24375 9642 24384
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9772 24404 9824 24410
rect 9772 24346 9824 24352
rect 9692 24041 9720 24346
rect 9770 24304 9826 24313
rect 9770 24239 9826 24248
rect 9784 24138 9812 24239
rect 9772 24132 9824 24138
rect 9772 24074 9824 24080
rect 9876 24070 9904 25842
rect 10060 25702 10088 28047
rect 10140 26444 10192 26450
rect 10140 26386 10192 26392
rect 10152 25786 10180 26386
rect 10244 26024 10272 29106
rect 10336 28121 10364 31078
rect 10876 30320 10928 30326
rect 10506 30288 10562 30297
rect 10876 30262 10928 30268
rect 10506 30223 10562 30232
rect 10520 29238 10548 30223
rect 10888 30122 10916 30262
rect 10876 30116 10928 30122
rect 10876 30058 10928 30064
rect 10692 29572 10744 29578
rect 10692 29514 10744 29520
rect 10508 29232 10560 29238
rect 10508 29174 10560 29180
rect 10704 29102 10732 29514
rect 10784 29504 10836 29510
rect 10784 29446 10836 29452
rect 10692 29096 10744 29102
rect 10692 29038 10744 29044
rect 10692 28960 10744 28966
rect 10796 28937 10824 29446
rect 10692 28902 10744 28908
rect 10782 28928 10838 28937
rect 10704 28642 10732 28902
rect 10782 28863 10838 28872
rect 10704 28614 10824 28642
rect 10692 28552 10744 28558
rect 10692 28494 10744 28500
rect 10600 28484 10652 28490
rect 10600 28426 10652 28432
rect 10414 28384 10470 28393
rect 10414 28319 10470 28328
rect 10322 28112 10378 28121
rect 10322 28047 10378 28056
rect 10428 27878 10456 28319
rect 10612 28257 10640 28426
rect 10598 28248 10654 28257
rect 10704 28218 10732 28494
rect 10796 28490 10824 28614
rect 10784 28484 10836 28490
rect 10784 28426 10836 28432
rect 10876 28484 10928 28490
rect 10876 28426 10928 28432
rect 10598 28183 10654 28192
rect 10692 28212 10744 28218
rect 10692 28154 10744 28160
rect 10416 27872 10468 27878
rect 10416 27814 10468 27820
rect 10416 27668 10468 27674
rect 10416 27610 10468 27616
rect 10322 26616 10378 26625
rect 10322 26551 10378 26560
rect 10336 26518 10364 26551
rect 10428 26518 10456 27610
rect 10324 26512 10376 26518
rect 10324 26454 10376 26460
rect 10416 26512 10468 26518
rect 10416 26454 10468 26460
rect 10324 26376 10376 26382
rect 10322 26344 10324 26353
rect 10376 26344 10378 26353
rect 10322 26279 10378 26288
rect 10244 25996 10364 26024
rect 10232 25900 10284 25906
rect 10232 25842 10284 25848
rect 10244 25786 10272 25842
rect 10152 25758 10272 25786
rect 10336 25770 10364 25996
rect 10324 25764 10376 25770
rect 10152 25702 10180 25758
rect 10324 25706 10376 25712
rect 10048 25696 10100 25702
rect 10048 25638 10100 25644
rect 10140 25696 10192 25702
rect 10140 25638 10192 25644
rect 10048 25492 10100 25498
rect 10048 25434 10100 25440
rect 10060 25158 10088 25434
rect 10048 25152 10100 25158
rect 10048 25094 10100 25100
rect 10048 24812 10100 24818
rect 10048 24754 10100 24760
rect 9956 24608 10008 24614
rect 9954 24576 9956 24585
rect 10008 24576 10010 24585
rect 9954 24511 10010 24520
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 9864 24064 9916 24070
rect 9678 24032 9734 24041
rect 9864 24006 9916 24012
rect 9968 24018 9996 24346
rect 10060 24274 10088 24754
rect 10152 24750 10180 25638
rect 10428 25294 10456 26454
rect 10508 25968 10560 25974
rect 10508 25910 10560 25916
rect 10520 25294 10548 25910
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 10232 25288 10284 25294
rect 10232 25230 10284 25236
rect 10416 25288 10468 25294
rect 10416 25230 10468 25236
rect 10508 25288 10560 25294
rect 10508 25230 10560 25236
rect 10140 24744 10192 24750
rect 10140 24686 10192 24692
rect 10048 24268 10100 24274
rect 10048 24210 10100 24216
rect 9968 23990 10088 24018
rect 9678 23967 9734 23976
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 9680 23792 9732 23798
rect 9680 23734 9732 23740
rect 9496 23520 9548 23526
rect 9496 23462 9548 23468
rect 9404 23044 9456 23050
rect 9404 22986 9456 22992
rect 9416 22710 9444 22986
rect 9404 22704 9456 22710
rect 9404 22646 9456 22652
rect 9126 22471 9182 22480
rect 9232 22494 9352 22522
rect 9404 22568 9456 22574
rect 9404 22510 9456 22516
rect 9508 22522 9536 23462
rect 9588 23248 9640 23254
rect 9588 23190 9640 23196
rect 9600 22642 9628 23190
rect 9588 22636 9640 22642
rect 9588 22578 9640 22584
rect 9036 21684 9088 21690
rect 9036 21626 9088 21632
rect 8850 21448 8906 21457
rect 8906 21406 9076 21434
rect 8850 21383 8906 21392
rect 8852 21344 8904 21350
rect 8852 21286 8904 21292
rect 8864 21146 8892 21286
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 9048 20913 9076 21406
rect 9128 21004 9180 21010
rect 9128 20946 9180 20952
rect 9034 20904 9090 20913
rect 8852 20868 8904 20874
rect 9034 20839 9090 20848
rect 8852 20810 8904 20816
rect 8864 20641 8892 20810
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8850 20632 8906 20641
rect 8850 20567 8906 20576
rect 8852 19916 8904 19922
rect 8852 19858 8904 19864
rect 8864 19417 8892 19858
rect 8956 19854 8984 20742
rect 9036 20528 9088 20534
rect 9036 20470 9088 20476
rect 9048 19854 9076 20470
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 8956 19514 8984 19790
rect 8944 19508 8996 19514
rect 8944 19450 8996 19456
rect 8850 19408 8906 19417
rect 8850 19343 8906 19352
rect 8864 18057 8892 19343
rect 8956 18766 8984 19450
rect 9048 18873 9076 19790
rect 9034 18864 9090 18873
rect 9034 18799 9090 18808
rect 8944 18760 8996 18766
rect 8944 18702 8996 18708
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 8942 18456 8998 18465
rect 8942 18391 8998 18400
rect 8956 18222 8984 18391
rect 9048 18290 9076 18566
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 8850 18048 8906 18057
rect 8850 17983 8906 17992
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8496 16782 8708 16810
rect 8772 16794 8800 17138
rect 8760 16788 8812 16794
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8220 16046 8248 16390
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 8208 16040 8260 16046
rect 8312 16028 8340 16662
rect 8392 16040 8444 16046
rect 8312 16000 8392 16028
rect 8208 15982 8260 15988
rect 8392 15982 8444 15988
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 8036 15026 8064 15982
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 8128 15162 8156 15438
rect 8404 15162 8432 15982
rect 8496 15366 8524 16782
rect 8760 16730 8812 16736
rect 8576 16720 8628 16726
rect 8574 16688 8576 16697
rect 8628 16688 8630 16697
rect 8574 16623 8630 16632
rect 8588 15502 8616 16623
rect 8864 16266 8892 17983
rect 8942 17776 8998 17785
rect 8942 17711 8998 17720
rect 8956 16590 8984 17711
rect 9048 17338 9076 18226
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8680 16238 8892 16266
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8116 15156 8168 15162
rect 8392 15156 8444 15162
rect 8116 15098 8168 15104
rect 8220 15116 8392 15144
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 7840 14884 7892 14890
rect 7840 14826 7892 14832
rect 7852 14618 7880 14826
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7760 14346 7788 14418
rect 7748 14340 7800 14346
rect 7748 14282 7800 14288
rect 7852 14006 7880 14554
rect 7944 14362 7972 14962
rect 8036 14482 8064 14962
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 7944 14334 8064 14362
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 7944 14113 7972 14214
rect 7930 14104 7986 14113
rect 7930 14039 7986 14048
rect 7840 14000 7892 14006
rect 7840 13942 7892 13948
rect 7930 13696 7986 13705
rect 7930 13631 7986 13640
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7944 12782 7972 13631
rect 8036 13394 8064 14334
rect 8128 13870 8156 15098
rect 8220 14550 8248 15116
rect 8392 15098 8444 15104
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8208 14544 8260 14550
rect 8496 14532 8524 14894
rect 8496 14504 8529 14532
rect 8208 14486 8260 14492
rect 8220 13938 8248 14486
rect 8501 14464 8529 14504
rect 8429 14436 8529 14464
rect 8429 14414 8457 14436
rect 8392 14408 8457 14414
rect 8444 14356 8457 14408
rect 8392 14350 8457 14356
rect 8404 14334 8457 14350
rect 8588 14372 8616 15438
rect 8680 14906 8708 16238
rect 8852 16176 8904 16182
rect 8758 16144 8814 16153
rect 8852 16118 8904 16124
rect 8758 16079 8760 16088
rect 8812 16079 8814 16088
rect 8760 16050 8812 16056
rect 8772 15706 8800 16050
rect 8864 15706 8892 16118
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 8864 15026 8892 15098
rect 8852 15020 8904 15026
rect 8852 14962 8904 14968
rect 8680 14878 8892 14906
rect 8760 14408 8812 14414
rect 8588 14356 8760 14372
rect 8588 14350 8812 14356
rect 8588 14344 8800 14350
rect 8588 13938 8616 14344
rect 8864 14090 8892 14878
rect 8680 14062 8892 14090
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 8588 13802 8616 13874
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8680 13682 8708 14062
rect 8850 13968 8906 13977
rect 8956 13954 8984 16526
rect 9048 16522 9076 17274
rect 9140 17202 9168 20946
rect 9232 20058 9260 22494
rect 9416 20992 9444 22510
rect 9508 22494 9628 22522
rect 9496 21480 9548 21486
rect 9496 21422 9548 21428
rect 9508 21078 9536 21422
rect 9496 21072 9548 21078
rect 9496 21014 9548 21020
rect 9324 20964 9444 20992
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 9324 19310 9352 20964
rect 9508 20942 9536 21014
rect 9496 20936 9548 20942
rect 9496 20878 9548 20884
rect 9404 20868 9456 20874
rect 9404 20810 9456 20816
rect 9416 20369 9444 20810
rect 9402 20360 9458 20369
rect 9402 20295 9458 20304
rect 9402 20088 9458 20097
rect 9402 20023 9404 20032
rect 9456 20023 9458 20032
rect 9404 19994 9456 20000
rect 9508 19938 9536 20878
rect 9600 20754 9628 22494
rect 9692 21962 9720 23734
rect 9784 23730 9812 23802
rect 9876 23730 9996 23746
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9876 23724 10008 23730
rect 9876 23718 9956 23724
rect 9784 23050 9812 23666
rect 9876 23118 9904 23718
rect 9956 23666 10008 23672
rect 10060 23610 10088 23990
rect 9968 23582 10088 23610
rect 10152 23594 10180 24686
rect 10140 23588 10192 23594
rect 9864 23112 9916 23118
rect 9864 23054 9916 23060
rect 9772 23044 9824 23050
rect 9772 22986 9824 22992
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9678 21856 9734 21865
rect 9678 21791 9734 21800
rect 9692 21418 9720 21791
rect 9680 21412 9732 21418
rect 9680 21354 9732 21360
rect 9784 21146 9812 22578
rect 9876 21690 9904 23054
rect 9968 22642 9996 23582
rect 10140 23530 10192 23536
rect 10244 23474 10272 25230
rect 10324 25220 10376 25226
rect 10324 25162 10376 25168
rect 10336 24614 10364 25162
rect 10612 24993 10640 25842
rect 10692 25832 10744 25838
rect 10692 25774 10744 25780
rect 10598 24984 10654 24993
rect 10598 24919 10654 24928
rect 10324 24608 10376 24614
rect 10324 24550 10376 24556
rect 10704 24426 10732 25774
rect 10796 24857 10824 28426
rect 10888 28218 10916 28426
rect 10876 28212 10928 28218
rect 10876 28154 10928 28160
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 10888 26586 10916 26930
rect 10980 26586 11008 31758
rect 11072 30190 11100 31962
rect 11152 31816 11204 31822
rect 11152 31758 11204 31764
rect 11164 31414 11192 31758
rect 12072 31476 12124 31482
rect 12072 31418 12124 31424
rect 11152 31408 11204 31414
rect 11152 31350 11204 31356
rect 11164 31113 11192 31350
rect 11150 31104 11206 31113
rect 11150 31039 11206 31048
rect 11888 30932 11940 30938
rect 11888 30874 11940 30880
rect 11060 30184 11112 30190
rect 11060 30126 11112 30132
rect 11152 29708 11204 29714
rect 11152 29650 11204 29656
rect 11060 29640 11112 29646
rect 11058 29608 11060 29617
rect 11112 29608 11114 29617
rect 11058 29543 11114 29552
rect 11060 29096 11112 29102
rect 11060 29038 11112 29044
rect 11072 28762 11100 29038
rect 11060 28756 11112 28762
rect 11060 28698 11112 28704
rect 11060 28076 11112 28082
rect 11060 28018 11112 28024
rect 11072 27606 11100 28018
rect 11060 27600 11112 27606
rect 11060 27542 11112 27548
rect 10876 26580 10928 26586
rect 10876 26522 10928 26528
rect 10968 26580 11020 26586
rect 10968 26522 11020 26528
rect 11164 26466 11192 29650
rect 11244 29640 11296 29646
rect 11244 29582 11296 29588
rect 11256 27334 11284 29582
rect 11796 29504 11848 29510
rect 11796 29446 11848 29452
rect 11808 29170 11836 29446
rect 11428 29164 11480 29170
rect 11428 29106 11480 29112
rect 11796 29164 11848 29170
rect 11796 29106 11848 29112
rect 11336 28756 11388 28762
rect 11336 28698 11388 28704
rect 11348 28529 11376 28698
rect 11440 28626 11468 29106
rect 11704 29028 11756 29034
rect 11704 28970 11756 28976
rect 11520 28688 11572 28694
rect 11520 28630 11572 28636
rect 11428 28620 11480 28626
rect 11428 28562 11480 28568
rect 11334 28520 11390 28529
rect 11334 28455 11390 28464
rect 11244 27328 11296 27334
rect 11244 27270 11296 27276
rect 10980 26438 11192 26466
rect 10876 26240 10928 26246
rect 10876 26182 10928 26188
rect 10888 26042 10916 26182
rect 10876 26036 10928 26042
rect 10876 25978 10928 25984
rect 10980 25922 11008 26438
rect 11152 26376 11204 26382
rect 11152 26318 11204 26324
rect 11164 26217 11192 26318
rect 11150 26208 11206 26217
rect 11150 26143 11206 26152
rect 10876 25900 10928 25906
rect 10980 25894 11100 25922
rect 10876 25842 10928 25848
rect 10888 25770 10916 25842
rect 10876 25764 10928 25770
rect 10876 25706 10928 25712
rect 10782 24848 10838 24857
rect 10782 24783 10838 24792
rect 10612 24398 10732 24426
rect 10416 24268 10468 24274
rect 10416 24210 10468 24216
rect 10324 24200 10376 24206
rect 10428 24177 10456 24210
rect 10324 24142 10376 24148
rect 10414 24168 10470 24177
rect 10336 24070 10364 24142
rect 10612 24138 10640 24398
rect 10690 24304 10746 24313
rect 10690 24239 10692 24248
rect 10744 24239 10746 24248
rect 10692 24210 10744 24216
rect 10414 24103 10470 24112
rect 10600 24132 10652 24138
rect 10600 24074 10652 24080
rect 10324 24064 10376 24070
rect 10324 24006 10376 24012
rect 10336 23866 10364 24006
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 10324 23724 10376 23730
rect 10324 23666 10376 23672
rect 10060 23446 10272 23474
rect 10060 22982 10088 23446
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 10048 22976 10100 22982
rect 10048 22918 10100 22924
rect 10244 22681 10272 23054
rect 10230 22672 10286 22681
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 10048 22636 10100 22642
rect 10048 22578 10100 22584
rect 10140 22636 10192 22642
rect 10230 22607 10286 22616
rect 10140 22578 10192 22584
rect 10060 22030 10088 22578
rect 10152 22166 10180 22578
rect 10336 22574 10364 23666
rect 10416 23112 10468 23118
rect 10416 23054 10468 23060
rect 10324 22568 10376 22574
rect 10324 22510 10376 22516
rect 10140 22160 10192 22166
rect 10140 22102 10192 22108
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9678 21040 9734 21049
rect 9678 20975 9734 20984
rect 9692 20942 9720 20975
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 9784 20754 9812 20878
rect 9600 20726 9812 20754
rect 9600 20641 9628 20726
rect 9586 20632 9642 20641
rect 9586 20567 9642 20576
rect 9876 20534 9904 21626
rect 10048 21616 10100 21622
rect 10048 21558 10100 21564
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9864 20528 9916 20534
rect 9600 20466 9812 20482
rect 9864 20470 9916 20476
rect 9588 20460 9824 20466
rect 9640 20454 9772 20460
rect 9588 20402 9640 20408
rect 9772 20402 9824 20408
rect 9968 20330 9996 21490
rect 10060 20466 10088 21558
rect 10048 20460 10100 20466
rect 10048 20402 10100 20408
rect 10046 20360 10102 20369
rect 9956 20324 10008 20330
rect 10046 20295 10102 20304
rect 9956 20266 10008 20272
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9784 19961 9812 20198
rect 9416 19910 9536 19938
rect 9586 19952 9642 19961
rect 9416 19786 9444 19910
rect 9586 19887 9642 19896
rect 9770 19952 9826 19961
rect 9770 19887 9772 19896
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 9404 19780 9456 19786
rect 9404 19722 9456 19728
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9220 18896 9272 18902
rect 9220 18838 9272 18844
rect 9232 18465 9260 18838
rect 9218 18456 9274 18465
rect 9218 18391 9274 18400
rect 9220 18284 9272 18290
rect 9324 18272 9352 19246
rect 9272 18244 9352 18272
rect 9220 18226 9272 18232
rect 9220 17604 9272 17610
rect 9220 17546 9272 17552
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9036 16516 9088 16522
rect 9036 16458 9088 16464
rect 9048 16114 9076 16458
rect 9140 16250 9168 17138
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 9128 16040 9180 16046
rect 9128 15982 9180 15988
rect 9036 15972 9088 15978
rect 9036 15914 9088 15920
rect 9048 15745 9076 15914
rect 9034 15736 9090 15745
rect 9034 15671 9090 15680
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 9048 14056 9076 15302
rect 9140 14793 9168 15982
rect 9232 15910 9260 17546
rect 9324 17338 9352 18244
rect 9508 17610 9536 19790
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9324 16658 9352 17274
rect 9496 17196 9548 17202
rect 9496 17138 9548 17144
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9324 15960 9352 16594
rect 9508 16454 9536 17138
rect 9496 16448 9548 16454
rect 9402 16416 9458 16425
rect 9496 16390 9548 16396
rect 9402 16351 9458 16360
rect 9416 16182 9444 16351
rect 9508 16250 9536 16390
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9404 16176 9456 16182
rect 9404 16118 9456 16124
rect 9404 15972 9456 15978
rect 9324 15932 9404 15960
rect 9404 15914 9456 15920
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 9508 15570 9536 16186
rect 9600 15994 9628 19887
rect 9824 19887 9826 19896
rect 9772 19858 9824 19864
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9692 18766 9720 19246
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9692 17882 9720 18294
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9784 17678 9812 19450
rect 9862 19000 9918 19009
rect 9862 18935 9864 18944
rect 9916 18935 9918 18944
rect 9864 18906 9916 18912
rect 9956 18896 10008 18902
rect 9876 18844 9956 18850
rect 9876 18838 10008 18844
rect 9876 18822 9996 18838
rect 9876 18766 9904 18822
rect 9864 18760 9916 18766
rect 9864 18702 9916 18708
rect 9772 17672 9824 17678
rect 9692 17632 9772 17660
rect 9692 16425 9720 17632
rect 9772 17614 9824 17620
rect 9876 17202 9904 18702
rect 9954 18320 10010 18329
rect 9954 18255 10010 18264
rect 9968 18222 9996 18255
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 9954 17912 10010 17921
rect 9954 17847 9956 17856
rect 10008 17847 10010 17856
rect 9956 17818 10008 17824
rect 9956 17536 10008 17542
rect 9956 17478 10008 17484
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9678 16416 9734 16425
rect 9678 16351 9734 16360
rect 9600 15966 9720 15994
rect 9692 15638 9720 15966
rect 9680 15632 9732 15638
rect 9680 15574 9732 15580
rect 9496 15564 9548 15570
rect 9496 15506 9548 15512
rect 9220 15088 9272 15094
rect 9220 15030 9272 15036
rect 9126 14784 9182 14793
rect 9126 14719 9182 14728
rect 9128 14544 9180 14550
rect 9128 14486 9180 14492
rect 9140 14249 9168 14486
rect 9232 14482 9260 15030
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9324 14414 9352 14962
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9508 14346 9536 14894
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 9692 14498 9720 15574
rect 9784 15502 9812 17138
rect 9876 16726 9904 17138
rect 9864 16720 9916 16726
rect 9864 16662 9916 16668
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9876 15026 9904 16662
rect 9968 16096 9996 17478
rect 10060 16572 10088 20295
rect 10152 19378 10180 22102
rect 10232 21344 10284 21350
rect 10230 21312 10232 21321
rect 10284 21312 10286 21321
rect 10230 21247 10286 21256
rect 10336 21010 10364 22510
rect 10428 22166 10456 23054
rect 10508 22432 10560 22438
rect 10508 22374 10560 22380
rect 10416 22160 10468 22166
rect 10416 22102 10468 22108
rect 10416 22024 10468 22030
rect 10416 21966 10468 21972
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10336 20466 10364 20946
rect 10428 20874 10456 21966
rect 10416 20868 10468 20874
rect 10416 20810 10468 20816
rect 10520 20505 10548 22374
rect 10506 20496 10562 20505
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10324 20460 10376 20466
rect 10506 20431 10562 20440
rect 10324 20402 10376 20408
rect 10244 20330 10272 20402
rect 10506 20360 10562 20369
rect 10232 20324 10284 20330
rect 10506 20295 10508 20304
rect 10232 20266 10284 20272
rect 10560 20295 10562 20304
rect 10508 20266 10560 20272
rect 10244 20058 10272 20266
rect 10232 20052 10284 20058
rect 10232 19994 10284 20000
rect 10506 19952 10562 19961
rect 10506 19887 10562 19896
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10428 19378 10456 19790
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 10152 18698 10180 19314
rect 10520 18970 10548 19887
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10140 18692 10192 18698
rect 10140 18634 10192 18640
rect 10232 18692 10284 18698
rect 10232 18634 10284 18640
rect 10244 18426 10272 18634
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10152 18222 10180 18362
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 10152 16794 10180 17138
rect 10244 17134 10272 18362
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10336 17882 10364 18226
rect 10416 18148 10468 18154
rect 10416 18090 10468 18096
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 10140 16584 10192 16590
rect 10060 16544 10140 16572
rect 10140 16526 10192 16532
rect 9968 16068 10088 16096
rect 9954 16008 10010 16017
rect 9954 15943 10010 15952
rect 9968 15910 9996 15943
rect 9956 15904 10008 15910
rect 10060 15881 10088 16068
rect 9956 15846 10008 15852
rect 10046 15872 10102 15881
rect 10046 15807 10102 15816
rect 10060 15450 10088 15807
rect 10152 15473 10180 16526
rect 10336 16114 10364 17818
rect 10428 17785 10456 18090
rect 10414 17776 10470 17785
rect 10414 17711 10470 17720
rect 10506 17640 10562 17649
rect 10506 17575 10562 17584
rect 10520 17202 10548 17575
rect 10612 17354 10640 24074
rect 10796 23866 10824 24783
rect 10888 24698 10916 25706
rect 11072 25378 11100 25894
rect 11072 25350 11192 25378
rect 10888 24670 11100 24698
rect 10876 24268 10928 24274
rect 10876 24210 10928 24216
rect 10888 23905 10916 24210
rect 10968 24064 11020 24070
rect 10968 24006 11020 24012
rect 10874 23896 10930 23905
rect 10784 23860 10836 23866
rect 10874 23831 10930 23840
rect 10784 23802 10836 23808
rect 10876 23792 10928 23798
rect 10876 23734 10928 23740
rect 10782 22944 10838 22953
rect 10782 22879 10838 22888
rect 10692 22636 10744 22642
rect 10692 22578 10744 22584
rect 10704 22234 10732 22578
rect 10796 22438 10824 22879
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10888 22250 10916 23734
rect 10980 23662 11008 24006
rect 10968 23656 11020 23662
rect 10968 23598 11020 23604
rect 11072 22409 11100 24670
rect 11058 22400 11114 22409
rect 11058 22335 11114 22344
rect 10692 22228 10744 22234
rect 10692 22170 10744 22176
rect 10796 22222 10916 22250
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10704 20874 10732 21490
rect 10692 20868 10744 20874
rect 10692 20810 10744 20816
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 10704 19514 10732 20334
rect 10796 20262 10824 22222
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 11072 22001 11100 22034
rect 11058 21992 11114 22001
rect 10876 21956 10928 21962
rect 11058 21927 11114 21936
rect 10876 21898 10928 21904
rect 10888 21078 10916 21898
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 10876 21072 10928 21078
rect 10876 21014 10928 21020
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10888 20074 10916 21014
rect 10980 20942 11008 21422
rect 10968 20936 11020 20942
rect 10968 20878 11020 20884
rect 10968 20800 11020 20806
rect 11072 20754 11100 21626
rect 11020 20748 11100 20754
rect 10968 20742 11100 20748
rect 10980 20726 11100 20742
rect 10968 20528 11020 20534
rect 10968 20470 11020 20476
rect 10796 20046 10916 20074
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10704 19378 10732 19450
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10796 18850 10824 20046
rect 10876 19984 10928 19990
rect 10876 19926 10928 19932
rect 10888 19378 10916 19926
rect 10980 19854 11008 20470
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 10796 18822 10916 18850
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10704 18358 10732 18702
rect 10692 18352 10744 18358
rect 10690 18320 10692 18329
rect 10744 18320 10746 18329
rect 10690 18255 10746 18264
rect 10612 17326 10824 17354
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10414 17096 10470 17105
rect 10414 17031 10470 17040
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10230 16008 10286 16017
rect 10230 15943 10232 15952
rect 10284 15943 10286 15952
rect 10232 15914 10284 15920
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10336 15570 10364 15846
rect 10428 15570 10456 17031
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10612 16522 10640 16594
rect 10600 16516 10652 16522
rect 10520 16476 10600 16504
rect 10520 16182 10548 16476
rect 10600 16458 10652 16464
rect 10598 16416 10654 16425
rect 10598 16351 10654 16360
rect 10508 16176 10560 16182
rect 10508 16118 10560 16124
rect 10612 16114 10640 16351
rect 10704 16289 10732 17138
rect 10690 16280 10746 16289
rect 10796 16250 10824 17326
rect 10690 16215 10746 16224
rect 10784 16244 10836 16250
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 10612 15706 10640 16050
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 9968 15422 10088 15450
rect 10138 15464 10194 15473
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9968 14958 9996 15422
rect 10138 15399 10194 15408
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 10060 15094 10088 15302
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9784 14618 9812 14758
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 9126 14240 9182 14249
rect 9126 14175 9182 14184
rect 9048 14028 9352 14056
rect 8956 13926 9260 13954
rect 8850 13903 8906 13912
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8588 13654 8708 13682
rect 8024 13388 8076 13394
rect 8024 13330 8076 13336
rect 8588 13326 8616 13654
rect 8666 13560 8722 13569
rect 8666 13495 8722 13504
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7760 12306 7788 12650
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 5460 11830 5488 12038
rect 5448 11824 5500 11830
rect 846 11792 902 11801
rect 5448 11766 5500 11772
rect 846 11727 848 11736
rect 900 11727 902 11736
rect 848 11698 900 11704
rect 7944 11694 7972 12718
rect 8036 12238 8064 12786
rect 8128 12782 8156 13126
rect 8680 12889 8708 13495
rect 8666 12880 8722 12889
rect 8666 12815 8722 12824
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8680 12306 8708 12815
rect 8772 12374 8800 13806
rect 8864 13462 8892 13903
rect 9232 13870 9260 13926
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9126 13560 9182 13569
rect 9126 13495 9182 13504
rect 9140 13462 9168 13495
rect 9324 13462 9352 14028
rect 9600 13938 9628 14486
rect 9692 14470 9812 14498
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9692 14113 9720 14350
rect 9678 14104 9734 14113
rect 9678 14039 9734 14048
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 8852 13456 8904 13462
rect 8852 13398 8904 13404
rect 9128 13456 9180 13462
rect 9128 13398 9180 13404
rect 9312 13456 9364 13462
rect 9312 13398 9364 13404
rect 9496 13456 9548 13462
rect 9496 13398 9548 13404
rect 8864 12850 8892 13398
rect 9404 13320 9456 13326
rect 9508 13308 9536 13398
rect 9600 13394 9628 13670
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9456 13280 9536 13308
rect 9404 13262 9456 13268
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 9508 12714 9536 13280
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9600 12714 9628 12854
rect 9692 12850 9720 14039
rect 9784 12850 9812 14470
rect 10152 13410 10180 15399
rect 9876 13382 10180 13410
rect 9876 13190 9904 13382
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9588 12708 9640 12714
rect 9588 12650 9640 12656
rect 9784 12442 9812 12786
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 8760 12368 8812 12374
rect 8760 12310 8812 12316
rect 8668 12300 8720 12306
rect 8668 12242 8720 12248
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 8300 12164 8352 12170
rect 8300 12106 8352 12112
rect 8312 11898 8340 12106
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 9968 11830 9996 13262
rect 10060 12986 10088 13262
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10336 12918 10364 15506
rect 10704 15162 10732 16215
rect 10784 16186 10836 16192
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10796 15745 10824 15982
rect 10888 15910 10916 18822
rect 10968 18692 11020 18698
rect 10968 18634 11020 18640
rect 10980 17882 11008 18634
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 10966 17776 11022 17785
rect 10966 17711 11022 17720
rect 10980 17066 11008 17711
rect 11058 17232 11114 17241
rect 11058 17167 11114 17176
rect 11072 17134 11100 17167
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10966 16960 11022 16969
rect 10966 16895 11022 16904
rect 10980 16658 11008 16895
rect 11072 16833 11100 17070
rect 11058 16824 11114 16833
rect 11058 16759 11114 16768
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 11164 16454 11192 25350
rect 11256 23322 11284 27270
rect 11440 26994 11468 28562
rect 11532 28422 11560 28630
rect 11520 28416 11572 28422
rect 11520 28358 11572 28364
rect 11612 28144 11664 28150
rect 11612 28086 11664 28092
rect 11520 27940 11572 27946
rect 11520 27882 11572 27888
rect 11428 26988 11480 26994
rect 11428 26930 11480 26936
rect 11428 26852 11480 26858
rect 11428 26794 11480 26800
rect 11336 26580 11388 26586
rect 11336 26522 11388 26528
rect 11244 23316 11296 23322
rect 11244 23258 11296 23264
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 11256 16674 11284 23054
rect 11348 22098 11376 26522
rect 11440 26450 11468 26794
rect 11428 26444 11480 26450
rect 11428 26386 11480 26392
rect 11336 22092 11388 22098
rect 11336 22034 11388 22040
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 11348 20602 11376 21898
rect 11440 21350 11468 26386
rect 11532 22137 11560 27882
rect 11624 26314 11652 28086
rect 11716 26858 11744 28970
rect 11796 28008 11848 28014
rect 11796 27950 11848 27956
rect 11704 26852 11756 26858
rect 11704 26794 11756 26800
rect 11704 26444 11756 26450
rect 11704 26386 11756 26392
rect 11612 26308 11664 26314
rect 11612 26250 11664 26256
rect 11624 25158 11652 26250
rect 11716 26081 11744 26386
rect 11702 26072 11758 26081
rect 11702 26007 11758 26016
rect 11704 25424 11756 25430
rect 11704 25366 11756 25372
rect 11612 25152 11664 25158
rect 11612 25094 11664 25100
rect 11612 24744 11664 24750
rect 11612 24686 11664 24692
rect 11624 24342 11652 24686
rect 11716 24410 11744 25366
rect 11808 24614 11836 27950
rect 11900 25702 11928 30874
rect 12084 30666 12112 31418
rect 12360 30938 12388 32438
rect 13544 32360 13596 32366
rect 13544 32302 13596 32308
rect 13634 32328 13690 32337
rect 13176 32224 13228 32230
rect 13176 32166 13228 32172
rect 12348 30932 12400 30938
rect 12348 30874 12400 30880
rect 12808 30796 12860 30802
rect 12808 30738 12860 30744
rect 12072 30660 12124 30666
rect 12072 30602 12124 30608
rect 11980 29300 12032 29306
rect 11980 29242 12032 29248
rect 11992 29209 12020 29242
rect 11978 29200 12034 29209
rect 11978 29135 12034 29144
rect 11978 26616 12034 26625
rect 11978 26551 12034 26560
rect 11992 26382 12020 26551
rect 11980 26376 12032 26382
rect 11980 26318 12032 26324
rect 11980 25900 12032 25906
rect 11980 25842 12032 25848
rect 11992 25786 12020 25842
rect 12084 25786 12112 30602
rect 12622 27568 12678 27577
rect 12622 27503 12678 27512
rect 12256 26784 12308 26790
rect 12256 26726 12308 26732
rect 12268 26382 12296 26726
rect 12636 26586 12664 27503
rect 12624 26580 12676 26586
rect 12624 26522 12676 26528
rect 12360 26450 12480 26466
rect 12348 26444 12480 26450
rect 12400 26438 12480 26444
rect 12348 26386 12400 26392
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 12452 26042 12480 26438
rect 12532 26240 12584 26246
rect 12532 26182 12584 26188
rect 12716 26240 12768 26246
rect 12716 26182 12768 26188
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12544 25974 12572 26182
rect 12532 25968 12584 25974
rect 12532 25910 12584 25916
rect 12256 25900 12308 25906
rect 12256 25842 12308 25848
rect 11992 25758 12112 25786
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 11796 24608 11848 24614
rect 11794 24576 11796 24585
rect 11848 24576 11850 24585
rect 11794 24511 11850 24520
rect 11704 24404 11756 24410
rect 11704 24346 11756 24352
rect 11612 24336 11664 24342
rect 11612 24278 11664 24284
rect 11796 24336 11848 24342
rect 11796 24278 11848 24284
rect 11704 23248 11756 23254
rect 11704 23190 11756 23196
rect 11716 22574 11744 23190
rect 11704 22568 11756 22574
rect 11704 22510 11756 22516
rect 11518 22128 11574 22137
rect 11518 22063 11574 22072
rect 11428 21344 11480 21350
rect 11428 21286 11480 21292
rect 11532 21146 11560 22063
rect 11610 21992 11666 22001
rect 11716 21962 11744 22510
rect 11610 21927 11666 21936
rect 11704 21956 11756 21962
rect 11624 21729 11652 21927
rect 11704 21898 11756 21904
rect 11610 21720 11666 21729
rect 11610 21655 11666 21664
rect 11612 21616 11664 21622
rect 11612 21558 11664 21564
rect 11520 21140 11572 21146
rect 11520 21082 11572 21088
rect 11624 21049 11652 21558
rect 11610 21040 11666 21049
rect 11610 20975 11666 20984
rect 11428 20800 11480 20806
rect 11428 20742 11480 20748
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 11348 17610 11376 20538
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 11440 17490 11468 20742
rect 11518 20224 11574 20233
rect 11518 20159 11574 20168
rect 11532 19922 11560 20159
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 11520 17604 11572 17610
rect 11520 17546 11572 17552
rect 11348 17462 11468 17490
rect 11348 17241 11376 17462
rect 11334 17232 11390 17241
rect 11334 17167 11390 17176
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11256 16646 11376 16674
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10980 15745 11008 16390
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 10782 15736 10838 15745
rect 10782 15671 10838 15680
rect 10966 15736 11022 15745
rect 10966 15671 11022 15680
rect 10876 15632 10928 15638
rect 11072 15620 11100 16118
rect 11164 15910 11192 16186
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 10876 15574 10928 15580
rect 10980 15592 11100 15620
rect 10888 15366 10916 15574
rect 10784 15360 10836 15366
rect 10782 15328 10784 15337
rect 10876 15360 10928 15366
rect 10836 15328 10838 15337
rect 10876 15302 10928 15308
rect 10782 15263 10838 15272
rect 10980 15178 11008 15592
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10796 15150 11008 15178
rect 11058 15192 11114 15201
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10520 14822 10548 14962
rect 10600 14952 10652 14958
rect 10796 14940 10824 15150
rect 11058 15127 11060 15136
rect 11112 15127 11114 15136
rect 11060 15098 11112 15104
rect 11164 15065 11192 15438
rect 11150 15056 11206 15065
rect 10876 15020 10928 15026
rect 11150 14991 11206 15000
rect 10876 14962 10928 14968
rect 10652 14912 10824 14940
rect 10600 14894 10652 14900
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10428 13530 10456 13874
rect 10600 13728 10652 13734
rect 10704 13716 10732 14912
rect 10888 14074 10916 14962
rect 11152 14884 11204 14890
rect 11152 14826 11204 14832
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10876 13728 10928 13734
rect 10704 13688 10876 13716
rect 10600 13670 10652 13676
rect 10876 13670 10928 13676
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10324 12912 10376 12918
rect 10324 12854 10376 12860
rect 10428 12434 10456 13126
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10520 12646 10548 12922
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10428 12406 10548 12434
rect 10520 12170 10548 12406
rect 10612 12238 10640 13670
rect 10888 13258 10916 13670
rect 10980 13462 11008 13806
rect 10968 13456 11020 13462
rect 10968 13398 11020 13404
rect 10980 13326 11008 13398
rect 10968 13320 11020 13326
rect 11164 13308 11192 14826
rect 10968 13262 11020 13268
rect 11072 13280 11192 13308
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10690 13152 10746 13161
rect 10690 13087 10746 13096
rect 10704 12850 10732 13087
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10784 12640 10836 12646
rect 10782 12608 10784 12617
rect 10836 12608 10838 12617
rect 10782 12543 10838 12552
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 11072 12170 11100 13280
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12850 11192 13126
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11164 12753 11192 12786
rect 11150 12744 11206 12753
rect 11150 12679 11206 12688
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 10520 11762 10548 12106
rect 11256 12102 11284 16526
rect 11348 15978 11376 16646
rect 11440 16522 11468 17138
rect 11428 16516 11480 16522
rect 11428 16458 11480 16464
rect 11440 16250 11468 16458
rect 11532 16425 11560 17546
rect 11624 16726 11652 20975
rect 11702 20768 11758 20777
rect 11702 20703 11758 20712
rect 11716 19174 11744 20703
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11702 18864 11758 18873
rect 11702 18799 11758 18808
rect 11716 18329 11744 18799
rect 11702 18320 11758 18329
rect 11702 18255 11758 18264
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11716 17678 11744 17818
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11716 16726 11744 17274
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11518 16416 11574 16425
rect 11518 16351 11574 16360
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11624 16114 11652 16186
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 11624 15638 11652 16050
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11808 15552 11836 24278
rect 11900 23361 11928 25638
rect 11980 24744 12032 24750
rect 11980 24686 12032 24692
rect 11992 23497 12020 24686
rect 11978 23488 12034 23497
rect 11978 23423 12034 23432
rect 11886 23352 11942 23361
rect 11886 23287 11942 23296
rect 12084 23118 12112 25758
rect 12268 25430 12296 25842
rect 12256 25424 12308 25430
rect 12256 25366 12308 25372
rect 12728 24206 12756 26182
rect 12820 25140 12848 30738
rect 12900 30592 12952 30598
rect 12900 30534 12952 30540
rect 12912 25906 12940 30534
rect 12992 29300 13044 29306
rect 13188 29288 13216 32166
rect 13556 32026 13584 32302
rect 13634 32263 13690 32272
rect 13648 32230 13676 32263
rect 13636 32224 13688 32230
rect 13636 32166 13688 32172
rect 13740 32042 13768 32710
rect 13544 32020 13596 32026
rect 13544 31962 13596 31968
rect 13648 32014 13768 32042
rect 13648 31890 13676 32014
rect 13636 31884 13688 31890
rect 13636 31826 13688 31832
rect 13648 31754 13676 31826
rect 13648 31726 13768 31754
rect 13450 31512 13506 31521
rect 13450 31447 13506 31456
rect 13360 30728 13412 30734
rect 13360 30670 13412 30676
rect 13044 29260 13216 29288
rect 12992 29242 13044 29248
rect 12992 29164 13044 29170
rect 12992 29106 13044 29112
rect 13004 27470 13032 29106
rect 13268 29096 13320 29102
rect 13266 29064 13268 29073
rect 13320 29064 13322 29073
rect 13266 28999 13322 29008
rect 13084 28960 13136 28966
rect 13082 28928 13084 28937
rect 13136 28928 13138 28937
rect 13082 28863 13138 28872
rect 13176 28688 13228 28694
rect 13176 28630 13228 28636
rect 13084 27940 13136 27946
rect 13084 27882 13136 27888
rect 13096 27538 13124 27882
rect 13084 27532 13136 27538
rect 13084 27474 13136 27480
rect 12992 27464 13044 27470
rect 12992 27406 13044 27412
rect 13004 27062 13032 27406
rect 13084 27396 13136 27402
rect 13084 27338 13136 27344
rect 12992 27056 13044 27062
rect 12992 26998 13044 27004
rect 13096 26042 13124 27338
rect 13084 26036 13136 26042
rect 13084 25978 13136 25984
rect 12900 25900 12952 25906
rect 12900 25842 12952 25848
rect 13084 25900 13136 25906
rect 13084 25842 13136 25848
rect 12992 25832 13044 25838
rect 12992 25774 13044 25780
rect 13004 25362 13032 25774
rect 12992 25356 13044 25362
rect 12992 25298 13044 25304
rect 12820 25112 12940 25140
rect 12808 24404 12860 24410
rect 12808 24346 12860 24352
rect 12716 24200 12768 24206
rect 12716 24142 12768 24148
rect 12716 23792 12768 23798
rect 12820 23780 12848 24346
rect 12912 24206 12940 25112
rect 12900 24200 12952 24206
rect 12898 24168 12900 24177
rect 12952 24168 12954 24177
rect 12898 24103 12954 24112
rect 12768 23752 12848 23780
rect 12716 23734 12768 23740
rect 12728 23322 12756 23734
rect 13096 23594 13124 25842
rect 13188 25702 13216 28630
rect 13268 28008 13320 28014
rect 13268 27950 13320 27956
rect 13280 27538 13308 27950
rect 13268 27532 13320 27538
rect 13268 27474 13320 27480
rect 13280 27130 13308 27474
rect 13268 27124 13320 27130
rect 13268 27066 13320 27072
rect 13266 27024 13322 27033
rect 13266 26959 13268 26968
rect 13320 26959 13322 26968
rect 13268 26930 13320 26936
rect 13176 25696 13228 25702
rect 13268 25696 13320 25702
rect 13176 25638 13228 25644
rect 13266 25664 13268 25673
rect 13320 25664 13322 25673
rect 13266 25599 13322 25608
rect 13372 24800 13400 30670
rect 13464 30190 13492 31447
rect 13636 30592 13688 30598
rect 13636 30534 13688 30540
rect 13452 30184 13504 30190
rect 13452 30126 13504 30132
rect 13648 29850 13676 30534
rect 13740 30122 13768 31726
rect 13820 30184 13872 30190
rect 13820 30126 13872 30132
rect 13728 30116 13780 30122
rect 13728 30058 13780 30064
rect 13740 30025 13768 30058
rect 13726 30016 13782 30025
rect 13726 29951 13782 29960
rect 13636 29844 13688 29850
rect 13636 29786 13688 29792
rect 13728 29844 13780 29850
rect 13728 29786 13780 29792
rect 13452 29776 13504 29782
rect 13452 29718 13504 29724
rect 13464 27878 13492 29718
rect 13648 29646 13676 29786
rect 13740 29714 13768 29786
rect 13728 29708 13780 29714
rect 13728 29650 13780 29656
rect 13636 29640 13688 29646
rect 13636 29582 13688 29588
rect 13544 29164 13596 29170
rect 13544 29106 13596 29112
rect 13636 29164 13688 29170
rect 13636 29106 13688 29112
rect 13556 29073 13584 29106
rect 13542 29064 13598 29073
rect 13542 28999 13598 29008
rect 13544 28076 13596 28082
rect 13544 28018 13596 28024
rect 13452 27872 13504 27878
rect 13452 27814 13504 27820
rect 13280 24772 13400 24800
rect 13174 24576 13230 24585
rect 13174 24511 13230 24520
rect 13188 24313 13216 24511
rect 13174 24304 13230 24313
rect 13174 24239 13230 24248
rect 13084 23588 13136 23594
rect 13084 23530 13136 23536
rect 12716 23316 12768 23322
rect 12900 23316 12952 23322
rect 12716 23258 12768 23264
rect 12820 23276 12900 23304
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 12256 23112 12308 23118
rect 12256 23054 12308 23060
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 11980 22976 12032 22982
rect 11980 22918 12032 22924
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 11900 21962 11928 22646
rect 11992 22030 12020 22918
rect 12164 22568 12216 22574
rect 12164 22510 12216 22516
rect 12176 22166 12204 22510
rect 12164 22160 12216 22166
rect 12164 22102 12216 22108
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 11888 21956 11940 21962
rect 11888 21898 11940 21904
rect 11900 21622 11928 21898
rect 11888 21616 11940 21622
rect 11888 21558 11940 21564
rect 11980 21412 12032 21418
rect 11980 21354 12032 21360
rect 11992 21321 12020 21354
rect 11978 21312 12034 21321
rect 11978 21247 12034 21256
rect 12084 21078 12112 21966
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 12072 21072 12124 21078
rect 12072 21014 12124 21020
rect 11888 20868 11940 20874
rect 11888 20810 11940 20816
rect 11900 20618 11928 20810
rect 11980 20800 12032 20806
rect 11978 20768 11980 20777
rect 12032 20768 12034 20777
rect 11978 20703 12034 20712
rect 11900 20590 12020 20618
rect 11888 20460 11940 20466
rect 11888 20402 11940 20408
rect 11900 18630 11928 20402
rect 11992 19281 12020 20590
rect 12084 19378 12112 21014
rect 12176 19854 12204 21490
rect 12268 21078 12296 23054
rect 12636 22982 12664 23054
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12438 22672 12494 22681
rect 12820 22642 12848 23276
rect 12900 23258 12952 23264
rect 13174 23216 13230 23225
rect 13174 23151 13230 23160
rect 13084 23044 13136 23050
rect 13084 22986 13136 22992
rect 12992 22976 13044 22982
rect 12992 22918 13044 22924
rect 12438 22607 12440 22616
rect 12492 22607 12494 22616
rect 12808 22636 12860 22642
rect 12440 22578 12492 22584
rect 12808 22578 12860 22584
rect 12716 22432 12768 22438
rect 12820 22420 12848 22578
rect 12768 22392 12848 22420
rect 12716 22374 12768 22380
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12452 21554 12480 21966
rect 12532 21956 12584 21962
rect 12584 21916 12664 21944
rect 12532 21898 12584 21904
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12530 21448 12586 21457
rect 12530 21383 12586 21392
rect 12346 21312 12402 21321
rect 12346 21247 12402 21256
rect 12256 21072 12308 21078
rect 12254 21040 12256 21049
rect 12308 21040 12310 21049
rect 12254 20975 12310 20984
rect 12256 20936 12308 20942
rect 12360 20924 12388 21247
rect 12544 21128 12572 21383
rect 12452 21100 12572 21128
rect 12452 21010 12480 21100
rect 12530 21040 12586 21049
rect 12440 21004 12492 21010
rect 12530 20975 12586 20984
rect 12440 20946 12492 20952
rect 12308 20896 12388 20924
rect 12256 20878 12308 20884
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 12176 19514 12204 19790
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 11978 19272 12034 19281
rect 11978 19207 12034 19216
rect 11980 18896 12032 18902
rect 11980 18838 12032 18844
rect 11888 18624 11940 18630
rect 11888 18566 11940 18572
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11900 18272 11928 18362
rect 11992 18290 12020 18838
rect 11980 18284 12032 18290
rect 11900 18244 11980 18272
rect 11900 17610 11928 18244
rect 11980 18226 12032 18232
rect 11980 17672 12032 17678
rect 12084 17660 12112 19314
rect 12164 19236 12216 19242
rect 12164 19178 12216 19184
rect 12176 18766 12204 19178
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 12176 18290 12204 18566
rect 12268 18306 12296 20878
rect 12440 20868 12492 20874
rect 12440 20810 12492 20816
rect 12452 20602 12480 20810
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12452 18834 12480 19450
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12348 18692 12400 18698
rect 12348 18634 12400 18640
rect 12360 18426 12388 18634
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12164 18284 12216 18290
rect 12268 18278 12480 18306
rect 12164 18226 12216 18232
rect 12176 18086 12204 18226
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12032 17632 12112 17660
rect 11980 17614 12032 17620
rect 11888 17604 11940 17610
rect 11888 17546 11940 17552
rect 11900 17218 11928 17546
rect 12084 17524 12112 17632
rect 12164 17536 12216 17542
rect 12084 17496 12164 17524
rect 12452 17490 12480 18278
rect 12164 17478 12216 17484
rect 12268 17462 12480 17490
rect 11900 17190 12020 17218
rect 11992 17184 12020 17190
rect 11992 17156 12204 17184
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 11900 16114 11928 17070
rect 11978 16416 12034 16425
rect 11978 16351 12034 16360
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11808 15524 11844 15552
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11624 14958 11652 15098
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11716 14890 11744 15438
rect 11816 15416 11844 15524
rect 11808 15388 11844 15416
rect 11808 15348 11836 15388
rect 11992 15366 12020 16351
rect 12176 16182 12204 17156
rect 12164 16176 12216 16182
rect 12164 16118 12216 16124
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 11980 15360 12032 15366
rect 11808 15320 11928 15348
rect 11900 15026 11928 15320
rect 11980 15302 12032 15308
rect 11992 15162 12020 15302
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11704 14884 11756 14890
rect 11704 14826 11756 14832
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11532 13462 11560 14758
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11520 13456 11572 13462
rect 11520 13398 11572 13404
rect 11532 13326 11560 13398
rect 11716 13326 11744 14418
rect 11794 13696 11850 13705
rect 11794 13631 11850 13640
rect 11808 13530 11836 13631
rect 11900 13530 11928 14962
rect 11992 14074 12020 14962
rect 12084 14822 12112 16050
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12176 15065 12204 15098
rect 12162 15056 12218 15065
rect 12162 14991 12218 15000
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 11978 13968 12034 13977
rect 11978 13903 11980 13912
rect 12032 13903 12034 13912
rect 11980 13874 12032 13880
rect 12084 13841 12112 14010
rect 12164 13864 12216 13870
rect 12070 13832 12126 13841
rect 12164 13806 12216 13812
rect 12070 13767 12126 13776
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 11992 13326 12020 13398
rect 12176 13326 12204 13806
rect 12268 13433 12296 17462
rect 12544 17320 12572 20975
rect 12636 20806 12664 21916
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12728 21554 12756 21830
rect 12820 21690 12848 21830
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 12820 21078 12848 21626
rect 12808 21072 12860 21078
rect 13004 21049 13032 22918
rect 13096 21321 13124 22986
rect 13188 22438 13216 23151
rect 13176 22432 13228 22438
rect 13176 22374 13228 22380
rect 13082 21312 13138 21321
rect 13082 21247 13138 21256
rect 13084 21140 13136 21146
rect 13188 21128 13216 22374
rect 13280 21554 13308 24772
rect 13360 24676 13412 24682
rect 13360 24618 13412 24624
rect 13372 24410 13400 24618
rect 13360 24404 13412 24410
rect 13360 24346 13412 24352
rect 13358 22808 13414 22817
rect 13358 22743 13360 22752
rect 13412 22743 13414 22752
rect 13360 22714 13412 22720
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13280 21457 13308 21490
rect 13266 21448 13322 21457
rect 13266 21383 13322 21392
rect 13372 21321 13400 22714
rect 13358 21312 13414 21321
rect 13358 21247 13414 21256
rect 13464 21146 13492 27814
rect 13556 23730 13584 28018
rect 13648 27962 13676 29106
rect 13740 29102 13768 29650
rect 13728 29096 13780 29102
rect 13728 29038 13780 29044
rect 13728 28688 13780 28694
rect 13832 28665 13860 30126
rect 14280 29640 14332 29646
rect 14280 29582 14332 29588
rect 14096 29504 14148 29510
rect 14096 29446 14148 29452
rect 13728 28630 13780 28636
rect 13818 28656 13874 28665
rect 13740 28257 13768 28630
rect 13818 28591 13874 28600
rect 13726 28248 13782 28257
rect 13726 28183 13782 28192
rect 13648 27934 13768 27962
rect 13636 27872 13688 27878
rect 13634 27840 13636 27849
rect 13688 27840 13690 27849
rect 13634 27775 13690 27784
rect 13634 27160 13690 27169
rect 13634 27095 13690 27104
rect 13648 27062 13676 27095
rect 13636 27056 13688 27062
rect 13636 26998 13688 27004
rect 13648 25906 13676 26998
rect 13740 26790 13768 27934
rect 13728 26784 13780 26790
rect 13728 26726 13780 26732
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13636 24948 13688 24954
rect 13636 24890 13688 24896
rect 13648 24818 13676 24890
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13634 24304 13690 24313
rect 13634 24239 13690 24248
rect 13648 23730 13676 24239
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 13636 23588 13688 23594
rect 13636 23530 13688 23536
rect 13544 22500 13596 22506
rect 13544 22442 13596 22448
rect 13556 22234 13584 22442
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 13136 21100 13216 21128
rect 13268 21140 13320 21146
rect 13084 21082 13136 21088
rect 13268 21082 13320 21088
rect 13452 21140 13504 21146
rect 13452 21082 13504 21088
rect 12808 21014 12860 21020
rect 12990 21040 13046 21049
rect 12990 20975 13046 20984
rect 12808 20936 12860 20942
rect 12728 20896 12808 20924
rect 12624 20800 12676 20806
rect 12622 20768 12624 20777
rect 12676 20768 12678 20777
rect 12622 20703 12678 20712
rect 12728 20058 12756 20896
rect 12808 20878 12860 20884
rect 12806 20768 12862 20777
rect 12806 20703 12862 20712
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 12728 19378 12756 19994
rect 12820 19514 12848 20703
rect 12898 19544 12954 19553
rect 12808 19508 12860 19514
rect 12898 19479 12954 19488
rect 12808 19450 12860 19456
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12714 19272 12770 19281
rect 12624 19236 12676 19242
rect 12714 19207 12770 19216
rect 12624 19178 12676 19184
rect 12636 18290 12664 19178
rect 12728 18834 12756 19207
rect 12820 18902 12848 19450
rect 12912 19009 12940 19479
rect 12898 19000 12954 19009
rect 12898 18935 12954 18944
rect 12808 18896 12860 18902
rect 12808 18838 12860 18844
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12716 18692 12768 18698
rect 12716 18634 12768 18640
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12452 17292 12572 17320
rect 12348 16108 12400 16114
rect 12348 16050 12400 16056
rect 12360 15434 12388 16050
rect 12348 15428 12400 15434
rect 12348 15370 12400 15376
rect 12452 14113 12480 17292
rect 12636 17270 12664 17818
rect 12728 17524 12756 18634
rect 12808 18216 12860 18222
rect 12808 18158 12860 18164
rect 12820 17649 12848 18158
rect 12912 17746 12940 18935
rect 13004 18222 13032 20975
rect 13176 20868 13228 20874
rect 13176 20810 13228 20816
rect 13188 20641 13216 20810
rect 13174 20632 13230 20641
rect 13280 20602 13308 21082
rect 13358 21040 13414 21049
rect 13358 20975 13414 20984
rect 13372 20942 13400 20975
rect 13556 20942 13584 21830
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 13452 20868 13504 20874
rect 13452 20810 13504 20816
rect 13464 20777 13492 20810
rect 13544 20800 13596 20806
rect 13450 20768 13506 20777
rect 13544 20742 13596 20748
rect 13450 20703 13506 20712
rect 13174 20567 13230 20576
rect 13268 20596 13320 20602
rect 13268 20538 13320 20544
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13176 20528 13228 20534
rect 13082 20496 13138 20505
rect 13176 20470 13228 20476
rect 13082 20431 13084 20440
rect 13136 20431 13138 20440
rect 13084 20402 13136 20408
rect 13084 19984 13136 19990
rect 13084 19926 13136 19932
rect 13096 19854 13124 19926
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 13004 18086 13032 18158
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 12990 17776 13046 17785
rect 12900 17740 12952 17746
rect 12990 17711 13046 17720
rect 12900 17682 12952 17688
rect 13004 17678 13032 17711
rect 12992 17672 13044 17678
rect 12806 17640 12862 17649
rect 12992 17614 13044 17620
rect 12806 17575 12862 17584
rect 12728 17496 12848 17524
rect 12624 17264 12676 17270
rect 12530 17232 12586 17241
rect 12624 17206 12676 17212
rect 12530 17167 12586 17176
rect 12438 14104 12494 14113
rect 12438 14039 12494 14048
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12254 13424 12310 13433
rect 12254 13359 12310 13368
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 11610 13016 11666 13025
rect 11610 12951 11612 12960
rect 11664 12951 11666 12960
rect 11612 12922 11664 12928
rect 11624 12481 11652 12922
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 11610 12472 11666 12481
rect 11610 12407 11666 12416
rect 12176 12306 12204 12786
rect 12268 12782 12296 13359
rect 12360 13326 12388 13738
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12452 12986 12480 14039
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12452 12850 12480 12922
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12256 12776 12308 12782
rect 12544 12753 12572 17167
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12636 15706 12664 16050
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12636 14618 12664 15642
rect 12728 15638 12756 16594
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 12820 15570 12848 17496
rect 12990 17232 13046 17241
rect 12990 17167 12992 17176
rect 13044 17167 13046 17176
rect 12992 17138 13044 17144
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12912 15881 12940 16934
rect 12992 16516 13044 16522
rect 12992 16458 13044 16464
rect 13004 16114 13032 16458
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13004 15978 13032 16050
rect 12992 15972 13044 15978
rect 12992 15914 13044 15920
rect 12898 15872 12954 15881
rect 12898 15807 12954 15816
rect 12900 15632 12952 15638
rect 12900 15574 12952 15580
rect 12992 15632 13044 15638
rect 12992 15574 13044 15580
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12912 15502 12940 15574
rect 12716 15496 12768 15502
rect 12714 15464 12716 15473
rect 12900 15496 12952 15502
rect 12768 15464 12770 15473
rect 13004 15473 13032 15574
rect 12900 15438 12952 15444
rect 12990 15464 13046 15473
rect 12714 15399 12770 15408
rect 12808 15428 12860 15434
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12728 14006 12756 15399
rect 12808 15370 12860 15376
rect 12820 15201 12848 15370
rect 12806 15192 12862 15201
rect 12806 15127 12862 15136
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12636 13394 12664 13466
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12728 13326 12756 13942
rect 12912 13938 12940 15438
rect 12990 15399 13046 15408
rect 13096 15094 13124 19790
rect 13188 18698 13216 20470
rect 13372 20058 13400 20538
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13266 19544 13322 19553
rect 13266 19479 13322 19488
rect 13280 19310 13308 19479
rect 13268 19304 13320 19310
rect 13268 19246 13320 19252
rect 13464 18902 13492 20703
rect 13556 19378 13584 20742
rect 13648 20398 13676 23530
rect 13740 22001 13768 26726
rect 13832 26382 13860 28591
rect 14004 26444 14056 26450
rect 14004 26386 14056 26392
rect 13820 26376 13872 26382
rect 13820 26318 13872 26324
rect 13832 24818 13860 26318
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13832 24410 13860 24754
rect 13912 24676 13964 24682
rect 13912 24618 13964 24624
rect 13820 24404 13872 24410
rect 13820 24346 13872 24352
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13832 23633 13860 24006
rect 13924 23905 13952 24618
rect 13910 23896 13966 23905
rect 13910 23831 13966 23840
rect 13912 23724 13964 23730
rect 13912 23666 13964 23672
rect 13818 23624 13874 23633
rect 13818 23559 13874 23568
rect 13820 22568 13872 22574
rect 13820 22510 13872 22516
rect 13832 22409 13860 22510
rect 13818 22400 13874 22409
rect 13818 22335 13874 22344
rect 13924 22166 13952 23666
rect 14016 22166 14044 26386
rect 14108 24274 14136 29446
rect 14292 28937 14320 29582
rect 14278 28928 14334 28937
rect 14278 28863 14334 28872
rect 14292 28082 14320 28863
rect 14280 28076 14332 28082
rect 14280 28018 14332 28024
rect 14280 25152 14332 25158
rect 14280 25094 14332 25100
rect 14188 24404 14240 24410
rect 14188 24346 14240 24352
rect 14200 24274 14228 24346
rect 14096 24268 14148 24274
rect 14096 24210 14148 24216
rect 14188 24268 14240 24274
rect 14188 24210 14240 24216
rect 14292 24177 14320 25094
rect 14384 24818 14412 34682
rect 22192 34604 22244 34610
rect 22192 34546 22244 34552
rect 22204 34066 22232 34546
rect 16304 34060 16356 34066
rect 16304 34002 16356 34008
rect 22192 34060 22244 34066
rect 22192 34002 22244 34008
rect 14832 32564 14884 32570
rect 14832 32506 14884 32512
rect 14554 31376 14610 31385
rect 14554 31311 14556 31320
rect 14608 31311 14610 31320
rect 14740 31340 14792 31346
rect 14556 31282 14608 31288
rect 14740 31282 14792 31288
rect 14568 30938 14596 31282
rect 14556 30932 14608 30938
rect 14556 30874 14608 30880
rect 14752 30666 14780 31282
rect 14464 30660 14516 30666
rect 14464 30602 14516 30608
rect 14740 30660 14792 30666
rect 14740 30602 14792 30608
rect 14476 30569 14504 30602
rect 14462 30560 14518 30569
rect 14462 30495 14518 30504
rect 14476 30394 14504 30495
rect 14464 30388 14516 30394
rect 14464 30330 14516 30336
rect 14556 30048 14608 30054
rect 14556 29990 14608 29996
rect 14464 29708 14516 29714
rect 14464 29650 14516 29656
rect 14476 28150 14504 29650
rect 14568 29646 14596 29990
rect 14556 29640 14608 29646
rect 14556 29582 14608 29588
rect 14740 29504 14792 29510
rect 14740 29446 14792 29452
rect 14464 28144 14516 28150
rect 14464 28086 14516 28092
rect 14556 27532 14608 27538
rect 14556 27474 14608 27480
rect 14464 26580 14516 26586
rect 14464 26522 14516 26528
rect 14372 24812 14424 24818
rect 14372 24754 14424 24760
rect 14384 24721 14412 24754
rect 14370 24712 14426 24721
rect 14370 24647 14426 24656
rect 14372 24608 14424 24614
rect 14372 24550 14424 24556
rect 14384 24410 14412 24550
rect 14372 24404 14424 24410
rect 14372 24346 14424 24352
rect 14278 24168 14334 24177
rect 14278 24103 14280 24112
rect 14332 24103 14334 24112
rect 14280 24074 14332 24080
rect 14096 24064 14148 24070
rect 14096 24006 14148 24012
rect 13912 22160 13964 22166
rect 13818 22128 13874 22137
rect 13912 22102 13964 22108
rect 14004 22160 14056 22166
rect 14004 22102 14056 22108
rect 13818 22063 13874 22072
rect 13726 21992 13782 22001
rect 13726 21927 13782 21936
rect 13832 21706 13860 22063
rect 13832 21678 13952 21706
rect 13728 21616 13780 21622
rect 13728 21558 13780 21564
rect 13740 20924 13768 21558
rect 13820 20936 13872 20942
rect 13740 20896 13820 20924
rect 13740 20466 13768 20896
rect 13820 20878 13872 20884
rect 13924 20466 13952 21678
rect 14108 21078 14136 24006
rect 14280 23860 14332 23866
rect 14280 23802 14332 23808
rect 14186 23352 14242 23361
rect 14186 23287 14242 23296
rect 14200 22817 14228 23287
rect 14186 22808 14242 22817
rect 14186 22743 14242 22752
rect 14200 22574 14228 22743
rect 14188 22568 14240 22574
rect 14188 22510 14240 22516
rect 14292 22420 14320 23802
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14384 22506 14412 22578
rect 14372 22500 14424 22506
rect 14372 22442 14424 22448
rect 14200 22392 14320 22420
rect 14096 21072 14148 21078
rect 14096 21014 14148 21020
rect 14004 21004 14056 21010
rect 14004 20946 14056 20952
rect 13728 20460 13780 20466
rect 13912 20460 13964 20466
rect 13780 20420 13860 20448
rect 13728 20402 13780 20408
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 13648 20058 13676 20334
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13832 19990 13860 20420
rect 13912 20402 13964 20408
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 13820 19984 13872 19990
rect 13820 19926 13872 19932
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13360 18896 13412 18902
rect 13360 18838 13412 18844
rect 13452 18896 13504 18902
rect 13452 18838 13504 18844
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 13176 18692 13228 18698
rect 13176 18634 13228 18640
rect 13188 18290 13216 18634
rect 13280 18426 13308 18770
rect 13372 18426 13400 18838
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13268 18420 13320 18426
rect 13268 18362 13320 18368
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 13464 18358 13492 18566
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 13372 17610 13400 18226
rect 13556 17882 13584 19314
rect 13740 19242 13768 19926
rect 13832 19786 13860 19926
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 13832 19378 13860 19722
rect 14016 19530 14044 20946
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 14108 19553 14136 20742
rect 13924 19502 14044 19530
rect 14094 19544 14150 19553
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 13544 17876 13596 17882
rect 13544 17818 13596 17824
rect 13360 17604 13412 17610
rect 13360 17546 13412 17552
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13188 17202 13216 17478
rect 13266 17368 13322 17377
rect 13266 17303 13322 17312
rect 13280 17202 13308 17303
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13280 15994 13308 17138
rect 13188 15966 13308 15994
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 13082 13968 13138 13977
rect 12900 13932 12952 13938
rect 13082 13903 13138 13912
rect 12900 13874 12952 13880
rect 12912 13326 12940 13874
rect 13096 13530 13124 13903
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12256 12718 12308 12724
rect 12530 12744 12586 12753
rect 12268 12442 12296 12718
rect 12530 12679 12586 12688
rect 12990 12744 13046 12753
rect 12990 12679 13046 12688
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 13004 12306 13032 12679
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 12900 12164 12952 12170
rect 13084 12164 13136 12170
rect 12952 12124 13084 12152
rect 12900 12106 12952 12112
rect 13084 12106 13136 12112
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 13188 11762 13216 15966
rect 13268 15904 13320 15910
rect 13266 15872 13268 15881
rect 13320 15872 13322 15881
rect 13266 15807 13322 15816
rect 13280 14521 13308 15807
rect 13266 14512 13322 14521
rect 13372 14482 13400 17546
rect 13542 17368 13598 17377
rect 13542 17303 13598 17312
rect 13556 17066 13584 17303
rect 13648 17184 13676 18702
rect 13924 18442 13952 19502
rect 14094 19479 14150 19488
rect 14108 19360 14136 19479
rect 13832 18414 13952 18442
rect 14016 19332 14136 19360
rect 13728 17808 13780 17814
rect 13726 17776 13728 17785
rect 13780 17776 13782 17785
rect 13726 17711 13782 17720
rect 13728 17196 13780 17202
rect 13648 17156 13728 17184
rect 13728 17138 13780 17144
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13740 15910 13768 17138
rect 13832 16833 13860 18414
rect 13912 18352 13964 18358
rect 13912 18294 13964 18300
rect 13924 17202 13952 18294
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 13818 16824 13874 16833
rect 13818 16759 13874 16768
rect 13924 16425 13952 17138
rect 13910 16416 13966 16425
rect 13910 16351 13966 16360
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13924 15434 13952 16351
rect 13728 15428 13780 15434
rect 13728 15370 13780 15376
rect 13912 15428 13964 15434
rect 13912 15370 13964 15376
rect 13740 15162 13768 15370
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13924 14482 13952 15370
rect 14016 15094 14044 19332
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 14108 18086 14136 18226
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 14108 16998 14136 17138
rect 14200 17066 14228 22392
rect 14280 22160 14332 22166
rect 14280 22102 14332 22108
rect 14188 17060 14240 17066
rect 14188 17002 14240 17008
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14108 15586 14136 16934
rect 14108 15558 14228 15586
rect 14200 15502 14228 15558
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 14004 15088 14056 15094
rect 14004 15030 14056 15036
rect 13266 14447 13322 14456
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 13832 13462 13860 13738
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13636 13320 13688 13326
rect 13266 13288 13322 13297
rect 13636 13262 13688 13268
rect 13266 13223 13322 13232
rect 13452 13252 13504 13258
rect 13280 12918 13308 13223
rect 13452 13194 13504 13200
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 13464 12753 13492 13194
rect 13648 13161 13676 13262
rect 13634 13152 13690 13161
rect 13634 13087 13690 13096
rect 13832 12850 13860 13398
rect 13924 13190 13952 13466
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 14016 12918 14044 15030
rect 14004 12912 14056 12918
rect 14004 12854 14056 12860
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13450 12744 13506 12753
rect 14108 12714 14136 15438
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 14200 13802 14228 14350
rect 14188 13796 14240 13802
rect 14188 13738 14240 13744
rect 14188 13456 14240 13462
rect 14188 13398 14240 13404
rect 13450 12679 13452 12688
rect 13504 12679 13506 12688
rect 14096 12708 14148 12714
rect 13452 12650 13504 12656
rect 14096 12650 14148 12656
rect 14200 12646 14228 13398
rect 14292 13190 14320 22102
rect 14384 21690 14412 22442
rect 14372 21684 14424 21690
rect 14372 21626 14424 21632
rect 14476 21457 14504 26522
rect 14568 26450 14596 27474
rect 14752 27112 14780 29446
rect 14660 27084 14780 27112
rect 14556 26444 14608 26450
rect 14556 26386 14608 26392
rect 14660 26314 14688 27084
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14648 26308 14700 26314
rect 14648 26250 14700 26256
rect 14556 24132 14608 24138
rect 14556 24074 14608 24080
rect 14568 23866 14596 24074
rect 14556 23860 14608 23866
rect 14556 23802 14608 23808
rect 14568 23594 14596 23802
rect 14556 23588 14608 23594
rect 14556 23530 14608 23536
rect 14660 23322 14688 26250
rect 14752 25906 14780 26930
rect 14844 26586 14872 32506
rect 15844 32428 15896 32434
rect 15844 32370 15896 32376
rect 15856 32201 15884 32370
rect 16028 32360 16080 32366
rect 16028 32302 16080 32308
rect 16120 32360 16172 32366
rect 16120 32302 16172 32308
rect 15936 32224 15988 32230
rect 15842 32192 15898 32201
rect 15936 32166 15988 32172
rect 15842 32127 15898 32136
rect 15200 31340 15252 31346
rect 15200 31282 15252 31288
rect 15476 31340 15528 31346
rect 15476 31282 15528 31288
rect 15212 30977 15240 31282
rect 15488 31249 15516 31282
rect 15474 31240 15530 31249
rect 15474 31175 15530 31184
rect 15292 31136 15344 31142
rect 15292 31078 15344 31084
rect 15198 30968 15254 30977
rect 15198 30903 15254 30912
rect 15212 29578 15240 30903
rect 15200 29572 15252 29578
rect 15200 29514 15252 29520
rect 14924 28416 14976 28422
rect 14924 28358 14976 28364
rect 14936 27878 14964 28358
rect 15014 28112 15070 28121
rect 15014 28047 15016 28056
rect 15068 28047 15070 28056
rect 15200 28076 15252 28082
rect 15016 28018 15068 28024
rect 15200 28018 15252 28024
rect 14924 27872 14976 27878
rect 14924 27814 14976 27820
rect 15016 27872 15068 27878
rect 15016 27814 15068 27820
rect 15028 26994 15056 27814
rect 15212 27538 15240 28018
rect 15200 27532 15252 27538
rect 15200 27474 15252 27480
rect 15108 27328 15160 27334
rect 15108 27270 15160 27276
rect 15120 27130 15148 27270
rect 15108 27124 15160 27130
rect 15108 27066 15160 27072
rect 15016 26988 15068 26994
rect 15016 26930 15068 26936
rect 15200 26988 15252 26994
rect 15200 26930 15252 26936
rect 15212 26625 15240 26930
rect 15198 26616 15254 26625
rect 14832 26580 14884 26586
rect 15198 26551 15254 26560
rect 14832 26522 14884 26528
rect 15304 26450 15332 31078
rect 15488 30433 15516 31175
rect 15660 30728 15712 30734
rect 15660 30670 15712 30676
rect 15474 30424 15530 30433
rect 15474 30359 15530 30368
rect 15474 30288 15530 30297
rect 15474 30223 15530 30232
rect 15488 28121 15516 30223
rect 15568 28212 15620 28218
rect 15568 28154 15620 28160
rect 15474 28112 15530 28121
rect 15474 28047 15476 28056
rect 15528 28047 15530 28056
rect 15476 28018 15528 28024
rect 15580 28014 15608 28154
rect 15568 28008 15620 28014
rect 15568 27950 15620 27956
rect 15384 27396 15436 27402
rect 15384 27338 15436 27344
rect 15292 26444 15344 26450
rect 15292 26386 15344 26392
rect 14924 26376 14976 26382
rect 14924 26318 14976 26324
rect 14830 26208 14886 26217
rect 14830 26143 14886 26152
rect 14844 25906 14872 26143
rect 14740 25900 14792 25906
rect 14740 25842 14792 25848
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 14648 23316 14700 23322
rect 14648 23258 14700 23264
rect 14646 22672 14702 22681
rect 14556 22636 14608 22642
rect 14646 22607 14702 22616
rect 14556 22578 14608 22584
rect 14568 22234 14596 22578
rect 14556 22228 14608 22234
rect 14556 22170 14608 22176
rect 14556 21956 14608 21962
rect 14556 21898 14608 21904
rect 14568 21622 14596 21898
rect 14556 21616 14608 21622
rect 14556 21558 14608 21564
rect 14462 21448 14518 21457
rect 14462 21383 14518 21392
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14476 20040 14504 20878
rect 14568 20602 14596 21558
rect 14660 21298 14688 22607
rect 14752 21978 14780 25842
rect 14936 24342 14964 26318
rect 15106 25800 15162 25809
rect 15106 25735 15108 25744
rect 15160 25735 15162 25744
rect 15108 25706 15160 25712
rect 15200 25696 15252 25702
rect 15396 25684 15424 27338
rect 15476 27056 15528 27062
rect 15476 26998 15528 27004
rect 15488 26586 15516 26998
rect 15476 26580 15528 26586
rect 15476 26522 15528 26528
rect 15476 26376 15528 26382
rect 15474 26344 15476 26353
rect 15528 26344 15530 26353
rect 15474 26279 15530 26288
rect 15252 25656 15424 25684
rect 15200 25638 15252 25644
rect 14924 24336 14976 24342
rect 14924 24278 14976 24284
rect 14832 24268 14884 24274
rect 14832 24210 14884 24216
rect 14844 24154 14872 24210
rect 15108 24200 15160 24206
rect 15106 24168 15108 24177
rect 15160 24168 15162 24177
rect 14844 24126 14964 24154
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 14844 22778 14872 23054
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 14936 22234 14964 24126
rect 15106 24103 15162 24112
rect 15016 23724 15068 23730
rect 15016 23666 15068 23672
rect 15028 22778 15056 23666
rect 15212 23610 15240 25638
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15488 23730 15516 24346
rect 15384 23724 15436 23730
rect 15384 23666 15436 23672
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15120 23582 15240 23610
rect 15120 23322 15148 23582
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 15212 23322 15240 23462
rect 15108 23316 15160 23322
rect 15108 23258 15160 23264
rect 15200 23316 15252 23322
rect 15200 23258 15252 23264
rect 15200 23112 15252 23118
rect 15198 23080 15200 23089
rect 15252 23080 15254 23089
rect 15198 23015 15254 23024
rect 15016 22772 15068 22778
rect 15016 22714 15068 22720
rect 14924 22228 14976 22234
rect 14924 22170 14976 22176
rect 14924 22024 14976 22030
rect 14922 21992 14924 22001
rect 15016 22024 15068 22030
rect 14976 21992 14978 22001
rect 14752 21962 14872 21978
rect 14752 21956 14884 21962
rect 14752 21950 14832 21956
rect 14752 21865 14780 21950
rect 15016 21966 15068 21972
rect 14922 21927 14978 21936
rect 14832 21898 14884 21904
rect 14738 21856 14794 21865
rect 14738 21791 14794 21800
rect 14936 21729 14964 21927
rect 14922 21720 14978 21729
rect 14922 21655 14978 21664
rect 14832 21480 14884 21486
rect 14832 21422 14884 21428
rect 14924 21480 14976 21486
rect 14924 21422 14976 21428
rect 14660 21270 14780 21298
rect 14648 21140 14700 21146
rect 14648 21082 14700 21088
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 14660 20262 14688 21082
rect 14752 20942 14780 21270
rect 14740 20936 14792 20942
rect 14740 20878 14792 20884
rect 14844 20806 14872 21422
rect 14936 21350 14964 21422
rect 15028 21350 15056 21966
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 15028 21078 15056 21286
rect 15016 21072 15068 21078
rect 15016 21014 15068 21020
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 15108 20868 15160 20874
rect 15108 20810 15160 20816
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14752 20058 14780 20402
rect 14740 20052 14792 20058
rect 14476 20012 14688 20040
rect 14476 19922 14504 20012
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 14370 19544 14426 19553
rect 14370 19479 14426 19488
rect 14384 19446 14412 19479
rect 14372 19440 14424 19446
rect 14372 19382 14424 19388
rect 14568 19310 14596 19858
rect 14660 19446 14688 20012
rect 14740 19994 14792 20000
rect 14844 19904 14872 20742
rect 14924 20256 14976 20262
rect 14924 20198 14976 20204
rect 14752 19876 14872 19904
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 14556 19304 14608 19310
rect 14556 19246 14608 19252
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14372 18692 14424 18698
rect 14372 18634 14424 18640
rect 14384 16998 14412 18634
rect 14476 17542 14504 18702
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14476 17270 14504 17478
rect 14464 17264 14516 17270
rect 14464 17206 14516 17212
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14384 15638 14412 16934
rect 14372 15632 14424 15638
rect 14372 15574 14424 15580
rect 14384 15434 14412 15574
rect 14372 15428 14424 15434
rect 14372 15370 14424 15376
rect 14568 15026 14596 19246
rect 14660 18766 14688 19382
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14752 18290 14780 19876
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14844 18766 14872 19314
rect 14936 18834 14964 20198
rect 15120 19922 15148 20810
rect 15108 19916 15160 19922
rect 15304 19904 15332 20878
rect 15396 20058 15424 23666
rect 15580 22234 15608 27950
rect 15672 27878 15700 30670
rect 15750 30288 15806 30297
rect 15856 30258 15884 32127
rect 15750 30223 15752 30232
rect 15804 30223 15806 30232
rect 15844 30252 15896 30258
rect 15752 30194 15804 30200
rect 15844 30194 15896 30200
rect 15752 30116 15804 30122
rect 15752 30058 15804 30064
rect 15660 27872 15712 27878
rect 15660 27814 15712 27820
rect 15660 26988 15712 26994
rect 15660 26930 15712 26936
rect 15672 26586 15700 26930
rect 15660 26580 15712 26586
rect 15660 26522 15712 26528
rect 15764 26246 15792 30058
rect 15948 28778 15976 32166
rect 16040 31278 16068 32302
rect 16132 31822 16160 32302
rect 16120 31816 16172 31822
rect 16120 31758 16172 31764
rect 16028 31272 16080 31278
rect 16028 31214 16080 31220
rect 16028 30048 16080 30054
rect 16028 29990 16080 29996
rect 16040 29850 16068 29990
rect 16028 29844 16080 29850
rect 16028 29786 16080 29792
rect 15948 28750 16252 28778
rect 16120 28688 16172 28694
rect 16120 28630 16172 28636
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 15856 27441 15884 28018
rect 16028 28008 16080 28014
rect 16028 27950 16080 27956
rect 15842 27432 15898 27441
rect 15842 27367 15898 27376
rect 15936 27396 15988 27402
rect 15936 27338 15988 27344
rect 15948 27033 15976 27338
rect 15934 27024 15990 27033
rect 15856 26982 15934 27010
rect 15752 26240 15804 26246
rect 15752 26182 15804 26188
rect 15752 25900 15804 25906
rect 15752 25842 15804 25848
rect 15660 25152 15712 25158
rect 15660 25094 15712 25100
rect 15672 24954 15700 25094
rect 15660 24948 15712 24954
rect 15660 24890 15712 24896
rect 15658 23896 15714 23905
rect 15658 23831 15660 23840
rect 15712 23831 15714 23840
rect 15660 23802 15712 23808
rect 15568 22228 15620 22234
rect 15568 22170 15620 22176
rect 15764 22030 15792 25842
rect 15856 22234 15884 26982
rect 15934 26959 15990 26968
rect 16040 26432 16068 27950
rect 16132 27878 16160 28630
rect 16120 27872 16172 27878
rect 16120 27814 16172 27820
rect 16132 27402 16160 27814
rect 16120 27396 16172 27402
rect 16120 27338 16172 27344
rect 15948 26404 16068 26432
rect 15948 24993 15976 26404
rect 16224 26194 16252 28750
rect 16316 28218 16344 34002
rect 21640 33992 21692 33998
rect 21640 33934 21692 33940
rect 21916 33992 21968 33998
rect 21916 33934 21968 33940
rect 17776 33652 17828 33658
rect 17776 33594 17828 33600
rect 17682 32056 17738 32065
rect 17224 32020 17276 32026
rect 17682 31991 17684 32000
rect 17224 31962 17276 31968
rect 17736 31991 17738 32000
rect 17684 31962 17736 31968
rect 17040 31952 17092 31958
rect 17040 31894 17092 31900
rect 16488 31272 16540 31278
rect 16488 31214 16540 31220
rect 16396 29640 16448 29646
rect 16396 29582 16448 29588
rect 16408 29034 16436 29582
rect 16396 29028 16448 29034
rect 16396 28970 16448 28976
rect 16304 28212 16356 28218
rect 16304 28154 16356 28160
rect 16396 27328 16448 27334
rect 16500 27316 16528 31214
rect 16762 30424 16818 30433
rect 16762 30359 16818 30368
rect 16776 29850 16804 30359
rect 16856 30116 16908 30122
rect 16856 30058 16908 30064
rect 16764 29844 16816 29850
rect 16764 29786 16816 29792
rect 16764 29708 16816 29714
rect 16764 29650 16816 29656
rect 16776 29617 16804 29650
rect 16762 29608 16818 29617
rect 16580 29572 16632 29578
rect 16762 29543 16764 29552
rect 16580 29514 16632 29520
rect 16816 29543 16818 29552
rect 16764 29514 16816 29520
rect 16592 28994 16620 29514
rect 16592 28966 16712 28994
rect 16684 28218 16712 28966
rect 16672 28212 16724 28218
rect 16672 28154 16724 28160
rect 16448 27288 16528 27316
rect 16396 27270 16448 27276
rect 16224 26166 16344 26194
rect 16210 26072 16266 26081
rect 16210 26007 16266 26016
rect 16028 25900 16080 25906
rect 16028 25842 16080 25848
rect 16040 25430 16068 25842
rect 16118 25528 16174 25537
rect 16118 25463 16174 25472
rect 16028 25424 16080 25430
rect 16028 25366 16080 25372
rect 15934 24984 15990 24993
rect 15934 24919 15990 24928
rect 15936 24812 15988 24818
rect 15936 24754 15988 24760
rect 15948 24274 15976 24754
rect 15936 24268 15988 24274
rect 15936 24210 15988 24216
rect 15844 22228 15896 22234
rect 15844 22170 15896 22176
rect 15844 22092 15896 22098
rect 15844 22034 15896 22040
rect 15752 22024 15804 22030
rect 15672 21984 15752 22012
rect 15476 21412 15528 21418
rect 15476 21354 15528 21360
rect 15488 21078 15516 21354
rect 15476 21072 15528 21078
rect 15476 21014 15528 21020
rect 15568 20528 15620 20534
rect 15568 20470 15620 20476
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15304 19876 15424 19904
rect 15108 19858 15160 19864
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15016 19780 15068 19786
rect 15016 19722 15068 19728
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 14922 18320 14978 18329
rect 14740 18284 14792 18290
rect 14922 18255 14924 18264
rect 14740 18226 14792 18232
rect 14976 18255 14978 18264
rect 14924 18226 14976 18232
rect 14924 17604 14976 17610
rect 14924 17546 14976 17552
rect 14646 16824 14702 16833
rect 14646 16759 14702 16768
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14568 13938 14596 14962
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14568 12986 14596 13874
rect 14660 13326 14688 16759
rect 14738 16008 14794 16017
rect 14738 15943 14794 15952
rect 14752 15502 14780 15943
rect 14936 15706 14964 17546
rect 15028 17202 15056 19722
rect 15106 19408 15162 19417
rect 15212 19378 15240 19790
rect 15106 19343 15162 19352
rect 15200 19372 15252 19378
rect 15120 19258 15148 19343
rect 15200 19314 15252 19320
rect 15292 19304 15344 19310
rect 15120 19230 15240 19258
rect 15292 19246 15344 19252
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 15120 18057 15148 18226
rect 15106 18048 15162 18057
rect 15106 17983 15162 17992
rect 15212 17882 15240 19230
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15212 17649 15240 17818
rect 15304 17678 15332 19246
rect 15396 18358 15424 19876
rect 15488 19378 15516 20334
rect 15580 19922 15608 20470
rect 15672 20466 15700 21984
rect 15752 21966 15804 21972
rect 15750 21448 15806 21457
rect 15750 21383 15806 21392
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 15672 19718 15700 20402
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 15476 19372 15528 19378
rect 15476 19314 15528 19320
rect 15488 18902 15516 19314
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15384 18352 15436 18358
rect 15384 18294 15436 18300
rect 15292 17672 15344 17678
rect 15198 17640 15254 17649
rect 15108 17604 15160 17610
rect 15292 17614 15344 17620
rect 15198 17575 15254 17584
rect 15108 17546 15160 17552
rect 15120 17513 15148 17546
rect 15106 17504 15162 17513
rect 15106 17439 15162 17448
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15028 16697 15056 17138
rect 15014 16688 15070 16697
rect 15764 16674 15792 21383
rect 15856 20466 15884 22034
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15856 19786 15884 20402
rect 15948 19854 15976 24210
rect 16040 21332 16068 25366
rect 16132 25226 16160 25463
rect 16120 25220 16172 25226
rect 16120 25162 16172 25168
rect 16224 24138 16252 26007
rect 16316 25498 16344 26166
rect 16304 25492 16356 25498
rect 16304 25434 16356 25440
rect 16302 25256 16358 25265
rect 16302 25191 16304 25200
rect 16356 25191 16358 25200
rect 16304 25162 16356 25168
rect 16408 24818 16436 27270
rect 16488 26376 16540 26382
rect 16488 26318 16540 26324
rect 16500 26042 16528 26318
rect 16488 26036 16540 26042
rect 16488 25978 16540 25984
rect 16488 25152 16540 25158
rect 16488 25094 16540 25100
rect 16500 24954 16528 25094
rect 16488 24948 16540 24954
rect 16488 24890 16540 24896
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 16500 24698 16528 24890
rect 16408 24670 16528 24698
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 16304 24404 16356 24410
rect 16304 24346 16356 24352
rect 16212 24132 16264 24138
rect 16212 24074 16264 24080
rect 16224 23118 16252 24074
rect 16212 23112 16264 23118
rect 16212 23054 16264 23060
rect 16316 22438 16344 24346
rect 16408 24274 16436 24670
rect 16488 24608 16540 24614
rect 16488 24550 16540 24556
rect 16500 24410 16528 24550
rect 16488 24404 16540 24410
rect 16488 24346 16540 24352
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 16592 24206 16620 24686
rect 16580 24200 16632 24206
rect 16580 24142 16632 24148
rect 16684 24138 16712 28154
rect 16764 24744 16816 24750
rect 16764 24686 16816 24692
rect 16672 24132 16724 24138
rect 16672 24074 16724 24080
rect 16578 24032 16634 24041
rect 16578 23967 16634 23976
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 16040 21304 16160 21332
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 16040 20058 16068 20538
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15844 19780 15896 19786
rect 15844 19722 15896 19728
rect 15948 19378 15976 19790
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 15936 19236 15988 19242
rect 15936 19178 15988 19184
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 15014 16623 15070 16632
rect 15292 16652 15344 16658
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14384 12442 14412 12922
rect 14568 12850 14596 12922
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14372 12436 14424 12442
rect 14660 12434 14688 13262
rect 14752 12850 14780 15302
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14844 14278 14872 14826
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14936 13938 14964 14962
rect 15028 14482 15056 16623
rect 15292 16594 15344 16600
rect 15488 16646 15792 16674
rect 15856 16658 15884 17070
rect 15844 16652 15896 16658
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15120 16046 15148 16390
rect 15198 16280 15254 16289
rect 15198 16215 15254 16224
rect 15212 16182 15240 16215
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 15120 15162 15148 15506
rect 15108 15156 15160 15162
rect 15108 15098 15160 15104
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15212 15042 15240 15098
rect 15120 15014 15240 15042
rect 15120 14890 15148 15014
rect 15108 14884 15160 14890
rect 15108 14826 15160 14832
rect 15198 14648 15254 14657
rect 15198 14583 15254 14592
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14832 12844 14884 12850
rect 14936 12832 14964 13874
rect 15120 13870 15148 14214
rect 15212 14006 15240 14583
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15016 13320 15068 13326
rect 15120 13308 15148 13806
rect 15068 13280 15148 13308
rect 15016 13262 15068 13268
rect 15028 12918 15056 13262
rect 15198 13152 15254 13161
rect 15198 13087 15254 13096
rect 15016 12912 15068 12918
rect 15016 12854 15068 12860
rect 14884 12804 14964 12832
rect 14832 12786 14884 12792
rect 14752 12753 14780 12786
rect 14738 12744 14794 12753
rect 14794 12702 14964 12730
rect 14738 12679 14794 12688
rect 14660 12406 14780 12434
rect 14372 12378 14424 12384
rect 14752 12306 14780 12406
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14936 12238 14964 12702
rect 15028 12442 15056 12854
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15212 12238 15240 13087
rect 15304 12850 15332 16594
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15396 15026 15424 16186
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15488 13462 15516 16646
rect 15844 16594 15896 16600
rect 15856 16250 15884 16594
rect 15948 16522 15976 19178
rect 16040 18426 16068 19994
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 16132 17762 16160 21304
rect 16316 20262 16344 22170
rect 16486 22128 16542 22137
rect 16486 22063 16488 22072
rect 16540 22063 16542 22072
rect 16488 22034 16540 22040
rect 16500 21962 16528 22034
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16486 20360 16542 20369
rect 16486 20295 16542 20304
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16316 17882 16344 20198
rect 16500 20058 16528 20295
rect 16488 20052 16540 20058
rect 16488 19994 16540 20000
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16396 19780 16448 19786
rect 16396 19722 16448 19728
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 16132 17734 16344 17762
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 16132 16590 16160 17614
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 15936 16516 15988 16522
rect 15936 16458 15988 16464
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15948 16114 15976 16458
rect 16040 16425 16068 16458
rect 16026 16416 16082 16425
rect 16026 16351 16082 16360
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15752 15972 15804 15978
rect 15752 15914 15804 15920
rect 15764 14822 15792 15914
rect 15856 15366 15884 16050
rect 15948 15638 15976 16050
rect 15936 15632 15988 15638
rect 15936 15574 15988 15580
rect 16040 15570 16068 16351
rect 16132 15978 16160 16526
rect 16210 16008 16266 16017
rect 16120 15972 16172 15978
rect 16210 15943 16212 15952
rect 16120 15914 16172 15920
rect 16264 15943 16266 15952
rect 16212 15914 16264 15920
rect 16120 15632 16172 15638
rect 16120 15574 16172 15580
rect 16028 15564 16080 15570
rect 16028 15506 16080 15512
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 15844 15360 15896 15366
rect 15844 15302 15896 15308
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15764 14482 15792 14758
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15672 13938 15700 14214
rect 15856 14074 15884 14962
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15948 13938 15976 15438
rect 16132 14414 16160 15574
rect 16212 15428 16264 15434
rect 16212 15370 16264 15376
rect 16224 14793 16252 15370
rect 16316 15366 16344 17734
rect 16408 16561 16436 19722
rect 16394 16552 16450 16561
rect 16394 16487 16450 16496
rect 16500 16402 16528 19790
rect 16592 19174 16620 23967
rect 16684 19446 16712 24074
rect 16672 19440 16724 19446
rect 16672 19382 16724 19388
rect 16580 19168 16632 19174
rect 16580 19110 16632 19116
rect 16592 18748 16620 19110
rect 16592 18720 16712 18748
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16592 17678 16620 18566
rect 16684 18222 16712 18720
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16500 16374 16620 16402
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16408 15502 16436 16050
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 16210 14784 16266 14793
rect 16210 14719 16266 14728
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16040 13938 16068 14350
rect 16224 13938 16252 14719
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 15672 13326 15700 13874
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 16040 13258 16068 13874
rect 16028 13252 16080 13258
rect 16028 13194 16080 13200
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15764 11898 15792 12786
rect 16040 12782 16068 13194
rect 16408 13161 16436 15438
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16394 13152 16450 13161
rect 16394 13087 16450 13096
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 16500 12617 16528 15302
rect 16592 14618 16620 16374
rect 16776 16250 16804 24686
rect 16868 24274 16896 30058
rect 17052 29578 17080 31894
rect 17130 31512 17186 31521
rect 17130 31447 17186 31456
rect 17040 29572 17092 29578
rect 17040 29514 17092 29520
rect 17052 29238 17080 29514
rect 17144 29322 17172 31447
rect 17236 30054 17264 31962
rect 17500 31680 17552 31686
rect 17500 31622 17552 31628
rect 17408 30252 17460 30258
rect 17408 30194 17460 30200
rect 17316 30184 17368 30190
rect 17316 30126 17368 30132
rect 17224 30048 17276 30054
rect 17224 29990 17276 29996
rect 17144 29294 17264 29322
rect 17040 29232 17092 29238
rect 17040 29174 17092 29180
rect 17132 29232 17184 29238
rect 17132 29174 17184 29180
rect 16948 29164 17000 29170
rect 16948 29106 17000 29112
rect 16960 27402 16988 29106
rect 16948 27396 17000 27402
rect 16948 27338 17000 27344
rect 16960 26518 16988 27338
rect 17040 26580 17092 26586
rect 17040 26522 17092 26528
rect 16948 26512 17000 26518
rect 16948 26454 17000 26460
rect 16948 24404 17000 24410
rect 16948 24346 17000 24352
rect 16856 24268 16908 24274
rect 16856 24210 16908 24216
rect 16868 22273 16896 24210
rect 16960 24070 16988 24346
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 16960 23866 16988 24006
rect 16948 23860 17000 23866
rect 16948 23802 17000 23808
rect 16948 22500 17000 22506
rect 16948 22442 17000 22448
rect 16854 22264 16910 22273
rect 16854 22199 16910 22208
rect 16868 22030 16896 22199
rect 16960 22166 16988 22442
rect 16948 22160 17000 22166
rect 16948 22102 17000 22108
rect 16856 22024 16908 22030
rect 16856 21966 16908 21972
rect 16948 21956 17000 21962
rect 16948 21898 17000 21904
rect 16960 21729 16988 21898
rect 16946 21720 17002 21729
rect 16946 21655 17002 21664
rect 16854 20632 16910 20641
rect 16854 20567 16910 20576
rect 16868 20330 16896 20567
rect 16856 20324 16908 20330
rect 16856 20266 16908 20272
rect 17052 19334 17080 26522
rect 17144 22234 17172 29174
rect 17236 28200 17264 29294
rect 17328 29073 17356 30126
rect 17420 29889 17448 30194
rect 17406 29880 17462 29889
rect 17406 29815 17462 29824
rect 17408 29572 17460 29578
rect 17408 29514 17460 29520
rect 17420 29238 17448 29514
rect 17408 29232 17460 29238
rect 17408 29174 17460 29180
rect 17314 29064 17370 29073
rect 17314 28999 17370 29008
rect 17236 28172 17356 28200
rect 17222 28112 17278 28121
rect 17222 28047 17278 28056
rect 17236 27713 17264 28047
rect 17222 27704 17278 27713
rect 17222 27639 17278 27648
rect 17224 27396 17276 27402
rect 17224 27338 17276 27344
rect 17236 26926 17264 27338
rect 17328 27282 17356 28172
rect 17408 28144 17460 28150
rect 17408 28086 17460 28092
rect 17420 27402 17448 28086
rect 17512 27538 17540 31622
rect 17684 30864 17736 30870
rect 17684 30806 17736 30812
rect 17592 30252 17644 30258
rect 17592 30194 17644 30200
rect 17604 30161 17632 30194
rect 17590 30152 17646 30161
rect 17696 30122 17724 30806
rect 17590 30087 17646 30096
rect 17684 30116 17736 30122
rect 17684 30058 17736 30064
rect 17590 29608 17646 29617
rect 17590 29543 17646 29552
rect 17604 29306 17632 29543
rect 17592 29300 17644 29306
rect 17592 29242 17644 29248
rect 17500 27532 17552 27538
rect 17500 27474 17552 27480
rect 17408 27396 17460 27402
rect 17408 27338 17460 27344
rect 17328 27254 17540 27282
rect 17224 26920 17276 26926
rect 17224 26862 17276 26868
rect 17236 26042 17264 26862
rect 17314 26616 17370 26625
rect 17314 26551 17370 26560
rect 17328 26518 17356 26551
rect 17316 26512 17368 26518
rect 17316 26454 17368 26460
rect 17406 26344 17462 26353
rect 17406 26279 17462 26288
rect 17224 26036 17276 26042
rect 17224 25978 17276 25984
rect 17316 25356 17368 25362
rect 17316 25298 17368 25304
rect 17224 24812 17276 24818
rect 17224 24754 17276 24760
rect 17236 24410 17264 24754
rect 17224 24404 17276 24410
rect 17224 24346 17276 24352
rect 17224 24268 17276 24274
rect 17224 24210 17276 24216
rect 17236 24070 17264 24210
rect 17224 24064 17276 24070
rect 17224 24006 17276 24012
rect 17132 22228 17184 22234
rect 17132 22170 17184 22176
rect 17144 21146 17172 22170
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 17236 20942 17264 21354
rect 17224 20936 17276 20942
rect 17222 20904 17224 20913
rect 17276 20904 17278 20913
rect 17222 20839 17278 20848
rect 17052 19306 17264 19334
rect 16856 19236 16908 19242
rect 16856 19178 16908 19184
rect 16868 18086 16896 19178
rect 17040 18964 17092 18970
rect 17040 18906 17092 18912
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16960 18426 16988 18702
rect 17052 18601 17080 18906
rect 17130 18864 17186 18873
rect 17130 18799 17186 18808
rect 17038 18592 17094 18601
rect 17038 18527 17094 18536
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 17144 18222 17172 18799
rect 17236 18766 17264 19306
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17132 18216 17184 18222
rect 17132 18158 17184 18164
rect 17236 18086 17264 18566
rect 17328 18290 17356 25298
rect 17420 19242 17448 26279
rect 17512 24206 17540 27254
rect 17592 26512 17644 26518
rect 17592 26454 17644 26460
rect 17604 24818 17632 26454
rect 17684 25424 17736 25430
rect 17684 25366 17736 25372
rect 17696 25294 17724 25366
rect 17684 25288 17736 25294
rect 17684 25230 17736 25236
rect 17682 24848 17738 24857
rect 17592 24812 17644 24818
rect 17682 24783 17684 24792
rect 17592 24754 17644 24760
rect 17736 24783 17738 24792
rect 17684 24754 17736 24760
rect 17696 24274 17724 24754
rect 17788 24682 17816 33594
rect 21652 33454 21680 33934
rect 21640 33448 21692 33454
rect 21640 33390 21692 33396
rect 21928 33386 21956 33934
rect 22664 33522 22692 35430
rect 23204 35080 23256 35086
rect 23204 35022 23256 35028
rect 23216 34678 23244 35022
rect 23296 35012 23348 35018
rect 23296 34954 23348 34960
rect 23204 34672 23256 34678
rect 23204 34614 23256 34620
rect 22836 34196 22888 34202
rect 22836 34138 22888 34144
rect 23112 34196 23164 34202
rect 23112 34138 23164 34144
rect 23204 34196 23256 34202
rect 23204 34138 23256 34144
rect 22744 33856 22796 33862
rect 22744 33798 22796 33804
rect 22652 33516 22704 33522
rect 22652 33458 22704 33464
rect 22756 33386 22784 33798
rect 21916 33380 21968 33386
rect 21916 33322 21968 33328
rect 22744 33380 22796 33386
rect 22744 33322 22796 33328
rect 21824 33040 21876 33046
rect 21824 32982 21876 32988
rect 20720 32972 20772 32978
rect 20720 32914 20772 32920
rect 18420 32904 18472 32910
rect 18420 32846 18472 32852
rect 17868 31816 17920 31822
rect 17868 31758 17920 31764
rect 17880 30054 17908 31758
rect 18432 31754 18460 32846
rect 19340 32564 19392 32570
rect 19340 32506 19392 32512
rect 19064 32428 19116 32434
rect 19064 32370 19116 32376
rect 18972 31816 19024 31822
rect 18972 31758 19024 31764
rect 18340 31726 18460 31754
rect 18236 30592 18288 30598
rect 18236 30534 18288 30540
rect 18248 30258 18276 30534
rect 18052 30252 18104 30258
rect 18052 30194 18104 30200
rect 18236 30252 18288 30258
rect 18236 30194 18288 30200
rect 18064 30161 18092 30194
rect 18050 30152 18106 30161
rect 18050 30087 18106 30096
rect 17868 30048 17920 30054
rect 17868 29990 17920 29996
rect 18144 30048 18196 30054
rect 18144 29990 18196 29996
rect 17880 27713 17908 29990
rect 18156 29646 18184 29990
rect 18144 29640 18196 29646
rect 18144 29582 18196 29588
rect 18052 29232 18104 29238
rect 18052 29174 18104 29180
rect 17960 28960 18012 28966
rect 17960 28902 18012 28908
rect 17972 27878 18000 28902
rect 18064 28490 18092 29174
rect 18144 29164 18196 29170
rect 18144 29106 18196 29112
rect 18052 28484 18104 28490
rect 18052 28426 18104 28432
rect 17960 27872 18012 27878
rect 17960 27814 18012 27820
rect 17866 27704 17922 27713
rect 17866 27639 17922 27648
rect 17880 27169 17908 27639
rect 17866 27160 17922 27169
rect 18064 27130 18092 28426
rect 17866 27095 17922 27104
rect 18052 27124 18104 27130
rect 18052 27066 18104 27072
rect 17960 26580 18012 26586
rect 18064 26568 18092 27066
rect 18156 26586 18184 29106
rect 18236 28484 18288 28490
rect 18236 28426 18288 28432
rect 18012 26540 18092 26568
rect 18144 26580 18196 26586
rect 17960 26522 18012 26528
rect 18144 26522 18196 26528
rect 17972 24750 18000 26522
rect 17960 24744 18012 24750
rect 17960 24686 18012 24692
rect 17776 24676 17828 24682
rect 17776 24618 17828 24624
rect 17868 24608 17920 24614
rect 17920 24568 18000 24596
rect 17868 24550 17920 24556
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 17776 24132 17828 24138
rect 17776 24074 17828 24080
rect 17590 21992 17646 22001
rect 17590 21927 17646 21936
rect 17500 21480 17552 21486
rect 17500 21422 17552 21428
rect 17512 20398 17540 21422
rect 17604 20942 17632 21927
rect 17684 21548 17736 21554
rect 17788 21536 17816 24074
rect 17736 21508 17816 21536
rect 17684 21490 17736 21496
rect 17696 20942 17724 21490
rect 17592 20936 17644 20942
rect 17590 20904 17592 20913
rect 17684 20936 17736 20942
rect 17644 20904 17646 20913
rect 17684 20878 17736 20884
rect 17590 20839 17646 20848
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17408 19236 17460 19242
rect 17408 19178 17460 19184
rect 17498 18864 17554 18873
rect 17498 18799 17554 18808
rect 17512 18630 17540 18799
rect 17788 18630 17816 20198
rect 17880 19718 17908 24142
rect 17972 22953 18000 24568
rect 18050 24576 18106 24585
rect 18156 24562 18184 26522
rect 18248 24818 18276 28426
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 18234 24712 18290 24721
rect 18234 24647 18236 24656
rect 18288 24647 18290 24656
rect 18236 24618 18288 24624
rect 18156 24534 18276 24562
rect 18050 24511 18106 24520
rect 18064 24392 18092 24511
rect 18248 24410 18276 24534
rect 18236 24404 18288 24410
rect 18064 24364 18184 24392
rect 18052 24268 18104 24274
rect 18052 24210 18104 24216
rect 17958 22944 18014 22953
rect 17958 22879 18014 22888
rect 18064 22098 18092 24210
rect 18156 22964 18184 24364
rect 18236 24346 18288 24352
rect 18340 24274 18368 31726
rect 18512 30796 18564 30802
rect 18512 30738 18564 30744
rect 18524 30394 18552 30738
rect 18786 30560 18842 30569
rect 18786 30495 18842 30504
rect 18800 30394 18828 30495
rect 18512 30388 18564 30394
rect 18512 30330 18564 30336
rect 18788 30388 18840 30394
rect 18788 30330 18840 30336
rect 18984 30326 19012 31758
rect 18696 30320 18748 30326
rect 18696 30262 18748 30268
rect 18972 30320 19024 30326
rect 18972 30262 19024 30268
rect 18708 30161 18736 30262
rect 18788 30252 18840 30258
rect 18788 30194 18840 30200
rect 18694 30152 18750 30161
rect 18604 30116 18656 30122
rect 18694 30087 18750 30096
rect 18604 30058 18656 30064
rect 18616 29578 18644 30058
rect 18800 30054 18828 30194
rect 18880 30184 18932 30190
rect 18880 30126 18932 30132
rect 18788 30048 18840 30054
rect 18788 29990 18840 29996
rect 18892 29889 18920 30126
rect 18878 29880 18934 29889
rect 18788 29844 18840 29850
rect 18878 29815 18934 29824
rect 18788 29786 18840 29792
rect 18694 29744 18750 29753
rect 18694 29679 18750 29688
rect 18708 29646 18736 29679
rect 18696 29640 18748 29646
rect 18696 29582 18748 29588
rect 18604 29572 18656 29578
rect 18604 29514 18656 29520
rect 18800 28994 18828 29786
rect 18984 29073 19012 30262
rect 19076 29850 19104 32370
rect 19352 31822 19380 32506
rect 19432 32428 19484 32434
rect 19432 32370 19484 32376
rect 19444 31929 19472 32370
rect 20732 32366 20760 32914
rect 21836 32434 21864 32982
rect 21916 32904 21968 32910
rect 21916 32846 21968 32852
rect 21824 32428 21876 32434
rect 21824 32370 21876 32376
rect 20720 32360 20772 32366
rect 20720 32302 20772 32308
rect 19524 32292 19576 32298
rect 19524 32234 19576 32240
rect 19430 31920 19486 31929
rect 19430 31855 19486 31864
rect 19340 31816 19392 31822
rect 19340 31758 19392 31764
rect 19246 30968 19302 30977
rect 19536 30938 19564 32234
rect 19982 31920 20038 31929
rect 19982 31855 20038 31864
rect 19996 31822 20024 31855
rect 19984 31816 20036 31822
rect 19984 31758 20036 31764
rect 19616 31680 19668 31686
rect 19614 31648 19616 31657
rect 19668 31648 19670 31657
rect 19614 31583 19670 31592
rect 20732 31414 20760 32302
rect 20812 31884 20864 31890
rect 20812 31826 20864 31832
rect 20720 31408 20772 31414
rect 20720 31350 20772 31356
rect 20076 31340 20128 31346
rect 20076 31282 20128 31288
rect 19892 31272 19944 31278
rect 19892 31214 19944 31220
rect 19616 31136 19668 31142
rect 19616 31078 19668 31084
rect 19246 30903 19302 30912
rect 19524 30932 19576 30938
rect 19156 30592 19208 30598
rect 19156 30534 19208 30540
rect 19168 30054 19196 30534
rect 19156 30048 19208 30054
rect 19156 29990 19208 29996
rect 19064 29844 19116 29850
rect 19064 29786 19116 29792
rect 19156 29844 19208 29850
rect 19156 29786 19208 29792
rect 19062 29744 19118 29753
rect 19168 29730 19196 29786
rect 19118 29702 19196 29730
rect 19260 29730 19288 30903
rect 19524 30874 19576 30880
rect 19432 30252 19484 30258
rect 19432 30194 19484 30200
rect 19524 30252 19576 30258
rect 19524 30194 19576 30200
rect 19260 29702 19334 29730
rect 19444 29714 19472 30194
rect 19536 30054 19564 30194
rect 19628 30054 19656 31078
rect 19800 30660 19852 30666
rect 19800 30602 19852 30608
rect 19524 30048 19576 30054
rect 19524 29990 19576 29996
rect 19616 30048 19668 30054
rect 19616 29990 19668 29996
rect 19062 29679 19118 29688
rect 18970 29064 19026 29073
rect 18970 28999 19026 29008
rect 18708 28966 18828 28994
rect 18420 28484 18472 28490
rect 18420 28426 18472 28432
rect 18432 26353 18460 28426
rect 18512 28416 18564 28422
rect 18512 28358 18564 28364
rect 18604 28416 18656 28422
rect 18604 28358 18656 28364
rect 18524 28082 18552 28358
rect 18512 28076 18564 28082
rect 18512 28018 18564 28024
rect 18616 26858 18644 28358
rect 18604 26852 18656 26858
rect 18604 26794 18656 26800
rect 18512 26784 18564 26790
rect 18512 26726 18564 26732
rect 18524 26382 18552 26726
rect 18512 26376 18564 26382
rect 18418 26344 18474 26353
rect 18512 26318 18564 26324
rect 18708 26330 18736 28966
rect 18788 28416 18840 28422
rect 19076 28393 19104 29679
rect 19306 29578 19334 29702
rect 19432 29708 19484 29714
rect 19432 29650 19484 29656
rect 19294 29572 19346 29578
rect 19294 29514 19346 29520
rect 19156 29504 19208 29510
rect 19156 29446 19208 29452
rect 18788 28358 18840 28364
rect 19062 28384 19118 28393
rect 18800 28218 18828 28358
rect 19062 28319 19118 28328
rect 18788 28212 18840 28218
rect 18788 28154 18840 28160
rect 18972 28212 19024 28218
rect 18972 28154 19024 28160
rect 18880 28076 18932 28082
rect 18880 28018 18932 28024
rect 18892 27674 18920 28018
rect 18984 27878 19012 28154
rect 19076 27962 19104 28319
rect 19168 28082 19196 29446
rect 19444 29306 19472 29650
rect 19432 29300 19484 29306
rect 19352 29260 19432 29288
rect 19248 29164 19300 29170
rect 19248 29106 19300 29112
rect 19260 29073 19288 29106
rect 19246 29064 19302 29073
rect 19352 29034 19380 29260
rect 19432 29242 19484 29248
rect 19432 29164 19484 29170
rect 19432 29106 19484 29112
rect 19246 28999 19302 29008
rect 19340 29028 19392 29034
rect 19340 28970 19392 28976
rect 19156 28076 19208 28082
rect 19156 28018 19208 28024
rect 19248 28076 19300 28082
rect 19248 28018 19300 28024
rect 19260 27962 19288 28018
rect 19076 27934 19288 27962
rect 18972 27872 19024 27878
rect 18972 27814 19024 27820
rect 19064 27872 19116 27878
rect 19064 27814 19116 27820
rect 18880 27668 18932 27674
rect 18880 27610 18932 27616
rect 18786 27296 18842 27305
rect 18786 27231 18842 27240
rect 18800 26450 18828 27231
rect 19076 26790 19104 27814
rect 19064 26784 19116 26790
rect 19064 26726 19116 26732
rect 19062 26616 19118 26625
rect 18880 26580 18932 26586
rect 19062 26551 19118 26560
rect 18880 26522 18932 26528
rect 18788 26444 18840 26450
rect 18788 26386 18840 26392
rect 18708 26302 18828 26330
rect 18418 26279 18474 26288
rect 18420 26240 18472 26246
rect 18420 26182 18472 26188
rect 18512 26240 18564 26246
rect 18512 26182 18564 26188
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 18156 22936 18368 22964
rect 18052 22092 18104 22098
rect 18340 22094 18368 22936
rect 18052 22034 18104 22040
rect 18156 22066 18368 22094
rect 18156 21978 18184 22066
rect 18064 21950 18184 21978
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 18064 19854 18092 21950
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 18156 21622 18184 21830
rect 18144 21616 18196 21622
rect 18144 21558 18196 21564
rect 18144 21140 18196 21146
rect 18144 21082 18196 21088
rect 18156 20777 18184 21082
rect 18142 20768 18198 20777
rect 18142 20703 18198 20712
rect 18248 20534 18276 21966
rect 18340 21962 18368 22066
rect 18328 21956 18380 21962
rect 18328 21898 18380 21904
rect 18326 21584 18382 21593
rect 18326 21519 18382 21528
rect 18340 20942 18368 21519
rect 18432 21010 18460 26182
rect 18524 26042 18552 26182
rect 18512 26036 18564 26042
rect 18512 25978 18564 25984
rect 18512 24812 18564 24818
rect 18512 24754 18564 24760
rect 18524 24585 18552 24754
rect 18604 24744 18656 24750
rect 18604 24686 18656 24692
rect 18510 24576 18566 24585
rect 18510 24511 18566 24520
rect 18512 24132 18564 24138
rect 18512 24074 18564 24080
rect 18524 23118 18552 24074
rect 18616 23662 18644 24686
rect 18696 24676 18748 24682
rect 18696 24618 18748 24624
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18602 23488 18658 23497
rect 18602 23423 18658 23432
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 18524 22642 18552 23054
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18512 21956 18564 21962
rect 18512 21898 18564 21904
rect 18420 21004 18472 21010
rect 18420 20946 18472 20952
rect 18328 20936 18380 20942
rect 18328 20878 18380 20884
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 18236 20528 18288 20534
rect 18236 20470 18288 20476
rect 18234 20360 18290 20369
rect 18234 20295 18290 20304
rect 18248 19854 18276 20295
rect 18052 19848 18104 19854
rect 18052 19790 18104 19796
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 17868 19712 17920 19718
rect 18248 19689 18276 19790
rect 17868 19654 17920 19660
rect 18234 19680 18290 19689
rect 18234 19615 18290 19624
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 18156 18426 18184 19178
rect 18144 18420 18196 18426
rect 18144 18362 18196 18368
rect 17868 18352 17920 18358
rect 17498 18320 17554 18329
rect 17316 18284 17368 18290
rect 17868 18294 17920 18300
rect 17498 18255 17554 18264
rect 17592 18284 17644 18290
rect 17316 18226 17368 18232
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 17040 17740 17092 17746
rect 17040 17682 17092 17688
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16868 17270 16896 17614
rect 16856 17264 16908 17270
rect 16856 17206 16908 17212
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16684 14890 16712 16050
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 16776 15201 16804 15438
rect 16762 15192 16818 15201
rect 16762 15127 16818 15136
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16670 14648 16726 14657
rect 16580 14612 16632 14618
rect 16670 14583 16726 14592
rect 16580 14554 16632 14560
rect 16684 14550 16712 14583
rect 16672 14544 16724 14550
rect 16672 14486 16724 14492
rect 16776 14414 16804 14894
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16868 14346 16896 17206
rect 17052 16726 17080 17682
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 17040 16720 17092 16726
rect 17040 16662 17092 16668
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 16868 14074 16896 14282
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16960 13802 16988 15982
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17052 14278 17080 15846
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 17144 14074 17172 17478
rect 17406 16824 17462 16833
rect 17406 16759 17462 16768
rect 17420 16726 17448 16759
rect 17408 16720 17460 16726
rect 17408 16662 17460 16668
rect 17224 16516 17276 16522
rect 17224 16458 17276 16464
rect 17236 15910 17264 16458
rect 17314 16144 17370 16153
rect 17314 16079 17316 16088
rect 17368 16079 17370 16088
rect 17316 16050 17368 16056
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17512 15366 17540 18255
rect 17592 18226 17644 18232
rect 17684 18284 17736 18290
rect 17684 18226 17736 18232
rect 17604 18086 17632 18226
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17592 16516 17644 16522
rect 17592 16458 17644 16464
rect 17604 16182 17632 16458
rect 17592 16176 17644 16182
rect 17592 16118 17644 16124
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17696 14906 17724 18226
rect 17776 18216 17828 18222
rect 17776 18158 17828 18164
rect 17788 17814 17816 18158
rect 17776 17808 17828 17814
rect 17776 17750 17828 17756
rect 17880 17542 17908 18294
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18050 18048 18106 18057
rect 18050 17983 18106 17992
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17788 17202 17816 17478
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17880 16726 17908 17478
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17868 16720 17920 16726
rect 17868 16662 17920 16668
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 17788 15638 17816 16186
rect 17972 15638 18000 17070
rect 17776 15632 17828 15638
rect 17776 15574 17828 15580
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 17972 15502 18000 15574
rect 18064 15502 18092 17983
rect 18142 15736 18198 15745
rect 18142 15671 18198 15680
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 18064 15201 18092 15438
rect 18156 15434 18184 15671
rect 18144 15428 18196 15434
rect 18144 15370 18196 15376
rect 18050 15192 18106 15201
rect 18050 15127 18106 15136
rect 17696 14878 17816 14906
rect 17406 14104 17462 14113
rect 17132 14068 17184 14074
rect 17406 14039 17462 14048
rect 17132 14010 17184 14016
rect 16948 13796 17000 13802
rect 16948 13738 17000 13744
rect 17144 13512 17172 14010
rect 17420 13938 17448 14039
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17420 13530 17448 13670
rect 17408 13524 17460 13530
rect 16960 13484 17356 13512
rect 16960 13326 16988 13484
rect 17328 13410 17356 13484
rect 17408 13466 17460 13472
rect 17328 13382 17448 13410
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 17222 13288 17278 13297
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 17132 13252 17184 13258
rect 17222 13223 17278 13232
rect 17132 13194 17184 13200
rect 16486 12608 16542 12617
rect 16486 12543 16542 12552
rect 17052 12434 17080 13194
rect 17144 12850 17172 13194
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17236 12714 17264 13223
rect 17420 12918 17448 13382
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17316 12912 17368 12918
rect 17316 12854 17368 12860
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 17224 12708 17276 12714
rect 17224 12650 17276 12656
rect 17328 12434 17356 12854
rect 17512 12850 17540 13262
rect 17604 12986 17632 13874
rect 17696 13433 17724 13874
rect 17788 13462 17816 14878
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17776 13456 17828 13462
rect 17682 13424 17738 13433
rect 17776 13398 17828 13404
rect 17682 13359 17738 13368
rect 17880 13002 17908 13806
rect 17972 13326 18000 13874
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 18248 13025 18276 18226
rect 18340 18034 18368 20742
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 18432 19514 18460 20402
rect 18524 20369 18552 21898
rect 18510 20360 18566 20369
rect 18510 20295 18566 20304
rect 18512 20256 18564 20262
rect 18512 20198 18564 20204
rect 18524 19990 18552 20198
rect 18512 19984 18564 19990
rect 18512 19926 18564 19932
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 18524 19553 18552 19790
rect 18510 19544 18566 19553
rect 18420 19508 18472 19514
rect 18510 19479 18566 19488
rect 18420 19450 18472 19456
rect 18616 19258 18644 23423
rect 18708 20874 18736 24618
rect 18800 24410 18828 26302
rect 18892 25838 18920 26522
rect 19076 26314 19104 26551
rect 19064 26308 19116 26314
rect 19064 26250 19116 26256
rect 18880 25832 18932 25838
rect 18880 25774 18932 25780
rect 18788 24404 18840 24410
rect 18788 24346 18840 24352
rect 19064 24336 19116 24342
rect 19064 24278 19116 24284
rect 18880 24132 18932 24138
rect 18880 24074 18932 24080
rect 18892 23322 18920 24074
rect 18880 23316 18932 23322
rect 18880 23258 18932 23264
rect 18892 23225 18920 23258
rect 18878 23216 18934 23225
rect 18878 23151 18934 23160
rect 18878 22808 18934 22817
rect 18878 22743 18934 22752
rect 18892 22094 18920 22743
rect 18892 22066 19012 22094
rect 18880 21956 18932 21962
rect 18880 21898 18932 21904
rect 18696 20868 18748 20874
rect 18696 20810 18748 20816
rect 18696 20392 18748 20398
rect 18696 20334 18748 20340
rect 18432 19230 18644 19258
rect 18708 19258 18736 20334
rect 18786 20088 18842 20097
rect 18786 20023 18842 20032
rect 18800 19378 18828 20023
rect 18892 19938 18920 21898
rect 18984 20398 19012 22066
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18970 20088 19026 20097
rect 18970 20023 18972 20032
rect 19024 20023 19026 20032
rect 18972 19994 19024 20000
rect 18892 19910 19012 19938
rect 18878 19408 18934 19417
rect 18788 19372 18840 19378
rect 18878 19343 18880 19352
rect 18788 19314 18840 19320
rect 18932 19343 18934 19352
rect 18880 19314 18932 19320
rect 18708 19230 18920 19258
rect 18432 18170 18460 19230
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18524 18358 18552 19110
rect 18512 18352 18564 18358
rect 18512 18294 18564 18300
rect 18616 18193 18644 19110
rect 18602 18184 18658 18193
rect 18432 18142 18552 18170
rect 18340 18006 18460 18034
rect 18326 16552 18382 16561
rect 18326 16487 18382 16496
rect 18340 15978 18368 16487
rect 18328 15972 18380 15978
rect 18328 15914 18380 15920
rect 18432 15881 18460 18006
rect 18418 15872 18474 15881
rect 18418 15807 18474 15816
rect 18432 15162 18460 15807
rect 18524 15609 18552 18142
rect 18602 18119 18658 18128
rect 18892 17241 18920 19230
rect 18878 17232 18934 17241
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18788 17196 18840 17202
rect 18878 17167 18934 17176
rect 18788 17138 18840 17144
rect 18708 16425 18736 17138
rect 18800 16998 18828 17138
rect 18788 16992 18840 16998
rect 18892 16969 18920 17167
rect 18788 16934 18840 16940
rect 18878 16960 18934 16969
rect 18878 16895 18934 16904
rect 18694 16416 18750 16425
rect 18694 16351 18750 16360
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18510 15600 18566 15609
rect 18510 15535 18566 15544
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18524 15094 18552 15438
rect 18512 15088 18564 15094
rect 18512 15030 18564 15036
rect 18616 14550 18644 15982
rect 18708 15502 18736 16351
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18696 15496 18748 15502
rect 18800 15473 18828 15846
rect 18892 15609 18920 16050
rect 18878 15600 18934 15609
rect 18878 15535 18934 15544
rect 18880 15496 18932 15502
rect 18696 15438 18748 15444
rect 18786 15464 18842 15473
rect 18708 15162 18736 15438
rect 18880 15438 18932 15444
rect 18786 15399 18842 15408
rect 18892 15201 18920 15438
rect 18878 15192 18934 15201
rect 18696 15156 18748 15162
rect 18878 15127 18934 15136
rect 18696 15098 18748 15104
rect 18604 14544 18656 14550
rect 18604 14486 18656 14492
rect 18616 13870 18644 14486
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18510 13424 18566 13433
rect 18510 13359 18566 13368
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18234 13016 18290 13025
rect 17592 12980 17644 12986
rect 17880 12974 18000 13002
rect 17592 12922 17644 12928
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 16960 12406 17356 12434
rect 16960 12170 16988 12406
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 17052 12102 17080 12310
rect 17328 12238 17356 12406
rect 17512 12238 17540 12786
rect 17972 12782 18000 12974
rect 18234 12951 18290 12960
rect 17960 12776 18012 12782
rect 17682 12744 17738 12753
rect 17960 12718 18012 12724
rect 17682 12679 17684 12688
rect 17736 12679 17738 12688
rect 17684 12650 17736 12656
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17500 12232 17552 12238
rect 17604 12220 17632 12378
rect 18248 12374 18276 12951
rect 18340 12918 18368 13126
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18524 12850 18552 13359
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18708 12714 18736 13874
rect 18788 13864 18840 13870
rect 18984 13818 19012 19910
rect 19076 17134 19104 24278
rect 19168 22030 19196 27934
rect 19338 27704 19394 27713
rect 19338 27639 19340 27648
rect 19392 27639 19394 27648
rect 19340 27610 19392 27616
rect 19444 26926 19472 29106
rect 19628 27674 19656 29990
rect 19812 29578 19840 30602
rect 19904 30258 19932 31214
rect 19984 31136 20036 31142
rect 19984 31078 20036 31084
rect 19996 30841 20024 31078
rect 19982 30832 20038 30841
rect 19982 30767 20038 30776
rect 19892 30252 19944 30258
rect 19892 30194 19944 30200
rect 19800 29572 19852 29578
rect 19800 29514 19852 29520
rect 19708 29504 19760 29510
rect 19708 29446 19760 29452
rect 19720 29345 19748 29446
rect 19706 29336 19762 29345
rect 19706 29271 19762 29280
rect 19812 28801 19840 29514
rect 19798 28792 19854 28801
rect 19798 28727 19854 28736
rect 19800 28144 19852 28150
rect 19800 28086 19852 28092
rect 19708 27872 19760 27878
rect 19708 27814 19760 27820
rect 19616 27668 19668 27674
rect 19616 27610 19668 27616
rect 19720 27606 19748 27814
rect 19708 27600 19760 27606
rect 19708 27542 19760 27548
rect 19812 27470 19840 28086
rect 19616 27464 19668 27470
rect 19616 27406 19668 27412
rect 19800 27464 19852 27470
rect 19800 27406 19852 27412
rect 19524 26988 19576 26994
rect 19524 26930 19576 26936
rect 19432 26920 19484 26926
rect 19432 26862 19484 26868
rect 19340 26580 19392 26586
rect 19340 26522 19392 26528
rect 19352 25974 19380 26522
rect 19340 25968 19392 25974
rect 19340 25910 19392 25916
rect 19536 25770 19564 26930
rect 19628 26450 19656 27406
rect 19706 27160 19762 27169
rect 19706 27095 19708 27104
rect 19760 27095 19762 27104
rect 19708 27066 19760 27072
rect 19616 26444 19668 26450
rect 19616 26386 19668 26392
rect 19708 26308 19760 26314
rect 19708 26250 19760 26256
rect 19524 25764 19576 25770
rect 19524 25706 19576 25712
rect 19522 25528 19578 25537
rect 19720 25498 19748 26250
rect 19522 25463 19524 25472
rect 19576 25463 19578 25472
rect 19708 25492 19760 25498
rect 19524 25434 19576 25440
rect 19708 25434 19760 25440
rect 19800 25492 19852 25498
rect 19800 25434 19852 25440
rect 19616 25424 19668 25430
rect 19338 25392 19394 25401
rect 19616 25366 19668 25372
rect 19338 25327 19394 25336
rect 19432 25356 19484 25362
rect 19352 25129 19380 25327
rect 19432 25298 19484 25304
rect 19338 25120 19394 25129
rect 19338 25055 19394 25064
rect 19340 24880 19392 24886
rect 19444 24868 19472 25298
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19392 24840 19472 24868
rect 19340 24822 19392 24828
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19352 23089 19380 23122
rect 19338 23080 19394 23089
rect 19338 23015 19394 23024
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19260 22030 19288 22918
rect 19340 22704 19392 22710
rect 19340 22646 19392 22652
rect 19352 22545 19380 22646
rect 19338 22536 19394 22545
rect 19338 22471 19394 22480
rect 19444 22420 19472 24006
rect 19536 23497 19564 25230
rect 19628 25158 19656 25366
rect 19812 25362 19840 25434
rect 19800 25356 19852 25362
rect 19800 25298 19852 25304
rect 19904 25242 19932 30194
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 19996 29306 20024 29582
rect 19984 29300 20036 29306
rect 19984 29242 20036 29248
rect 19996 27962 20024 29242
rect 20088 28422 20116 31282
rect 20720 31136 20772 31142
rect 20720 31078 20772 31084
rect 20444 30592 20496 30598
rect 20442 30560 20444 30569
rect 20496 30560 20498 30569
rect 20442 30495 20498 30504
rect 20536 29708 20588 29714
rect 20536 29650 20588 29656
rect 20168 29504 20220 29510
rect 20168 29446 20220 29452
rect 20180 28966 20208 29446
rect 20168 28960 20220 28966
rect 20168 28902 20220 28908
rect 20180 28422 20208 28902
rect 20260 28484 20312 28490
rect 20260 28426 20312 28432
rect 20076 28416 20128 28422
rect 20076 28358 20128 28364
rect 20168 28416 20220 28422
rect 20168 28358 20220 28364
rect 20088 28150 20116 28358
rect 20076 28144 20128 28150
rect 20076 28086 20128 28092
rect 19996 27934 20116 27962
rect 19982 27432 20038 27441
rect 19982 27367 19984 27376
rect 20036 27367 20038 27376
rect 19984 27338 20036 27344
rect 19984 25424 20036 25430
rect 19984 25366 20036 25372
rect 19720 25214 19932 25242
rect 19616 25152 19668 25158
rect 19616 25094 19668 25100
rect 19614 24984 19670 24993
rect 19614 24919 19670 24928
rect 19628 24818 19656 24919
rect 19720 24818 19748 25214
rect 19890 25120 19946 25129
rect 19890 25055 19946 25064
rect 19616 24812 19668 24818
rect 19616 24754 19668 24760
rect 19708 24812 19760 24818
rect 19708 24754 19760 24760
rect 19708 24608 19760 24614
rect 19708 24550 19760 24556
rect 19720 24070 19748 24550
rect 19800 24404 19852 24410
rect 19800 24346 19852 24352
rect 19812 24274 19840 24346
rect 19800 24268 19852 24274
rect 19800 24210 19852 24216
rect 19708 24064 19760 24070
rect 19708 24006 19760 24012
rect 19522 23488 19578 23497
rect 19522 23423 19578 23432
rect 19706 23488 19762 23497
rect 19706 23423 19762 23432
rect 19352 22392 19472 22420
rect 19156 22024 19208 22030
rect 19156 21966 19208 21972
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 19248 21140 19300 21146
rect 19248 21082 19300 21088
rect 19156 19712 19208 19718
rect 19156 19654 19208 19660
rect 19168 19156 19196 19654
rect 19260 19514 19288 21082
rect 19352 20534 19380 22392
rect 19616 22160 19668 22166
rect 19616 22102 19668 22108
rect 19524 22024 19576 22030
rect 19524 21966 19576 21972
rect 19536 21350 19564 21966
rect 19628 21350 19656 22102
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19616 21344 19668 21350
rect 19616 21286 19668 21292
rect 19720 21146 19748 23423
rect 19798 22808 19854 22817
rect 19798 22743 19854 22752
rect 19812 22642 19840 22743
rect 19800 22636 19852 22642
rect 19800 22578 19852 22584
rect 19708 21140 19760 21146
rect 19708 21082 19760 21088
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19248 19168 19300 19174
rect 19168 19128 19248 19156
rect 19248 19110 19300 19116
rect 19260 18902 19288 19110
rect 19248 18896 19300 18902
rect 19248 18838 19300 18844
rect 19156 18760 19208 18766
rect 19208 18720 19288 18748
rect 19156 18702 19208 18708
rect 19260 18290 19288 18720
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19154 17232 19210 17241
rect 19154 17167 19156 17176
rect 19208 17167 19210 17176
rect 19156 17138 19208 17144
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 19076 15638 19104 15846
rect 19064 15632 19116 15638
rect 19064 15574 19116 15580
rect 19168 13938 19196 16934
rect 19260 15745 19288 18226
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 19352 17610 19380 18022
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19338 17096 19394 17105
rect 19338 17031 19394 17040
rect 19352 16998 19380 17031
rect 19444 16998 19472 20878
rect 19904 20806 19932 25055
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19892 20800 19944 20806
rect 19892 20742 19944 20748
rect 19536 20602 19564 20742
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19536 19378 19564 20538
rect 19996 20466 20024 25366
rect 20088 24596 20116 27934
rect 20166 25392 20222 25401
rect 20166 25327 20222 25336
rect 20180 24818 20208 25327
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20168 24608 20220 24614
rect 20088 24568 20168 24596
rect 20168 24550 20220 24556
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 20088 23866 20116 24346
rect 20076 23860 20128 23866
rect 20180 23848 20208 24550
rect 20272 24410 20300 28426
rect 20548 28082 20576 29650
rect 20626 29608 20682 29617
rect 20626 29543 20628 29552
rect 20680 29543 20682 29552
rect 20628 29514 20680 29520
rect 20536 28076 20588 28082
rect 20536 28018 20588 28024
rect 20444 27872 20496 27878
rect 20444 27814 20496 27820
rect 20456 27538 20484 27814
rect 20444 27532 20496 27538
rect 20444 27474 20496 27480
rect 20444 26784 20496 26790
rect 20444 26726 20496 26732
rect 20456 26382 20484 26726
rect 20444 26376 20496 26382
rect 20444 26318 20496 26324
rect 20548 26234 20576 28018
rect 20732 27554 20760 31078
rect 20640 27526 20760 27554
rect 20640 26994 20668 27526
rect 20720 27328 20772 27334
rect 20720 27270 20772 27276
rect 20628 26988 20680 26994
rect 20628 26930 20680 26936
rect 20640 26761 20668 26930
rect 20626 26752 20682 26761
rect 20626 26687 20682 26696
rect 20732 26382 20760 27270
rect 20628 26376 20680 26382
rect 20628 26318 20680 26324
rect 20720 26376 20772 26382
rect 20720 26318 20772 26324
rect 20456 26206 20576 26234
rect 20352 25356 20404 25362
rect 20352 25298 20404 25304
rect 20260 24404 20312 24410
rect 20260 24346 20312 24352
rect 20180 23820 20300 23848
rect 20076 23802 20128 23808
rect 20168 23724 20220 23730
rect 20168 23666 20220 23672
rect 20180 23526 20208 23666
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 19892 20460 19944 20466
rect 19892 20402 19944 20408
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19628 19922 19656 20198
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19522 19272 19578 19281
rect 19522 19207 19524 19216
rect 19576 19207 19578 19216
rect 19524 19178 19576 19184
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19536 16658 19564 18566
rect 19628 18426 19656 19314
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19614 18320 19670 18329
rect 19614 18255 19616 18264
rect 19668 18255 19670 18264
rect 19616 18226 19668 18232
rect 19628 17678 19656 18226
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19628 17338 19656 17614
rect 19616 17332 19668 17338
rect 19616 17274 19668 17280
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19246 15736 19302 15745
rect 19246 15671 19302 15680
rect 19432 15428 19484 15434
rect 19432 15370 19484 15376
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 19260 14550 19288 14962
rect 19444 14890 19472 15370
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19432 14884 19484 14890
rect 19432 14826 19484 14832
rect 19248 14544 19300 14550
rect 19248 14486 19300 14492
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 18788 13806 18840 13812
rect 18800 12986 18828 13806
rect 18892 13790 19012 13818
rect 18892 12986 18920 13790
rect 19168 13258 19196 13874
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 18800 12850 18828 12922
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18892 12646 18920 12922
rect 19260 12850 19288 14214
rect 19536 12850 19564 14894
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19628 14006 19656 14350
rect 19616 14000 19668 14006
rect 19616 13942 19668 13948
rect 19720 13938 19748 20402
rect 19800 19916 19852 19922
rect 19800 19858 19852 19864
rect 19812 18465 19840 19858
rect 19798 18456 19854 18465
rect 19798 18391 19854 18400
rect 19812 18290 19840 18391
rect 19800 18284 19852 18290
rect 19800 18226 19852 18232
rect 19904 18086 19932 20402
rect 19984 20324 20036 20330
rect 19984 20266 20036 20272
rect 19996 19378 20024 20266
rect 20088 19922 20116 21286
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 20180 19802 20208 23462
rect 20088 19774 20208 19802
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19996 18766 20024 19314
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 19892 18080 19944 18086
rect 19798 18048 19854 18057
rect 19892 18022 19944 18028
rect 19798 17983 19854 17992
rect 19812 17746 19840 17983
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19812 16794 19840 16934
rect 19800 16788 19852 16794
rect 19800 16730 19852 16736
rect 19996 15337 20024 18158
rect 20088 16250 20116 19774
rect 20166 19544 20222 19553
rect 20166 19479 20168 19488
rect 20220 19479 20222 19488
rect 20168 19450 20220 19456
rect 20168 19304 20220 19310
rect 20166 19272 20168 19281
rect 20220 19272 20222 19281
rect 20166 19207 20222 19216
rect 20166 19000 20222 19009
rect 20166 18935 20222 18944
rect 20180 18222 20208 18935
rect 20168 18216 20220 18222
rect 20168 18158 20220 18164
rect 20272 17678 20300 23820
rect 20364 23186 20392 25298
rect 20456 24834 20484 26206
rect 20640 25498 20668 26318
rect 20824 26234 20852 31826
rect 21928 31822 21956 32846
rect 22008 32768 22060 32774
rect 22008 32710 22060 32716
rect 22020 31822 22048 32710
rect 22284 32224 22336 32230
rect 22284 32166 22336 32172
rect 22558 32192 22614 32201
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 22008 31816 22060 31822
rect 22008 31758 22060 31764
rect 22296 31754 22324 32166
rect 22558 32127 22614 32136
rect 22572 31793 22600 32127
rect 22744 31816 22796 31822
rect 22558 31784 22614 31793
rect 22296 31726 22416 31754
rect 22192 31476 22244 31482
rect 22192 31418 22244 31424
rect 22204 31226 22232 31418
rect 22296 31346 22324 31726
rect 22388 31686 22416 31726
rect 22468 31748 22520 31754
rect 22744 31758 22796 31764
rect 22558 31719 22614 31728
rect 22468 31690 22520 31696
rect 22376 31680 22428 31686
rect 22376 31622 22428 31628
rect 22480 31634 22508 31690
rect 22480 31606 22600 31634
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22468 31272 22520 31278
rect 22204 31198 22324 31226
rect 22468 31214 22520 31220
rect 22100 31136 22152 31142
rect 21730 31104 21786 31113
rect 22100 31078 22152 31084
rect 21730 31039 21786 31048
rect 21640 30320 21692 30326
rect 21640 30262 21692 30268
rect 20916 29850 21036 29866
rect 20904 29844 21036 29850
rect 20956 29838 21036 29844
rect 20904 29786 20956 29792
rect 21008 29764 21036 29838
rect 21088 29776 21140 29782
rect 21008 29736 21088 29764
rect 21088 29718 21140 29724
rect 20904 29708 20956 29714
rect 20904 29650 20956 29656
rect 21456 29708 21508 29714
rect 21456 29650 21508 29656
rect 20916 27062 20944 29650
rect 21088 29640 21140 29646
rect 21086 29608 21088 29617
rect 21140 29608 21142 29617
rect 21086 29543 21142 29552
rect 21088 27328 21140 27334
rect 21088 27270 21140 27276
rect 20904 27056 20956 27062
rect 20956 27016 21036 27044
rect 20904 26998 20956 27004
rect 20902 26752 20958 26761
rect 20902 26687 20958 26696
rect 20916 26586 20944 26687
rect 20904 26580 20956 26586
rect 20904 26522 20956 26528
rect 20824 26206 20944 26234
rect 20720 25900 20772 25906
rect 20720 25842 20772 25848
rect 20732 25809 20760 25842
rect 20718 25800 20774 25809
rect 20718 25735 20774 25744
rect 20916 25684 20944 26206
rect 20732 25656 20944 25684
rect 20628 25492 20680 25498
rect 20628 25434 20680 25440
rect 20536 25424 20588 25430
rect 20588 25372 20668 25378
rect 20536 25366 20668 25372
rect 20548 25350 20668 25366
rect 20536 25220 20588 25226
rect 20536 25162 20588 25168
rect 20548 24954 20576 25162
rect 20536 24948 20588 24954
rect 20536 24890 20588 24896
rect 20456 24806 20576 24834
rect 20640 24818 20668 25350
rect 20548 23644 20576 24806
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 20456 23616 20576 23644
rect 20352 23180 20404 23186
rect 20352 23122 20404 23128
rect 20364 22710 20392 23122
rect 20352 22704 20404 22710
rect 20352 22646 20404 22652
rect 20456 22166 20484 23616
rect 20628 23112 20680 23118
rect 20534 23080 20590 23089
rect 20628 23054 20680 23060
rect 20534 23015 20536 23024
rect 20588 23015 20590 23024
rect 20536 22986 20588 22992
rect 20536 22432 20588 22438
rect 20536 22374 20588 22380
rect 20444 22160 20496 22166
rect 20444 22102 20496 22108
rect 20548 20602 20576 22374
rect 20640 22137 20668 23054
rect 20626 22128 20682 22137
rect 20626 22063 20682 22072
rect 20628 21888 20680 21894
rect 20732 21876 20760 25656
rect 21008 23866 21036 27016
rect 21100 26518 21128 27270
rect 21180 26920 21232 26926
rect 21180 26862 21232 26868
rect 21088 26512 21140 26518
rect 21088 26454 21140 26460
rect 21088 25356 21140 25362
rect 21088 25298 21140 25304
rect 20996 23860 21048 23866
rect 20996 23802 21048 23808
rect 20996 23112 21048 23118
rect 20916 23072 20996 23100
rect 20812 22976 20864 22982
rect 20916 22953 20944 23072
rect 20996 23054 21048 23060
rect 20812 22918 20864 22924
rect 20902 22944 20958 22953
rect 20824 22817 20852 22918
rect 20902 22879 20958 22888
rect 20810 22808 20866 22817
rect 20810 22743 20866 22752
rect 20812 22636 20864 22642
rect 20916 22624 20944 22879
rect 20864 22596 20944 22624
rect 20812 22578 20864 22584
rect 20996 22568 21048 22574
rect 20996 22510 21048 22516
rect 20812 22432 20864 22438
rect 20812 22374 20864 22380
rect 20824 22234 20852 22374
rect 20812 22228 20864 22234
rect 20864 22188 20944 22216
rect 20812 22170 20864 22176
rect 20810 22128 20866 22137
rect 20810 22063 20866 22072
rect 20680 21848 20760 21876
rect 20628 21830 20680 21836
rect 20824 21690 20852 22063
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 20628 21548 20680 21554
rect 20628 21490 20680 21496
rect 20640 20874 20668 21490
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20628 20868 20680 20874
rect 20628 20810 20680 20816
rect 20536 20596 20588 20602
rect 20536 20538 20588 20544
rect 20352 20392 20404 20398
rect 20352 20334 20404 20340
rect 20364 19258 20392 20334
rect 20732 19514 20760 21422
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20824 21146 20852 21286
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20916 21010 20944 22188
rect 21008 21350 21036 22510
rect 21100 22273 21128 25298
rect 21192 24614 21220 26862
rect 21364 26376 21416 26382
rect 21364 26318 21416 26324
rect 21272 24744 21324 24750
rect 21272 24686 21324 24692
rect 21180 24608 21232 24614
rect 21180 24550 21232 24556
rect 21192 24138 21220 24550
rect 21180 24132 21232 24138
rect 21180 24074 21232 24080
rect 21178 23760 21234 23769
rect 21178 23695 21234 23704
rect 21086 22264 21142 22273
rect 21192 22234 21220 23695
rect 21086 22199 21142 22208
rect 21180 22228 21232 22234
rect 21180 22170 21232 22176
rect 21192 22094 21220 22170
rect 21284 22098 21312 24686
rect 21100 22066 21220 22094
rect 21272 22092 21324 22098
rect 21100 22001 21128 22066
rect 21272 22034 21324 22040
rect 21180 22024 21232 22030
rect 21086 21992 21142 22001
rect 21180 21966 21232 21972
rect 21086 21927 21142 21936
rect 21192 21536 21220 21966
rect 21272 21548 21324 21554
rect 21192 21508 21272 21536
rect 20996 21344 21048 21350
rect 20996 21286 21048 21292
rect 21086 21312 21142 21321
rect 20904 21004 20956 21010
rect 20904 20946 20956 20952
rect 20812 20800 20864 20806
rect 20812 20742 20864 20748
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20732 19378 20760 19450
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20628 19304 20680 19310
rect 20364 19230 20484 19258
rect 20628 19246 20680 19252
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 20272 17202 20300 17614
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 20076 16244 20128 16250
rect 20076 16186 20128 16192
rect 20088 16114 20116 16186
rect 20350 16144 20406 16153
rect 20076 16108 20128 16114
rect 20350 16079 20352 16088
rect 20076 16050 20128 16056
rect 20404 16079 20406 16088
rect 20352 16050 20404 16056
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 20180 15706 20208 15846
rect 20168 15700 20220 15706
rect 20168 15642 20220 15648
rect 19982 15328 20038 15337
rect 19982 15263 20038 15272
rect 19892 15088 19944 15094
rect 19892 15030 19944 15036
rect 19800 14408 19852 14414
rect 19800 14350 19852 14356
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19616 12912 19668 12918
rect 19616 12854 19668 12860
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19248 12708 19300 12714
rect 19248 12650 19300 12656
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 19260 12238 19288 12650
rect 19536 12238 19564 12786
rect 19628 12238 19656 12854
rect 19812 12374 19840 14350
rect 19904 12850 19932 15030
rect 19984 14884 20036 14890
rect 19984 14826 20036 14832
rect 19996 14618 20024 14826
rect 20350 14648 20406 14657
rect 19984 14612 20036 14618
rect 20350 14583 20406 14592
rect 19984 14554 20036 14560
rect 20260 14544 20312 14550
rect 20088 14492 20260 14498
rect 20088 14486 20312 14492
rect 20088 14470 20300 14486
rect 20364 14482 20392 14583
rect 20352 14476 20404 14482
rect 20088 14414 20116 14470
rect 20352 14418 20404 14424
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20180 13841 20208 14350
rect 20352 14340 20404 14346
rect 20456 14328 20484 19230
rect 20640 18970 20668 19246
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 20732 18465 20760 18634
rect 20718 18456 20774 18465
rect 20718 18391 20774 18400
rect 20536 16516 20588 16522
rect 20536 16458 20588 16464
rect 20548 16250 20576 16458
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20536 14408 20588 14414
rect 20404 14300 20484 14328
rect 20534 14376 20536 14385
rect 20588 14376 20590 14385
rect 20534 14311 20590 14320
rect 20352 14282 20404 14288
rect 20166 13832 20222 13841
rect 20166 13767 20222 13776
rect 20364 13705 20392 14282
rect 20350 13696 20406 13705
rect 20350 13631 20406 13640
rect 20076 13252 20128 13258
rect 20076 13194 20128 13200
rect 20088 12986 20116 13194
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20732 12918 20760 14826
rect 20824 14822 20852 20742
rect 20916 20466 20944 20946
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 21008 20262 21036 21286
rect 21086 21247 21142 21256
rect 20996 20256 21048 20262
rect 20996 20198 21048 20204
rect 20994 19952 21050 19961
rect 20994 19887 21050 19896
rect 21008 19718 21036 19887
rect 20996 19712 21048 19718
rect 20996 19654 21048 19660
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 20916 18426 20944 18634
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 21100 18329 21128 21247
rect 21192 20942 21220 21508
rect 21272 21490 21324 21496
rect 21180 20936 21232 20942
rect 21180 20878 21232 20884
rect 21192 20466 21220 20878
rect 21376 20806 21404 26318
rect 21468 25362 21496 29650
rect 21652 29102 21680 30262
rect 21640 29096 21692 29102
rect 21640 29038 21692 29044
rect 21640 28212 21692 28218
rect 21640 28154 21692 28160
rect 21652 27878 21680 28154
rect 21548 27872 21600 27878
rect 21548 27814 21600 27820
rect 21640 27872 21692 27878
rect 21640 27814 21692 27820
rect 21456 25356 21508 25362
rect 21456 25298 21508 25304
rect 21560 24274 21588 27814
rect 21744 27520 21772 31039
rect 21824 30592 21876 30598
rect 21824 30534 21876 30540
rect 21836 29850 21864 30534
rect 21916 30184 21968 30190
rect 21916 30126 21968 30132
rect 21928 29850 21956 30126
rect 21824 29844 21876 29850
rect 21824 29786 21876 29792
rect 21916 29844 21968 29850
rect 21916 29786 21968 29792
rect 21836 29238 21864 29786
rect 22008 29504 22060 29510
rect 22008 29446 22060 29452
rect 21824 29232 21876 29238
rect 21824 29174 21876 29180
rect 21914 29200 21970 29209
rect 21914 29135 21970 29144
rect 21928 29102 21956 29135
rect 21916 29096 21968 29102
rect 21916 29038 21968 29044
rect 21824 28960 21876 28966
rect 21824 28902 21876 28908
rect 21836 28762 21864 28902
rect 21824 28756 21876 28762
rect 21824 28698 21876 28704
rect 21836 27713 21864 28698
rect 22020 27946 22048 29446
rect 21916 27940 21968 27946
rect 21916 27882 21968 27888
rect 22008 27940 22060 27946
rect 22008 27882 22060 27888
rect 21822 27704 21878 27713
rect 21928 27674 21956 27882
rect 21822 27639 21878 27648
rect 21916 27668 21968 27674
rect 21916 27610 21968 27616
rect 21744 27492 22048 27520
rect 21732 27396 21784 27402
rect 21732 27338 21784 27344
rect 21916 27396 21968 27402
rect 21916 27338 21968 27344
rect 21456 24268 21508 24274
rect 21456 24210 21508 24216
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 21468 22642 21496 24210
rect 21548 22704 21600 22710
rect 21548 22646 21600 22652
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 21364 20800 21416 20806
rect 21364 20742 21416 20748
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 21364 20392 21416 20398
rect 21364 20334 21416 20340
rect 21270 19952 21326 19961
rect 21270 19887 21326 19896
rect 21178 19272 21234 19281
rect 21178 19207 21234 19216
rect 21192 18902 21220 19207
rect 21284 19174 21312 19887
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21180 18896 21232 18902
rect 21180 18838 21232 18844
rect 21086 18320 21142 18329
rect 21086 18255 21142 18264
rect 21100 16794 21128 18255
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 20994 15872 21050 15881
rect 20994 15807 21050 15816
rect 21008 15473 21036 15807
rect 20994 15464 21050 15473
rect 20994 15399 21050 15408
rect 21192 15162 21220 16526
rect 21376 15881 21404 20334
rect 21468 20330 21496 22578
rect 21560 22234 21588 22646
rect 21548 22228 21600 22234
rect 21548 22170 21600 22176
rect 21640 22092 21692 22098
rect 21640 22034 21692 22040
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21560 21078 21588 21286
rect 21548 21072 21600 21078
rect 21548 21014 21600 21020
rect 21548 20936 21600 20942
rect 21548 20878 21600 20884
rect 21560 20466 21588 20878
rect 21548 20460 21600 20466
rect 21548 20402 21600 20408
rect 21456 20324 21508 20330
rect 21456 20266 21508 20272
rect 21548 19440 21600 19446
rect 21548 19382 21600 19388
rect 21456 19236 21508 19242
rect 21456 19178 21508 19184
rect 21468 18358 21496 19178
rect 21560 18766 21588 19382
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 21548 18624 21600 18630
rect 21548 18566 21600 18572
rect 21456 18352 21508 18358
rect 21456 18294 21508 18300
rect 21560 18222 21588 18566
rect 21548 18216 21600 18222
rect 21548 18158 21600 18164
rect 21652 16046 21680 22034
rect 21744 21010 21772 27338
rect 21824 26444 21876 26450
rect 21824 26386 21876 26392
rect 21836 26042 21864 26386
rect 21824 26036 21876 26042
rect 21824 25978 21876 25984
rect 21824 22432 21876 22438
rect 21824 22374 21876 22380
rect 21836 21894 21864 22374
rect 21824 21888 21876 21894
rect 21824 21830 21876 21836
rect 21732 21004 21784 21010
rect 21732 20946 21784 20952
rect 21824 20800 21876 20806
rect 21824 20742 21876 20748
rect 21732 19168 21784 19174
rect 21732 19110 21784 19116
rect 21744 18970 21772 19110
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21836 18766 21864 20742
rect 21928 19258 21956 27338
rect 22020 20398 22048 27492
rect 22112 26586 22140 31078
rect 22192 29164 22244 29170
rect 22192 29106 22244 29112
rect 22204 28490 22232 29106
rect 22192 28484 22244 28490
rect 22192 28426 22244 28432
rect 22204 28393 22232 28426
rect 22190 28384 22246 28393
rect 22190 28319 22246 28328
rect 22192 27464 22244 27470
rect 22192 27406 22244 27412
rect 22204 27130 22232 27406
rect 22192 27124 22244 27130
rect 22192 27066 22244 27072
rect 22190 27024 22246 27033
rect 22190 26959 22246 26968
rect 22204 26586 22232 26959
rect 22100 26580 22152 26586
rect 22100 26522 22152 26528
rect 22192 26580 22244 26586
rect 22192 26522 22244 26528
rect 22100 26444 22152 26450
rect 22100 26386 22152 26392
rect 22112 25838 22140 26386
rect 22100 25832 22152 25838
rect 22100 25774 22152 25780
rect 22296 25226 22324 31198
rect 22376 31136 22428 31142
rect 22376 31078 22428 31084
rect 22388 30054 22416 31078
rect 22480 30841 22508 31214
rect 22572 30938 22600 31606
rect 22756 31482 22784 31758
rect 22744 31476 22796 31482
rect 22744 31418 22796 31424
rect 22560 30932 22612 30938
rect 22560 30874 22612 30880
rect 22466 30832 22522 30841
rect 22466 30767 22522 30776
rect 22572 30394 22600 30874
rect 22744 30728 22796 30734
rect 22744 30670 22796 30676
rect 22468 30388 22520 30394
rect 22468 30330 22520 30336
rect 22560 30388 22612 30394
rect 22560 30330 22612 30336
rect 22376 30048 22428 30054
rect 22376 29990 22428 29996
rect 22374 29880 22430 29889
rect 22374 29815 22430 29824
rect 22388 27334 22416 29815
rect 22480 29492 22508 30330
rect 22652 30252 22704 30258
rect 22652 30194 22704 30200
rect 22664 30025 22692 30194
rect 22650 30016 22706 30025
rect 22650 29951 22706 29960
rect 22652 29504 22704 29510
rect 22480 29464 22652 29492
rect 22652 29446 22704 29452
rect 22468 28960 22520 28966
rect 22468 28902 22520 28908
rect 22376 27328 22428 27334
rect 22376 27270 22428 27276
rect 22376 26920 22428 26926
rect 22376 26862 22428 26868
rect 22388 25702 22416 26862
rect 22376 25696 22428 25702
rect 22376 25638 22428 25644
rect 22376 25492 22428 25498
rect 22376 25434 22428 25440
rect 22284 25220 22336 25226
rect 22204 25180 22284 25208
rect 22098 24576 22154 24585
rect 22098 24511 22154 24520
rect 22112 24313 22140 24511
rect 22098 24304 22154 24313
rect 22098 24239 22154 24248
rect 22100 23520 22152 23526
rect 22100 23462 22152 23468
rect 22112 22710 22140 23462
rect 22204 23254 22232 25180
rect 22284 25162 22336 25168
rect 22284 24268 22336 24274
rect 22284 24210 22336 24216
rect 22296 24041 22324 24210
rect 22282 24032 22338 24041
rect 22282 23967 22338 23976
rect 22282 23624 22338 23633
rect 22282 23559 22284 23568
rect 22336 23559 22338 23568
rect 22284 23530 22336 23536
rect 22282 23488 22338 23497
rect 22282 23423 22338 23432
rect 22192 23248 22244 23254
rect 22192 23190 22244 23196
rect 22100 22704 22152 22710
rect 22100 22646 22152 22652
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 22204 22080 22232 22578
rect 22296 22438 22324 23423
rect 22388 23338 22416 25434
rect 22480 23497 22508 28902
rect 22560 27668 22612 27674
rect 22560 27610 22612 27616
rect 22572 26790 22600 27610
rect 22560 26784 22612 26790
rect 22560 26726 22612 26732
rect 22572 25498 22600 26726
rect 22664 25906 22692 29446
rect 22756 29238 22784 30670
rect 22744 29232 22796 29238
rect 22744 29174 22796 29180
rect 22848 28762 22876 34138
rect 23124 33658 23152 34138
rect 23112 33652 23164 33658
rect 23112 33594 23164 33600
rect 23216 33522 23244 34138
rect 23308 33658 23336 34954
rect 23400 34202 23428 37130
rect 23676 35154 23704 37130
rect 23664 35148 23716 35154
rect 23664 35090 23716 35096
rect 23572 35012 23624 35018
rect 23572 34954 23624 34960
rect 23584 34746 23612 34954
rect 23676 34746 23704 35090
rect 24124 34944 24176 34950
rect 24124 34886 24176 34892
rect 23572 34740 23624 34746
rect 23572 34682 23624 34688
rect 23664 34740 23716 34746
rect 23664 34682 23716 34688
rect 23664 34604 23716 34610
rect 23664 34546 23716 34552
rect 23676 34202 23704 34546
rect 24136 34202 24164 34886
rect 25608 34746 25636 37130
rect 26976 35012 27028 35018
rect 26976 34954 27028 34960
rect 25596 34740 25648 34746
rect 25596 34682 25648 34688
rect 25608 34610 25636 34682
rect 24308 34604 24360 34610
rect 24308 34546 24360 34552
rect 25596 34604 25648 34610
rect 25596 34546 25648 34552
rect 24320 34202 24348 34546
rect 25504 34400 25556 34406
rect 25504 34342 25556 34348
rect 23388 34196 23440 34202
rect 23388 34138 23440 34144
rect 23664 34196 23716 34202
rect 23664 34138 23716 34144
rect 24124 34196 24176 34202
rect 24124 34138 24176 34144
rect 24308 34196 24360 34202
rect 24308 34138 24360 34144
rect 25516 33998 25544 34342
rect 23388 33992 23440 33998
rect 23388 33934 23440 33940
rect 24584 33992 24636 33998
rect 24584 33934 24636 33940
rect 24768 33992 24820 33998
rect 24768 33934 24820 33940
rect 25504 33992 25556 33998
rect 25504 33934 25556 33940
rect 23400 33658 23428 33934
rect 23480 33924 23532 33930
rect 23480 33866 23532 33872
rect 23296 33652 23348 33658
rect 23296 33594 23348 33600
rect 23388 33652 23440 33658
rect 23388 33594 23440 33600
rect 23204 33516 23256 33522
rect 23204 33458 23256 33464
rect 22928 33448 22980 33454
rect 22928 33390 22980 33396
rect 22836 28756 22888 28762
rect 22836 28698 22888 28704
rect 22836 28008 22888 28014
rect 22836 27950 22888 27956
rect 22848 25945 22876 27950
rect 22940 27606 22968 33390
rect 23388 32972 23440 32978
rect 23388 32914 23440 32920
rect 23112 32564 23164 32570
rect 23112 32506 23164 32512
rect 23020 32496 23072 32502
rect 23020 32438 23072 32444
rect 23032 32298 23060 32438
rect 23020 32292 23072 32298
rect 23020 32234 23072 32240
rect 23032 32026 23060 32234
rect 23020 32020 23072 32026
rect 23020 31962 23072 31968
rect 23020 31816 23072 31822
rect 23020 31758 23072 31764
rect 23032 30802 23060 31758
rect 23020 30796 23072 30802
rect 23020 30738 23072 30744
rect 23020 30252 23072 30258
rect 23020 30194 23072 30200
rect 23032 29510 23060 30194
rect 23020 29504 23072 29510
rect 23020 29446 23072 29452
rect 23124 28994 23152 32506
rect 23296 32428 23348 32434
rect 23296 32370 23348 32376
rect 23204 32224 23256 32230
rect 23204 32166 23256 32172
rect 23216 32026 23244 32166
rect 23308 32065 23336 32370
rect 23294 32056 23350 32065
rect 23204 32020 23256 32026
rect 23294 31991 23350 32000
rect 23204 31962 23256 31968
rect 23400 31754 23428 32914
rect 23492 32570 23520 33866
rect 24596 33590 24624 33934
rect 24584 33584 24636 33590
rect 24584 33526 24636 33532
rect 23572 33380 23624 33386
rect 23572 33322 23624 33328
rect 23584 32570 23612 33322
rect 24780 33289 24808 33934
rect 26148 33924 26200 33930
rect 26148 33866 26200 33872
rect 26160 33658 26188 33866
rect 26608 33856 26660 33862
rect 26608 33798 26660 33804
rect 26148 33652 26200 33658
rect 26148 33594 26200 33600
rect 26620 33454 26648 33798
rect 26516 33448 26568 33454
rect 26516 33390 26568 33396
rect 26608 33448 26660 33454
rect 26608 33390 26660 33396
rect 24766 33280 24822 33289
rect 24766 33215 24822 33224
rect 26148 32768 26200 32774
rect 26148 32710 26200 32716
rect 23480 32564 23532 32570
rect 23480 32506 23532 32512
rect 23572 32564 23624 32570
rect 23572 32506 23624 32512
rect 23756 32360 23808 32366
rect 23756 32302 23808 32308
rect 24032 32360 24084 32366
rect 24032 32302 24084 32308
rect 23768 32026 23796 32302
rect 23940 32224 23992 32230
rect 23940 32166 23992 32172
rect 23952 32026 23980 32166
rect 23756 32020 23808 32026
rect 23756 31962 23808 31968
rect 23940 32020 23992 32026
rect 23940 31962 23992 31968
rect 23940 31816 23992 31822
rect 23938 31784 23940 31793
rect 23992 31784 23994 31793
rect 23308 31726 23428 31754
rect 23480 31748 23532 31754
rect 23308 31278 23336 31726
rect 23938 31719 23994 31728
rect 23480 31690 23532 31696
rect 23388 31340 23440 31346
rect 23388 31282 23440 31288
rect 23296 31272 23348 31278
rect 23296 31214 23348 31220
rect 23204 29504 23256 29510
rect 23204 29446 23256 29452
rect 23032 28966 23152 28994
rect 23216 28966 23244 29446
rect 23308 29170 23336 31214
rect 23400 30161 23428 31282
rect 23492 30938 23520 31690
rect 23572 31340 23624 31346
rect 23572 31282 23624 31288
rect 23584 30938 23612 31282
rect 23480 30932 23532 30938
rect 23480 30874 23532 30880
rect 23572 30932 23624 30938
rect 23572 30874 23624 30880
rect 23480 30252 23532 30258
rect 23480 30194 23532 30200
rect 23386 30152 23442 30161
rect 23492 30122 23520 30194
rect 23386 30087 23442 30096
rect 23480 30116 23532 30122
rect 23480 30058 23532 30064
rect 23388 30048 23440 30054
rect 23388 29990 23440 29996
rect 23296 29164 23348 29170
rect 23296 29106 23348 29112
rect 23400 29034 23428 29990
rect 23492 29170 23520 30058
rect 23480 29164 23532 29170
rect 23480 29106 23532 29112
rect 23296 29028 23348 29034
rect 23296 28970 23348 28976
rect 23388 29028 23440 29034
rect 23388 28970 23440 28976
rect 22928 27600 22980 27606
rect 22928 27542 22980 27548
rect 22834 25936 22890 25945
rect 22652 25900 22704 25906
rect 22834 25871 22890 25880
rect 22652 25842 22704 25848
rect 22560 25492 22612 25498
rect 22560 25434 22612 25440
rect 22560 24812 22612 24818
rect 22560 24754 22612 24760
rect 22572 24449 22600 24754
rect 22558 24440 22614 24449
rect 22558 24375 22614 24384
rect 22664 24324 22692 25842
rect 22836 25696 22888 25702
rect 22836 25638 22888 25644
rect 22848 24614 22876 25638
rect 22928 24812 22980 24818
rect 22928 24754 22980 24760
rect 22744 24608 22796 24614
rect 22744 24550 22796 24556
rect 22836 24608 22888 24614
rect 22940 24585 22968 24754
rect 22836 24550 22888 24556
rect 22926 24576 22982 24585
rect 22572 24296 22692 24324
rect 22466 23488 22522 23497
rect 22466 23423 22522 23432
rect 22388 23310 22508 23338
rect 22284 22432 22336 22438
rect 22284 22374 22336 22380
rect 22376 22432 22428 22438
rect 22376 22374 22428 22380
rect 22388 22273 22416 22374
rect 22374 22264 22430 22273
rect 22374 22199 22430 22208
rect 22204 22052 22324 22080
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 22008 20392 22060 20398
rect 22008 20334 22060 20340
rect 22112 19786 22140 20402
rect 22100 19780 22152 19786
rect 22100 19722 22152 19728
rect 22192 19780 22244 19786
rect 22192 19722 22244 19728
rect 22008 19712 22060 19718
rect 22008 19654 22060 19660
rect 22098 19680 22154 19689
rect 22020 19378 22048 19654
rect 22098 19615 22154 19624
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 21928 19230 22048 19258
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 21928 18834 21956 19110
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 21824 18760 21876 18766
rect 21824 18702 21876 18708
rect 22020 16250 22048 19230
rect 22112 19174 22140 19615
rect 22204 19378 22232 19722
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22296 19334 22324 22052
rect 22480 19334 22508 23310
rect 22572 23202 22600 24296
rect 22652 24132 22704 24138
rect 22652 24074 22704 24080
rect 22664 23769 22692 24074
rect 22650 23760 22706 23769
rect 22650 23695 22706 23704
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22664 23322 22692 23598
rect 22652 23316 22704 23322
rect 22652 23258 22704 23264
rect 22572 23174 22692 23202
rect 22664 20466 22692 23174
rect 22652 20460 22704 20466
rect 22652 20402 22704 20408
rect 22652 20256 22704 20262
rect 22650 20224 22652 20233
rect 22704 20224 22706 20233
rect 22650 20159 22706 20168
rect 22664 19553 22692 20159
rect 22650 19544 22706 19553
rect 22650 19479 22706 19488
rect 22296 19306 22416 19334
rect 22480 19306 22600 19334
rect 22284 19236 22336 19242
rect 22284 19178 22336 19184
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22296 19009 22324 19178
rect 22282 19000 22338 19009
rect 22282 18935 22338 18944
rect 22100 18896 22152 18902
rect 22100 18838 22152 18844
rect 22112 18698 22140 18838
rect 22190 18728 22246 18737
rect 22100 18692 22152 18698
rect 22388 18714 22416 19306
rect 22466 19000 22522 19009
rect 22466 18935 22522 18944
rect 22190 18663 22246 18672
rect 22296 18686 22416 18714
rect 22100 18634 22152 18640
rect 22204 18290 22232 18663
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22190 17912 22246 17921
rect 22190 17847 22246 17856
rect 22204 17678 22232 17847
rect 22192 17672 22244 17678
rect 22192 17614 22244 17620
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22112 17338 22140 17478
rect 22100 17332 22152 17338
rect 22100 17274 22152 17280
rect 22204 16590 22232 17478
rect 22296 16794 22324 18686
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22388 18290 22416 18566
rect 22480 18465 22508 18935
rect 22466 18456 22522 18465
rect 22466 18391 22522 18400
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22376 18080 22428 18086
rect 22376 18022 22428 18028
rect 22388 17678 22416 18022
rect 22376 17672 22428 17678
rect 22376 17614 22428 17620
rect 22374 17504 22430 17513
rect 22374 17439 22430 17448
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22296 16658 22324 16730
rect 22284 16652 22336 16658
rect 22284 16594 22336 16600
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 22008 16244 22060 16250
rect 22008 16186 22060 16192
rect 21640 16040 21692 16046
rect 21640 15982 21692 15988
rect 22098 16008 22154 16017
rect 21362 15872 21418 15881
rect 21362 15807 21418 15816
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 21652 14890 21680 15982
rect 22098 15943 22154 15952
rect 22112 15910 22140 15943
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 22112 15609 22140 15846
rect 22098 15600 22154 15609
rect 22098 15535 22154 15544
rect 22098 15328 22154 15337
rect 22098 15263 22154 15272
rect 21640 14884 21692 14890
rect 21640 14826 21692 14832
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 22112 14550 22140 15263
rect 22100 14544 22152 14550
rect 22100 14486 22152 14492
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 22006 14376 22062 14385
rect 21744 13870 21772 14350
rect 22006 14311 22062 14320
rect 22020 14278 22048 14311
rect 21916 14272 21968 14278
rect 21916 14214 21968 14220
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 21928 13988 21956 14214
rect 22204 14006 22232 16390
rect 22296 16182 22324 16458
rect 22284 16176 22336 16182
rect 22284 16118 22336 16124
rect 22388 16114 22416 17439
rect 22480 16182 22508 18226
rect 22572 17762 22600 19306
rect 22650 18184 22706 18193
rect 22650 18119 22652 18128
rect 22704 18119 22706 18128
rect 22652 18090 22704 18096
rect 22572 17734 22692 17762
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22572 16794 22600 17614
rect 22560 16788 22612 16794
rect 22560 16730 22612 16736
rect 22664 16674 22692 17734
rect 22756 17202 22784 24550
rect 22926 24511 22982 24520
rect 22836 24404 22888 24410
rect 23032 24392 23060 28966
rect 23204 28960 23256 28966
rect 23204 28902 23256 28908
rect 23308 28762 23336 28970
rect 23296 28756 23348 28762
rect 23296 28698 23348 28704
rect 23204 28620 23256 28626
rect 23204 28562 23256 28568
rect 23112 28552 23164 28558
rect 23112 28494 23164 28500
rect 22888 24364 23060 24392
rect 22836 24346 22888 24352
rect 22848 24313 22876 24346
rect 23124 24342 23152 28494
rect 23216 26926 23244 28562
rect 23308 27860 23336 28698
rect 23386 28656 23442 28665
rect 23386 28591 23388 28600
rect 23440 28591 23442 28600
rect 23388 28562 23440 28568
rect 23388 28484 23440 28490
rect 23388 28426 23440 28432
rect 23400 27985 23428 28426
rect 23480 28008 23532 28014
rect 23386 27976 23442 27985
rect 23480 27950 23532 27956
rect 23386 27911 23442 27920
rect 23388 27872 23440 27878
rect 23308 27832 23388 27860
rect 23388 27814 23440 27820
rect 23296 27396 23348 27402
rect 23296 27338 23348 27344
rect 23204 26920 23256 26926
rect 23204 26862 23256 26868
rect 23308 26858 23336 27338
rect 23296 26852 23348 26858
rect 23296 26794 23348 26800
rect 23492 26625 23520 27950
rect 23478 26616 23534 26625
rect 23204 26580 23256 26586
rect 23478 26551 23534 26560
rect 23204 26522 23256 26528
rect 23216 25702 23244 26522
rect 23480 26240 23532 26246
rect 23480 26182 23532 26188
rect 23492 25906 23520 26182
rect 23296 25900 23348 25906
rect 23296 25842 23348 25848
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 23204 25696 23256 25702
rect 23204 25638 23256 25644
rect 23204 25152 23256 25158
rect 23204 25094 23256 25100
rect 23112 24336 23164 24342
rect 22834 24304 22890 24313
rect 22834 24239 22890 24248
rect 23018 24304 23074 24313
rect 23112 24278 23164 24284
rect 23018 24239 23074 24248
rect 23032 24206 23060 24239
rect 22836 24200 22888 24206
rect 22836 24142 22888 24148
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 22848 22642 22876 24142
rect 23124 23746 23152 24278
rect 23216 24274 23244 25094
rect 23204 24268 23256 24274
rect 23204 24210 23256 24216
rect 23124 23718 23244 23746
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 22940 23225 22968 23462
rect 22926 23216 22982 23225
rect 22926 23151 22982 23160
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 23112 21480 23164 21486
rect 23112 21422 23164 21428
rect 23124 21010 23152 21422
rect 23112 21004 23164 21010
rect 23112 20946 23164 20952
rect 22834 20904 22890 20913
rect 22834 20839 22890 20848
rect 22848 18465 22876 20839
rect 23112 20596 23164 20602
rect 23112 20538 23164 20544
rect 23020 20392 23072 20398
rect 23020 20334 23072 20340
rect 22928 19304 22980 19310
rect 22928 19246 22980 19252
rect 22834 18456 22890 18465
rect 22834 18391 22890 18400
rect 22940 18358 22968 19246
rect 22928 18352 22980 18358
rect 22928 18294 22980 18300
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22848 17882 22876 18226
rect 22928 18216 22980 18222
rect 22928 18158 22980 18164
rect 22836 17876 22888 17882
rect 22836 17818 22888 17824
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22756 16810 22784 17138
rect 22756 16782 22876 16810
rect 22664 16646 22784 16674
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22468 16176 22520 16182
rect 22468 16118 22520 16124
rect 22664 16114 22692 16526
rect 22756 16454 22784 16646
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22756 16250 22784 16390
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22652 16108 22704 16114
rect 22704 16068 22784 16096
rect 22652 16050 22704 16056
rect 22282 16008 22338 16017
rect 22282 15943 22338 15952
rect 22296 15706 22324 15943
rect 22284 15700 22336 15706
rect 22284 15642 22336 15648
rect 22388 15502 22416 16050
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 22466 15872 22522 15881
rect 22466 15807 22522 15816
rect 22480 15570 22508 15807
rect 22572 15706 22600 15982
rect 22756 15978 22784 16068
rect 22652 15972 22704 15978
rect 22652 15914 22704 15920
rect 22744 15972 22796 15978
rect 22744 15914 22796 15920
rect 22664 15881 22692 15914
rect 22650 15872 22706 15881
rect 22650 15807 22706 15816
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22468 15564 22520 15570
rect 22468 15506 22520 15512
rect 22376 15496 22428 15502
rect 22282 15464 22338 15473
rect 22376 15438 22428 15444
rect 22282 15399 22284 15408
rect 22336 15399 22338 15408
rect 22284 15370 22336 15376
rect 22466 14512 22522 14521
rect 22466 14447 22522 14456
rect 22560 14476 22612 14482
rect 22480 14346 22508 14447
rect 22560 14418 22612 14424
rect 22468 14340 22520 14346
rect 22468 14282 22520 14288
rect 22008 14000 22060 14006
rect 21928 13960 22008 13988
rect 22008 13942 22060 13948
rect 22192 14000 22244 14006
rect 22572 13954 22600 14418
rect 22848 14006 22876 16782
rect 22940 14618 22968 18158
rect 23032 18086 23060 20334
rect 23124 20330 23152 20538
rect 23112 20324 23164 20330
rect 23112 20266 23164 20272
rect 23112 19780 23164 19786
rect 23112 19722 23164 19728
rect 23124 19689 23152 19722
rect 23110 19680 23166 19689
rect 23110 19615 23166 19624
rect 23112 19440 23164 19446
rect 23112 19382 23164 19388
rect 23020 18080 23072 18086
rect 23020 18022 23072 18028
rect 23032 17746 23060 18022
rect 23020 17740 23072 17746
rect 23020 17682 23072 17688
rect 23018 17640 23074 17649
rect 23018 17575 23020 17584
rect 23072 17575 23074 17584
rect 23020 17546 23072 17552
rect 23124 17338 23152 19382
rect 23216 17762 23244 23718
rect 23308 22681 23336 25842
rect 23584 25786 23612 30874
rect 23756 30728 23808 30734
rect 23756 30670 23808 30676
rect 23768 26586 23796 30670
rect 23940 30660 23992 30666
rect 23940 30602 23992 30608
rect 23848 30320 23900 30326
rect 23848 30262 23900 30268
rect 23860 29306 23888 30262
rect 23952 30122 23980 30602
rect 24044 30410 24072 32302
rect 25688 32292 25740 32298
rect 25688 32234 25740 32240
rect 24122 32192 24178 32201
rect 24122 32127 24178 32136
rect 24136 31822 24164 32127
rect 24124 31816 24176 31822
rect 24124 31758 24176 31764
rect 24492 30932 24544 30938
rect 24492 30874 24544 30880
rect 24044 30382 24164 30410
rect 24504 30394 24532 30874
rect 24768 30728 24820 30734
rect 24768 30670 24820 30676
rect 24780 30569 24808 30670
rect 25504 30592 25556 30598
rect 24766 30560 24822 30569
rect 25504 30534 25556 30540
rect 24766 30495 24822 30504
rect 24032 30252 24084 30258
rect 24032 30194 24084 30200
rect 23940 30116 23992 30122
rect 23940 30058 23992 30064
rect 24044 29345 24072 30194
rect 24030 29336 24086 29345
rect 23848 29300 23900 29306
rect 24030 29271 24086 29280
rect 23848 29242 23900 29248
rect 24136 29073 24164 30382
rect 24308 30388 24360 30394
rect 24308 30330 24360 30336
rect 24492 30388 24544 30394
rect 24492 30330 24544 30336
rect 24216 30320 24268 30326
rect 24216 30262 24268 30268
rect 24228 30190 24256 30262
rect 24216 30184 24268 30190
rect 24216 30126 24268 30132
rect 24228 29714 24256 30126
rect 24216 29708 24268 29714
rect 24216 29650 24268 29656
rect 24122 29064 24178 29073
rect 24122 28999 24178 29008
rect 24124 28076 24176 28082
rect 24124 28018 24176 28024
rect 24216 28076 24268 28082
rect 24216 28018 24268 28024
rect 23940 26852 23992 26858
rect 23940 26794 23992 26800
rect 23756 26580 23808 26586
rect 23756 26522 23808 26528
rect 23768 26314 23796 26522
rect 23952 26518 23980 26794
rect 23940 26512 23992 26518
rect 23940 26454 23992 26460
rect 24032 26512 24084 26518
rect 24032 26454 24084 26460
rect 23756 26308 23808 26314
rect 23756 26250 23808 26256
rect 23756 25968 23808 25974
rect 23808 25928 23980 25956
rect 23756 25910 23808 25916
rect 23664 25900 23716 25906
rect 23664 25842 23716 25848
rect 23492 25758 23612 25786
rect 23388 25356 23440 25362
rect 23388 25298 23440 25304
rect 23400 24993 23428 25298
rect 23386 24984 23442 24993
rect 23386 24919 23442 24928
rect 23388 24064 23440 24070
rect 23388 24006 23440 24012
rect 23400 23186 23428 24006
rect 23388 23180 23440 23186
rect 23388 23122 23440 23128
rect 23492 23118 23520 25758
rect 23676 25673 23704 25842
rect 23756 25696 23808 25702
rect 23662 25664 23718 25673
rect 23756 25638 23808 25644
rect 23662 25599 23718 25608
rect 23768 25498 23796 25638
rect 23756 25492 23808 25498
rect 23756 25434 23808 25440
rect 23572 25288 23624 25294
rect 23572 25230 23624 25236
rect 23584 25129 23612 25230
rect 23570 25120 23626 25129
rect 23570 25055 23626 25064
rect 23846 24576 23902 24585
rect 23846 24511 23902 24520
rect 23754 24440 23810 24449
rect 23860 24410 23888 24511
rect 23754 24375 23810 24384
rect 23848 24404 23900 24410
rect 23572 24268 23624 24274
rect 23572 24210 23624 24216
rect 23584 23662 23612 24210
rect 23572 23656 23624 23662
rect 23572 23598 23624 23604
rect 23768 23594 23796 24375
rect 23848 24346 23900 24352
rect 23848 24132 23900 24138
rect 23848 24074 23900 24080
rect 23756 23588 23808 23594
rect 23756 23530 23808 23536
rect 23756 23316 23808 23322
rect 23756 23258 23808 23264
rect 23480 23112 23532 23118
rect 23664 23112 23716 23118
rect 23480 23054 23532 23060
rect 23584 23072 23664 23100
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23492 22681 23520 22918
rect 23294 22672 23350 22681
rect 23294 22607 23350 22616
rect 23478 22672 23534 22681
rect 23478 22607 23534 22616
rect 23308 20942 23336 22607
rect 23584 22409 23612 23072
rect 23664 23054 23716 23060
rect 23664 22976 23716 22982
rect 23664 22918 23716 22924
rect 23676 22778 23704 22918
rect 23664 22772 23716 22778
rect 23664 22714 23716 22720
rect 23570 22400 23626 22409
rect 23570 22335 23626 22344
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 23296 20936 23348 20942
rect 23296 20878 23348 20884
rect 23294 20768 23350 20777
rect 23294 20703 23350 20712
rect 23308 18426 23336 20703
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 23400 20233 23428 20402
rect 23386 20224 23442 20233
rect 23386 20159 23442 20168
rect 23492 19854 23520 21286
rect 23584 19854 23612 22335
rect 23768 21457 23796 23258
rect 23860 22982 23888 24074
rect 23848 22976 23900 22982
rect 23848 22918 23900 22924
rect 23846 22808 23902 22817
rect 23846 22743 23902 22752
rect 23860 21554 23888 22743
rect 23952 22681 23980 25928
rect 23938 22672 23994 22681
rect 23938 22607 23994 22616
rect 23940 22432 23992 22438
rect 23940 22374 23992 22380
rect 23952 21622 23980 22374
rect 23940 21616 23992 21622
rect 23940 21558 23992 21564
rect 23848 21548 23900 21554
rect 23848 21490 23900 21496
rect 23754 21448 23810 21457
rect 23754 21383 23810 21392
rect 23848 21412 23900 21418
rect 23848 21354 23900 21360
rect 23664 20868 23716 20874
rect 23664 20810 23716 20816
rect 23676 20602 23704 20810
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 23756 20460 23808 20466
rect 23756 20402 23808 20408
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23572 19848 23624 19854
rect 23572 19790 23624 19796
rect 23388 19780 23440 19786
rect 23388 19722 23440 19728
rect 23400 19446 23428 19722
rect 23676 19514 23704 20198
rect 23768 19854 23796 20402
rect 23860 20262 23888 21354
rect 24044 21350 24072 26454
rect 24136 24410 24164 28018
rect 24228 26790 24256 28018
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 24214 26616 24270 26625
rect 24214 26551 24270 26560
rect 24124 24404 24176 24410
rect 24124 24346 24176 24352
rect 24136 24070 24164 24346
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 24124 23792 24176 23798
rect 24124 23734 24176 23740
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 23938 20632 23994 20641
rect 23938 20567 23994 20576
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23848 20052 23900 20058
rect 23848 19994 23900 20000
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 23664 19508 23716 19514
rect 23664 19450 23716 19456
rect 23388 19440 23440 19446
rect 23388 19382 23440 19388
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23492 18834 23520 18906
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23296 18420 23348 18426
rect 23296 18362 23348 18368
rect 23388 18216 23440 18222
rect 23388 18158 23440 18164
rect 23400 18057 23428 18158
rect 23492 18086 23520 18770
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23480 18080 23532 18086
rect 23386 18048 23442 18057
rect 23480 18022 23532 18028
rect 23386 17983 23442 17992
rect 23584 17882 23612 18226
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23216 17734 23336 17762
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 23124 16794 23152 17274
rect 23216 17270 23244 17614
rect 23204 17264 23256 17270
rect 23204 17206 23256 17212
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 23018 16416 23074 16425
rect 23018 16351 23074 16360
rect 23032 15910 23060 16351
rect 23020 15904 23072 15910
rect 23020 15846 23072 15852
rect 23204 15904 23256 15910
rect 23204 15846 23256 15852
rect 23032 15026 23060 15846
rect 23216 15502 23244 15846
rect 23204 15496 23256 15502
rect 23204 15438 23256 15444
rect 23308 15434 23336 17734
rect 23388 16108 23440 16114
rect 23388 16050 23440 16056
rect 23296 15428 23348 15434
rect 23296 15370 23348 15376
rect 23400 15337 23428 16050
rect 23386 15328 23442 15337
rect 23386 15263 23442 15272
rect 23676 15026 23704 19450
rect 23756 18080 23808 18086
rect 23860 18068 23888 19994
rect 23808 18040 23888 18068
rect 23756 18022 23808 18028
rect 23768 15366 23796 18022
rect 23952 15994 23980 20567
rect 24032 20460 24084 20466
rect 24032 20402 24084 20408
rect 24044 19310 24072 20402
rect 24136 20398 24164 23734
rect 24228 22094 24256 26551
rect 24320 22522 24348 30330
rect 24492 30116 24544 30122
rect 24492 30058 24544 30064
rect 24504 29782 24532 30058
rect 24492 29776 24544 29782
rect 24492 29718 24544 29724
rect 24400 29708 24452 29714
rect 24400 29650 24452 29656
rect 24412 29510 24440 29650
rect 24400 29504 24452 29510
rect 24400 29446 24452 29452
rect 24582 29336 24638 29345
rect 24582 29271 24638 29280
rect 24492 28008 24544 28014
rect 24492 27950 24544 27956
rect 24400 27328 24452 27334
rect 24504 27316 24532 27950
rect 24452 27288 24532 27316
rect 24400 27270 24452 27276
rect 24412 27062 24440 27270
rect 24400 27056 24452 27062
rect 24400 26998 24452 27004
rect 24596 26874 24624 29271
rect 24766 29200 24822 29209
rect 24766 29135 24822 29144
rect 24860 29164 24912 29170
rect 24676 27328 24728 27334
rect 24676 27270 24728 27276
rect 24688 27130 24716 27270
rect 24676 27124 24728 27130
rect 24676 27066 24728 27072
rect 24780 26994 24808 29135
rect 24860 29106 24912 29112
rect 24872 28082 24900 29106
rect 25042 29064 25098 29073
rect 25042 28999 25098 29008
rect 25056 28966 25084 28999
rect 24952 28960 25004 28966
rect 24952 28902 25004 28908
rect 25044 28960 25096 28966
rect 25044 28902 25096 28908
rect 24964 28490 24992 28902
rect 25516 28626 25544 30534
rect 25504 28620 25556 28626
rect 25504 28562 25556 28568
rect 24952 28484 25004 28490
rect 24952 28426 25004 28432
rect 25596 28484 25648 28490
rect 25596 28426 25648 28432
rect 24860 28076 24912 28082
rect 24860 28018 24912 28024
rect 25044 28076 25096 28082
rect 25044 28018 25096 28024
rect 24676 26988 24728 26994
rect 24676 26930 24728 26936
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24504 26846 24624 26874
rect 24400 25832 24452 25838
rect 24398 25800 24400 25809
rect 24452 25800 24454 25809
rect 24398 25735 24454 25744
rect 24504 25702 24532 26846
rect 24584 26784 24636 26790
rect 24584 26726 24636 26732
rect 24400 25696 24452 25702
rect 24400 25638 24452 25644
rect 24492 25696 24544 25702
rect 24492 25638 24544 25644
rect 24412 24954 24440 25638
rect 24400 24948 24452 24954
rect 24400 24890 24452 24896
rect 24398 24576 24454 24585
rect 24398 24511 24454 24520
rect 24412 24177 24440 24511
rect 24398 24168 24454 24177
rect 24398 24103 24454 24112
rect 24504 24070 24532 25638
rect 24400 24064 24452 24070
rect 24400 24006 24452 24012
rect 24492 24064 24544 24070
rect 24492 24006 24544 24012
rect 24412 23526 24440 24006
rect 24492 23724 24544 23730
rect 24492 23666 24544 23672
rect 24400 23520 24452 23526
rect 24400 23462 24452 23468
rect 24412 22642 24440 23462
rect 24504 22710 24532 23666
rect 24492 22704 24544 22710
rect 24492 22646 24544 22652
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24320 22494 24532 22522
rect 24228 22066 24348 22094
rect 24216 22024 24268 22030
rect 24216 21966 24268 21972
rect 24228 21350 24256 21966
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 24228 20777 24256 21286
rect 24214 20768 24270 20777
rect 24214 20703 24270 20712
rect 24216 20596 24268 20602
rect 24216 20538 24268 20544
rect 24228 20505 24256 20538
rect 24214 20496 24270 20505
rect 24214 20431 24270 20440
rect 24124 20392 24176 20398
rect 24124 20334 24176 20340
rect 24320 20058 24348 22066
rect 24398 21992 24454 22001
rect 24504 21978 24532 22494
rect 24596 22098 24624 26726
rect 24688 25809 24716 26930
rect 24952 26920 25004 26926
rect 24952 26862 25004 26868
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 24872 25974 24900 26318
rect 24860 25968 24912 25974
rect 24860 25910 24912 25916
rect 24964 25906 24992 26862
rect 25056 26042 25084 28018
rect 25412 27532 25464 27538
rect 25412 27474 25464 27480
rect 25320 27464 25372 27470
rect 25320 27406 25372 27412
rect 25136 26852 25188 26858
rect 25136 26794 25188 26800
rect 25044 26036 25096 26042
rect 25044 25978 25096 25984
rect 24768 25900 24820 25906
rect 24768 25842 24820 25848
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 24674 25800 24730 25809
rect 24674 25735 24730 25744
rect 24780 25430 24808 25842
rect 25044 25696 25096 25702
rect 25042 25664 25044 25673
rect 25096 25664 25098 25673
rect 25042 25599 25098 25608
rect 24860 25492 24912 25498
rect 24860 25434 24912 25440
rect 25044 25492 25096 25498
rect 25044 25434 25096 25440
rect 24768 25424 24820 25430
rect 24768 25366 24820 25372
rect 24674 25120 24730 25129
rect 24674 25055 24730 25064
rect 24688 24274 24716 25055
rect 24780 24886 24808 25366
rect 24872 24954 24900 25434
rect 24952 25288 25004 25294
rect 24952 25230 25004 25236
rect 24860 24948 24912 24954
rect 24860 24890 24912 24896
rect 24768 24880 24820 24886
rect 24768 24822 24820 24828
rect 24768 24336 24820 24342
rect 24768 24278 24820 24284
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 24780 24177 24808 24278
rect 24860 24200 24912 24206
rect 24766 24168 24822 24177
rect 24860 24142 24912 24148
rect 24766 24103 24822 24112
rect 24768 24064 24820 24070
rect 24768 24006 24820 24012
rect 24780 23508 24808 24006
rect 24688 23480 24808 23508
rect 24688 22166 24716 23480
rect 24872 23186 24900 24142
rect 24964 24070 24992 25230
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 24952 23792 25004 23798
rect 24952 23734 25004 23740
rect 24964 23633 24992 23734
rect 24950 23624 25006 23633
rect 24950 23559 25006 23568
rect 24860 23180 24912 23186
rect 24860 23122 24912 23128
rect 24952 23180 25004 23186
rect 24952 23122 25004 23128
rect 24872 22574 24900 23122
rect 24964 22953 24992 23122
rect 24950 22944 25006 22953
rect 24950 22879 25006 22888
rect 24860 22568 24912 22574
rect 24860 22510 24912 22516
rect 24676 22160 24728 22166
rect 24676 22102 24728 22108
rect 24584 22092 24636 22098
rect 24584 22034 24636 22040
rect 25056 21978 25084 25434
rect 25148 24138 25176 26794
rect 25228 26784 25280 26790
rect 25332 26772 25360 27406
rect 25280 26744 25360 26772
rect 25228 26726 25280 26732
rect 25332 26586 25360 26744
rect 25424 26586 25452 27474
rect 25608 27130 25636 28426
rect 25596 27124 25648 27130
rect 25596 27066 25648 27072
rect 25504 26920 25556 26926
rect 25504 26862 25556 26868
rect 25320 26580 25372 26586
rect 25320 26522 25372 26528
rect 25412 26580 25464 26586
rect 25412 26522 25464 26528
rect 25320 26376 25372 26382
rect 25318 26344 25320 26353
rect 25372 26344 25374 26353
rect 25318 26279 25374 26288
rect 25412 26036 25464 26042
rect 25412 25978 25464 25984
rect 25318 25664 25374 25673
rect 25318 25599 25374 25608
rect 25332 25294 25360 25599
rect 25424 25537 25452 25978
rect 25410 25528 25466 25537
rect 25516 25498 25544 26862
rect 25608 26790 25636 27066
rect 25596 26784 25648 26790
rect 25596 26726 25648 26732
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 25608 26042 25636 26318
rect 25596 26036 25648 26042
rect 25596 25978 25648 25984
rect 25596 25832 25648 25838
rect 25596 25774 25648 25780
rect 25608 25498 25636 25774
rect 25410 25463 25466 25472
rect 25504 25492 25556 25498
rect 25424 25378 25452 25463
rect 25504 25434 25556 25440
rect 25596 25492 25648 25498
rect 25596 25434 25648 25440
rect 25424 25350 25544 25378
rect 25320 25288 25372 25294
rect 25240 25236 25320 25242
rect 25240 25230 25372 25236
rect 25240 25214 25360 25230
rect 25240 25158 25268 25214
rect 25228 25152 25280 25158
rect 25228 25094 25280 25100
rect 25320 25152 25372 25158
rect 25320 25094 25372 25100
rect 25412 25152 25464 25158
rect 25412 25094 25464 25100
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 25136 24132 25188 24138
rect 25136 24074 25188 24080
rect 25136 23792 25188 23798
rect 25240 23769 25268 24210
rect 25136 23734 25188 23740
rect 25226 23760 25282 23769
rect 25148 23322 25176 23734
rect 25226 23695 25282 23704
rect 25228 23588 25280 23594
rect 25332 23576 25360 25094
rect 25280 23548 25360 23576
rect 25228 23530 25280 23536
rect 25136 23316 25188 23322
rect 25136 23258 25188 23264
rect 25228 23248 25280 23254
rect 25134 23216 25190 23225
rect 25228 23190 25280 23196
rect 25134 23151 25190 23160
rect 25148 22234 25176 23151
rect 25240 22642 25268 23190
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 25240 22234 25268 22578
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 25228 22228 25280 22234
rect 25228 22170 25280 22176
rect 25136 22024 25188 22030
rect 24504 21950 24624 21978
rect 24398 21927 24400 21936
rect 24452 21927 24454 21936
rect 24400 21898 24452 21904
rect 24492 21888 24544 21894
rect 24412 21836 24492 21842
rect 24412 21830 24544 21836
rect 24412 21814 24532 21830
rect 24412 21554 24440 21814
rect 24490 21720 24546 21729
rect 24490 21655 24546 21664
rect 24400 21548 24452 21554
rect 24400 21490 24452 21496
rect 24400 21412 24452 21418
rect 24400 21354 24452 21360
rect 24412 20942 24440 21354
rect 24504 21049 24532 21655
rect 24596 21622 24624 21950
rect 24860 21956 24912 21962
rect 24860 21898 24912 21904
rect 24964 21950 25084 21978
rect 25134 21992 25136 22001
rect 25188 21992 25190 22001
rect 24872 21865 24900 21898
rect 24858 21856 24914 21865
rect 24858 21791 24914 21800
rect 24688 21644 24900 21672
rect 24584 21616 24636 21622
rect 24584 21558 24636 21564
rect 24688 21554 24716 21644
rect 24872 21554 24900 21644
rect 24676 21548 24728 21554
rect 24676 21490 24728 21496
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 24584 21480 24636 21486
rect 24584 21422 24636 21428
rect 24674 21448 24730 21457
rect 24596 21146 24624 21422
rect 24674 21383 24730 21392
rect 24768 21412 24820 21418
rect 24584 21140 24636 21146
rect 24584 21082 24636 21088
rect 24490 21040 24546 21049
rect 24490 20975 24546 20984
rect 24584 21004 24636 21010
rect 24584 20946 24636 20952
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 24490 20768 24546 20777
rect 24490 20703 24546 20712
rect 24308 20052 24360 20058
rect 24308 19994 24360 20000
rect 24124 19916 24176 19922
rect 24124 19858 24176 19864
rect 24032 19304 24084 19310
rect 24032 19246 24084 19252
rect 24032 18760 24084 18766
rect 24032 18702 24084 18708
rect 24044 18426 24072 18702
rect 24032 18420 24084 18426
rect 24032 18362 24084 18368
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 24044 17921 24072 18226
rect 24030 17912 24086 17921
rect 24030 17847 24032 17856
rect 24084 17847 24086 17856
rect 24032 17818 24084 17824
rect 24032 17060 24084 17066
rect 24032 17002 24084 17008
rect 24044 16833 24072 17002
rect 24030 16824 24086 16833
rect 24030 16759 24086 16768
rect 24136 16522 24164 19858
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 24308 17128 24360 17134
rect 24308 17070 24360 17076
rect 24320 16794 24348 17070
rect 24308 16788 24360 16794
rect 24308 16730 24360 16736
rect 24320 16658 24348 16730
rect 24308 16652 24360 16658
rect 24308 16594 24360 16600
rect 24124 16516 24176 16522
rect 24124 16458 24176 16464
rect 23952 15966 24072 15994
rect 23848 15700 23900 15706
rect 23848 15642 23900 15648
rect 23756 15360 23808 15366
rect 23756 15302 23808 15308
rect 23860 15162 23888 15642
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 23848 15156 23900 15162
rect 23848 15098 23900 15104
rect 23020 15020 23072 15026
rect 23020 14962 23072 14968
rect 23572 15020 23624 15026
rect 23572 14962 23624 14968
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23584 14906 23612 14962
rect 23768 14958 23796 15098
rect 23756 14952 23808 14958
rect 23584 14878 23704 14906
rect 23756 14894 23808 14900
rect 23676 14822 23704 14878
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 23664 14816 23716 14822
rect 23664 14758 23716 14764
rect 23584 14618 23612 14758
rect 22928 14612 22980 14618
rect 22928 14554 22980 14560
rect 23572 14612 23624 14618
rect 23572 14554 23624 14560
rect 23020 14408 23072 14414
rect 23020 14350 23072 14356
rect 22192 13942 22244 13948
rect 22480 13938 22600 13954
rect 22836 14000 22888 14006
rect 22836 13942 22888 13948
rect 22468 13932 22600 13938
rect 22520 13926 22600 13932
rect 22468 13874 22520 13880
rect 21732 13864 21784 13870
rect 21732 13806 21784 13812
rect 22284 13796 22336 13802
rect 22284 13738 22336 13744
rect 22296 13569 22324 13738
rect 22282 13560 22338 13569
rect 22480 13530 22508 13874
rect 22282 13495 22284 13504
rect 22336 13495 22338 13504
rect 22468 13524 22520 13530
rect 22284 13466 22336 13472
rect 22468 13466 22520 13472
rect 22100 13456 22152 13462
rect 22100 13398 22152 13404
rect 22112 13190 22140 13398
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 23032 12986 23060 14350
rect 23110 14104 23166 14113
rect 23110 14039 23112 14048
rect 23164 14039 23166 14048
rect 23112 14010 23164 14016
rect 23202 13288 23258 13297
rect 23202 13223 23258 13232
rect 23480 13252 23532 13258
rect 23216 12986 23244 13223
rect 23480 13194 23532 13200
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 20720 12912 20772 12918
rect 20720 12854 20772 12860
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19800 12368 19852 12374
rect 19800 12310 19852 12316
rect 17684 12232 17736 12238
rect 17604 12192 17684 12220
rect 17500 12174 17552 12180
rect 17684 12174 17736 12180
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 19524 12232 19576 12238
rect 19524 12174 19576 12180
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19904 12170 19932 12786
rect 20732 12646 20760 12854
rect 23216 12850 23244 12922
rect 23492 12850 23520 13194
rect 23768 12986 23796 14894
rect 24044 14482 24072 15966
rect 24136 15910 24164 16458
rect 24124 15904 24176 15910
rect 24124 15846 24176 15852
rect 24216 15360 24268 15366
rect 24216 15302 24268 15308
rect 24124 14816 24176 14822
rect 24124 14758 24176 14764
rect 24136 14482 24164 14758
rect 24228 14521 24256 15302
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24320 14618 24348 14962
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 24214 14512 24270 14521
rect 24032 14476 24084 14482
rect 24032 14418 24084 14424
rect 24124 14476 24176 14482
rect 24214 14447 24270 14456
rect 24124 14418 24176 14424
rect 23846 13696 23902 13705
rect 23846 13631 23902 13640
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 23860 12850 23888 13631
rect 24412 13569 24440 17274
rect 24398 13560 24454 13569
rect 24398 13495 24454 13504
rect 23938 13016 23994 13025
rect 23938 12951 23994 12960
rect 23952 12850 23980 12951
rect 24412 12889 24440 13495
rect 24504 12986 24532 20703
rect 24596 19922 24624 20946
rect 24584 19916 24636 19922
rect 24584 19858 24636 19864
rect 24584 19780 24636 19786
rect 24584 19722 24636 19728
rect 24596 19514 24624 19722
rect 24584 19508 24636 19514
rect 24584 19450 24636 19456
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24596 16998 24624 17478
rect 24584 16992 24636 16998
rect 24584 16934 24636 16940
rect 24688 14414 24716 21383
rect 24768 21354 24820 21360
rect 24860 21412 24912 21418
rect 24860 21354 24912 21360
rect 24780 17338 24808 21354
rect 24872 21146 24900 21354
rect 24860 21140 24912 21146
rect 24860 21082 24912 21088
rect 24858 21040 24914 21049
rect 24858 20975 24914 20984
rect 24872 20942 24900 20975
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24860 20596 24912 20602
rect 24860 20538 24912 20544
rect 24872 20330 24900 20538
rect 24860 20324 24912 20330
rect 24860 20266 24912 20272
rect 24964 20210 24992 21950
rect 25134 21927 25190 21936
rect 25228 21956 25280 21962
rect 25228 21898 25280 21904
rect 25044 21888 25096 21894
rect 25044 21830 25096 21836
rect 25056 20330 25084 21830
rect 25134 21176 25190 21185
rect 25134 21111 25190 21120
rect 25148 20806 25176 21111
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 25044 20324 25096 20330
rect 25044 20266 25096 20272
rect 24964 20182 25084 20210
rect 24858 19272 24914 19281
rect 24858 19207 24914 19216
rect 24872 18834 24900 19207
rect 24860 18828 24912 18834
rect 24860 18770 24912 18776
rect 24860 18420 24912 18426
rect 24860 18362 24912 18368
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 24872 17218 24900 18362
rect 24952 17808 25004 17814
rect 24952 17750 25004 17756
rect 24780 17202 24900 17218
rect 24768 17196 24900 17202
rect 24820 17190 24900 17196
rect 24768 17138 24820 17144
rect 24860 17128 24912 17134
rect 24780 17076 24860 17082
rect 24780 17070 24912 17076
rect 24780 17054 24900 17070
rect 24780 16969 24808 17054
rect 24766 16960 24822 16969
rect 24766 16895 24822 16904
rect 24964 16522 24992 17750
rect 25056 17082 25084 20182
rect 25148 19174 25176 20334
rect 25136 19168 25188 19174
rect 25136 19110 25188 19116
rect 25240 17678 25268 21898
rect 25332 21010 25360 23548
rect 25320 21004 25372 21010
rect 25320 20946 25372 20952
rect 25320 20868 25372 20874
rect 25320 20810 25372 20816
rect 25228 17672 25280 17678
rect 25228 17614 25280 17620
rect 25332 17134 25360 20810
rect 25424 19990 25452 25094
rect 25516 20346 25544 25350
rect 25596 24336 25648 24342
rect 25594 24304 25596 24313
rect 25648 24304 25650 24313
rect 25594 24239 25650 24248
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25608 22438 25636 23666
rect 25596 22432 25648 22438
rect 25596 22374 25648 22380
rect 25700 22094 25728 32234
rect 26056 32224 26108 32230
rect 26056 32166 26108 32172
rect 26068 32026 26096 32166
rect 26056 32020 26108 32026
rect 26056 31962 26108 31968
rect 26160 31754 26188 32710
rect 26240 32360 26292 32366
rect 26240 32302 26292 32308
rect 26148 31748 26200 31754
rect 26148 31690 26200 31696
rect 25778 31648 25834 31657
rect 25778 31583 25834 31592
rect 25792 27614 25820 31583
rect 25964 31272 26016 31278
rect 25964 31214 26016 31220
rect 26148 31272 26200 31278
rect 26148 31214 26200 31220
rect 25872 31136 25924 31142
rect 25872 31078 25924 31084
rect 25884 30054 25912 31078
rect 25976 30870 26004 31214
rect 26056 31136 26108 31142
rect 26056 31078 26108 31084
rect 25964 30864 26016 30870
rect 25964 30806 26016 30812
rect 26068 30666 26096 31078
rect 26160 30938 26188 31214
rect 26252 31142 26280 32302
rect 26422 32192 26478 32201
rect 26422 32127 26478 32136
rect 26436 31890 26464 32127
rect 26528 32026 26556 33390
rect 26608 32428 26660 32434
rect 26608 32370 26660 32376
rect 26620 32026 26648 32370
rect 26516 32020 26568 32026
rect 26516 31962 26568 31968
rect 26608 32020 26660 32026
rect 26608 31962 26660 31968
rect 26424 31884 26476 31890
rect 26424 31826 26476 31832
rect 26620 31278 26648 31962
rect 26988 31822 27016 34954
rect 27080 34202 27108 37130
rect 28184 34746 28212 37130
rect 28172 34740 28224 34746
rect 28172 34682 28224 34688
rect 27528 34672 27580 34678
rect 27528 34614 27580 34620
rect 27068 34196 27120 34202
rect 27068 34138 27120 34144
rect 27080 33522 27108 34138
rect 27540 33998 27568 34614
rect 27712 34604 27764 34610
rect 27712 34546 27764 34552
rect 27528 33992 27580 33998
rect 27528 33934 27580 33940
rect 27068 33516 27120 33522
rect 27068 33458 27120 33464
rect 27436 33380 27488 33386
rect 27436 33322 27488 33328
rect 27252 32360 27304 32366
rect 27252 32302 27304 32308
rect 26976 31816 27028 31822
rect 26976 31758 27028 31764
rect 26608 31272 26660 31278
rect 26608 31214 26660 31220
rect 26700 31272 26752 31278
rect 26700 31214 26752 31220
rect 26332 31204 26384 31210
rect 26332 31146 26384 31152
rect 26240 31136 26292 31142
rect 26240 31078 26292 31084
rect 26148 30932 26200 30938
rect 26148 30874 26200 30880
rect 26056 30660 26108 30666
rect 26056 30602 26108 30608
rect 25964 30388 26016 30394
rect 25964 30330 26016 30336
rect 25872 30048 25924 30054
rect 25872 29990 25924 29996
rect 25976 29753 26004 30330
rect 26160 29850 26188 30874
rect 26344 30598 26372 31146
rect 26712 30841 26740 31214
rect 26698 30832 26754 30841
rect 26608 30796 26660 30802
rect 26698 30767 26754 30776
rect 26608 30738 26660 30744
rect 26332 30592 26384 30598
rect 26332 30534 26384 30540
rect 26240 30048 26292 30054
rect 26240 29990 26292 29996
rect 26148 29844 26200 29850
rect 26148 29786 26200 29792
rect 25962 29744 26018 29753
rect 25962 29679 26018 29688
rect 26252 29646 26280 29990
rect 26240 29640 26292 29646
rect 26240 29582 26292 29588
rect 25872 29504 25924 29510
rect 25872 29446 25924 29452
rect 25884 29238 25912 29446
rect 25872 29232 25924 29238
rect 25872 29174 25924 29180
rect 26148 28620 26200 28626
rect 26148 28562 26200 28568
rect 26160 28490 26188 28562
rect 26148 28484 26200 28490
rect 26148 28426 26200 28432
rect 26252 27962 26280 29582
rect 26516 29572 26568 29578
rect 26516 29514 26568 29520
rect 26332 28960 26384 28966
rect 26332 28902 26384 28908
rect 26344 28801 26372 28902
rect 26330 28792 26386 28801
rect 26330 28727 26386 28736
rect 26252 27934 26464 27962
rect 26240 27872 26292 27878
rect 26332 27872 26384 27878
rect 26240 27814 26292 27820
rect 26330 27840 26332 27849
rect 26384 27840 26386 27849
rect 25792 27586 25912 27614
rect 25780 26784 25832 26790
rect 25780 26726 25832 26732
rect 25792 26353 25820 26726
rect 25778 26344 25834 26353
rect 25778 26279 25834 26288
rect 25780 25288 25832 25294
rect 25780 25230 25832 25236
rect 25792 24750 25820 25230
rect 25884 24993 25912 27586
rect 26252 27538 26280 27814
rect 26330 27775 26386 27784
rect 26240 27532 26292 27538
rect 26240 27474 26292 27480
rect 26436 27402 26464 27934
rect 26240 27396 26292 27402
rect 26240 27338 26292 27344
rect 26424 27396 26476 27402
rect 26424 27338 26476 27344
rect 26056 27124 26108 27130
rect 26056 27066 26108 27072
rect 25964 27056 26016 27062
rect 25964 26998 26016 27004
rect 25976 26450 26004 26998
rect 25964 26444 26016 26450
rect 25964 26386 26016 26392
rect 25870 24984 25926 24993
rect 25870 24919 25926 24928
rect 25780 24744 25832 24750
rect 25780 24686 25832 24692
rect 25792 24313 25820 24686
rect 25778 24304 25834 24313
rect 25778 24239 25834 24248
rect 25976 24188 26004 26386
rect 26068 25838 26096 27066
rect 26252 26790 26280 27338
rect 26424 26988 26476 26994
rect 26344 26948 26424 26976
rect 26240 26784 26292 26790
rect 26240 26726 26292 26732
rect 26238 26344 26294 26353
rect 26238 26279 26294 26288
rect 26252 25906 26280 26279
rect 26240 25900 26292 25906
rect 26240 25842 26292 25848
rect 26056 25832 26108 25838
rect 26056 25774 26108 25780
rect 26068 25158 26096 25774
rect 26148 25220 26200 25226
rect 26148 25162 26200 25168
rect 26056 25152 26108 25158
rect 26056 25094 26108 25100
rect 26054 24848 26110 24857
rect 26160 24834 26188 25162
rect 26240 25152 26292 25158
rect 26238 25120 26240 25129
rect 26292 25120 26294 25129
rect 26238 25055 26294 25064
rect 26344 24886 26372 26948
rect 26424 26930 26476 26936
rect 26424 26512 26476 26518
rect 26424 26454 26476 26460
rect 26332 24880 26384 24886
rect 26160 24806 26280 24834
rect 26436 24857 26464 26454
rect 26528 25362 26556 29514
rect 26620 28082 26648 30738
rect 26976 30660 27028 30666
rect 26976 30602 27028 30608
rect 27068 30660 27120 30666
rect 27068 30602 27120 30608
rect 26790 30288 26846 30297
rect 26790 30223 26846 30232
rect 26700 29640 26752 29646
rect 26700 29582 26752 29588
rect 26712 29481 26740 29582
rect 26698 29472 26754 29481
rect 26698 29407 26754 29416
rect 26804 29170 26832 30223
rect 26884 29844 26936 29850
rect 26884 29786 26936 29792
rect 26792 29164 26844 29170
rect 26792 29106 26844 29112
rect 26700 28960 26752 28966
rect 26700 28902 26752 28908
rect 26792 28960 26844 28966
rect 26792 28902 26844 28908
rect 26712 28558 26740 28902
rect 26700 28552 26752 28558
rect 26700 28494 26752 28500
rect 26608 28076 26660 28082
rect 26608 28018 26660 28024
rect 26712 28014 26740 28494
rect 26804 28422 26832 28902
rect 26792 28416 26844 28422
rect 26792 28358 26844 28364
rect 26792 28212 26844 28218
rect 26792 28154 26844 28160
rect 26700 28008 26752 28014
rect 26700 27950 26752 27956
rect 26608 27872 26660 27878
rect 26608 27814 26660 27820
rect 26620 27674 26648 27814
rect 26608 27668 26660 27674
rect 26608 27610 26660 27616
rect 26700 27668 26752 27674
rect 26700 27610 26752 27616
rect 26606 27432 26662 27441
rect 26606 27367 26662 27376
rect 26620 26858 26648 27367
rect 26712 27130 26740 27610
rect 26804 27606 26832 28154
rect 26896 27674 26924 29786
rect 26884 27668 26936 27674
rect 26884 27610 26936 27616
rect 26792 27600 26844 27606
rect 26792 27542 26844 27548
rect 26792 27464 26844 27470
rect 26792 27406 26844 27412
rect 26882 27432 26938 27441
rect 26700 27124 26752 27130
rect 26700 27066 26752 27072
rect 26608 26852 26660 26858
rect 26608 26794 26660 26800
rect 26606 26616 26662 26625
rect 26606 26551 26608 26560
rect 26660 26551 26662 26560
rect 26608 26522 26660 26528
rect 26804 26382 26832 27406
rect 26882 27367 26938 27376
rect 26896 27169 26924 27367
rect 26882 27160 26938 27169
rect 26882 27095 26938 27104
rect 26792 26376 26844 26382
rect 26844 26336 26924 26364
rect 26792 26318 26844 26324
rect 26608 25900 26660 25906
rect 26608 25842 26660 25848
rect 26792 25900 26844 25906
rect 26792 25842 26844 25848
rect 26516 25356 26568 25362
rect 26516 25298 26568 25304
rect 26516 24948 26568 24954
rect 26516 24890 26568 24896
rect 26332 24822 26384 24828
rect 26422 24848 26478 24857
rect 26054 24783 26110 24792
rect 26068 24682 26096 24783
rect 26056 24676 26108 24682
rect 26056 24618 26108 24624
rect 25608 22066 25728 22094
rect 25792 24160 26004 24188
rect 25608 20466 25636 22066
rect 25686 21992 25742 22001
rect 25686 21927 25742 21936
rect 25700 21894 25728 21927
rect 25688 21888 25740 21894
rect 25688 21830 25740 21836
rect 25792 20874 25820 24160
rect 26056 24132 26108 24138
rect 26056 24074 26108 24080
rect 26068 24018 26096 24074
rect 25976 23990 26096 24018
rect 25870 23760 25926 23769
rect 25870 23695 25872 23704
rect 25924 23695 25926 23704
rect 25872 23666 25924 23672
rect 25870 23488 25926 23497
rect 25870 23423 25926 23432
rect 25780 20868 25832 20874
rect 25780 20810 25832 20816
rect 25596 20460 25648 20466
rect 25596 20402 25648 20408
rect 25516 20318 25820 20346
rect 25504 20052 25556 20058
rect 25504 19994 25556 20000
rect 25596 20052 25648 20058
rect 25596 19994 25648 20000
rect 25412 19984 25464 19990
rect 25412 19926 25464 19932
rect 25410 18728 25466 18737
rect 25410 18663 25466 18672
rect 25424 18465 25452 18663
rect 25410 18456 25466 18465
rect 25410 18391 25466 18400
rect 25424 18290 25452 18391
rect 25412 18284 25464 18290
rect 25412 18226 25464 18232
rect 25412 18080 25464 18086
rect 25410 18048 25412 18057
rect 25464 18048 25466 18057
rect 25410 17983 25466 17992
rect 25320 17128 25372 17134
rect 25056 17054 25176 17082
rect 25320 17070 25372 17076
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 25056 16658 25084 16934
rect 25148 16726 25176 17054
rect 25136 16720 25188 16726
rect 25136 16662 25188 16668
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 25136 16584 25188 16590
rect 25136 16526 25188 16532
rect 24952 16516 25004 16522
rect 24952 16458 25004 16464
rect 24964 16182 24992 16458
rect 25148 16250 25176 16526
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 24952 16176 25004 16182
rect 24952 16118 25004 16124
rect 25228 15972 25280 15978
rect 25228 15914 25280 15920
rect 25240 15366 25268 15914
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25240 14958 25268 15302
rect 25228 14952 25280 14958
rect 25228 14894 25280 14900
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 25332 13870 25360 17070
rect 25516 16794 25544 19994
rect 25608 19854 25636 19994
rect 25686 19952 25742 19961
rect 25686 19887 25688 19896
rect 25740 19887 25742 19896
rect 25688 19858 25740 19864
rect 25792 19854 25820 20318
rect 25884 20058 25912 23423
rect 25976 23254 26004 23990
rect 26148 23792 26200 23798
rect 26068 23752 26148 23780
rect 25964 23248 26016 23254
rect 25964 23190 26016 23196
rect 25976 22098 26004 23190
rect 26068 23050 26096 23752
rect 26148 23734 26200 23740
rect 26252 23497 26280 24806
rect 26422 24783 26478 24792
rect 26332 24744 26384 24750
rect 26332 24686 26384 24692
rect 26344 24313 26372 24686
rect 26528 24614 26556 24890
rect 26620 24857 26648 25842
rect 26698 25120 26754 25129
rect 26698 25055 26754 25064
rect 26606 24848 26662 24857
rect 26606 24783 26662 24792
rect 26516 24608 26568 24614
rect 26516 24550 26568 24556
rect 26330 24304 26386 24313
rect 26330 24239 26386 24248
rect 26344 24070 26372 24239
rect 26424 24132 26476 24138
rect 26424 24074 26476 24080
rect 26332 24064 26384 24070
rect 26332 24006 26384 24012
rect 26436 23746 26464 24074
rect 26712 23905 26740 25055
rect 26804 24993 26832 25842
rect 26790 24984 26846 24993
rect 26790 24919 26846 24928
rect 26792 24744 26844 24750
rect 26792 24686 26844 24692
rect 26698 23896 26754 23905
rect 26698 23831 26754 23840
rect 26344 23718 26464 23746
rect 26514 23760 26570 23769
rect 26238 23488 26294 23497
rect 26238 23423 26294 23432
rect 26056 23044 26108 23050
rect 26056 22986 26108 22992
rect 26148 23044 26200 23050
rect 26148 22986 26200 22992
rect 26160 22642 26188 22986
rect 26148 22636 26200 22642
rect 26148 22578 26200 22584
rect 26240 22636 26292 22642
rect 26240 22578 26292 22584
rect 26056 22568 26108 22574
rect 26056 22510 26108 22516
rect 26146 22536 26202 22545
rect 26068 22234 26096 22510
rect 26146 22471 26202 22480
rect 26056 22228 26108 22234
rect 26056 22170 26108 22176
rect 26160 22098 26188 22471
rect 26252 22409 26280 22578
rect 26344 22574 26372 23718
rect 26514 23695 26570 23704
rect 26700 23724 26752 23730
rect 26424 23656 26476 23662
rect 26424 23598 26476 23604
rect 26436 22658 26464 23598
rect 26528 23594 26556 23695
rect 26700 23666 26752 23672
rect 26608 23656 26660 23662
rect 26608 23598 26660 23604
rect 26516 23588 26568 23594
rect 26516 23530 26568 23536
rect 26516 23316 26568 23322
rect 26516 23258 26568 23264
rect 26528 23050 26556 23258
rect 26620 23254 26648 23598
rect 26608 23248 26660 23254
rect 26608 23190 26660 23196
rect 26712 23100 26740 23666
rect 26804 23254 26832 24686
rect 26896 24138 26924 26336
rect 26988 25158 27016 30602
rect 27080 30569 27108 30602
rect 27066 30560 27122 30569
rect 27066 30495 27122 30504
rect 27158 28792 27214 28801
rect 27158 28727 27214 28736
rect 27068 28144 27120 28150
rect 27068 28086 27120 28092
rect 27080 27878 27108 28086
rect 27172 27985 27200 28727
rect 27264 28558 27292 32302
rect 27344 30932 27396 30938
rect 27344 30874 27396 30880
rect 27252 28552 27304 28558
rect 27252 28494 27304 28500
rect 27252 28076 27304 28082
rect 27252 28018 27304 28024
rect 27158 27976 27214 27985
rect 27158 27911 27214 27920
rect 27068 27872 27120 27878
rect 27068 27814 27120 27820
rect 27160 27872 27212 27878
rect 27160 27814 27212 27820
rect 27068 27056 27120 27062
rect 27068 26998 27120 27004
rect 26976 25152 27028 25158
rect 26976 25094 27028 25100
rect 26976 24676 27028 24682
rect 26976 24618 27028 24624
rect 26884 24132 26936 24138
rect 26884 24074 26936 24080
rect 26988 23866 27016 24618
rect 26976 23860 27028 23866
rect 26976 23802 27028 23808
rect 26882 23760 26938 23769
rect 26882 23695 26938 23704
rect 26976 23724 27028 23730
rect 26896 23662 26924 23695
rect 26976 23666 27028 23672
rect 26884 23656 26936 23662
rect 26884 23598 26936 23604
rect 26884 23316 26936 23322
rect 26884 23258 26936 23264
rect 26792 23248 26844 23254
rect 26792 23190 26844 23196
rect 26896 23118 26924 23258
rect 26884 23112 26936 23118
rect 26712 23072 26832 23100
rect 26516 23044 26568 23050
rect 26516 22986 26568 22992
rect 26436 22642 26556 22658
rect 26436 22636 26568 22642
rect 26436 22630 26516 22636
rect 26516 22578 26568 22584
rect 26332 22568 26384 22574
rect 26332 22510 26384 22516
rect 26804 22488 26832 23072
rect 26988 23100 27016 23666
rect 27080 23322 27108 26998
rect 27172 24682 27200 27814
rect 27264 26790 27292 28018
rect 27252 26784 27304 26790
rect 27252 26726 27304 26732
rect 27264 26625 27292 26726
rect 27250 26616 27306 26625
rect 27250 26551 27306 26560
rect 27160 24676 27212 24682
rect 27160 24618 27212 24624
rect 27252 24608 27304 24614
rect 27252 24550 27304 24556
rect 27160 24132 27212 24138
rect 27160 24074 27212 24080
rect 27172 23526 27200 24074
rect 27160 23520 27212 23526
rect 27160 23462 27212 23468
rect 27068 23316 27120 23322
rect 27068 23258 27120 23264
rect 27160 23112 27212 23118
rect 26988 23072 27160 23100
rect 26884 23054 26936 23060
rect 27160 23054 27212 23060
rect 26884 22976 26936 22982
rect 26884 22918 26936 22924
rect 26896 22642 26924 22918
rect 27066 22808 27122 22817
rect 27066 22743 27122 22752
rect 26884 22636 26936 22642
rect 26884 22578 26936 22584
rect 26528 22460 26832 22488
rect 26882 22536 26938 22545
rect 26882 22471 26938 22480
rect 26332 22432 26384 22438
rect 26238 22400 26294 22409
rect 26384 22392 26464 22420
rect 26332 22374 26384 22380
rect 26238 22335 26294 22344
rect 26436 22166 26464 22392
rect 26332 22160 26384 22166
rect 26332 22102 26384 22108
rect 26424 22160 26476 22166
rect 26424 22102 26476 22108
rect 25964 22092 26016 22098
rect 25964 22034 26016 22040
rect 26148 22092 26200 22098
rect 26148 22034 26200 22040
rect 25964 21956 26016 21962
rect 25964 21898 26016 21904
rect 25976 21593 26004 21898
rect 25962 21584 26018 21593
rect 25962 21519 26018 21528
rect 26146 21584 26202 21593
rect 26146 21519 26202 21528
rect 25964 21480 26016 21486
rect 25964 21422 26016 21428
rect 25976 20262 26004 21422
rect 26160 21321 26188 21519
rect 26146 21312 26202 21321
rect 26146 21247 26202 21256
rect 26344 20942 26372 22102
rect 26422 21176 26478 21185
rect 26422 21111 26478 21120
rect 26332 20936 26384 20942
rect 26332 20878 26384 20884
rect 26054 20632 26110 20641
rect 26054 20567 26110 20576
rect 26068 20466 26096 20567
rect 26056 20460 26108 20466
rect 26056 20402 26108 20408
rect 26332 20460 26384 20466
rect 26332 20402 26384 20408
rect 26148 20392 26200 20398
rect 26148 20334 26200 20340
rect 25964 20256 26016 20262
rect 25964 20198 26016 20204
rect 26056 20256 26108 20262
rect 26056 20198 26108 20204
rect 25872 20052 25924 20058
rect 25872 19994 25924 20000
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25608 18426 25636 19790
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25596 18420 25648 18426
rect 25596 18362 25648 18368
rect 25700 18170 25728 19110
rect 25608 18142 25728 18170
rect 25504 16788 25556 16794
rect 25504 16730 25556 16736
rect 25412 16652 25464 16658
rect 25412 16594 25464 16600
rect 25424 14793 25452 16594
rect 25516 16114 25544 16730
rect 25608 16114 25636 18142
rect 25688 18080 25740 18086
rect 25688 18022 25740 18028
rect 25700 17678 25728 18022
rect 25688 17672 25740 17678
rect 25688 17614 25740 17620
rect 25792 16590 25820 19790
rect 25964 19372 26016 19378
rect 25964 19314 26016 19320
rect 25976 17882 26004 19314
rect 25964 17876 26016 17882
rect 25964 17818 26016 17824
rect 25872 16720 25924 16726
rect 25872 16662 25924 16668
rect 25780 16584 25832 16590
rect 25780 16526 25832 16532
rect 25504 16108 25556 16114
rect 25504 16050 25556 16056
rect 25596 16108 25648 16114
rect 25596 16050 25648 16056
rect 25410 14784 25466 14793
rect 25410 14719 25466 14728
rect 25320 13864 25372 13870
rect 25320 13806 25372 13812
rect 24492 12980 24544 12986
rect 24492 12922 24544 12928
rect 24398 12880 24454 12889
rect 23204 12844 23256 12850
rect 23204 12786 23256 12792
rect 23480 12844 23532 12850
rect 23480 12786 23532 12792
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 23940 12844 23992 12850
rect 25424 12850 25452 14719
rect 24398 12815 24454 12824
rect 25412 12844 25464 12850
rect 23940 12786 23992 12792
rect 20720 12640 20772 12646
rect 23204 12640 23256 12646
rect 20720 12582 20772 12588
rect 23202 12608 23204 12617
rect 23256 12608 23258 12617
rect 23202 12543 23258 12552
rect 17408 12164 17460 12170
rect 17408 12106 17460 12112
rect 19892 12164 19944 12170
rect 19892 12106 19944 12112
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 15856 11694 15884 11834
rect 17420 11762 17448 12106
rect 23860 11898 23888 12786
rect 24412 12646 24440 12815
rect 25412 12786 25464 12792
rect 25516 12714 25544 16050
rect 25596 15700 25648 15706
rect 25596 15642 25648 15648
rect 25608 15473 25636 15642
rect 25594 15464 25650 15473
rect 25594 15399 25650 15408
rect 25688 15360 25740 15366
rect 25688 15302 25740 15308
rect 25596 14544 25648 14550
rect 25596 14486 25648 14492
rect 25608 13938 25636 14486
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25700 13734 25728 15302
rect 25688 13728 25740 13734
rect 25688 13670 25740 13676
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 25504 12708 25556 12714
rect 25504 12650 25556 12656
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 25700 12481 25728 12786
rect 25792 12782 25820 16526
rect 25884 15978 25912 16662
rect 25964 16516 26016 16522
rect 25964 16458 26016 16464
rect 25872 15972 25924 15978
rect 25872 15914 25924 15920
rect 25872 13932 25924 13938
rect 25976 13920 26004 16458
rect 25924 13892 26004 13920
rect 25872 13874 25924 13880
rect 25884 13258 25912 13874
rect 26068 13530 26096 20198
rect 26160 18290 26188 20334
rect 26344 20058 26372 20402
rect 26436 20398 26464 21111
rect 26528 20874 26556 22460
rect 26790 22400 26846 22409
rect 26790 22335 26846 22344
rect 26804 22234 26832 22335
rect 26792 22228 26844 22234
rect 26792 22170 26844 22176
rect 26608 22160 26660 22166
rect 26608 22102 26660 22108
rect 26516 20868 26568 20874
rect 26516 20810 26568 20816
rect 26528 20602 26556 20810
rect 26620 20602 26648 22102
rect 26792 22024 26844 22030
rect 26792 21966 26844 21972
rect 26804 20777 26832 21966
rect 26790 20768 26846 20777
rect 26790 20703 26846 20712
rect 26516 20596 26568 20602
rect 26516 20538 26568 20544
rect 26608 20596 26660 20602
rect 26608 20538 26660 20544
rect 26424 20392 26476 20398
rect 26424 20334 26476 20340
rect 26528 20058 26556 20538
rect 26792 20460 26844 20466
rect 26792 20402 26844 20408
rect 26332 20052 26384 20058
rect 26332 19994 26384 20000
rect 26516 20052 26568 20058
rect 26516 19994 26568 20000
rect 26424 19916 26476 19922
rect 26424 19858 26476 19864
rect 26332 19712 26384 19718
rect 26332 19654 26384 19660
rect 26240 19304 26292 19310
rect 26240 19246 26292 19252
rect 26252 18358 26280 19246
rect 26240 18352 26292 18358
rect 26240 18294 26292 18300
rect 26148 18284 26200 18290
rect 26148 18226 26200 18232
rect 26146 17912 26202 17921
rect 26146 17847 26202 17856
rect 26240 17876 26292 17882
rect 26160 17746 26188 17847
rect 26240 17818 26292 17824
rect 26148 17740 26200 17746
rect 26148 17682 26200 17688
rect 26252 17270 26280 17818
rect 26344 17678 26372 19654
rect 26332 17672 26384 17678
rect 26332 17614 26384 17620
rect 26436 17542 26464 19858
rect 26804 19854 26832 20402
rect 26792 19848 26844 19854
rect 26792 19790 26844 19796
rect 26516 19712 26568 19718
rect 26514 19680 26516 19689
rect 26896 19700 26924 22471
rect 26976 21888 27028 21894
rect 26976 21830 27028 21836
rect 26988 21554 27016 21830
rect 26976 21548 27028 21554
rect 26976 21490 27028 21496
rect 27080 21418 27108 22743
rect 27172 22098 27200 23054
rect 27264 22234 27292 24550
rect 27356 22710 27384 30874
rect 27448 30818 27476 33322
rect 27540 31686 27568 33934
rect 27724 33658 27752 34546
rect 28448 34400 28500 34406
rect 28448 34342 28500 34348
rect 27804 33924 27856 33930
rect 27804 33866 27856 33872
rect 27712 33652 27764 33658
rect 27712 33594 27764 33600
rect 27816 33114 27844 33866
rect 27896 33516 27948 33522
rect 27896 33458 27948 33464
rect 27988 33516 28040 33522
rect 27988 33458 28040 33464
rect 28264 33516 28316 33522
rect 28264 33458 28316 33464
rect 27804 33108 27856 33114
rect 27804 33050 27856 33056
rect 27908 32910 27936 33458
rect 27804 32904 27856 32910
rect 27804 32846 27856 32852
rect 27896 32904 27948 32910
rect 27896 32846 27948 32852
rect 27620 32836 27672 32842
rect 27620 32778 27672 32784
rect 27632 31754 27660 32778
rect 27816 32230 27844 32846
rect 27908 32774 27936 32846
rect 27896 32768 27948 32774
rect 27896 32710 27948 32716
rect 27804 32224 27856 32230
rect 27804 32166 27856 32172
rect 27632 31726 27844 31754
rect 27528 31680 27580 31686
rect 27528 31622 27580 31628
rect 27448 30790 27568 30818
rect 27436 30728 27488 30734
rect 27436 30670 27488 30676
rect 27448 29850 27476 30670
rect 27436 29844 27488 29850
rect 27436 29786 27488 29792
rect 27436 28756 27488 28762
rect 27436 28698 27488 28704
rect 27448 28218 27476 28698
rect 27540 28218 27568 30790
rect 27712 30184 27764 30190
rect 27712 30126 27764 30132
rect 27724 29714 27752 30126
rect 27712 29708 27764 29714
rect 27712 29650 27764 29656
rect 27712 28416 27764 28422
rect 27712 28358 27764 28364
rect 27436 28212 27488 28218
rect 27436 28154 27488 28160
rect 27528 28212 27580 28218
rect 27528 28154 27580 28160
rect 27724 28082 27752 28358
rect 27712 28076 27764 28082
rect 27712 28018 27764 28024
rect 27436 27940 27488 27946
rect 27436 27882 27488 27888
rect 27448 27130 27476 27882
rect 27618 27704 27674 27713
rect 27618 27639 27674 27648
rect 27528 27532 27580 27538
rect 27528 27474 27580 27480
rect 27436 27124 27488 27130
rect 27436 27066 27488 27072
rect 27540 26858 27568 27474
rect 27632 27062 27660 27639
rect 27816 27606 27844 31726
rect 27894 31648 27950 31657
rect 27894 31583 27950 31592
rect 27908 31113 27936 31583
rect 27894 31104 27950 31113
rect 27894 31039 27950 31048
rect 28000 30938 28028 33458
rect 28276 33046 28304 33458
rect 28460 33454 28488 34342
rect 29656 34066 29684 37130
rect 29644 34060 29696 34066
rect 29644 34002 29696 34008
rect 29000 33856 29052 33862
rect 29000 33798 29052 33804
rect 28448 33448 28500 33454
rect 28448 33390 28500 33396
rect 29012 33114 29040 33798
rect 30484 33658 30512 37130
rect 30472 33652 30524 33658
rect 30472 33594 30524 33600
rect 30484 33522 30512 33594
rect 29552 33516 29604 33522
rect 29552 33458 29604 33464
rect 30472 33516 30524 33522
rect 30472 33458 30524 33464
rect 29564 33114 29592 33458
rect 30656 33448 30708 33454
rect 30656 33390 30708 33396
rect 30196 33312 30248 33318
rect 30196 33254 30248 33260
rect 29000 33108 29052 33114
rect 29000 33050 29052 33056
rect 29552 33108 29604 33114
rect 29552 33050 29604 33056
rect 28264 33040 28316 33046
rect 28264 32982 28316 32988
rect 28276 32910 28304 32982
rect 30208 32910 30236 33254
rect 30668 32910 30696 33390
rect 32232 33114 32260 37130
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 31576 33108 31628 33114
rect 31576 33050 31628 33056
rect 32220 33108 32272 33114
rect 32220 33050 32272 33056
rect 28264 32904 28316 32910
rect 28264 32846 28316 32852
rect 29736 32904 29788 32910
rect 29736 32846 29788 32852
rect 29828 32904 29880 32910
rect 29828 32846 29880 32852
rect 29920 32904 29972 32910
rect 29920 32846 29972 32852
rect 30196 32904 30248 32910
rect 30196 32846 30248 32852
rect 30656 32904 30708 32910
rect 30656 32846 30708 32852
rect 29748 32774 29776 32846
rect 29736 32768 29788 32774
rect 29736 32710 29788 32716
rect 28356 32428 28408 32434
rect 28356 32370 28408 32376
rect 28540 32428 28592 32434
rect 28540 32370 28592 32376
rect 29000 32428 29052 32434
rect 29000 32370 29052 32376
rect 29644 32428 29696 32434
rect 29644 32370 29696 32376
rect 28368 32065 28396 32370
rect 28078 32056 28134 32065
rect 28354 32056 28410 32065
rect 28134 32014 28304 32042
rect 28078 31991 28134 32000
rect 28170 31920 28226 31929
rect 28170 31855 28226 31864
rect 28080 31680 28132 31686
rect 28080 31622 28132 31628
rect 28092 31346 28120 31622
rect 28080 31340 28132 31346
rect 28080 31282 28132 31288
rect 27988 30932 28040 30938
rect 27988 30874 28040 30880
rect 27988 30728 28040 30734
rect 27988 30670 28040 30676
rect 28000 29782 28028 30670
rect 27988 29776 28040 29782
rect 27988 29718 28040 29724
rect 28000 29238 28028 29718
rect 28078 29472 28134 29481
rect 28078 29407 28134 29416
rect 27988 29232 28040 29238
rect 27988 29174 28040 29180
rect 28092 29034 28120 29407
rect 28080 29028 28132 29034
rect 28080 28970 28132 28976
rect 27896 28552 27948 28558
rect 27896 28494 27948 28500
rect 27804 27600 27856 27606
rect 27804 27542 27856 27548
rect 27712 27464 27764 27470
rect 27908 27452 27936 28494
rect 27988 28416 28040 28422
rect 27988 28358 28040 28364
rect 28000 28121 28028 28358
rect 27986 28112 28042 28121
rect 27986 28047 28042 28056
rect 27986 27704 28042 27713
rect 27986 27639 28042 27648
rect 27764 27424 27936 27452
rect 27712 27406 27764 27412
rect 27620 27056 27672 27062
rect 27620 26998 27672 27004
rect 27528 26852 27580 26858
rect 27528 26794 27580 26800
rect 27436 26444 27488 26450
rect 27436 26386 27488 26392
rect 27448 26353 27476 26386
rect 27434 26344 27490 26353
rect 27434 26279 27490 26288
rect 27526 26072 27582 26081
rect 27526 26007 27582 26016
rect 27434 25528 27490 25537
rect 27434 25463 27490 25472
rect 27448 25265 27476 25463
rect 27434 25256 27490 25265
rect 27434 25191 27490 25200
rect 27540 25158 27568 26007
rect 27620 25696 27672 25702
rect 27620 25638 27672 25644
rect 27632 25265 27660 25638
rect 27618 25256 27674 25265
rect 27618 25191 27674 25200
rect 27436 25152 27488 25158
rect 27436 25094 27488 25100
rect 27528 25152 27580 25158
rect 27528 25094 27580 25100
rect 27448 23866 27476 25094
rect 27528 24336 27580 24342
rect 27526 24304 27528 24313
rect 27620 24336 27672 24342
rect 27580 24304 27582 24313
rect 27620 24278 27672 24284
rect 27526 24239 27582 24248
rect 27632 24206 27660 24278
rect 27620 24200 27672 24206
rect 27620 24142 27672 24148
rect 27436 23860 27488 23866
rect 27436 23802 27488 23808
rect 27528 23792 27580 23798
rect 27528 23734 27580 23740
rect 27436 23724 27488 23730
rect 27436 23666 27488 23672
rect 27448 23526 27476 23666
rect 27436 23520 27488 23526
rect 27436 23462 27488 23468
rect 27540 23322 27568 23734
rect 27528 23316 27580 23322
rect 27528 23258 27580 23264
rect 27344 22704 27396 22710
rect 27344 22646 27396 22652
rect 27344 22568 27396 22574
rect 27344 22510 27396 22516
rect 27252 22228 27304 22234
rect 27252 22170 27304 22176
rect 27160 22092 27212 22098
rect 27160 22034 27212 22040
rect 27068 21412 27120 21418
rect 27068 21354 27120 21360
rect 26976 21140 27028 21146
rect 26976 21082 27028 21088
rect 26988 20777 27016 21082
rect 27068 20936 27120 20942
rect 27068 20878 27120 20884
rect 27080 20806 27108 20878
rect 27068 20800 27120 20806
rect 26974 20768 27030 20777
rect 27068 20742 27120 20748
rect 26974 20703 27030 20712
rect 26976 20256 27028 20262
rect 26976 20198 27028 20204
rect 26568 19680 26570 19689
rect 26514 19615 26570 19624
rect 26712 19672 26924 19700
rect 26516 18284 26568 18290
rect 26516 18226 26568 18232
rect 26424 17536 26476 17542
rect 26424 17478 26476 17484
rect 26240 17264 26292 17270
rect 26240 17206 26292 17212
rect 26528 17202 26556 18226
rect 26712 17762 26740 19672
rect 26988 19378 27016 20198
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 27080 19174 27108 20742
rect 27068 19168 27120 19174
rect 26974 19136 27030 19145
rect 27068 19110 27120 19116
rect 26974 19071 27030 19080
rect 26988 18358 27016 19071
rect 27066 18456 27122 18465
rect 27066 18391 27122 18400
rect 26976 18352 27028 18358
rect 26976 18294 27028 18300
rect 27080 18222 27108 18391
rect 27068 18216 27120 18222
rect 27068 18158 27120 18164
rect 26884 18080 26936 18086
rect 26884 18022 26936 18028
rect 26620 17734 26740 17762
rect 26790 17776 26846 17785
rect 26332 17196 26384 17202
rect 26332 17138 26384 17144
rect 26516 17196 26568 17202
rect 26516 17138 26568 17144
rect 26344 16658 26372 17138
rect 26332 16652 26384 16658
rect 26332 16594 26384 16600
rect 26148 16516 26200 16522
rect 26148 16458 26200 16464
rect 26160 15366 26188 16458
rect 26332 16176 26384 16182
rect 26332 16118 26384 16124
rect 26344 15910 26372 16118
rect 26422 16008 26478 16017
rect 26422 15943 26478 15952
rect 26332 15904 26384 15910
rect 26332 15846 26384 15852
rect 26344 15502 26372 15846
rect 26436 15609 26464 15943
rect 26528 15910 26556 17138
rect 26620 16250 26648 17734
rect 26790 17711 26846 17720
rect 26804 17610 26832 17711
rect 26792 17604 26844 17610
rect 26792 17546 26844 17552
rect 26700 17536 26752 17542
rect 26700 17478 26752 17484
rect 26712 17270 26740 17478
rect 26792 17332 26844 17338
rect 26792 17274 26844 17280
rect 26700 17264 26752 17270
rect 26700 17206 26752 17212
rect 26804 17082 26832 17274
rect 26712 17054 26832 17082
rect 26608 16244 26660 16250
rect 26608 16186 26660 16192
rect 26712 16130 26740 17054
rect 26896 16998 26924 18022
rect 26976 17876 27028 17882
rect 26976 17818 27028 17824
rect 26988 17377 27016 17818
rect 26974 17368 27030 17377
rect 26974 17303 27030 17312
rect 27080 17218 27108 18158
rect 27172 17338 27200 22034
rect 27356 21350 27384 22510
rect 27436 22432 27488 22438
rect 27436 22374 27488 22380
rect 27344 21344 27396 21350
rect 27344 21286 27396 21292
rect 27250 20632 27306 20641
rect 27250 20567 27306 20576
rect 27264 19922 27292 20567
rect 27252 19916 27304 19922
rect 27252 19858 27304 19864
rect 27448 19689 27476 22374
rect 27620 20800 27672 20806
rect 27724 20777 27752 27406
rect 27804 27124 27856 27130
rect 27804 27066 27856 27072
rect 27816 24886 27844 27066
rect 28000 26897 28028 27639
rect 27986 26888 28042 26897
rect 27986 26823 28042 26832
rect 27804 24880 27856 24886
rect 27804 24822 27856 24828
rect 27816 24120 27844 24822
rect 27896 24676 27948 24682
rect 27896 24618 27948 24624
rect 27908 24410 27936 24618
rect 27896 24404 27948 24410
rect 27896 24346 27948 24352
rect 28080 24336 28132 24342
rect 28078 24304 28080 24313
rect 28132 24304 28134 24313
rect 28078 24239 28134 24248
rect 27988 24200 28040 24206
rect 27988 24142 28040 24148
rect 27896 24132 27948 24138
rect 27816 24092 27896 24120
rect 27896 24074 27948 24080
rect 27802 23760 27858 23769
rect 27802 23695 27804 23704
rect 27856 23695 27858 23704
rect 27804 23666 27856 23672
rect 27802 23488 27858 23497
rect 27802 23423 27858 23432
rect 27816 23050 27844 23423
rect 27908 23322 27936 24074
rect 27896 23316 27948 23322
rect 27896 23258 27948 23264
rect 27804 23044 27856 23050
rect 27804 22986 27856 22992
rect 27816 22953 27844 22986
rect 27802 22944 27858 22953
rect 27802 22879 27858 22888
rect 28000 22234 28028 24142
rect 28184 23497 28212 31855
rect 28276 31113 28304 32014
rect 28354 31991 28410 32000
rect 28356 31748 28408 31754
rect 28356 31690 28408 31696
rect 28368 31346 28396 31690
rect 28552 31521 28580 32370
rect 28816 31816 28868 31822
rect 28816 31758 28868 31764
rect 28538 31512 28594 31521
rect 28538 31447 28594 31456
rect 28552 31414 28580 31447
rect 28540 31408 28592 31414
rect 28540 31350 28592 31356
rect 28356 31340 28408 31346
rect 28356 31282 28408 31288
rect 28262 31104 28318 31113
rect 28262 31039 28318 31048
rect 28368 30954 28396 31282
rect 28276 30926 28396 30954
rect 28722 30968 28778 30977
rect 28276 30870 28304 30926
rect 28722 30903 28724 30912
rect 28776 30903 28778 30912
rect 28724 30874 28776 30880
rect 28264 30864 28316 30870
rect 28264 30806 28316 30812
rect 28276 29238 28304 30806
rect 28448 30592 28500 30598
rect 28448 30534 28500 30540
rect 28356 29572 28408 29578
rect 28356 29514 28408 29520
rect 28368 29306 28396 29514
rect 28356 29300 28408 29306
rect 28356 29242 28408 29248
rect 28264 29232 28316 29238
rect 28264 29174 28316 29180
rect 28356 29164 28408 29170
rect 28356 29106 28408 29112
rect 28264 28484 28316 28490
rect 28264 28426 28316 28432
rect 28276 28393 28304 28426
rect 28262 28384 28318 28393
rect 28262 28319 28318 28328
rect 28276 26790 28304 28319
rect 28368 28257 28396 29106
rect 28460 28490 28488 30534
rect 28630 30152 28686 30161
rect 28630 30087 28686 30096
rect 28644 29578 28672 30087
rect 28724 29844 28776 29850
rect 28724 29786 28776 29792
rect 28632 29572 28684 29578
rect 28632 29514 28684 29520
rect 28540 29096 28592 29102
rect 28540 29038 28592 29044
rect 28448 28484 28500 28490
rect 28448 28426 28500 28432
rect 28354 28248 28410 28257
rect 28354 28183 28410 28192
rect 28460 26994 28488 28426
rect 28448 26988 28500 26994
rect 28448 26930 28500 26936
rect 28552 26897 28580 29038
rect 28632 28960 28684 28966
rect 28632 28902 28684 28908
rect 28644 28393 28672 28902
rect 28736 28422 28764 29786
rect 28828 28762 28856 31758
rect 28908 31136 28960 31142
rect 28908 31078 28960 31084
rect 28920 30734 28948 31078
rect 28908 30728 28960 30734
rect 28908 30670 28960 30676
rect 29012 29238 29040 32370
rect 29368 31272 29420 31278
rect 29368 31214 29420 31220
rect 29380 30258 29408 31214
rect 29092 30252 29144 30258
rect 29092 30194 29144 30200
rect 29368 30252 29420 30258
rect 29368 30194 29420 30200
rect 29104 29782 29132 30194
rect 29276 30184 29328 30190
rect 29276 30126 29328 30132
rect 29092 29776 29144 29782
rect 29092 29718 29144 29724
rect 29184 29776 29236 29782
rect 29184 29718 29236 29724
rect 29196 29306 29224 29718
rect 29288 29306 29316 30126
rect 29460 30048 29512 30054
rect 29460 29990 29512 29996
rect 29552 30048 29604 30054
rect 29552 29990 29604 29996
rect 29184 29300 29236 29306
rect 29184 29242 29236 29248
rect 29276 29300 29328 29306
rect 29472 29288 29500 29990
rect 29564 29889 29592 29990
rect 29550 29880 29606 29889
rect 29550 29815 29606 29824
rect 29550 29744 29606 29753
rect 29550 29679 29606 29688
rect 29564 29578 29592 29679
rect 29552 29572 29604 29578
rect 29552 29514 29604 29520
rect 29552 29300 29604 29306
rect 29472 29260 29552 29288
rect 29276 29242 29328 29248
rect 29552 29242 29604 29248
rect 29000 29232 29052 29238
rect 29000 29174 29052 29180
rect 29276 29164 29328 29170
rect 29276 29106 29328 29112
rect 29552 29164 29604 29170
rect 29552 29106 29604 29112
rect 28908 29028 28960 29034
rect 28960 28988 29040 29016
rect 28908 28970 28960 28976
rect 28906 28792 28962 28801
rect 28816 28756 28868 28762
rect 28906 28727 28962 28736
rect 28816 28698 28868 28704
rect 28920 28694 28948 28727
rect 29012 28694 29040 28988
rect 28908 28688 28960 28694
rect 28908 28630 28960 28636
rect 29000 28688 29052 28694
rect 29000 28630 29052 28636
rect 28816 28620 28868 28626
rect 28816 28562 28868 28568
rect 28828 28472 28856 28562
rect 28828 28444 28948 28472
rect 28724 28416 28776 28422
rect 28630 28384 28686 28393
rect 28724 28358 28776 28364
rect 28630 28319 28686 28328
rect 28736 28082 28764 28358
rect 28816 28144 28868 28150
rect 28816 28086 28868 28092
rect 28920 28098 28948 28444
rect 29000 28416 29052 28422
rect 29000 28358 29052 28364
rect 29012 28218 29040 28358
rect 29090 28248 29146 28257
rect 29000 28212 29052 28218
rect 29288 28234 29316 29106
rect 29460 29096 29512 29102
rect 29366 29064 29422 29073
rect 29460 29038 29512 29044
rect 29366 28999 29422 29008
rect 29380 28966 29408 28999
rect 29368 28960 29420 28966
rect 29368 28902 29420 28908
rect 29368 28416 29420 28422
rect 29368 28358 29420 28364
rect 29090 28183 29146 28192
rect 29196 28206 29316 28234
rect 29000 28154 29052 28160
rect 29104 28098 29132 28183
rect 28724 28076 28776 28082
rect 28724 28018 28776 28024
rect 28538 26888 28594 26897
rect 28356 26852 28408 26858
rect 28538 26823 28594 26832
rect 28356 26794 28408 26800
rect 28264 26784 28316 26790
rect 28264 26726 28316 26732
rect 28276 25702 28304 26726
rect 28264 25696 28316 25702
rect 28264 25638 28316 25644
rect 28264 24608 28316 24614
rect 28264 24550 28316 24556
rect 28276 24410 28304 24550
rect 28264 24404 28316 24410
rect 28264 24346 28316 24352
rect 28368 24206 28396 26794
rect 28630 25936 28686 25945
rect 28630 25871 28686 25880
rect 28540 25696 28592 25702
rect 28540 25638 28592 25644
rect 28448 25220 28500 25226
rect 28448 25162 28500 25168
rect 28460 24886 28488 25162
rect 28448 24880 28500 24886
rect 28448 24822 28500 24828
rect 28552 24206 28580 25638
rect 28644 25430 28672 25871
rect 28632 25424 28684 25430
rect 28632 25366 28684 25372
rect 28356 24200 28408 24206
rect 28356 24142 28408 24148
rect 28540 24200 28592 24206
rect 28540 24142 28592 24148
rect 28264 23520 28316 23526
rect 28170 23488 28226 23497
rect 28316 23480 28580 23508
rect 28264 23462 28316 23468
rect 28170 23423 28226 23432
rect 28080 23044 28132 23050
rect 28080 22986 28132 22992
rect 27804 22228 27856 22234
rect 27804 22170 27856 22176
rect 27988 22228 28040 22234
rect 27988 22170 28040 22176
rect 27816 21486 27844 22170
rect 27986 22128 28042 22137
rect 28092 22114 28120 22986
rect 28262 22672 28318 22681
rect 28262 22607 28318 22616
rect 28172 22228 28224 22234
rect 28172 22170 28224 22176
rect 28042 22086 28120 22114
rect 27986 22063 27988 22072
rect 28040 22063 28042 22072
rect 27988 22034 28040 22040
rect 28080 22024 28132 22030
rect 28078 21992 28080 22001
rect 28132 21992 28134 22001
rect 28078 21927 28134 21936
rect 27804 21480 27856 21486
rect 27804 21422 27856 21428
rect 27894 21040 27950 21049
rect 27894 20975 27950 20984
rect 27804 20936 27856 20942
rect 27804 20878 27856 20884
rect 27620 20742 27672 20748
rect 27710 20768 27766 20777
rect 27632 20262 27660 20742
rect 27710 20703 27766 20712
rect 27620 20256 27672 20262
rect 27620 20198 27672 20204
rect 27434 19680 27490 19689
rect 27434 19615 27490 19624
rect 27342 19408 27398 19417
rect 27342 19343 27398 19352
rect 27252 18148 27304 18154
rect 27252 18090 27304 18096
rect 27264 17814 27292 18090
rect 27252 17808 27304 17814
rect 27252 17750 27304 17756
rect 27252 17536 27304 17542
rect 27252 17478 27304 17484
rect 27160 17332 27212 17338
rect 27160 17274 27212 17280
rect 26988 17190 27108 17218
rect 26884 16992 26936 16998
rect 26884 16934 26936 16940
rect 26792 16788 26844 16794
rect 26792 16730 26844 16736
rect 26620 16102 26740 16130
rect 26516 15904 26568 15910
rect 26516 15846 26568 15852
rect 26422 15600 26478 15609
rect 26422 15535 26478 15544
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 26240 15428 26292 15434
rect 26240 15370 26292 15376
rect 26148 15360 26200 15366
rect 26148 15302 26200 15308
rect 26252 15162 26280 15370
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26148 15020 26200 15026
rect 26148 14962 26200 14968
rect 26160 14006 26188 14962
rect 26148 14000 26200 14006
rect 26148 13942 26200 13948
rect 26056 13524 26108 13530
rect 26056 13466 26108 13472
rect 25872 13252 25924 13258
rect 25872 13194 25924 13200
rect 26054 13016 26110 13025
rect 26160 12986 26188 13942
rect 26252 13938 26280 15098
rect 26436 15026 26464 15535
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 26330 14920 26386 14929
rect 26330 14855 26386 14864
rect 26344 14822 26372 14855
rect 26332 14816 26384 14822
rect 26332 14758 26384 14764
rect 26424 14408 26476 14414
rect 26424 14350 26476 14356
rect 26240 13932 26292 13938
rect 26240 13874 26292 13880
rect 26332 13864 26384 13870
rect 26332 13806 26384 13812
rect 26344 13326 26372 13806
rect 26436 13734 26464 14350
rect 26528 13977 26556 15846
rect 26620 15314 26648 16102
rect 26698 15872 26754 15881
rect 26698 15807 26754 15816
rect 26712 15502 26740 15807
rect 26700 15496 26752 15502
rect 26700 15438 26752 15444
rect 26698 15328 26754 15337
rect 26620 15286 26698 15314
rect 26698 15263 26754 15272
rect 26514 13968 26570 13977
rect 26514 13903 26516 13912
rect 26568 13903 26570 13912
rect 26608 13932 26660 13938
rect 26516 13874 26568 13880
rect 26608 13874 26660 13880
rect 26424 13728 26476 13734
rect 26424 13670 26476 13676
rect 26620 13530 26648 13874
rect 26712 13734 26740 15263
rect 26804 13938 26832 16730
rect 26884 16720 26936 16726
rect 26884 16662 26936 16668
rect 26896 16522 26924 16662
rect 26884 16516 26936 16522
rect 26884 16458 26936 16464
rect 26882 16280 26938 16289
rect 26882 16215 26938 16224
rect 26896 15881 26924 16215
rect 26882 15872 26938 15881
rect 26882 15807 26938 15816
rect 26988 15434 27016 17190
rect 27160 17128 27212 17134
rect 27080 17076 27160 17082
rect 27080 17070 27212 17076
rect 27080 17054 27200 17070
rect 26976 15428 27028 15434
rect 26976 15370 27028 15376
rect 27080 15366 27108 17054
rect 27160 16992 27212 16998
rect 27160 16934 27212 16940
rect 27068 15360 27120 15366
rect 27068 15302 27120 15308
rect 26884 15088 26936 15094
rect 26884 15030 26936 15036
rect 26896 14822 26924 15030
rect 27080 14822 27108 15302
rect 26884 14816 26936 14822
rect 26884 14758 26936 14764
rect 27068 14816 27120 14822
rect 27068 14758 27120 14764
rect 27172 13938 27200 16934
rect 26792 13932 26844 13938
rect 26792 13874 26844 13880
rect 27160 13932 27212 13938
rect 27160 13874 27212 13880
rect 26700 13728 26752 13734
rect 26700 13670 26752 13676
rect 27172 13530 27200 13874
rect 26608 13524 26660 13530
rect 26608 13466 26660 13472
rect 27160 13524 27212 13530
rect 27160 13466 27212 13472
rect 26620 13394 26648 13466
rect 26608 13388 26660 13394
rect 26608 13330 26660 13336
rect 26332 13320 26384 13326
rect 26332 13262 26384 13268
rect 26054 12951 26110 12960
rect 26148 12980 26200 12986
rect 26068 12782 26096 12951
rect 26148 12922 26200 12928
rect 25780 12776 25832 12782
rect 25780 12718 25832 12724
rect 26056 12776 26108 12782
rect 26056 12718 26108 12724
rect 25686 12472 25742 12481
rect 27264 12434 27292 17478
rect 27356 16726 27384 19343
rect 27344 16720 27396 16726
rect 27344 16662 27396 16668
rect 27342 16552 27398 16561
rect 27342 16487 27398 16496
rect 27356 16289 27384 16487
rect 27342 16280 27398 16289
rect 27342 16215 27398 16224
rect 27342 15192 27398 15201
rect 27342 15127 27344 15136
rect 27396 15127 27398 15136
rect 27344 15098 27396 15104
rect 27344 14952 27396 14958
rect 27344 14894 27396 14900
rect 27356 14482 27384 14894
rect 27344 14476 27396 14482
rect 27344 14418 27396 14424
rect 27448 14414 27476 19615
rect 27816 19378 27844 20878
rect 27908 20777 27936 20975
rect 27894 20768 27950 20777
rect 27894 20703 27950 20712
rect 27986 20632 28042 20641
rect 27986 20567 27988 20576
rect 28040 20567 28042 20576
rect 27988 20538 28040 20544
rect 28092 20466 28120 21927
rect 28184 21593 28212 22170
rect 28170 21584 28226 21593
rect 28170 21519 28226 21528
rect 28276 21468 28304 22607
rect 28446 22264 28502 22273
rect 28446 22199 28448 22208
rect 28500 22199 28502 22208
rect 28448 22170 28500 22176
rect 28354 21992 28410 22001
rect 28354 21927 28410 21936
rect 28184 21440 28304 21468
rect 28080 20460 28132 20466
rect 28080 20402 28132 20408
rect 27804 19372 27856 19378
rect 27804 19314 27856 19320
rect 27988 19372 28040 19378
rect 27988 19314 28040 19320
rect 27896 19304 27948 19310
rect 27802 19272 27858 19281
rect 27896 19246 27948 19252
rect 27802 19207 27858 19216
rect 27528 18964 27580 18970
rect 27528 18906 27580 18912
rect 27540 17882 27568 18906
rect 27620 18148 27672 18154
rect 27620 18090 27672 18096
rect 27528 17876 27580 17882
rect 27528 17818 27580 17824
rect 27632 17746 27660 18090
rect 27712 18080 27764 18086
rect 27816 18057 27844 19207
rect 27908 18970 27936 19246
rect 27896 18964 27948 18970
rect 27896 18906 27948 18912
rect 27896 18420 27948 18426
rect 27896 18362 27948 18368
rect 27712 18022 27764 18028
rect 27802 18048 27858 18057
rect 27620 17740 27672 17746
rect 27620 17682 27672 17688
rect 27528 17672 27580 17678
rect 27528 17614 27580 17620
rect 27540 17241 27568 17614
rect 27724 17270 27752 18022
rect 27802 17983 27858 17992
rect 27712 17264 27764 17270
rect 27526 17232 27582 17241
rect 27712 17206 27764 17212
rect 27526 17167 27582 17176
rect 27816 17082 27844 17983
rect 27632 17054 27844 17082
rect 27528 16108 27580 16114
rect 27528 16050 27580 16056
rect 27540 15366 27568 16050
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27436 14408 27488 14414
rect 27436 14350 27488 14356
rect 27540 13938 27568 15302
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 25686 12407 25742 12416
rect 27172 12406 27292 12434
rect 27172 12345 27200 12406
rect 27158 12336 27214 12345
rect 27158 12271 27214 12280
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 27632 10985 27660 17054
rect 27908 16833 27936 18362
rect 28000 18034 28028 19314
rect 28092 19310 28120 20402
rect 28080 19304 28132 19310
rect 28080 19246 28132 19252
rect 28000 18006 28120 18034
rect 27986 17912 28042 17921
rect 27986 17847 28042 17856
rect 28000 17814 28028 17847
rect 27988 17808 28040 17814
rect 27988 17750 28040 17756
rect 28092 17678 28120 18006
rect 28184 17882 28212 21440
rect 28264 20460 28316 20466
rect 28264 20402 28316 20408
rect 28276 18766 28304 20402
rect 28264 18760 28316 18766
rect 28264 18702 28316 18708
rect 28276 18290 28304 18702
rect 28264 18284 28316 18290
rect 28264 18226 28316 18232
rect 28172 17876 28224 17882
rect 28172 17818 28224 17824
rect 28172 17740 28224 17746
rect 28172 17682 28224 17688
rect 27988 17672 28040 17678
rect 27988 17614 28040 17620
rect 28080 17672 28132 17678
rect 28080 17614 28132 17620
rect 28000 16998 28028 17614
rect 28078 17232 28134 17241
rect 28078 17167 28080 17176
rect 28132 17167 28134 17176
rect 28080 17138 28132 17144
rect 27988 16992 28040 16998
rect 27988 16934 28040 16940
rect 27894 16824 27950 16833
rect 28184 16794 28212 17682
rect 28368 17241 28396 21927
rect 28446 21040 28502 21049
rect 28446 20975 28502 20984
rect 28460 18222 28488 20975
rect 28552 18766 28580 23480
rect 28644 22273 28672 25366
rect 28630 22264 28686 22273
rect 28630 22199 28686 22208
rect 28736 20534 28764 28018
rect 28828 27849 28856 28086
rect 28920 28070 29132 28098
rect 28908 27872 28960 27878
rect 28814 27840 28870 27849
rect 28908 27814 28960 27820
rect 28814 27775 28870 27784
rect 28816 27464 28868 27470
rect 28816 27406 28868 27412
rect 28828 25537 28856 27406
rect 28920 26625 28948 27814
rect 29092 27328 29144 27334
rect 29092 27270 29144 27276
rect 28998 27160 29054 27169
rect 28998 27095 29054 27104
rect 29012 26858 29040 27095
rect 29000 26852 29052 26858
rect 29000 26794 29052 26800
rect 28906 26616 28962 26625
rect 28906 26551 28962 26560
rect 28814 25528 28870 25537
rect 28814 25463 28870 25472
rect 28920 25412 28948 26551
rect 29104 25537 29132 27270
rect 29196 25906 29224 28206
rect 29380 27849 29408 28358
rect 29472 28218 29500 29038
rect 29460 28212 29512 28218
rect 29460 28154 29512 28160
rect 29366 27840 29422 27849
rect 29366 27775 29422 27784
rect 29564 27614 29592 29106
rect 29656 29050 29684 32370
rect 29748 32366 29776 32710
rect 29840 32570 29868 32846
rect 29828 32564 29880 32570
rect 29828 32506 29880 32512
rect 29736 32360 29788 32366
rect 29736 32302 29788 32308
rect 29736 32224 29788 32230
rect 29736 32166 29788 32172
rect 29748 31958 29776 32166
rect 29736 31952 29788 31958
rect 29736 31894 29788 31900
rect 29932 30598 29960 32846
rect 30288 32836 30340 32842
rect 30288 32778 30340 32784
rect 31024 32836 31076 32842
rect 31024 32778 31076 32784
rect 30300 31414 30328 32778
rect 31036 32570 31064 32778
rect 31024 32564 31076 32570
rect 31024 32506 31076 32512
rect 31392 32496 31444 32502
rect 31392 32438 31444 32444
rect 30380 32360 30432 32366
rect 30380 32302 30432 32308
rect 30392 32201 30420 32302
rect 30378 32192 30434 32201
rect 30378 32127 30434 32136
rect 31404 31890 31432 32438
rect 31588 32366 31616 33050
rect 36084 32836 36136 32842
rect 36084 32778 36136 32784
rect 32128 32768 32180 32774
rect 32128 32710 32180 32716
rect 32140 32434 32168 32710
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 32128 32428 32180 32434
rect 32128 32370 32180 32376
rect 31576 32360 31628 32366
rect 31576 32302 31628 32308
rect 32128 32292 32180 32298
rect 32128 32234 32180 32240
rect 30932 31884 30984 31890
rect 30932 31826 30984 31832
rect 31392 31884 31444 31890
rect 31392 31826 31444 31832
rect 30378 31784 30434 31793
rect 30434 31728 30604 31754
rect 30378 31726 30604 31728
rect 30378 31719 30434 31726
rect 30288 31408 30340 31414
rect 30288 31350 30340 31356
rect 29920 30592 29972 30598
rect 30300 30569 30328 31350
rect 30576 31226 30604 31726
rect 30576 31198 30880 31226
rect 30562 31104 30618 31113
rect 30562 31039 30618 31048
rect 29920 30534 29972 30540
rect 30286 30560 30342 30569
rect 30286 30495 30342 30504
rect 30196 30252 30248 30258
rect 30196 30194 30248 30200
rect 30380 30252 30432 30258
rect 30380 30194 30432 30200
rect 29828 30184 29880 30190
rect 30104 30184 30156 30190
rect 29828 30126 29880 30132
rect 30102 30152 30104 30161
rect 30156 30152 30158 30161
rect 29736 29776 29788 29782
rect 29736 29718 29788 29724
rect 29748 29238 29776 29718
rect 29840 29714 29868 30126
rect 30102 30087 30158 30096
rect 29920 30048 29972 30054
rect 29920 29990 29972 29996
rect 29828 29708 29880 29714
rect 29828 29650 29880 29656
rect 29736 29232 29788 29238
rect 29736 29174 29788 29180
rect 29656 29022 29776 29050
rect 29932 29034 29960 29990
rect 30208 29866 30236 30194
rect 30288 30116 30340 30122
rect 30288 30058 30340 30064
rect 30300 30025 30328 30058
rect 30286 30016 30342 30025
rect 30286 29951 30342 29960
rect 30012 29844 30064 29850
rect 30208 29838 30328 29866
rect 30392 29850 30420 30194
rect 30576 30190 30604 31039
rect 30748 30252 30800 30258
rect 30748 30194 30800 30200
rect 30564 30184 30616 30190
rect 30564 30126 30616 30132
rect 30472 30048 30524 30054
rect 30472 29990 30524 29996
rect 30012 29786 30064 29792
rect 30024 29492 30052 29786
rect 30300 29730 30328 29838
rect 30380 29844 30432 29850
rect 30380 29786 30432 29792
rect 30300 29714 30420 29730
rect 30300 29708 30432 29714
rect 30300 29702 30380 29708
rect 30380 29650 30432 29656
rect 30104 29504 30156 29510
rect 30024 29464 30104 29492
rect 30024 29345 30052 29464
rect 30104 29446 30156 29452
rect 30010 29336 30066 29345
rect 30010 29271 30066 29280
rect 29748 28948 29776 29022
rect 29920 29028 29972 29034
rect 29920 28970 29972 28976
rect 29288 27586 29592 27614
rect 29656 28920 29776 28948
rect 29828 28960 29880 28966
rect 29184 25900 29236 25906
rect 29184 25842 29236 25848
rect 29090 25528 29146 25537
rect 29090 25463 29146 25472
rect 28828 25384 28948 25412
rect 28828 24868 28856 25384
rect 28908 25220 28960 25226
rect 28908 25162 28960 25168
rect 29092 25220 29144 25226
rect 29092 25162 29144 25168
rect 28920 24993 28948 25162
rect 28906 24984 28962 24993
rect 28906 24919 28962 24928
rect 28828 24840 28948 24868
rect 28816 23724 28868 23730
rect 28816 23666 28868 23672
rect 28724 20528 28776 20534
rect 28724 20470 28776 20476
rect 28828 20058 28856 23666
rect 28816 20052 28868 20058
rect 28816 19994 28868 20000
rect 28920 19938 28948 24840
rect 29104 24138 29132 25162
rect 29092 24132 29144 24138
rect 29092 24074 29144 24080
rect 29104 23905 29132 24074
rect 29090 23896 29146 23905
rect 29000 23860 29052 23866
rect 29090 23831 29146 23840
rect 29000 23802 29052 23808
rect 29012 23254 29040 23802
rect 29196 23610 29224 25842
rect 29288 24410 29316 27586
rect 29460 27532 29512 27538
rect 29460 27474 29512 27480
rect 29368 27328 29420 27334
rect 29368 27270 29420 27276
rect 29380 26994 29408 27270
rect 29368 26988 29420 26994
rect 29368 26930 29420 26936
rect 29276 24404 29328 24410
rect 29276 24346 29328 24352
rect 29104 23582 29224 23610
rect 29000 23248 29052 23254
rect 29000 23190 29052 23196
rect 29104 23186 29132 23582
rect 29184 23520 29236 23526
rect 29184 23462 29236 23468
rect 29092 23180 29144 23186
rect 29092 23122 29144 23128
rect 29000 23044 29052 23050
rect 29000 22986 29052 22992
rect 29012 22574 29040 22986
rect 29092 22704 29144 22710
rect 29092 22646 29144 22652
rect 29000 22568 29052 22574
rect 29000 22510 29052 22516
rect 29000 22432 29052 22438
rect 28998 22400 29000 22409
rect 29052 22400 29054 22409
rect 28998 22335 29054 22344
rect 29104 22273 29132 22646
rect 29196 22438 29224 23462
rect 29276 23180 29328 23186
rect 29276 23122 29328 23128
rect 29288 22642 29316 23122
rect 29380 22710 29408 26930
rect 29472 26518 29500 27474
rect 29552 27396 29604 27402
rect 29552 27338 29604 27344
rect 29460 26512 29512 26518
rect 29460 26454 29512 26460
rect 29564 26314 29592 27338
rect 29552 26308 29604 26314
rect 29552 26250 29604 26256
rect 29552 25696 29604 25702
rect 29552 25638 29604 25644
rect 29564 25294 29592 25638
rect 29552 25288 29604 25294
rect 29552 25230 29604 25236
rect 29460 24948 29512 24954
rect 29460 24890 29512 24896
rect 29368 22704 29420 22710
rect 29368 22646 29420 22652
rect 29276 22636 29328 22642
rect 29276 22578 29328 22584
rect 29366 22536 29422 22545
rect 29276 22500 29328 22506
rect 29366 22471 29422 22480
rect 29276 22442 29328 22448
rect 29184 22432 29236 22438
rect 29184 22374 29236 22380
rect 29090 22264 29146 22273
rect 29090 22199 29146 22208
rect 29000 22024 29052 22030
rect 29000 21966 29052 21972
rect 29012 20466 29040 21966
rect 29104 20602 29132 22199
rect 29182 21720 29238 21729
rect 29182 21655 29238 21664
rect 29092 20596 29144 20602
rect 29092 20538 29144 20544
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 29092 20392 29144 20398
rect 29090 20360 29092 20369
rect 29144 20360 29146 20369
rect 29090 20295 29146 20304
rect 29000 20256 29052 20262
rect 29000 20198 29052 20204
rect 29012 20097 29040 20198
rect 28998 20088 29054 20097
rect 28998 20023 29054 20032
rect 28644 19910 28948 19938
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 28540 18624 28592 18630
rect 28540 18566 28592 18572
rect 28552 18358 28580 18566
rect 28540 18352 28592 18358
rect 28540 18294 28592 18300
rect 28448 18216 28500 18222
rect 28448 18158 28500 18164
rect 28538 18048 28594 18057
rect 28538 17983 28594 17992
rect 28448 17536 28500 17542
rect 28448 17478 28500 17484
rect 28354 17232 28410 17241
rect 28354 17167 28410 17176
rect 28460 16794 28488 17478
rect 27894 16759 27950 16768
rect 28172 16788 28224 16794
rect 28172 16730 28224 16736
rect 28448 16788 28500 16794
rect 28448 16730 28500 16736
rect 28552 16658 28580 17983
rect 28644 17746 28672 19910
rect 28908 19848 28960 19854
rect 28908 19790 28960 19796
rect 28814 19000 28870 19009
rect 28920 18970 28948 19790
rect 29104 19786 29132 20295
rect 29000 19780 29052 19786
rect 29000 19722 29052 19728
rect 29092 19780 29144 19786
rect 29092 19722 29144 19728
rect 29012 19310 29040 19722
rect 29000 19304 29052 19310
rect 29000 19246 29052 19252
rect 28814 18935 28870 18944
rect 28908 18964 28960 18970
rect 28828 18850 28856 18935
rect 28908 18906 28960 18912
rect 28828 18822 28948 18850
rect 28920 18766 28948 18822
rect 28816 18760 28868 18766
rect 28816 18702 28868 18708
rect 28908 18760 28960 18766
rect 28908 18702 28960 18708
rect 28724 18624 28776 18630
rect 28724 18566 28776 18572
rect 28736 18154 28764 18566
rect 28724 18148 28776 18154
rect 28724 18090 28776 18096
rect 28632 17740 28684 17746
rect 28632 17682 28684 17688
rect 28828 17626 28856 18702
rect 29012 18426 29040 19246
rect 29090 19136 29146 19145
rect 29090 19071 29146 19080
rect 29104 18766 29132 19071
rect 29196 18766 29224 21655
rect 29288 21049 29316 22442
rect 29380 21457 29408 22471
rect 29366 21448 29422 21457
rect 29366 21383 29422 21392
rect 29274 21040 29330 21049
rect 29274 20975 29330 20984
rect 29276 20460 29328 20466
rect 29276 20402 29328 20408
rect 29288 20262 29316 20402
rect 29276 20256 29328 20262
rect 29276 20198 29328 20204
rect 29368 20256 29420 20262
rect 29368 20198 29420 20204
rect 29274 20088 29330 20097
rect 29274 20023 29330 20032
rect 29288 19689 29316 20023
rect 29380 19922 29408 20198
rect 29368 19916 29420 19922
rect 29368 19858 29420 19864
rect 29274 19680 29330 19689
rect 29274 19615 29330 19624
rect 29092 18760 29144 18766
rect 29092 18702 29144 18708
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 29000 18420 29052 18426
rect 29000 18362 29052 18368
rect 29104 18170 29132 18702
rect 29368 18692 29420 18698
rect 29368 18634 29420 18640
rect 29274 18592 29330 18601
rect 29274 18527 29330 18536
rect 29288 18358 29316 18527
rect 29276 18352 29328 18358
rect 29276 18294 29328 18300
rect 29380 18222 29408 18634
rect 29368 18216 29420 18222
rect 29104 18142 29224 18170
rect 29368 18158 29420 18164
rect 29196 18086 29224 18142
rect 29184 18080 29236 18086
rect 29184 18022 29236 18028
rect 29366 17912 29422 17921
rect 29366 17847 29422 17856
rect 29380 17678 29408 17847
rect 28736 17598 28856 17626
rect 29368 17672 29420 17678
rect 29368 17614 29420 17620
rect 29472 17626 29500 24890
rect 29552 24200 29604 24206
rect 29552 24142 29604 24148
rect 29564 23866 29592 24142
rect 29552 23860 29604 23866
rect 29552 23802 29604 23808
rect 29552 23724 29604 23730
rect 29552 23666 29604 23672
rect 29564 23254 29592 23666
rect 29656 23526 29684 28920
rect 29828 28902 29880 28908
rect 29736 28756 29788 28762
rect 29736 28698 29788 28704
rect 29748 27538 29776 28698
rect 29840 28393 29868 28902
rect 30288 28552 30340 28558
rect 30288 28494 30340 28500
rect 29826 28384 29882 28393
rect 29826 28319 29882 28328
rect 30196 28144 30248 28150
rect 30196 28086 30248 28092
rect 29920 28076 29972 28082
rect 29920 28018 29972 28024
rect 29736 27532 29788 27538
rect 29736 27474 29788 27480
rect 29736 26240 29788 26246
rect 29736 26182 29788 26188
rect 29748 25294 29776 26182
rect 29828 25492 29880 25498
rect 29828 25434 29880 25440
rect 29736 25288 29788 25294
rect 29736 25230 29788 25236
rect 29840 24993 29868 25434
rect 29932 25430 29960 28018
rect 30010 27976 30066 27985
rect 30010 27911 30066 27920
rect 29920 25424 29972 25430
rect 29920 25366 29972 25372
rect 30024 25242 30052 27911
rect 30102 26072 30158 26081
rect 30102 26007 30158 26016
rect 30116 25498 30144 26007
rect 30104 25492 30156 25498
rect 30104 25434 30156 25440
rect 30104 25356 30156 25362
rect 30104 25298 30156 25304
rect 29932 25214 30052 25242
rect 29826 24984 29882 24993
rect 29826 24919 29882 24928
rect 29828 24404 29880 24410
rect 29828 24346 29880 24352
rect 29734 24304 29790 24313
rect 29734 24239 29790 24248
rect 29748 23905 29776 24239
rect 29734 23896 29790 23905
rect 29734 23831 29790 23840
rect 29840 23780 29868 24346
rect 29932 23866 29960 25214
rect 30012 25152 30064 25158
rect 30012 25094 30064 25100
rect 29920 23860 29972 23866
rect 29920 23802 29972 23808
rect 29748 23752 29868 23780
rect 29644 23520 29696 23526
rect 29644 23462 29696 23468
rect 29552 23248 29604 23254
rect 29552 23190 29604 23196
rect 29644 23248 29696 23254
rect 29644 23190 29696 23196
rect 29552 22704 29604 22710
rect 29552 22646 29604 22652
rect 29564 18834 29592 22646
rect 29552 18828 29604 18834
rect 29552 18770 29604 18776
rect 29564 18290 29592 18770
rect 29552 18284 29604 18290
rect 29552 18226 29604 18232
rect 29656 17660 29684 23190
rect 29748 22506 29776 23752
rect 29920 23724 29972 23730
rect 29920 23666 29972 23672
rect 29828 23520 29880 23526
rect 29826 23488 29828 23497
rect 29880 23488 29882 23497
rect 29826 23423 29882 23432
rect 29840 23254 29868 23423
rect 29828 23248 29880 23254
rect 29828 23190 29880 23196
rect 29828 22704 29880 22710
rect 29828 22646 29880 22652
rect 29736 22500 29788 22506
rect 29736 22442 29788 22448
rect 29734 21448 29790 21457
rect 29734 21383 29736 21392
rect 29788 21383 29790 21392
rect 29736 21354 29788 21360
rect 29736 20868 29788 20874
rect 29736 20810 29788 20816
rect 29748 20534 29776 20810
rect 29736 20528 29788 20534
rect 29736 20470 29788 20476
rect 29736 20324 29788 20330
rect 29736 20266 29788 20272
rect 29748 19553 29776 20266
rect 29840 19922 29868 22646
rect 29828 19916 29880 19922
rect 29828 19858 29880 19864
rect 29932 19802 29960 23666
rect 30024 21350 30052 25094
rect 30116 24954 30144 25298
rect 30104 24948 30156 24954
rect 30104 24890 30156 24896
rect 30104 24268 30156 24274
rect 30104 24210 30156 24216
rect 30116 24070 30144 24210
rect 30104 24064 30156 24070
rect 30104 24006 30156 24012
rect 30104 23860 30156 23866
rect 30104 23802 30156 23808
rect 30012 21344 30064 21350
rect 30012 21286 30064 21292
rect 30010 20632 30066 20641
rect 30010 20567 30066 20576
rect 30024 20330 30052 20567
rect 30012 20324 30064 20330
rect 30012 20266 30064 20272
rect 29840 19774 29960 19802
rect 30012 19780 30064 19786
rect 29734 19544 29790 19553
rect 29734 19479 29790 19488
rect 29734 18048 29790 18057
rect 29734 17983 29790 17992
rect 29748 17882 29776 17983
rect 29840 17882 29868 19774
rect 30012 19722 30064 19728
rect 29920 19508 29972 19514
rect 29920 19450 29972 19456
rect 29736 17876 29788 17882
rect 29736 17818 29788 17824
rect 29828 17876 29880 17882
rect 29828 17818 29880 17824
rect 29736 17672 29788 17678
rect 29550 17640 29606 17649
rect 29472 17598 29550 17626
rect 28540 16652 28592 16658
rect 28540 16594 28592 16600
rect 28264 16516 28316 16522
rect 28264 16458 28316 16464
rect 28080 16244 28132 16250
rect 28080 16186 28132 16192
rect 28092 15706 28120 16186
rect 28276 15706 28304 16458
rect 28080 15700 28132 15706
rect 28080 15642 28132 15648
rect 28264 15700 28316 15706
rect 28264 15642 28316 15648
rect 27804 15428 27856 15434
rect 27804 15370 27856 15376
rect 27816 15162 27844 15370
rect 27804 15156 27856 15162
rect 27804 15098 27856 15104
rect 28736 15026 28764 17598
rect 29550 17575 29552 17584
rect 29604 17575 29606 17584
rect 29656 17632 29736 17660
rect 29552 17546 29604 17552
rect 28816 17536 28868 17542
rect 28816 17478 28868 17484
rect 27712 15020 27764 15026
rect 27712 14962 27764 14968
rect 28724 15020 28776 15026
rect 28724 14962 28776 14968
rect 27724 14657 27752 14962
rect 27804 14952 27856 14958
rect 27804 14894 27856 14900
rect 27816 14822 27844 14894
rect 27804 14816 27856 14822
rect 27802 14784 27804 14793
rect 27856 14784 27858 14793
rect 27802 14719 27858 14728
rect 27710 14648 27766 14657
rect 27710 14583 27766 14592
rect 28828 14346 28856 17478
rect 29656 17202 29684 17632
rect 29736 17614 29788 17620
rect 29644 17196 29696 17202
rect 29644 17138 29696 17144
rect 29552 17128 29604 17134
rect 29840 17082 29868 17818
rect 29552 17070 29604 17076
rect 29368 16992 29420 16998
rect 29368 16934 29420 16940
rect 29460 16992 29512 16998
rect 29460 16934 29512 16940
rect 29380 16726 29408 16934
rect 29368 16720 29420 16726
rect 29368 16662 29420 16668
rect 29000 16584 29052 16590
rect 28906 16552 28962 16561
rect 29000 16526 29052 16532
rect 28906 16487 28962 16496
rect 28920 16454 28948 16487
rect 28908 16448 28960 16454
rect 28908 16390 28960 16396
rect 29012 16250 29040 16526
rect 29368 16516 29420 16522
rect 29368 16458 29420 16464
rect 29184 16448 29236 16454
rect 29184 16390 29236 16396
rect 29000 16244 29052 16250
rect 29000 16186 29052 16192
rect 29092 15700 29144 15706
rect 29092 15642 29144 15648
rect 28816 14340 28868 14346
rect 28816 14282 28868 14288
rect 28078 14104 28134 14113
rect 28078 14039 28080 14048
rect 28132 14039 28134 14048
rect 29000 14068 29052 14074
rect 28080 14010 28132 14016
rect 29000 14010 29052 14016
rect 28908 14000 28960 14006
rect 28828 13960 28908 13988
rect 28540 13932 28592 13938
rect 28540 13874 28592 13880
rect 27712 13864 27764 13870
rect 27712 13806 27764 13812
rect 27724 12306 27752 13806
rect 28552 13326 28580 13874
rect 28828 13802 28856 13960
rect 28908 13942 28960 13948
rect 28816 13796 28868 13802
rect 28816 13738 28868 13744
rect 28908 13796 28960 13802
rect 28908 13738 28960 13744
rect 28540 13320 28592 13326
rect 28540 13262 28592 13268
rect 28828 13258 28856 13738
rect 28920 13394 28948 13738
rect 29012 13530 29040 14010
rect 29000 13524 29052 13530
rect 29000 13466 29052 13472
rect 28908 13388 28960 13394
rect 28908 13330 28960 13336
rect 28356 13252 28408 13258
rect 28356 13194 28408 13200
rect 28816 13252 28868 13258
rect 28816 13194 28868 13200
rect 28368 13161 28396 13194
rect 28354 13152 28410 13161
rect 28354 13087 28410 13096
rect 27712 12300 27764 12306
rect 27712 12242 27764 12248
rect 29104 12209 29132 15642
rect 29196 15570 29224 16390
rect 29380 16046 29408 16458
rect 29368 16040 29420 16046
rect 29368 15982 29420 15988
rect 29184 15564 29236 15570
rect 29184 15506 29236 15512
rect 29472 15094 29500 16934
rect 29564 16017 29592 17070
rect 29748 17054 29868 17082
rect 29748 16998 29776 17054
rect 29736 16992 29788 16998
rect 29736 16934 29788 16940
rect 29932 16522 29960 19450
rect 29920 16516 29972 16522
rect 29920 16458 29972 16464
rect 29642 16416 29698 16425
rect 29642 16351 29698 16360
rect 29656 16114 29684 16351
rect 29644 16108 29696 16114
rect 29644 16050 29696 16056
rect 29828 16108 29880 16114
rect 29828 16050 29880 16056
rect 29550 16008 29606 16017
rect 29550 15943 29606 15952
rect 29734 16008 29790 16017
rect 29734 15943 29790 15952
rect 29748 15910 29776 15943
rect 29736 15904 29788 15910
rect 29736 15846 29788 15852
rect 29550 15600 29606 15609
rect 29550 15535 29606 15544
rect 29564 15502 29592 15535
rect 29552 15496 29604 15502
rect 29552 15438 29604 15444
rect 29644 15496 29696 15502
rect 29644 15438 29696 15444
rect 29564 15094 29592 15438
rect 29460 15088 29512 15094
rect 29460 15030 29512 15036
rect 29552 15088 29604 15094
rect 29552 15030 29604 15036
rect 29656 13394 29684 15438
rect 29644 13388 29696 13394
rect 29644 13330 29696 13336
rect 29460 13252 29512 13258
rect 29460 13194 29512 13200
rect 29472 12918 29500 13194
rect 29748 12918 29776 15846
rect 29840 13569 29868 16050
rect 29932 15706 29960 16458
rect 29920 15700 29972 15706
rect 29920 15642 29972 15648
rect 29826 13560 29882 13569
rect 30024 13530 30052 19722
rect 30116 18970 30144 23802
rect 30208 21434 30236 28086
rect 30300 25362 30328 28494
rect 30484 28218 30512 29990
rect 30564 29776 30616 29782
rect 30564 29718 30616 29724
rect 30576 29510 30604 29718
rect 30760 29617 30788 30194
rect 30746 29608 30802 29617
rect 30746 29543 30802 29552
rect 30564 29504 30616 29510
rect 30564 29446 30616 29452
rect 30656 29504 30708 29510
rect 30656 29446 30708 29452
rect 30564 29164 30616 29170
rect 30564 29106 30616 29112
rect 30472 28212 30524 28218
rect 30472 28154 30524 28160
rect 30380 28144 30432 28150
rect 30380 28086 30432 28092
rect 30392 26586 30420 28086
rect 30472 27600 30524 27606
rect 30472 27542 30524 27548
rect 30380 26580 30432 26586
rect 30380 26522 30432 26528
rect 30378 25664 30434 25673
rect 30378 25599 30434 25608
rect 30288 25356 30340 25362
rect 30288 25298 30340 25304
rect 30300 23730 30328 25298
rect 30392 24993 30420 25599
rect 30378 24984 30434 24993
rect 30378 24919 30434 24928
rect 30288 23724 30340 23730
rect 30288 23666 30340 23672
rect 30208 21406 30328 21434
rect 30196 21344 30248 21350
rect 30196 21286 30248 21292
rect 30208 21010 30236 21286
rect 30196 21004 30248 21010
rect 30196 20946 30248 20952
rect 30196 20528 30248 20534
rect 30196 20470 30248 20476
rect 30208 19718 30236 20470
rect 30300 20346 30328 21406
rect 30484 21350 30512 27542
rect 30576 22166 30604 29106
rect 30564 22160 30616 22166
rect 30564 22102 30616 22108
rect 30564 21548 30616 21554
rect 30564 21490 30616 21496
rect 30472 21344 30524 21350
rect 30472 21286 30524 21292
rect 30576 21146 30604 21490
rect 30564 21140 30616 21146
rect 30564 21082 30616 21088
rect 30300 20318 30420 20346
rect 30288 20256 30340 20262
rect 30288 20198 30340 20204
rect 30300 19990 30328 20198
rect 30288 19984 30340 19990
rect 30288 19926 30340 19932
rect 30392 19836 30420 20318
rect 30564 20052 30616 20058
rect 30564 19994 30616 20000
rect 30300 19808 30420 19836
rect 30196 19712 30248 19718
rect 30196 19654 30248 19660
rect 30104 18964 30156 18970
rect 30104 18906 30156 18912
rect 30300 17678 30328 19808
rect 30472 19780 30524 19786
rect 30472 19722 30524 19728
rect 30288 17672 30340 17678
rect 30288 17614 30340 17620
rect 30194 17368 30250 17377
rect 30194 17303 30250 17312
rect 30208 17066 30236 17303
rect 30300 17134 30328 17614
rect 30288 17128 30340 17134
rect 30288 17070 30340 17076
rect 30196 17060 30248 17066
rect 30196 17002 30248 17008
rect 30104 16040 30156 16046
rect 30104 15982 30156 15988
rect 30116 15910 30144 15982
rect 30104 15904 30156 15910
rect 30104 15846 30156 15852
rect 30288 14340 30340 14346
rect 30288 14282 30340 14288
rect 30300 13802 30328 14282
rect 30484 14278 30512 19722
rect 30576 19689 30604 19994
rect 30562 19680 30618 19689
rect 30562 19615 30618 19624
rect 30668 18698 30696 29446
rect 30746 29064 30802 29073
rect 30746 28999 30802 29008
rect 30760 28558 30788 28999
rect 30748 28552 30800 28558
rect 30748 28494 30800 28500
rect 30748 26376 30800 26382
rect 30748 26318 30800 26324
rect 30760 25673 30788 26318
rect 30746 25664 30802 25673
rect 30746 25599 30802 25608
rect 30748 24676 30800 24682
rect 30748 24618 30800 24624
rect 30760 24410 30788 24618
rect 30748 24404 30800 24410
rect 30748 24346 30800 24352
rect 30746 24168 30802 24177
rect 30746 24103 30802 24112
rect 30760 23730 30788 24103
rect 30852 23769 30880 31198
rect 30944 29753 30972 31826
rect 31024 31816 31076 31822
rect 31024 31758 31076 31764
rect 31484 31816 31536 31822
rect 31484 31758 31536 31764
rect 30930 29744 30986 29753
rect 30930 29679 30986 29688
rect 30944 29170 30972 29679
rect 30932 29164 30984 29170
rect 30932 29106 30984 29112
rect 30932 27396 30984 27402
rect 30932 27338 30984 27344
rect 30944 26353 30972 27338
rect 31036 26790 31064 31758
rect 31496 31657 31524 31758
rect 31482 31648 31538 31657
rect 31482 31583 31538 31592
rect 31496 31346 31524 31583
rect 31116 31340 31168 31346
rect 31116 31282 31168 31288
rect 31484 31340 31536 31346
rect 31484 31282 31536 31288
rect 31128 30870 31156 31282
rect 31116 30864 31168 30870
rect 31116 30806 31168 30812
rect 31116 30592 31168 30598
rect 31116 30534 31168 30540
rect 31128 30122 31156 30534
rect 31668 30320 31720 30326
rect 31666 30288 31668 30297
rect 31852 30320 31904 30326
rect 31720 30288 31722 30297
rect 31484 30252 31536 30258
rect 31852 30262 31904 30268
rect 31666 30223 31722 30232
rect 31760 30252 31812 30258
rect 31484 30194 31536 30200
rect 31760 30194 31812 30200
rect 31116 30116 31168 30122
rect 31116 30058 31168 30064
rect 31390 29744 31446 29753
rect 31390 29679 31392 29688
rect 31444 29679 31446 29688
rect 31392 29650 31444 29656
rect 31116 29640 31168 29646
rect 31114 29608 31116 29617
rect 31168 29608 31170 29617
rect 31114 29543 31170 29552
rect 31300 29232 31352 29238
rect 31206 29200 31262 29209
rect 31116 29164 31168 29170
rect 31300 29174 31352 29180
rect 31206 29135 31262 29144
rect 31116 29106 31168 29112
rect 31128 28762 31156 29106
rect 31220 29102 31248 29135
rect 31208 29096 31260 29102
rect 31208 29038 31260 29044
rect 31116 28756 31168 28762
rect 31116 28698 31168 28704
rect 31312 28694 31340 29174
rect 31300 28688 31352 28694
rect 31300 28630 31352 28636
rect 31404 28490 31432 29650
rect 31496 29073 31524 30194
rect 31574 30152 31630 30161
rect 31574 30087 31630 30096
rect 31588 29628 31616 30087
rect 31668 29844 31720 29850
rect 31772 29832 31800 30194
rect 31864 29850 31892 30262
rect 32140 30122 32168 32234
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34428 32020 34480 32026
rect 34428 31962 34480 31968
rect 32772 31884 32824 31890
rect 32772 31826 32824 31832
rect 32784 31362 32812 31826
rect 33324 31748 33376 31754
rect 33324 31690 33376 31696
rect 32784 31346 32904 31362
rect 32784 31340 32916 31346
rect 32784 31334 32864 31340
rect 32220 30932 32272 30938
rect 32220 30874 32272 30880
rect 32128 30116 32180 30122
rect 32128 30058 32180 30064
rect 31944 30048 31996 30054
rect 31944 29990 31996 29996
rect 31720 29804 31800 29832
rect 31852 29844 31904 29850
rect 31668 29786 31720 29792
rect 31852 29786 31904 29792
rect 31668 29640 31720 29646
rect 31588 29600 31668 29628
rect 31720 29600 31800 29628
rect 31668 29582 31720 29588
rect 31666 29336 31722 29345
rect 31666 29271 31722 29280
rect 31482 29064 31538 29073
rect 31482 28999 31538 29008
rect 31576 29028 31628 29034
rect 31576 28970 31628 28976
rect 31392 28484 31444 28490
rect 31220 28444 31392 28472
rect 31024 26784 31076 26790
rect 31024 26726 31076 26732
rect 31022 26480 31078 26489
rect 31022 26415 31078 26424
rect 30930 26344 30986 26353
rect 31036 26314 31064 26415
rect 30930 26279 30986 26288
rect 31024 26308 31076 26314
rect 31024 26250 31076 26256
rect 30932 26240 30984 26246
rect 30932 26182 30984 26188
rect 30944 25294 30972 26182
rect 31116 25492 31168 25498
rect 31116 25434 31168 25440
rect 30932 25288 30984 25294
rect 30932 25230 30984 25236
rect 31128 24818 31156 25434
rect 31116 24812 31168 24818
rect 31116 24754 31168 24760
rect 31024 24676 31076 24682
rect 31024 24618 31076 24624
rect 30932 24268 30984 24274
rect 30932 24210 30984 24216
rect 30838 23760 30894 23769
rect 30748 23724 30800 23730
rect 30838 23695 30894 23704
rect 30748 23666 30800 23672
rect 30944 23526 30972 24210
rect 30932 23520 30984 23526
rect 30932 23462 30984 23468
rect 31036 23322 31064 24618
rect 31024 23316 31076 23322
rect 31024 23258 31076 23264
rect 31024 23044 31076 23050
rect 31024 22986 31076 22992
rect 31036 22642 31064 22986
rect 31024 22636 31076 22642
rect 31024 22578 31076 22584
rect 30932 22568 30984 22574
rect 30932 22510 30984 22516
rect 30944 22438 30972 22510
rect 30932 22432 30984 22438
rect 30932 22374 30984 22380
rect 31128 22250 31156 24754
rect 31220 23254 31248 28444
rect 31392 28426 31444 28432
rect 31484 27328 31536 27334
rect 31484 27270 31536 27276
rect 31496 27062 31524 27270
rect 31484 27056 31536 27062
rect 31484 26998 31536 27004
rect 31392 26784 31444 26790
rect 31392 26726 31444 26732
rect 31300 26580 31352 26586
rect 31300 26522 31352 26528
rect 31208 23248 31260 23254
rect 31208 23190 31260 23196
rect 31312 23168 31340 26522
rect 31404 25430 31432 26726
rect 31484 25832 31536 25838
rect 31484 25774 31536 25780
rect 31392 25424 31444 25430
rect 31392 25366 31444 25372
rect 31496 25294 31524 25774
rect 31484 25288 31536 25294
rect 31484 25230 31536 25236
rect 31392 25220 31444 25226
rect 31392 25162 31444 25168
rect 31404 23338 31432 25162
rect 31482 25120 31538 25129
rect 31482 25055 31538 25064
rect 31496 23730 31524 25055
rect 31484 23724 31536 23730
rect 31484 23666 31536 23672
rect 31588 23526 31616 28970
rect 31680 28762 31708 29271
rect 31772 29073 31800 29600
rect 31956 29306 31984 29990
rect 32036 29776 32088 29782
rect 32036 29718 32088 29724
rect 32048 29510 32076 29718
rect 32128 29640 32180 29646
rect 32128 29582 32180 29588
rect 32036 29504 32088 29510
rect 32036 29446 32088 29452
rect 31944 29300 31996 29306
rect 31944 29242 31996 29248
rect 31758 29064 31814 29073
rect 31758 28999 31814 29008
rect 31668 28756 31720 28762
rect 31668 28698 31720 28704
rect 31668 27600 31720 27606
rect 31772 27588 31800 28999
rect 31720 27560 31800 27588
rect 31668 27542 31720 27548
rect 31956 27520 31984 29242
rect 32048 27674 32076 29446
rect 32140 29209 32168 29582
rect 32126 29200 32182 29209
rect 32126 29135 32182 29144
rect 32036 27668 32088 27674
rect 32036 27610 32088 27616
rect 31772 27492 31984 27520
rect 31668 27464 31720 27470
rect 31668 27406 31720 27412
rect 31680 26353 31708 27406
rect 31772 26790 31800 27492
rect 32128 27464 32180 27470
rect 32048 27424 32128 27452
rect 32048 27384 32076 27424
rect 32128 27406 32180 27412
rect 31864 27356 32076 27384
rect 31760 26784 31812 26790
rect 31760 26726 31812 26732
rect 31864 26382 31892 27356
rect 32128 27328 32180 27334
rect 32126 27296 32128 27305
rect 32180 27296 32182 27305
rect 32126 27231 32182 27240
rect 32128 26988 32180 26994
rect 32128 26930 32180 26936
rect 32036 26920 32088 26926
rect 32036 26862 32088 26868
rect 32048 26586 32076 26862
rect 32036 26580 32088 26586
rect 32036 26522 32088 26528
rect 31944 26444 31996 26450
rect 31944 26386 31996 26392
rect 31852 26376 31904 26382
rect 31666 26344 31722 26353
rect 31852 26318 31904 26324
rect 31666 26279 31722 26288
rect 31760 26308 31812 26314
rect 31680 24818 31708 26279
rect 31760 26250 31812 26256
rect 31772 25362 31800 26250
rect 31956 25974 31984 26386
rect 32036 26308 32088 26314
rect 32036 26250 32088 26256
rect 32048 26042 32076 26250
rect 32036 26036 32088 26042
rect 32036 25978 32088 25984
rect 31944 25968 31996 25974
rect 31944 25910 31996 25916
rect 32036 25832 32088 25838
rect 32036 25774 32088 25780
rect 31944 25764 31996 25770
rect 31944 25706 31996 25712
rect 31760 25356 31812 25362
rect 31760 25298 31812 25304
rect 31772 24954 31800 25298
rect 31850 25120 31906 25129
rect 31850 25055 31906 25064
rect 31760 24948 31812 24954
rect 31760 24890 31812 24896
rect 31668 24812 31720 24818
rect 31668 24754 31720 24760
rect 31666 24576 31722 24585
rect 31666 24511 31722 24520
rect 31680 24274 31708 24511
rect 31760 24404 31812 24410
rect 31760 24346 31812 24352
rect 31668 24268 31720 24274
rect 31668 24210 31720 24216
rect 31680 24177 31708 24210
rect 31666 24168 31722 24177
rect 31666 24103 31722 24112
rect 31666 23896 31722 23905
rect 31666 23831 31722 23840
rect 31576 23520 31628 23526
rect 31576 23462 31628 23468
rect 31404 23310 31616 23338
rect 31312 23140 31524 23168
rect 31208 23112 31260 23118
rect 31208 23054 31260 23060
rect 31220 22642 31248 23054
rect 31392 23044 31444 23050
rect 31392 22986 31444 22992
rect 31208 22636 31260 22642
rect 31208 22578 31260 22584
rect 31300 22636 31352 22642
rect 31300 22578 31352 22584
rect 30944 22222 31156 22250
rect 30748 21548 30800 21554
rect 30748 21490 30800 21496
rect 30840 21548 30892 21554
rect 30840 21490 30892 21496
rect 30760 18766 30788 21490
rect 30852 20942 30880 21490
rect 30944 21486 30972 22222
rect 31220 22166 31248 22578
rect 31312 22438 31340 22578
rect 31404 22438 31432 22986
rect 31496 22710 31524 23140
rect 31484 22704 31536 22710
rect 31484 22646 31536 22652
rect 31496 22438 31524 22646
rect 31300 22432 31352 22438
rect 31300 22374 31352 22380
rect 31392 22432 31444 22438
rect 31392 22374 31444 22380
rect 31484 22432 31536 22438
rect 31484 22374 31536 22380
rect 31116 22160 31168 22166
rect 31116 22102 31168 22108
rect 31208 22160 31260 22166
rect 31208 22102 31260 22108
rect 31024 22092 31076 22098
rect 31024 22034 31076 22040
rect 31036 21690 31064 22034
rect 31024 21684 31076 21690
rect 31024 21626 31076 21632
rect 30932 21480 30984 21486
rect 30932 21422 30984 21428
rect 31036 21350 31064 21626
rect 31024 21344 31076 21350
rect 31024 21286 31076 21292
rect 30840 20936 30892 20942
rect 30840 20878 30892 20884
rect 31024 20800 31076 20806
rect 31024 20742 31076 20748
rect 30930 20632 30986 20641
rect 30930 20567 30986 20576
rect 30840 20256 30892 20262
rect 30840 20198 30892 20204
rect 30748 18760 30800 18766
rect 30748 18702 30800 18708
rect 30656 18692 30708 18698
rect 30656 18634 30708 18640
rect 30760 18426 30788 18702
rect 30748 18420 30800 18426
rect 30748 18362 30800 18368
rect 30852 16658 30880 20198
rect 30944 19417 30972 20567
rect 30930 19408 30986 19417
rect 30930 19343 30986 19352
rect 30840 16652 30892 16658
rect 30840 16594 30892 16600
rect 30852 16250 30880 16594
rect 30840 16244 30892 16250
rect 30840 16186 30892 16192
rect 30748 16176 30800 16182
rect 30748 16118 30800 16124
rect 30760 15366 30788 16118
rect 30748 15360 30800 15366
rect 30748 15302 30800 15308
rect 30656 14952 30708 14958
rect 30654 14920 30656 14929
rect 30708 14920 30710 14929
rect 30654 14855 30710 14864
rect 30760 14396 30788 15302
rect 30838 15192 30894 15201
rect 30838 15127 30894 15136
rect 30852 15026 30880 15127
rect 30840 15020 30892 15026
rect 30840 14962 30892 14968
rect 30944 14822 30972 19343
rect 31036 18834 31064 20742
rect 31024 18828 31076 18834
rect 31024 18770 31076 18776
rect 31022 18456 31078 18465
rect 31022 18391 31078 18400
rect 31036 17542 31064 18391
rect 31128 17678 31156 22102
rect 31208 21548 31260 21554
rect 31208 21490 31260 21496
rect 31220 18952 31248 21490
rect 31312 19378 31340 22374
rect 31404 20641 31432 22374
rect 31484 22160 31536 22166
rect 31484 22102 31536 22108
rect 31390 20632 31446 20641
rect 31390 20567 31446 20576
rect 31392 20052 31444 20058
rect 31392 19994 31444 20000
rect 31404 19553 31432 19994
rect 31390 19544 31446 19553
rect 31390 19479 31446 19488
rect 31300 19372 31352 19378
rect 31300 19314 31352 19320
rect 31496 19174 31524 22102
rect 31588 21554 31616 23310
rect 31576 21548 31628 21554
rect 31576 21490 31628 21496
rect 31574 20632 31630 20641
rect 31574 20567 31630 20576
rect 31588 20369 31616 20567
rect 31574 20360 31630 20369
rect 31574 20295 31630 20304
rect 31680 20262 31708 23831
rect 31772 22817 31800 24346
rect 31864 24274 31892 25055
rect 31956 24857 31984 25706
rect 32048 25498 32076 25774
rect 32036 25492 32088 25498
rect 32036 25434 32088 25440
rect 31942 24848 31998 24857
rect 31942 24783 31998 24792
rect 31944 24744 31996 24750
rect 31944 24686 31996 24692
rect 31956 24410 31984 24686
rect 32036 24608 32088 24614
rect 32036 24550 32088 24556
rect 31944 24404 31996 24410
rect 31944 24346 31996 24352
rect 31852 24268 31904 24274
rect 31852 24210 31904 24216
rect 31942 24168 31998 24177
rect 31942 24103 31998 24112
rect 31852 23860 31904 23866
rect 31852 23802 31904 23808
rect 31864 23594 31892 23802
rect 31956 23633 31984 24103
rect 31942 23624 31998 23633
rect 31852 23588 31904 23594
rect 31942 23559 31998 23568
rect 31852 23530 31904 23536
rect 31944 23520 31996 23526
rect 31944 23462 31996 23468
rect 31852 22976 31904 22982
rect 31852 22918 31904 22924
rect 31758 22808 31814 22817
rect 31864 22778 31892 22918
rect 31758 22743 31814 22752
rect 31852 22772 31904 22778
rect 31852 22714 31904 22720
rect 31956 22681 31984 23462
rect 31942 22672 31998 22681
rect 31942 22607 31998 22616
rect 32048 22556 32076 24550
rect 32140 24342 32168 26930
rect 32232 25378 32260 30874
rect 32784 30598 32812 31334
rect 32864 31282 32916 31288
rect 33140 31340 33192 31346
rect 33140 31282 33192 31288
rect 32862 31240 32918 31249
rect 32862 31175 32918 31184
rect 32956 31204 33008 31210
rect 32876 31142 32904 31175
rect 32956 31146 33008 31152
rect 32864 31136 32916 31142
rect 32864 31078 32916 31084
rect 32312 30592 32364 30598
rect 32312 30534 32364 30540
rect 32772 30592 32824 30598
rect 32772 30534 32824 30540
rect 32324 26625 32352 30534
rect 32404 30252 32456 30258
rect 32680 30252 32732 30258
rect 32456 30212 32536 30240
rect 32404 30194 32456 30200
rect 32404 29776 32456 29782
rect 32404 29718 32456 29724
rect 32416 29617 32444 29718
rect 32402 29608 32458 29617
rect 32508 29578 32536 30212
rect 32680 30194 32732 30200
rect 32586 30016 32642 30025
rect 32586 29951 32642 29960
rect 32402 29543 32458 29552
rect 32496 29572 32548 29578
rect 32496 29514 32548 29520
rect 32404 27532 32456 27538
rect 32404 27474 32456 27480
rect 32310 26616 32366 26625
rect 32310 26551 32366 26560
rect 32324 26314 32352 26551
rect 32312 26308 32364 26314
rect 32312 26250 32364 26256
rect 32310 26208 32366 26217
rect 32310 26143 32366 26152
rect 32324 25702 32352 26143
rect 32312 25696 32364 25702
rect 32312 25638 32364 25644
rect 32232 25350 32352 25378
rect 32220 25288 32272 25294
rect 32220 25230 32272 25236
rect 32232 24721 32260 25230
rect 32324 24954 32352 25350
rect 32312 24948 32364 24954
rect 32312 24890 32364 24896
rect 32218 24712 32274 24721
rect 32218 24647 32274 24656
rect 32312 24676 32364 24682
rect 32232 24342 32260 24647
rect 32312 24618 32364 24624
rect 32324 24585 32352 24618
rect 32310 24576 32366 24585
rect 32310 24511 32366 24520
rect 32128 24336 32180 24342
rect 32128 24278 32180 24284
rect 32220 24336 32272 24342
rect 32220 24278 32272 24284
rect 32310 24304 32366 24313
rect 32310 24239 32366 24248
rect 32324 24206 32352 24239
rect 32312 24200 32364 24206
rect 32218 24168 32274 24177
rect 32312 24142 32364 24148
rect 32218 24103 32274 24112
rect 32232 23662 32260 24103
rect 32312 23860 32364 23866
rect 32312 23802 32364 23808
rect 32220 23656 32272 23662
rect 32220 23598 32272 23604
rect 32128 22976 32180 22982
rect 32128 22918 32180 22924
rect 31956 22528 32076 22556
rect 31852 20324 31904 20330
rect 31852 20266 31904 20272
rect 31668 20256 31720 20262
rect 31668 20198 31720 20204
rect 31576 19916 31628 19922
rect 31576 19858 31628 19864
rect 31392 19168 31444 19174
rect 31484 19168 31536 19174
rect 31392 19110 31444 19116
rect 31482 19136 31484 19145
rect 31536 19136 31538 19145
rect 31220 18924 31340 18952
rect 31206 18864 31262 18873
rect 31206 18799 31262 18808
rect 31220 18290 31248 18799
rect 31208 18284 31260 18290
rect 31208 18226 31260 18232
rect 31208 17740 31260 17746
rect 31208 17682 31260 17688
rect 31116 17672 31168 17678
rect 31116 17614 31168 17620
rect 31024 17536 31076 17542
rect 31024 17478 31076 17484
rect 31220 15366 31248 17682
rect 31312 16590 31340 18924
rect 31404 18290 31432 19110
rect 31482 19071 31538 19080
rect 31484 18692 31536 18698
rect 31484 18634 31536 18640
rect 31392 18284 31444 18290
rect 31392 18226 31444 18232
rect 31404 17882 31432 18226
rect 31392 17876 31444 17882
rect 31392 17818 31444 17824
rect 31392 17672 31444 17678
rect 31392 17614 31444 17620
rect 31404 17202 31432 17614
rect 31392 17196 31444 17202
rect 31392 17138 31444 17144
rect 31496 17066 31524 18634
rect 31484 17060 31536 17066
rect 31484 17002 31536 17008
rect 31392 16720 31444 16726
rect 31392 16662 31444 16668
rect 31300 16584 31352 16590
rect 31300 16526 31352 16532
rect 31404 16425 31432 16662
rect 31390 16416 31446 16425
rect 31390 16351 31446 16360
rect 31208 15360 31260 15366
rect 31208 15302 31260 15308
rect 31300 15156 31352 15162
rect 31300 15098 31352 15104
rect 31022 15056 31078 15065
rect 31022 14991 31078 15000
rect 31116 15020 31168 15026
rect 31036 14958 31064 14991
rect 31116 14962 31168 14968
rect 31208 15020 31260 15026
rect 31208 14962 31260 14968
rect 31024 14952 31076 14958
rect 31024 14894 31076 14900
rect 30932 14816 30984 14822
rect 30932 14758 30984 14764
rect 30930 14648 30986 14657
rect 31128 14618 31156 14962
rect 31220 14890 31248 14962
rect 31312 14890 31340 15098
rect 31392 14952 31444 14958
rect 31392 14894 31444 14900
rect 31208 14884 31260 14890
rect 31208 14826 31260 14832
rect 31300 14884 31352 14890
rect 31300 14826 31352 14832
rect 30930 14583 30932 14592
rect 30984 14583 30986 14592
rect 31116 14612 31168 14618
rect 30932 14554 30984 14560
rect 31116 14554 31168 14560
rect 30840 14408 30892 14414
rect 30760 14368 30840 14396
rect 30840 14350 30892 14356
rect 30472 14272 30524 14278
rect 30472 14214 30524 14220
rect 30288 13796 30340 13802
rect 30288 13738 30340 13744
rect 30930 13696 30986 13705
rect 30930 13631 30986 13640
rect 29826 13495 29882 13504
rect 30012 13524 30064 13530
rect 30012 13466 30064 13472
rect 30944 13258 30972 13631
rect 31022 13560 31078 13569
rect 31022 13495 31078 13504
rect 31036 13394 31064 13495
rect 31024 13388 31076 13394
rect 31024 13330 31076 13336
rect 30932 13252 30984 13258
rect 30932 13194 30984 13200
rect 29460 12912 29512 12918
rect 29460 12854 29512 12860
rect 29736 12912 29788 12918
rect 29736 12854 29788 12860
rect 30288 12912 30340 12918
rect 30288 12854 30340 12860
rect 30300 12442 30328 12854
rect 30944 12850 30972 13194
rect 30932 12844 30984 12850
rect 30932 12786 30984 12792
rect 31036 12646 31064 13330
rect 31404 13326 31432 14894
rect 31392 13320 31444 13326
rect 31392 13262 31444 13268
rect 31116 13252 31168 13258
rect 31116 13194 31168 13200
rect 31128 12918 31156 13194
rect 31496 12986 31524 17002
rect 31588 15162 31616 19858
rect 31864 19242 31892 20266
rect 31668 19236 31720 19242
rect 31668 19178 31720 19184
rect 31852 19236 31904 19242
rect 31852 19178 31904 19184
rect 31680 18601 31708 19178
rect 31864 18970 31892 19178
rect 31852 18964 31904 18970
rect 31852 18906 31904 18912
rect 31760 18828 31812 18834
rect 31760 18770 31812 18776
rect 31666 18592 31722 18601
rect 31666 18527 31722 18536
rect 31668 18284 31720 18290
rect 31668 18226 31720 18232
rect 31680 18086 31708 18226
rect 31668 18080 31720 18086
rect 31668 18022 31720 18028
rect 31772 17746 31800 18770
rect 31956 18601 31984 22528
rect 32036 22432 32088 22438
rect 32036 22374 32088 22380
rect 32048 21894 32076 22374
rect 32036 21888 32088 21894
rect 32036 21830 32088 21836
rect 32036 21684 32088 21690
rect 32036 21626 32088 21632
rect 31942 18592 31998 18601
rect 31864 18550 31942 18578
rect 31760 17740 31812 17746
rect 31760 17682 31812 17688
rect 31668 17604 31720 17610
rect 31668 17546 31720 17552
rect 31680 17338 31708 17546
rect 31668 17332 31720 17338
rect 31668 17274 31720 17280
rect 31668 16992 31720 16998
rect 31668 16934 31720 16940
rect 31680 16794 31708 16934
rect 31668 16788 31720 16794
rect 31668 16730 31720 16736
rect 31760 16652 31812 16658
rect 31760 16594 31812 16600
rect 31772 15638 31800 16594
rect 31864 15706 31892 18550
rect 31942 18527 31998 18536
rect 31942 17912 31998 17921
rect 31942 17847 31998 17856
rect 31956 17678 31984 17847
rect 31944 17672 31996 17678
rect 31944 17614 31996 17620
rect 32048 17626 32076 21626
rect 32140 19514 32168 22918
rect 32232 21865 32260 23598
rect 32218 21856 32274 21865
rect 32218 21791 32274 21800
rect 32324 21690 32352 23802
rect 32416 23662 32444 27474
rect 32508 26994 32536 29514
rect 32600 27538 32628 29951
rect 32692 29646 32720 30194
rect 32680 29640 32732 29646
rect 32680 29582 32732 29588
rect 32862 29472 32918 29481
rect 32862 29407 32918 29416
rect 32876 28490 32904 29407
rect 32864 28484 32916 28490
rect 32864 28426 32916 28432
rect 32680 28416 32732 28422
rect 32678 28384 32680 28393
rect 32732 28384 32734 28393
rect 32678 28319 32734 28328
rect 32772 28008 32824 28014
rect 32772 27950 32824 27956
rect 32784 27713 32812 27950
rect 32770 27704 32826 27713
rect 32876 27674 32904 28426
rect 32770 27639 32826 27648
rect 32864 27668 32916 27674
rect 32864 27610 32916 27616
rect 32588 27532 32640 27538
rect 32588 27474 32640 27480
rect 32588 27328 32640 27334
rect 32588 27270 32640 27276
rect 32864 27328 32916 27334
rect 32864 27270 32916 27276
rect 32600 26994 32628 27270
rect 32496 26988 32548 26994
rect 32496 26930 32548 26936
rect 32588 26988 32640 26994
rect 32588 26930 32640 26936
rect 32508 26330 32536 26930
rect 32770 26888 32826 26897
rect 32770 26823 32826 26832
rect 32588 26784 32640 26790
rect 32588 26726 32640 26732
rect 32600 26518 32628 26726
rect 32784 26586 32812 26823
rect 32772 26580 32824 26586
rect 32772 26522 32824 26528
rect 32588 26512 32640 26518
rect 32588 26454 32640 26460
rect 32680 26376 32732 26382
rect 32508 26302 32628 26330
rect 32680 26318 32732 26324
rect 32496 24812 32548 24818
rect 32496 24754 32548 24760
rect 32508 24274 32536 24754
rect 32496 24268 32548 24274
rect 32496 24210 32548 24216
rect 32600 24154 32628 26302
rect 32508 24126 32628 24154
rect 32404 23656 32456 23662
rect 32404 23598 32456 23604
rect 32508 22094 32536 24126
rect 32588 23724 32640 23730
rect 32588 23666 32640 23672
rect 32600 23254 32628 23666
rect 32588 23248 32640 23254
rect 32588 23190 32640 23196
rect 32600 22545 32628 23190
rect 32586 22536 32642 22545
rect 32586 22471 32642 22480
rect 32692 22273 32720 26318
rect 32772 26036 32824 26042
rect 32772 25978 32824 25984
rect 32784 25226 32812 25978
rect 32876 25906 32904 27270
rect 32864 25900 32916 25906
rect 32864 25842 32916 25848
rect 32772 25220 32824 25226
rect 32772 25162 32824 25168
rect 32772 24948 32824 24954
rect 32772 24890 32824 24896
rect 32784 24682 32812 24890
rect 32968 24818 32996 31146
rect 33152 30954 33180 31282
rect 33060 30938 33180 30954
rect 33048 30932 33180 30938
rect 33100 30926 33180 30932
rect 33048 30874 33100 30880
rect 33140 30864 33192 30870
rect 33140 30806 33192 30812
rect 33152 30666 33180 30806
rect 33336 30734 33364 31690
rect 33784 31476 33836 31482
rect 33784 31418 33836 31424
rect 33416 31340 33468 31346
rect 33416 31282 33468 31288
rect 33428 31142 33456 31282
rect 33600 31204 33652 31210
rect 33600 31146 33652 31152
rect 33692 31204 33744 31210
rect 33692 31146 33744 31152
rect 33416 31136 33468 31142
rect 33416 31078 33468 31084
rect 33232 30728 33284 30734
rect 33232 30670 33284 30676
rect 33324 30728 33376 30734
rect 33428 30705 33456 31078
rect 33508 30932 33560 30938
rect 33508 30874 33560 30880
rect 33324 30670 33376 30676
rect 33414 30696 33470 30705
rect 33140 30660 33192 30666
rect 33140 30602 33192 30608
rect 33138 28792 33194 28801
rect 33138 28727 33194 28736
rect 33152 28694 33180 28727
rect 33140 28688 33192 28694
rect 33140 28630 33192 28636
rect 33140 27872 33192 27878
rect 33140 27814 33192 27820
rect 33048 27532 33100 27538
rect 33048 27474 33100 27480
rect 33060 27334 33088 27474
rect 33048 27328 33100 27334
rect 33048 27270 33100 27276
rect 32956 24812 33008 24818
rect 32956 24754 33008 24760
rect 32772 24676 32824 24682
rect 32772 24618 32824 24624
rect 32784 23497 32812 24618
rect 32956 24608 33008 24614
rect 32956 24550 33008 24556
rect 32968 23497 32996 24550
rect 33060 23526 33088 27270
rect 33152 26790 33180 27814
rect 33244 27470 33272 30670
rect 33414 30631 33470 30640
rect 33520 30598 33548 30874
rect 33508 30592 33560 30598
rect 33508 30534 33560 30540
rect 33416 30320 33468 30326
rect 33416 30262 33468 30268
rect 33324 28688 33376 28694
rect 33324 28630 33376 28636
rect 33336 27614 33364 28630
rect 33428 27985 33456 30262
rect 33520 28490 33548 30534
rect 33508 28484 33560 28490
rect 33508 28426 33560 28432
rect 33414 27976 33470 27985
rect 33414 27911 33470 27920
rect 33336 27586 33548 27614
rect 33324 27532 33376 27538
rect 33324 27474 33376 27480
rect 33232 27464 33284 27470
rect 33232 27406 33284 27412
rect 33140 26784 33192 26790
rect 33140 26726 33192 26732
rect 33152 26586 33180 26726
rect 33140 26580 33192 26586
rect 33140 26522 33192 26528
rect 33244 26466 33272 27406
rect 33152 26450 33272 26466
rect 33140 26444 33272 26450
rect 33192 26438 33272 26444
rect 33140 26386 33192 26392
rect 33232 26376 33284 26382
rect 33232 26318 33284 26324
rect 33140 25832 33192 25838
rect 33140 25774 33192 25780
rect 33048 23520 33100 23526
rect 32770 23488 32826 23497
rect 32770 23423 32826 23432
rect 32954 23488 33010 23497
rect 33048 23462 33100 23468
rect 32954 23423 33010 23432
rect 32864 23316 32916 23322
rect 32864 23258 32916 23264
rect 32772 23180 32824 23186
rect 32772 23122 32824 23128
rect 32678 22264 32734 22273
rect 32678 22199 32734 22208
rect 32508 22066 32628 22094
rect 32496 21956 32548 21962
rect 32496 21898 32548 21904
rect 32312 21684 32364 21690
rect 32312 21626 32364 21632
rect 32312 21548 32364 21554
rect 32312 21490 32364 21496
rect 32324 21457 32352 21490
rect 32404 21480 32456 21486
rect 32310 21448 32366 21457
rect 32404 21422 32456 21428
rect 32310 21383 32366 21392
rect 32312 21344 32364 21350
rect 32312 21286 32364 21292
rect 32218 20768 32274 20777
rect 32218 20703 32274 20712
rect 32232 19922 32260 20703
rect 32220 19916 32272 19922
rect 32220 19858 32272 19864
rect 32232 19786 32260 19858
rect 32220 19780 32272 19786
rect 32220 19722 32272 19728
rect 32324 19553 32352 21286
rect 32416 20534 32444 21422
rect 32404 20528 32456 20534
rect 32404 20470 32456 20476
rect 32310 19544 32366 19553
rect 32128 19508 32180 19514
rect 32310 19479 32366 19488
rect 32404 19508 32456 19514
rect 32128 19450 32180 19456
rect 32404 19450 32456 19456
rect 32220 19304 32272 19310
rect 32218 19272 32220 19281
rect 32272 19272 32274 19281
rect 32218 19207 32274 19216
rect 32128 19168 32180 19174
rect 32126 19136 32128 19145
rect 32180 19136 32182 19145
rect 32126 19071 32182 19080
rect 32312 18624 32364 18630
rect 32312 18566 32364 18572
rect 32324 18290 32352 18566
rect 32312 18284 32364 18290
rect 32312 18226 32364 18232
rect 32312 18080 32364 18086
rect 32218 18048 32274 18057
rect 32312 18022 32364 18028
rect 32218 17983 32274 17992
rect 32232 17762 32260 17983
rect 32324 17882 32352 18022
rect 32312 17876 32364 17882
rect 32312 17818 32364 17824
rect 32232 17734 32352 17762
rect 32416 17746 32444 19450
rect 32048 17598 32260 17626
rect 32128 17536 32180 17542
rect 32128 17478 32180 17484
rect 31944 17332 31996 17338
rect 31944 17274 31996 17280
rect 31956 16794 31984 17274
rect 32140 17270 32168 17478
rect 32128 17264 32180 17270
rect 32128 17206 32180 17212
rect 31944 16788 31996 16794
rect 31944 16730 31996 16736
rect 32036 16720 32088 16726
rect 32036 16662 32088 16668
rect 32048 16590 32076 16662
rect 32036 16584 32088 16590
rect 32036 16526 32088 16532
rect 31852 15700 31904 15706
rect 31852 15642 31904 15648
rect 31760 15632 31812 15638
rect 31760 15574 31812 15580
rect 32232 15434 32260 17598
rect 32324 17270 32352 17734
rect 32404 17740 32456 17746
rect 32404 17682 32456 17688
rect 32312 17264 32364 17270
rect 32312 17206 32364 17212
rect 32402 16824 32458 16833
rect 32508 16794 32536 21898
rect 32600 21729 32628 22066
rect 32586 21720 32642 21729
rect 32586 21655 32642 21664
rect 32680 20528 32732 20534
rect 32680 20470 32732 20476
rect 32692 19922 32720 20470
rect 32680 19916 32732 19922
rect 32680 19858 32732 19864
rect 32784 19802 32812 23122
rect 32876 22080 32904 23258
rect 32956 23044 33008 23050
rect 32956 22986 33008 22992
rect 32968 22778 32996 22986
rect 32956 22772 33008 22778
rect 32956 22714 33008 22720
rect 32968 22574 32996 22714
rect 32956 22568 33008 22574
rect 32956 22510 33008 22516
rect 33046 22536 33102 22545
rect 33046 22471 33102 22480
rect 33060 22234 33088 22471
rect 33048 22228 33100 22234
rect 33048 22170 33100 22176
rect 32876 22052 32996 22080
rect 32862 21992 32918 22001
rect 32862 21927 32918 21936
rect 32692 19774 32812 19802
rect 32588 18760 32640 18766
rect 32588 18702 32640 18708
rect 32600 18426 32628 18702
rect 32588 18420 32640 18426
rect 32588 18362 32640 18368
rect 32586 17912 32642 17921
rect 32586 17847 32642 17856
rect 32600 17678 32628 17847
rect 32588 17672 32640 17678
rect 32588 17614 32640 17620
rect 32600 17513 32628 17614
rect 32586 17504 32642 17513
rect 32586 17439 32642 17448
rect 32402 16759 32458 16768
rect 32496 16788 32548 16794
rect 32416 16726 32444 16759
rect 32496 16730 32548 16736
rect 32404 16720 32456 16726
rect 32404 16662 32456 16668
rect 32312 16652 32364 16658
rect 32312 16594 32364 16600
rect 32324 15910 32352 16594
rect 32402 16280 32458 16289
rect 32402 16215 32404 16224
rect 32456 16215 32458 16224
rect 32588 16244 32640 16250
rect 32404 16186 32456 16192
rect 32588 16186 32640 16192
rect 32416 16046 32444 16186
rect 32600 16153 32628 16186
rect 32586 16144 32642 16153
rect 32586 16079 32588 16088
rect 32640 16079 32642 16088
rect 32588 16050 32640 16056
rect 32404 16040 32456 16046
rect 32404 15982 32456 15988
rect 32312 15904 32364 15910
rect 32312 15846 32364 15852
rect 32588 15904 32640 15910
rect 32588 15846 32640 15852
rect 32600 15706 32628 15846
rect 32588 15700 32640 15706
rect 32588 15642 32640 15648
rect 32692 15638 32720 19774
rect 32772 19712 32824 19718
rect 32772 19654 32824 19660
rect 32784 18290 32812 19654
rect 32772 18284 32824 18290
rect 32772 18226 32824 18232
rect 32772 15904 32824 15910
rect 32772 15846 32824 15852
rect 32680 15632 32732 15638
rect 32680 15574 32732 15580
rect 32220 15428 32272 15434
rect 32220 15370 32272 15376
rect 31576 15156 31628 15162
rect 31628 15116 31708 15144
rect 31576 15098 31628 15104
rect 31574 15056 31630 15065
rect 31574 14991 31576 15000
rect 31628 14991 31630 15000
rect 31576 14962 31628 14968
rect 31576 14816 31628 14822
rect 31574 14784 31576 14793
rect 31628 14784 31630 14793
rect 31574 14719 31630 14728
rect 31576 14476 31628 14482
rect 31576 14418 31628 14424
rect 31588 13394 31616 14418
rect 31680 14006 31708 15116
rect 31760 15020 31812 15026
rect 31760 14962 31812 14968
rect 31772 14550 31800 14962
rect 31852 14816 31904 14822
rect 31852 14758 31904 14764
rect 31760 14544 31812 14550
rect 31760 14486 31812 14492
rect 31864 14346 31892 14758
rect 32692 14657 32720 15574
rect 32784 15502 32812 15846
rect 32876 15745 32904 21927
rect 32968 19786 32996 22052
rect 33048 21956 33100 21962
rect 33048 21898 33100 21904
rect 33060 21690 33088 21898
rect 33048 21684 33100 21690
rect 33048 21626 33100 21632
rect 33048 21480 33100 21486
rect 33048 21422 33100 21428
rect 33060 21350 33088 21422
rect 33048 21344 33100 21350
rect 33048 21286 33100 21292
rect 33152 19854 33180 25774
rect 33244 23798 33272 26318
rect 33336 24682 33364 27474
rect 33414 27296 33470 27305
rect 33414 27231 33470 27240
rect 33428 27130 33456 27231
rect 33416 27124 33468 27130
rect 33416 27066 33468 27072
rect 33416 26444 33468 26450
rect 33416 26386 33468 26392
rect 33428 25702 33456 26386
rect 33416 25696 33468 25702
rect 33416 25638 33468 25644
rect 33416 25492 33468 25498
rect 33416 25434 33468 25440
rect 33324 24676 33376 24682
rect 33324 24618 33376 24624
rect 33324 24404 33376 24410
rect 33324 24346 33376 24352
rect 33336 23866 33364 24346
rect 33324 23860 33376 23866
rect 33324 23802 33376 23808
rect 33232 23792 33284 23798
rect 33232 23734 33284 23740
rect 33244 23118 33272 23734
rect 33232 23112 33284 23118
rect 33232 23054 33284 23060
rect 33428 22778 33456 25434
rect 33520 23118 33548 27586
rect 33612 25702 33640 31146
rect 33704 30802 33732 31146
rect 33796 30802 33824 31418
rect 34440 30938 34468 31962
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 34612 31340 34664 31346
rect 34612 31282 34664 31288
rect 34428 30932 34480 30938
rect 34428 30874 34480 30880
rect 33692 30796 33744 30802
rect 33692 30738 33744 30744
rect 33784 30796 33836 30802
rect 33784 30738 33836 30744
rect 34520 30728 34572 30734
rect 34520 30670 34572 30676
rect 33692 30660 33744 30666
rect 33692 30602 33744 30608
rect 33784 30660 33836 30666
rect 33784 30602 33836 30608
rect 33704 30394 33732 30602
rect 33692 30388 33744 30394
rect 33692 30330 33744 30336
rect 33796 30274 33824 30602
rect 33704 30246 33824 30274
rect 33600 25696 33652 25702
rect 33600 25638 33652 25644
rect 33704 25498 33732 30246
rect 33784 30184 33836 30190
rect 33784 30126 33836 30132
rect 33692 25492 33744 25498
rect 33692 25434 33744 25440
rect 33692 25356 33744 25362
rect 33692 25298 33744 25304
rect 33600 24880 33652 24886
rect 33600 24822 33652 24828
rect 33612 24449 33640 24822
rect 33704 24818 33732 25298
rect 33692 24812 33744 24818
rect 33692 24754 33744 24760
rect 33692 24676 33744 24682
rect 33692 24618 33744 24624
rect 33598 24440 33654 24449
rect 33598 24375 33654 24384
rect 33612 23662 33640 24375
rect 33600 23656 33652 23662
rect 33600 23598 33652 23604
rect 33600 23316 33652 23322
rect 33600 23258 33652 23264
rect 33508 23112 33560 23118
rect 33508 23054 33560 23060
rect 33416 22772 33468 22778
rect 33416 22714 33468 22720
rect 33324 22704 33376 22710
rect 33324 22646 33376 22652
rect 33232 22228 33284 22234
rect 33232 22170 33284 22176
rect 33244 22001 33272 22170
rect 33230 21992 33286 22001
rect 33230 21927 33286 21936
rect 33230 21720 33286 21729
rect 33230 21655 33232 21664
rect 33284 21655 33286 21664
rect 33232 21626 33284 21632
rect 33230 21312 33286 21321
rect 33230 21247 33286 21256
rect 33140 19848 33192 19854
rect 33140 19790 33192 19796
rect 32956 19780 33008 19786
rect 32956 19722 33008 19728
rect 32968 18358 32996 19722
rect 33048 19712 33100 19718
rect 33048 19654 33100 19660
rect 32956 18352 33008 18358
rect 32956 18294 33008 18300
rect 32968 17882 32996 18294
rect 33060 18154 33088 19654
rect 33140 18216 33192 18222
rect 33140 18158 33192 18164
rect 33048 18148 33100 18154
rect 33048 18090 33100 18096
rect 32956 17876 33008 17882
rect 32956 17818 33008 17824
rect 33152 17746 33180 18158
rect 33244 17762 33272 21247
rect 33336 18222 33364 22646
rect 33416 22500 33468 22506
rect 33416 22442 33468 22448
rect 33428 21078 33456 22442
rect 33520 22234 33548 23054
rect 33508 22228 33560 22234
rect 33508 22170 33560 22176
rect 33612 22001 33640 23258
rect 33704 22030 33732 24618
rect 33796 24614 33824 30126
rect 33968 29844 34020 29850
rect 33968 29786 34020 29792
rect 33876 29164 33928 29170
rect 33876 29106 33928 29112
rect 33888 29073 33916 29106
rect 33874 29064 33930 29073
rect 33874 28999 33930 29008
rect 33876 28960 33928 28966
rect 33876 28902 33928 28908
rect 33888 28490 33916 28902
rect 33876 28484 33928 28490
rect 33876 28426 33928 28432
rect 33980 28370 34008 29786
rect 34532 29594 34560 30670
rect 34440 29566 34560 29594
rect 34440 29186 34468 29566
rect 34440 29170 34560 29186
rect 34440 29164 34572 29170
rect 34440 29158 34520 29164
rect 34520 29106 34572 29112
rect 34152 29028 34204 29034
rect 34532 28994 34560 29106
rect 34152 28970 34204 28976
rect 34164 28665 34192 28970
rect 34440 28966 34560 28994
rect 34336 28960 34388 28966
rect 34336 28902 34388 28908
rect 34348 28762 34376 28902
rect 34336 28756 34388 28762
rect 34336 28698 34388 28704
rect 34150 28656 34206 28665
rect 34060 28620 34112 28626
rect 34150 28591 34206 28600
rect 34060 28562 34112 28568
rect 33888 28342 34008 28370
rect 33888 24886 33916 28342
rect 33968 28212 34020 28218
rect 33968 28154 34020 28160
rect 33876 24880 33928 24886
rect 33876 24822 33928 24828
rect 33784 24608 33836 24614
rect 33784 24550 33836 24556
rect 33874 24576 33930 24585
rect 33874 24511 33930 24520
rect 33888 24410 33916 24511
rect 33876 24404 33928 24410
rect 33876 24346 33928 24352
rect 33980 24274 34008 28154
rect 34072 28150 34100 28562
rect 34336 28416 34388 28422
rect 34336 28358 34388 28364
rect 34060 28144 34112 28150
rect 34060 28086 34112 28092
rect 34060 28008 34112 28014
rect 34060 27950 34112 27956
rect 34072 27674 34100 27950
rect 34060 27668 34112 27674
rect 34060 27610 34112 27616
rect 34072 25242 34100 27610
rect 34348 27538 34376 28358
rect 34336 27532 34388 27538
rect 34336 27474 34388 27480
rect 34348 27334 34376 27474
rect 34440 27402 34468 28966
rect 34624 28626 34652 31282
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35992 30728 36044 30734
rect 35992 30670 36044 30676
rect 34796 30660 34848 30666
rect 34796 30602 34848 30608
rect 34702 30424 34758 30433
rect 34702 30359 34758 30368
rect 34716 29578 34744 30359
rect 34808 30054 34836 30602
rect 35348 30592 35400 30598
rect 35348 30534 35400 30540
rect 34796 30048 34848 30054
rect 34796 29990 34848 29996
rect 34704 29572 34756 29578
rect 34704 29514 34756 29520
rect 34716 29170 34744 29514
rect 34808 29306 34836 29990
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35070 29336 35126 29345
rect 34796 29300 34848 29306
rect 35070 29271 35126 29280
rect 34796 29242 34848 29248
rect 35084 29238 35112 29271
rect 35072 29232 35124 29238
rect 35072 29174 35124 29180
rect 34704 29164 34756 29170
rect 34704 29106 34756 29112
rect 34796 29096 34848 29102
rect 34702 29064 34758 29073
rect 35256 29096 35308 29102
rect 34796 29038 34848 29044
rect 34886 29064 34942 29073
rect 34702 28999 34758 29008
rect 34716 28937 34744 28999
rect 34702 28928 34758 28937
rect 34702 28863 34758 28872
rect 34612 28620 34664 28626
rect 34612 28562 34664 28568
rect 34612 28484 34664 28490
rect 34612 28426 34664 28432
rect 34518 28248 34574 28257
rect 34518 28183 34574 28192
rect 34428 27396 34480 27402
rect 34428 27338 34480 27344
rect 34336 27328 34388 27334
rect 34336 27270 34388 27276
rect 34532 27130 34560 28183
rect 34520 27124 34572 27130
rect 34520 27066 34572 27072
rect 34244 26988 34296 26994
rect 34244 26930 34296 26936
rect 34336 26988 34388 26994
rect 34336 26930 34388 26936
rect 34152 25696 34204 25702
rect 34256 25673 34284 26930
rect 34152 25638 34204 25644
rect 34242 25664 34298 25673
rect 34164 25498 34192 25638
rect 34242 25599 34298 25608
rect 34242 25528 34298 25537
rect 34152 25492 34204 25498
rect 34242 25463 34298 25472
rect 34152 25434 34204 25440
rect 34072 25214 34192 25242
rect 34060 25152 34112 25158
rect 34060 25094 34112 25100
rect 33876 24268 33928 24274
rect 33876 24210 33928 24216
rect 33968 24268 34020 24274
rect 33968 24210 34020 24216
rect 33784 23520 33836 23526
rect 33784 23462 33836 23468
rect 33796 23050 33824 23462
rect 33784 23044 33836 23050
rect 33784 22986 33836 22992
rect 33692 22024 33744 22030
rect 33598 21992 33654 22001
rect 33692 21966 33744 21972
rect 33598 21927 33654 21936
rect 33506 21720 33562 21729
rect 33506 21655 33562 21664
rect 33520 21554 33548 21655
rect 33508 21548 33560 21554
rect 33508 21490 33560 21496
rect 33704 21350 33732 21966
rect 33692 21344 33744 21350
rect 33692 21286 33744 21292
rect 33416 21072 33468 21078
rect 33416 21014 33468 21020
rect 33692 21004 33744 21010
rect 33692 20946 33744 20952
rect 33600 20596 33652 20602
rect 33600 20538 33652 20544
rect 33612 20058 33640 20538
rect 33600 20052 33652 20058
rect 33600 19994 33652 20000
rect 33416 19848 33468 19854
rect 33416 19790 33468 19796
rect 33508 19848 33560 19854
rect 33508 19790 33560 19796
rect 33324 18216 33376 18222
rect 33324 18158 33376 18164
rect 33428 17882 33456 19790
rect 33520 19446 33548 19790
rect 33508 19440 33560 19446
rect 33508 19382 33560 19388
rect 33508 19168 33560 19174
rect 33508 19110 33560 19116
rect 33416 17876 33468 17882
rect 33416 17818 33468 17824
rect 33140 17740 33192 17746
rect 33244 17734 33364 17762
rect 33140 17682 33192 17688
rect 33232 17672 33284 17678
rect 33232 17614 33284 17620
rect 33140 16992 33192 16998
rect 33140 16934 33192 16940
rect 32956 16244 33008 16250
rect 32956 16186 33008 16192
rect 32968 16153 32996 16186
rect 32954 16144 33010 16153
rect 32954 16079 33010 16088
rect 32862 15736 32918 15745
rect 32862 15671 32864 15680
rect 32916 15671 32918 15680
rect 32864 15642 32916 15648
rect 33048 15632 33100 15638
rect 33048 15574 33100 15580
rect 33060 15502 33088 15574
rect 32772 15496 32824 15502
rect 32956 15496 33008 15502
rect 32772 15438 32824 15444
rect 32862 15464 32918 15473
rect 32956 15438 33008 15444
rect 33048 15496 33100 15502
rect 33048 15438 33100 15444
rect 32862 15399 32864 15408
rect 32916 15399 32918 15408
rect 32864 15370 32916 15376
rect 32968 15162 32996 15438
rect 32956 15156 33008 15162
rect 32956 15098 33008 15104
rect 33152 15026 33180 16934
rect 33244 16590 33272 17614
rect 33336 17218 33364 17734
rect 33336 17190 33456 17218
rect 33322 17096 33378 17105
rect 33322 17031 33378 17040
rect 33232 16584 33284 16590
rect 33232 16526 33284 16532
rect 33230 16280 33286 16289
rect 33230 16215 33286 16224
rect 33244 15638 33272 16215
rect 33336 15706 33364 17031
rect 33428 16794 33456 17190
rect 33416 16788 33468 16794
rect 33416 16730 33468 16736
rect 33416 16584 33468 16590
rect 33416 16526 33468 16532
rect 33428 16425 33456 16526
rect 33414 16416 33470 16425
rect 33414 16351 33470 16360
rect 33520 15706 33548 19110
rect 33612 17610 33640 19994
rect 33600 17604 33652 17610
rect 33600 17546 33652 17552
rect 33612 15910 33640 17546
rect 33704 16182 33732 20946
rect 33796 18086 33824 22986
rect 33888 20602 33916 24210
rect 33968 23656 34020 23662
rect 33968 23598 34020 23604
rect 33980 23118 34008 23598
rect 33968 23112 34020 23118
rect 33968 23054 34020 23060
rect 33968 22772 34020 22778
rect 33968 22714 34020 22720
rect 33980 21706 34008 22714
rect 34072 21962 34100 25094
rect 34164 24954 34192 25214
rect 34152 24948 34204 24954
rect 34152 24890 34204 24896
rect 34256 24290 34284 25463
rect 34348 24410 34376 26930
rect 34520 26920 34572 26926
rect 34520 26862 34572 26868
rect 34532 26790 34560 26862
rect 34520 26784 34572 26790
rect 34520 26726 34572 26732
rect 34428 25900 34480 25906
rect 34428 25842 34480 25848
rect 34440 24993 34468 25842
rect 34520 25696 34572 25702
rect 34520 25638 34572 25644
rect 34532 25362 34560 25638
rect 34520 25356 34572 25362
rect 34520 25298 34572 25304
rect 34426 24984 34482 24993
rect 34426 24919 34482 24928
rect 34336 24404 34388 24410
rect 34336 24346 34388 24352
rect 34428 24404 34480 24410
rect 34428 24346 34480 24352
rect 34440 24290 34468 24346
rect 34256 24262 34468 24290
rect 34152 24064 34204 24070
rect 34152 24006 34204 24012
rect 34164 23662 34192 24006
rect 34152 23656 34204 23662
rect 34152 23598 34204 23604
rect 34152 23180 34204 23186
rect 34152 23122 34204 23128
rect 34164 22166 34192 23122
rect 34256 22273 34284 24262
rect 34426 24032 34482 24041
rect 34426 23967 34482 23976
rect 34440 23798 34468 23967
rect 34532 23905 34560 25298
rect 34624 24177 34652 28426
rect 34716 27878 34744 28863
rect 34704 27872 34756 27878
rect 34704 27814 34756 27820
rect 34702 27704 34758 27713
rect 34702 27639 34704 27648
rect 34756 27639 34758 27648
rect 34704 27610 34756 27616
rect 34808 26994 34836 29038
rect 35360 29084 35388 30534
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 36004 30326 36032 30670
rect 35992 30320 36044 30326
rect 35992 30262 36044 30268
rect 36004 29714 36032 30262
rect 35992 29708 36044 29714
rect 35992 29650 36044 29656
rect 36096 29646 36124 32778
rect 37464 32564 37516 32570
rect 37464 32506 37516 32512
rect 37096 32360 37148 32366
rect 37096 32302 37148 32308
rect 36360 32224 36412 32230
rect 36360 32166 36412 32172
rect 36174 31376 36230 31385
rect 36174 31311 36230 31320
rect 36188 30734 36216 31311
rect 36268 31204 36320 31210
rect 36268 31146 36320 31152
rect 36176 30728 36228 30734
rect 36176 30670 36228 30676
rect 36084 29640 36136 29646
rect 36084 29582 36136 29588
rect 35440 29504 35492 29510
rect 35440 29446 35492 29452
rect 35452 29238 35480 29446
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 35716 29300 35768 29306
rect 35716 29242 35768 29248
rect 35440 29232 35492 29238
rect 35440 29174 35492 29180
rect 35440 29096 35492 29102
rect 35360 29056 35440 29084
rect 35256 29038 35308 29044
rect 35440 29038 35492 29044
rect 34886 28999 34942 29008
rect 34900 28966 34928 28999
rect 34888 28960 34940 28966
rect 34888 28902 34940 28908
rect 35268 28914 35296 29038
rect 35624 29028 35676 29034
rect 35544 28976 35624 28994
rect 35544 28970 35676 28976
rect 35544 28966 35664 28970
rect 35268 28886 35480 28914
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35348 28756 35400 28762
rect 35348 28698 35400 28704
rect 35360 28422 35388 28698
rect 35348 28416 35400 28422
rect 35348 28358 35400 28364
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35164 27668 35216 27674
rect 35164 27610 35216 27616
rect 35176 26994 35204 27610
rect 35360 27538 35388 28358
rect 35348 27532 35400 27538
rect 35348 27474 35400 27480
rect 35452 27418 35480 28886
rect 35544 28422 35572 28966
rect 35728 28558 35756 29242
rect 35808 29232 35860 29238
rect 35808 29174 35860 29180
rect 35820 28558 35848 29174
rect 36096 28762 36124 29582
rect 36280 29102 36308 31146
rect 36268 29096 36320 29102
rect 36268 29038 36320 29044
rect 36176 29028 36228 29034
rect 36176 28970 36228 28976
rect 36084 28756 36136 28762
rect 36084 28698 36136 28704
rect 35716 28552 35768 28558
rect 35622 28520 35678 28529
rect 35716 28494 35768 28500
rect 35808 28552 35860 28558
rect 35808 28494 35860 28500
rect 35622 28455 35624 28464
rect 35676 28455 35678 28464
rect 35992 28484 36044 28490
rect 35624 28426 35676 28432
rect 35992 28426 36044 28432
rect 35532 28416 35584 28422
rect 35532 28358 35584 28364
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 35808 27940 35860 27946
rect 35808 27882 35860 27888
rect 35530 27704 35586 27713
rect 35530 27639 35532 27648
rect 35584 27639 35586 27648
rect 35532 27610 35584 27616
rect 35360 27390 35480 27418
rect 35254 27296 35310 27305
rect 35254 27231 35310 27240
rect 35268 27062 35296 27231
rect 35256 27056 35308 27062
rect 35256 26998 35308 27004
rect 34796 26988 34848 26994
rect 34796 26930 34848 26936
rect 35164 26988 35216 26994
rect 35164 26930 35216 26936
rect 34704 26240 34756 26246
rect 34704 26182 34756 26188
rect 34610 24168 34666 24177
rect 34610 24103 34666 24112
rect 34612 24064 34664 24070
rect 34612 24006 34664 24012
rect 34518 23896 34574 23905
rect 34518 23831 34574 23840
rect 34428 23792 34480 23798
rect 34428 23734 34480 23740
rect 34624 23730 34652 24006
rect 34336 23724 34388 23730
rect 34336 23666 34388 23672
rect 34520 23724 34572 23730
rect 34520 23666 34572 23672
rect 34612 23724 34664 23730
rect 34612 23666 34664 23672
rect 34242 22264 34298 22273
rect 34242 22199 34298 22208
rect 34152 22160 34204 22166
rect 34152 22102 34204 22108
rect 34242 21992 34298 22001
rect 34060 21956 34112 21962
rect 34060 21898 34112 21904
rect 34164 21950 34242 21978
rect 33980 21678 34100 21706
rect 34072 21321 34100 21678
rect 34058 21312 34114 21321
rect 34058 21247 34114 21256
rect 33966 21176 34022 21185
rect 33966 21111 34022 21120
rect 34060 21140 34112 21146
rect 33980 21078 34008 21111
rect 34060 21082 34112 21088
rect 33968 21072 34020 21078
rect 33968 21014 34020 21020
rect 33876 20596 33928 20602
rect 33876 20538 33928 20544
rect 33876 20256 33928 20262
rect 33876 20198 33928 20204
rect 33888 20058 33916 20198
rect 33966 20088 34022 20097
rect 33876 20052 33928 20058
rect 33966 20023 34022 20032
rect 33876 19994 33928 20000
rect 33888 19417 33916 19994
rect 33980 19825 34008 20023
rect 34072 19922 34100 21082
rect 34060 19916 34112 19922
rect 34060 19858 34112 19864
rect 33966 19816 34022 19825
rect 33966 19751 33968 19760
rect 34020 19751 34022 19760
rect 33968 19722 34020 19728
rect 34060 19712 34112 19718
rect 34060 19654 34112 19660
rect 34072 19446 34100 19654
rect 34164 19446 34192 21950
rect 34242 21927 34298 21936
rect 34242 21856 34298 21865
rect 34242 21791 34298 21800
rect 34256 19802 34284 21791
rect 34348 21049 34376 23666
rect 34532 23610 34560 23666
rect 34440 23582 34560 23610
rect 34440 23361 34468 23582
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 34426 23352 34482 23361
rect 34532 23322 34560 23462
rect 34426 23287 34482 23296
rect 34520 23316 34572 23322
rect 34520 23258 34572 23264
rect 34612 23316 34664 23322
rect 34612 23258 34664 23264
rect 34518 23216 34574 23225
rect 34518 23151 34574 23160
rect 34532 22794 34560 23151
rect 34624 22982 34652 23258
rect 34612 22976 34664 22982
rect 34612 22918 34664 22924
rect 34532 22766 34652 22794
rect 34518 22400 34574 22409
rect 34518 22335 34574 22344
rect 34532 22234 34560 22335
rect 34520 22228 34572 22234
rect 34440 22188 34520 22216
rect 34334 21040 34390 21049
rect 34334 20975 34390 20984
rect 34440 20466 34468 22188
rect 34520 22170 34572 22176
rect 34520 21956 34572 21962
rect 34520 21898 34572 21904
rect 34428 20460 34480 20466
rect 34428 20402 34480 20408
rect 34532 19922 34560 21898
rect 34624 20942 34652 22766
rect 34716 22080 34744 26182
rect 34808 26042 34836 26930
rect 34888 26852 34940 26858
rect 35072 26852 35124 26858
rect 34940 26812 35072 26840
rect 34888 26794 34940 26800
rect 35072 26794 35124 26800
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35162 26072 35218 26081
rect 34796 26036 34848 26042
rect 35162 26007 35218 26016
rect 34796 25978 34848 25984
rect 35176 25838 35204 26007
rect 35164 25832 35216 25838
rect 35164 25774 35216 25780
rect 34794 25664 34850 25673
rect 34794 25599 34850 25608
rect 34808 24324 34836 25599
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35164 25492 35216 25498
rect 35164 25434 35216 25440
rect 34888 25288 34940 25294
rect 34888 25230 34940 25236
rect 34900 24857 34928 25230
rect 35176 24954 35204 25434
rect 35164 24948 35216 24954
rect 35164 24890 35216 24896
rect 34886 24848 34942 24857
rect 34886 24783 34942 24792
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34980 24336 35032 24342
rect 34808 24296 34980 24324
rect 34980 24278 35032 24284
rect 34980 24200 35032 24206
rect 34980 24142 35032 24148
rect 34992 24041 35020 24142
rect 34978 24032 35034 24041
rect 34978 23967 35034 23976
rect 34796 23724 34848 23730
rect 34796 23666 34848 23672
rect 34808 23100 34836 23666
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34888 23248 34940 23254
rect 34886 23216 34888 23225
rect 34940 23216 34942 23225
rect 34886 23151 34942 23160
rect 34888 23112 34940 23118
rect 34808 23072 34888 23100
rect 34888 23054 34940 23060
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35164 22228 35216 22234
rect 35164 22170 35216 22176
rect 34716 22052 34836 22080
rect 34704 21956 34756 21962
rect 34704 21898 34756 21904
rect 34612 20936 34664 20942
rect 34612 20878 34664 20884
rect 34612 20392 34664 20398
rect 34610 20360 34612 20369
rect 34664 20360 34666 20369
rect 34610 20295 34666 20304
rect 34624 19922 34652 20295
rect 34520 19916 34572 19922
rect 34520 19858 34572 19864
rect 34612 19916 34664 19922
rect 34612 19858 34664 19864
rect 34428 19848 34480 19854
rect 34256 19774 34376 19802
rect 34428 19790 34480 19796
rect 34518 19816 34574 19825
rect 34244 19712 34296 19718
rect 34244 19654 34296 19660
rect 34060 19440 34112 19446
rect 33874 19408 33930 19417
rect 34060 19382 34112 19388
rect 34152 19440 34204 19446
rect 34152 19382 34204 19388
rect 33874 19343 33930 19352
rect 34060 18624 34112 18630
rect 34060 18566 34112 18572
rect 34072 18290 34100 18566
rect 34060 18284 34112 18290
rect 34060 18226 34112 18232
rect 34060 18148 34112 18154
rect 34060 18090 34112 18096
rect 33784 18080 33836 18086
rect 33784 18022 33836 18028
rect 33968 18080 34020 18086
rect 33968 18022 34020 18028
rect 33876 17876 33928 17882
rect 33876 17818 33928 17824
rect 33782 17776 33838 17785
rect 33782 17711 33838 17720
rect 33796 17678 33824 17711
rect 33784 17672 33836 17678
rect 33784 17614 33836 17620
rect 33888 17610 33916 17818
rect 33980 17678 34008 18022
rect 34072 17882 34100 18090
rect 34164 18086 34192 19382
rect 34256 19378 34284 19654
rect 34244 19372 34296 19378
rect 34244 19314 34296 19320
rect 34242 18456 34298 18465
rect 34242 18391 34298 18400
rect 34256 18290 34284 18391
rect 34244 18284 34296 18290
rect 34244 18226 34296 18232
rect 34152 18080 34204 18086
rect 34152 18022 34204 18028
rect 34256 17882 34284 18226
rect 34060 17876 34112 17882
rect 34060 17818 34112 17824
rect 34244 17876 34296 17882
rect 34244 17818 34296 17824
rect 33968 17672 34020 17678
rect 33968 17614 34020 17620
rect 33876 17604 33928 17610
rect 33876 17546 33928 17552
rect 34072 17338 34100 17818
rect 34152 17536 34204 17542
rect 34152 17478 34204 17484
rect 34060 17332 34112 17338
rect 34060 17274 34112 17280
rect 34164 17105 34192 17478
rect 34150 17096 34206 17105
rect 34150 17031 34206 17040
rect 34060 16788 34112 16794
rect 34060 16730 34112 16736
rect 33692 16176 33744 16182
rect 33692 16118 33744 16124
rect 33600 15904 33652 15910
rect 33600 15846 33652 15852
rect 33324 15700 33376 15706
rect 33324 15642 33376 15648
rect 33508 15700 33560 15706
rect 33508 15642 33560 15648
rect 33232 15632 33284 15638
rect 33232 15574 33284 15580
rect 33140 15020 33192 15026
rect 33140 14962 33192 14968
rect 32678 14648 32734 14657
rect 32678 14583 32734 14592
rect 31852 14340 31904 14346
rect 31852 14282 31904 14288
rect 31668 14000 31720 14006
rect 31668 13942 31720 13948
rect 32312 14000 32364 14006
rect 32312 13942 32364 13948
rect 32324 13802 32352 13942
rect 33244 13938 33272 15574
rect 33324 15496 33376 15502
rect 33600 15496 33652 15502
rect 33324 15438 33376 15444
rect 33598 15464 33600 15473
rect 33652 15464 33654 15473
rect 33336 14006 33364 15438
rect 33598 15399 33654 15408
rect 33784 15428 33836 15434
rect 33784 15370 33836 15376
rect 33796 15162 33824 15370
rect 33784 15156 33836 15162
rect 33784 15098 33836 15104
rect 33508 15088 33560 15094
rect 33508 15030 33560 15036
rect 33690 15056 33746 15065
rect 33520 14929 33548 15030
rect 33690 14991 33692 15000
rect 33744 14991 33746 15000
rect 33692 14962 33744 14968
rect 33506 14920 33562 14929
rect 33506 14855 33562 14864
rect 33704 14482 33732 14962
rect 33692 14476 33744 14482
rect 33692 14418 33744 14424
rect 33324 14000 33376 14006
rect 33324 13942 33376 13948
rect 33232 13932 33284 13938
rect 33232 13874 33284 13880
rect 34072 13870 34100 16730
rect 34256 15502 34284 17818
rect 34348 16046 34376 19774
rect 34440 17678 34468 19790
rect 34518 19751 34574 19760
rect 34532 18170 34560 19751
rect 34716 19514 34744 21898
rect 34808 20262 34836 22052
rect 35070 21720 35126 21729
rect 35070 21655 35126 21664
rect 35084 21622 35112 21655
rect 35072 21616 35124 21622
rect 35072 21558 35124 21564
rect 35176 21486 35204 22170
rect 35256 22160 35308 22166
rect 35256 22102 35308 22108
rect 35268 21554 35296 22102
rect 35360 21690 35388 27390
rect 35820 27334 35848 27882
rect 35808 27328 35860 27334
rect 35808 27270 35860 27276
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35438 27160 35494 27169
rect 35594 27163 35902 27172
rect 35438 27095 35494 27104
rect 35452 26994 35480 27095
rect 35440 26988 35492 26994
rect 35440 26930 35492 26936
rect 35440 26784 35492 26790
rect 35440 26726 35492 26732
rect 35452 26246 35480 26726
rect 35530 26616 35586 26625
rect 35530 26551 35532 26560
rect 35584 26551 35586 26560
rect 35532 26522 35584 26528
rect 35440 26240 35492 26246
rect 35440 26182 35492 26188
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 35440 25696 35492 25702
rect 35440 25638 35492 25644
rect 35452 24818 35480 25638
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 35532 24880 35584 24886
rect 35532 24822 35584 24828
rect 35440 24812 35492 24818
rect 35440 24754 35492 24760
rect 35544 24206 35572 24822
rect 36004 24750 36032 28426
rect 36084 27396 36136 27402
rect 36084 27338 36136 27344
rect 36096 26081 36124 27338
rect 36082 26072 36138 26081
rect 36082 26007 36138 26016
rect 36084 25900 36136 25906
rect 36084 25842 36136 25848
rect 35992 24744 36044 24750
rect 35992 24686 36044 24692
rect 35716 24608 35768 24614
rect 35716 24550 35768 24556
rect 35624 24404 35676 24410
rect 35624 24346 35676 24352
rect 35636 24206 35664 24346
rect 35728 24274 35756 24550
rect 35716 24268 35768 24274
rect 35716 24210 35768 24216
rect 35440 24200 35492 24206
rect 35440 24142 35492 24148
rect 35532 24200 35584 24206
rect 35532 24142 35584 24148
rect 35624 24200 35676 24206
rect 35624 24142 35676 24148
rect 35452 23186 35480 24142
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 36004 23798 36032 24686
rect 36096 24206 36124 25842
rect 36188 25294 36216 28970
rect 36268 28960 36320 28966
rect 36268 28902 36320 28908
rect 36176 25288 36228 25294
rect 36176 25230 36228 25236
rect 36280 24682 36308 28902
rect 36268 24676 36320 24682
rect 36268 24618 36320 24624
rect 36084 24200 36136 24206
rect 36084 24142 36136 24148
rect 36268 24200 36320 24206
rect 36268 24142 36320 24148
rect 35992 23792 36044 23798
rect 35992 23734 36044 23740
rect 35440 23180 35492 23186
rect 35440 23122 35492 23128
rect 35624 23112 35676 23118
rect 35624 23054 35676 23060
rect 35440 23044 35492 23050
rect 35440 22986 35492 22992
rect 35452 22234 35480 22986
rect 35636 22982 35664 23054
rect 35624 22976 35676 22982
rect 35624 22918 35676 22924
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 35624 22636 35676 22642
rect 35624 22578 35676 22584
rect 35532 22500 35584 22506
rect 35532 22442 35584 22448
rect 35440 22228 35492 22234
rect 35440 22170 35492 22176
rect 35544 22098 35572 22442
rect 35532 22092 35584 22098
rect 35532 22034 35584 22040
rect 35440 22024 35492 22030
rect 35440 21966 35492 21972
rect 35530 21992 35586 22001
rect 35348 21684 35400 21690
rect 35348 21626 35400 21632
rect 35256 21548 35308 21554
rect 35256 21490 35308 21496
rect 35164 21480 35216 21486
rect 35164 21422 35216 21428
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34888 21140 34940 21146
rect 34888 21082 34940 21088
rect 34900 20874 34928 21082
rect 35360 21010 35388 21626
rect 35348 21004 35400 21010
rect 35348 20946 35400 20952
rect 35452 20913 35480 21966
rect 35636 21978 35664 22578
rect 36096 22166 36124 24142
rect 36176 23112 36228 23118
rect 36176 23054 36228 23060
rect 36084 22160 36136 22166
rect 36084 22102 36136 22108
rect 35586 21950 35664 21978
rect 35530 21927 35532 21936
rect 35584 21927 35586 21936
rect 35532 21898 35584 21904
rect 35992 21888 36044 21894
rect 35992 21830 36044 21836
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 35532 21480 35584 21486
rect 35532 21422 35584 21428
rect 35544 21146 35572 21422
rect 36004 21146 36032 21830
rect 35532 21140 35584 21146
rect 35532 21082 35584 21088
rect 35992 21140 36044 21146
rect 35992 21082 36044 21088
rect 36188 21026 36216 23054
rect 36280 21146 36308 24142
rect 36372 22710 36400 32166
rect 36544 31272 36596 31278
rect 36544 31214 36596 31220
rect 36452 28416 36504 28422
rect 36452 28358 36504 28364
rect 36464 25770 36492 28358
rect 36556 28150 36584 31214
rect 37004 30048 37056 30054
rect 37004 29990 37056 29996
rect 36728 28620 36780 28626
rect 36728 28562 36780 28568
rect 36740 28150 36768 28562
rect 37016 28558 37044 29990
rect 37004 28552 37056 28558
rect 37004 28494 37056 28500
rect 36544 28144 36596 28150
rect 36544 28086 36596 28092
rect 36728 28144 36780 28150
rect 36728 28086 36780 28092
rect 36912 28008 36964 28014
rect 36912 27950 36964 27956
rect 36544 27872 36596 27878
rect 36544 27814 36596 27820
rect 36452 25764 36504 25770
rect 36452 25706 36504 25712
rect 36452 25492 36504 25498
rect 36452 25434 36504 25440
rect 36464 25401 36492 25434
rect 36450 25392 36506 25401
rect 36556 25378 36584 27814
rect 36728 27464 36780 27470
rect 36634 27432 36690 27441
rect 36728 27406 36780 27412
rect 36634 27367 36690 27376
rect 36648 26042 36676 27367
rect 36636 26036 36688 26042
rect 36636 25978 36688 25984
rect 36556 25350 36676 25378
rect 36450 25327 36506 25336
rect 36648 25294 36676 25350
rect 36636 25288 36688 25294
rect 36464 25236 36636 25242
rect 36464 25230 36688 25236
rect 36464 25214 36676 25230
rect 36464 23526 36492 25214
rect 36740 25140 36768 27406
rect 36924 26790 36952 27950
rect 36912 26784 36964 26790
rect 36648 25112 36768 25140
rect 36832 26744 36912 26772
rect 36544 24064 36596 24070
rect 36544 24006 36596 24012
rect 36452 23520 36504 23526
rect 36452 23462 36504 23468
rect 36556 22778 36584 24006
rect 36544 22772 36596 22778
rect 36544 22714 36596 22720
rect 36360 22704 36412 22710
rect 36360 22646 36412 22652
rect 36372 22234 36400 22646
rect 36450 22536 36506 22545
rect 36450 22471 36506 22480
rect 36360 22228 36412 22234
rect 36360 22170 36412 22176
rect 36464 21894 36492 22471
rect 36452 21888 36504 21894
rect 36452 21830 36504 21836
rect 36268 21140 36320 21146
rect 36268 21082 36320 21088
rect 36004 20998 36216 21026
rect 36360 21072 36412 21078
rect 36360 21014 36412 21020
rect 36542 21040 36598 21049
rect 35438 20904 35494 20913
rect 34888 20868 34940 20874
rect 34888 20810 34940 20816
rect 35348 20868 35400 20874
rect 35438 20839 35494 20848
rect 35348 20810 35400 20816
rect 34796 20256 34848 20262
rect 34796 20198 34848 20204
rect 34704 19508 34756 19514
rect 34704 19450 34756 19456
rect 34702 18320 34758 18329
rect 34702 18255 34704 18264
rect 34756 18255 34758 18264
rect 34704 18226 34756 18232
rect 34532 18142 34652 18170
rect 34520 18080 34572 18086
rect 34518 18048 34520 18057
rect 34572 18048 34574 18057
rect 34518 17983 34574 17992
rect 34428 17672 34480 17678
rect 34428 17614 34480 17620
rect 34336 16040 34388 16046
rect 34336 15982 34388 15988
rect 34348 15706 34376 15982
rect 34336 15700 34388 15706
rect 34336 15642 34388 15648
rect 34244 15496 34296 15502
rect 34244 15438 34296 15444
rect 34060 13864 34112 13870
rect 34060 13806 34112 13812
rect 32312 13796 32364 13802
rect 32312 13738 32364 13744
rect 34440 13433 34468 17614
rect 34624 14074 34652 18142
rect 34704 18080 34756 18086
rect 34704 18022 34756 18028
rect 34716 15570 34744 18022
rect 34808 16776 34836 20198
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34980 18692 35032 18698
rect 34980 18634 35032 18640
rect 34888 18216 34940 18222
rect 34888 18158 34940 18164
rect 34900 18086 34928 18158
rect 34992 18086 35020 18634
rect 35360 18329 35388 20810
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 35440 20052 35492 20058
rect 35440 19994 35492 20000
rect 35532 20052 35584 20058
rect 35532 19994 35584 20000
rect 35452 19854 35480 19994
rect 35440 19848 35492 19854
rect 35440 19790 35492 19796
rect 35346 18320 35402 18329
rect 35346 18255 35402 18264
rect 35348 18148 35400 18154
rect 35348 18090 35400 18096
rect 34888 18080 34940 18086
rect 34888 18022 34940 18028
rect 34980 18080 35032 18086
rect 34980 18022 35032 18028
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35360 17785 35388 18090
rect 35346 17776 35402 17785
rect 35164 17740 35216 17746
rect 35346 17711 35402 17720
rect 35164 17682 35216 17688
rect 35176 17610 35204 17682
rect 35360 17678 35388 17711
rect 35348 17672 35400 17678
rect 35348 17614 35400 17620
rect 35072 17604 35124 17610
rect 35072 17546 35124 17552
rect 35164 17604 35216 17610
rect 35164 17546 35216 17552
rect 35084 17377 35112 17546
rect 35348 17536 35400 17542
rect 35452 17490 35480 19790
rect 35544 19786 35572 19994
rect 35532 19780 35584 19786
rect 35532 19722 35584 19728
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 35400 17484 35480 17490
rect 35348 17478 35480 17484
rect 35360 17462 35480 17478
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35070 17368 35126 17377
rect 35594 17371 35902 17380
rect 35070 17303 35126 17312
rect 35716 17264 35768 17270
rect 35346 17232 35402 17241
rect 35544 17212 35716 17218
rect 35544 17206 35768 17212
rect 35544 17202 35756 17206
rect 35346 17167 35402 17176
rect 35532 17196 35756 17202
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34808 16748 34928 16776
rect 34900 16114 34928 16748
rect 35360 16114 35388 17167
rect 35584 17190 35756 17196
rect 35900 17196 35952 17202
rect 35532 17138 35584 17144
rect 35900 17138 35952 17144
rect 35440 17128 35492 17134
rect 35440 17070 35492 17076
rect 35716 17128 35768 17134
rect 35716 17070 35768 17076
rect 34888 16108 34940 16114
rect 34888 16050 34940 16056
rect 35348 16108 35400 16114
rect 35348 16050 35400 16056
rect 34796 16040 34848 16046
rect 34796 15982 34848 15988
rect 34808 15706 34836 15982
rect 35452 15978 35480 17070
rect 35728 16998 35756 17070
rect 35716 16992 35768 16998
rect 35716 16934 35768 16940
rect 35912 16794 35940 17138
rect 35900 16788 35952 16794
rect 35900 16730 35952 16736
rect 36004 16538 36032 20998
rect 36176 20936 36228 20942
rect 36176 20878 36228 20884
rect 36268 20936 36320 20942
rect 36268 20878 36320 20884
rect 36188 20602 36216 20878
rect 36176 20596 36228 20602
rect 36176 20538 36228 20544
rect 36176 20392 36228 20398
rect 36176 20334 36228 20340
rect 36084 17604 36136 17610
rect 36084 17546 36136 17552
rect 36096 17338 36124 17546
rect 36084 17332 36136 17338
rect 36084 17274 36136 17280
rect 36004 16510 36124 16538
rect 35992 16448 36044 16454
rect 35992 16390 36044 16396
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 36004 16130 36032 16390
rect 35820 16114 36032 16130
rect 35808 16108 36032 16114
rect 35860 16102 36032 16108
rect 35808 16050 35860 16056
rect 35440 15972 35492 15978
rect 35440 15914 35492 15920
rect 35808 15904 35860 15910
rect 35808 15846 35860 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34796 15700 34848 15706
rect 34796 15642 34848 15648
rect 34704 15564 34756 15570
rect 34704 15506 34756 15512
rect 34796 15564 34848 15570
rect 34796 15506 34848 15512
rect 34808 14385 34836 15506
rect 35820 15434 35848 15846
rect 35808 15428 35860 15434
rect 35808 15370 35860 15376
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34794 14376 34850 14385
rect 34794 14311 34850 14320
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 34612 14068 34664 14074
rect 34612 14010 34664 14016
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 36096 13530 36124 16510
rect 36188 15162 36216 20334
rect 36280 17882 36308 20878
rect 36372 20262 36400 21014
rect 36542 20975 36598 20984
rect 36360 20256 36412 20262
rect 36360 20198 36412 20204
rect 36556 19310 36584 20975
rect 36544 19304 36596 19310
rect 36544 19246 36596 19252
rect 36544 18896 36596 18902
rect 36544 18838 36596 18844
rect 36268 17876 36320 17882
rect 36268 17818 36320 17824
rect 36556 17814 36584 18838
rect 36648 18358 36676 25112
rect 36728 24676 36780 24682
rect 36728 24618 36780 24624
rect 36740 24018 36768 24618
rect 36832 24206 36860 26744
rect 36912 26726 36964 26732
rect 36912 26444 36964 26450
rect 36912 26386 36964 26392
rect 36924 26246 36952 26386
rect 36912 26240 36964 26246
rect 36912 26182 36964 26188
rect 36912 26036 36964 26042
rect 36912 25978 36964 25984
rect 36924 25362 36952 25978
rect 36912 25356 36964 25362
rect 36912 25298 36964 25304
rect 37016 24290 37044 28494
rect 37108 28014 37136 32302
rect 37476 31754 37504 32506
rect 39026 32328 39082 32337
rect 39026 32263 39082 32272
rect 37476 31726 37872 31754
rect 37738 30016 37794 30025
rect 37738 29951 37794 29960
rect 37370 29744 37426 29753
rect 37370 29679 37426 29688
rect 37384 29238 37412 29679
rect 37648 29572 37700 29578
rect 37648 29514 37700 29520
rect 37372 29232 37424 29238
rect 37372 29174 37424 29180
rect 37188 29096 37240 29102
rect 37188 29038 37240 29044
rect 37200 28762 37228 29038
rect 37660 29034 37688 29514
rect 37648 29028 37700 29034
rect 37648 28970 37700 28976
rect 37188 28756 37240 28762
rect 37188 28698 37240 28704
rect 37096 28008 37148 28014
rect 37096 27950 37148 27956
rect 37200 27674 37228 28698
rect 37464 28484 37516 28490
rect 37464 28426 37516 28432
rect 37476 27878 37504 28426
rect 37556 28144 37608 28150
rect 37608 28092 37688 28098
rect 37556 28086 37688 28092
rect 37568 28070 37688 28086
rect 37464 27872 37516 27878
rect 37464 27814 37516 27820
rect 37188 27668 37240 27674
rect 37188 27610 37240 27616
rect 37372 27668 37424 27674
rect 37372 27610 37424 27616
rect 37384 27130 37412 27610
rect 37372 27124 37424 27130
rect 37372 27066 37424 27072
rect 37476 27010 37504 27814
rect 37556 27464 37608 27470
rect 37556 27406 37608 27412
rect 37384 26982 37504 27010
rect 37188 26920 37240 26926
rect 37186 26888 37188 26897
rect 37240 26888 37242 26897
rect 37186 26823 37242 26832
rect 37200 26586 37228 26823
rect 37188 26580 37240 26586
rect 37188 26522 37240 26528
rect 37096 26036 37148 26042
rect 37096 25978 37148 25984
rect 36924 24262 37044 24290
rect 36820 24200 36872 24206
rect 36820 24142 36872 24148
rect 36740 23990 36860 24018
rect 36726 23760 36782 23769
rect 36726 23695 36728 23704
rect 36780 23695 36782 23704
rect 36728 23666 36780 23672
rect 36728 23520 36780 23526
rect 36728 23462 36780 23468
rect 36636 18352 36688 18358
rect 36636 18294 36688 18300
rect 36544 17808 36596 17814
rect 36544 17750 36596 17756
rect 36452 17672 36504 17678
rect 36372 17632 36452 17660
rect 36372 17270 36400 17632
rect 36452 17614 36504 17620
rect 36556 17490 36584 17750
rect 36740 17746 36768 23462
rect 36832 22438 36860 23990
rect 36924 23118 36952 24262
rect 37004 24132 37056 24138
rect 37004 24074 37056 24080
rect 36912 23112 36964 23118
rect 36912 23054 36964 23060
rect 36820 22432 36872 22438
rect 36820 22374 36872 22380
rect 36818 21584 36874 21593
rect 36818 21519 36874 21528
rect 36832 20534 36860 21519
rect 36820 20528 36872 20534
rect 36820 20470 36872 20476
rect 36912 20392 36964 20398
rect 36912 20334 36964 20340
rect 36924 19334 36952 20334
rect 37016 20058 37044 24074
rect 37108 23322 37136 25978
rect 37096 23316 37148 23322
rect 37096 23258 37148 23264
rect 37108 21078 37136 23258
rect 37200 23118 37228 26522
rect 37278 25800 37334 25809
rect 37278 25735 37280 25744
rect 37332 25735 37334 25744
rect 37280 25706 37332 25712
rect 37280 23316 37332 23322
rect 37280 23258 37332 23264
rect 37292 23225 37320 23258
rect 37278 23216 37334 23225
rect 37278 23151 37334 23160
rect 37188 23112 37240 23118
rect 37188 23054 37240 23060
rect 37096 21072 37148 21078
rect 37096 21014 37148 21020
rect 37096 20460 37148 20466
rect 37096 20402 37148 20408
rect 37004 20052 37056 20058
rect 37004 19994 37056 20000
rect 37108 19961 37136 20402
rect 37200 20398 37228 23054
rect 37384 22094 37412 26982
rect 37464 26376 37516 26382
rect 37464 26318 37516 26324
rect 37476 26042 37504 26318
rect 37464 26036 37516 26042
rect 37464 25978 37516 25984
rect 37464 25900 37516 25906
rect 37464 25842 37516 25848
rect 37476 25702 37504 25842
rect 37464 25696 37516 25702
rect 37464 25638 37516 25644
rect 37476 24993 37504 25638
rect 37568 25498 37596 27406
rect 37660 26353 37688 28070
rect 37646 26344 37702 26353
rect 37646 26279 37702 26288
rect 37556 25492 37608 25498
rect 37556 25434 37608 25440
rect 37462 24984 37518 24993
rect 37462 24919 37518 24928
rect 37556 23656 37608 23662
rect 37462 23624 37518 23633
rect 37556 23598 37608 23604
rect 37462 23559 37518 23568
rect 37476 23322 37504 23559
rect 37464 23316 37516 23322
rect 37464 23258 37516 23264
rect 37476 23118 37504 23258
rect 37568 23186 37596 23598
rect 37556 23180 37608 23186
rect 37556 23122 37608 23128
rect 37464 23112 37516 23118
rect 37464 23054 37516 23060
rect 37660 22094 37688 26279
rect 37752 25430 37780 29951
rect 37740 25424 37792 25430
rect 37740 25366 37792 25372
rect 37740 24200 37792 24206
rect 37740 24142 37792 24148
rect 37292 22066 37412 22094
rect 37568 22066 37688 22094
rect 37292 21622 37320 22066
rect 37280 21616 37332 21622
rect 37280 21558 37332 21564
rect 37372 21616 37424 21622
rect 37372 21558 37424 21564
rect 37462 21584 37518 21593
rect 37384 21350 37412 21558
rect 37462 21519 37464 21528
rect 37516 21519 37518 21528
rect 37464 21490 37516 21496
rect 37568 21350 37596 22066
rect 37752 21486 37780 24142
rect 37740 21480 37792 21486
rect 37740 21422 37792 21428
rect 37372 21344 37424 21350
rect 37372 21286 37424 21292
rect 37556 21344 37608 21350
rect 37556 21286 37608 21292
rect 37188 20392 37240 20398
rect 37188 20334 37240 20340
rect 37188 20052 37240 20058
rect 37188 19994 37240 20000
rect 37094 19952 37150 19961
rect 37094 19887 37150 19896
rect 36832 19306 36952 19334
rect 36728 17740 36780 17746
rect 36728 17682 36780 17688
rect 36464 17462 36584 17490
rect 36360 17264 36412 17270
rect 36360 17206 36412 17212
rect 36464 17134 36492 17462
rect 36634 17232 36690 17241
rect 36634 17167 36636 17176
rect 36688 17167 36690 17176
rect 36636 17138 36688 17144
rect 36452 17128 36504 17134
rect 36544 17128 36596 17134
rect 36452 17070 36504 17076
rect 36542 17096 36544 17105
rect 36596 17096 36598 17105
rect 36542 17031 36598 17040
rect 36728 17060 36780 17066
rect 36728 17002 36780 17008
rect 36544 16244 36596 16250
rect 36544 16186 36596 16192
rect 36556 16046 36584 16186
rect 36634 16144 36690 16153
rect 36634 16079 36690 16088
rect 36648 16046 36676 16079
rect 36544 16040 36596 16046
rect 36544 15982 36596 15988
rect 36636 16040 36688 16046
rect 36636 15982 36688 15988
rect 36740 15978 36768 17002
rect 36832 16522 36860 19306
rect 37004 18760 37056 18766
rect 36910 18728 36966 18737
rect 37004 18702 37056 18708
rect 37096 18760 37148 18766
rect 37096 18702 37148 18708
rect 36910 18663 36966 18672
rect 36924 18290 36952 18663
rect 36912 18284 36964 18290
rect 36912 18226 36964 18232
rect 37016 17542 37044 18702
rect 37108 18426 37136 18702
rect 37200 18630 37228 19994
rect 37464 19712 37516 19718
rect 37464 19654 37516 19660
rect 37476 18970 37504 19654
rect 37464 18964 37516 18970
rect 37464 18906 37516 18912
rect 37280 18828 37332 18834
rect 37280 18770 37332 18776
rect 37188 18624 37240 18630
rect 37188 18566 37240 18572
rect 37096 18420 37148 18426
rect 37096 18362 37148 18368
rect 37200 17882 37228 18566
rect 37292 18222 37320 18770
rect 37476 18290 37504 18906
rect 37372 18284 37424 18290
rect 37372 18226 37424 18232
rect 37464 18284 37516 18290
rect 37464 18226 37516 18232
rect 37280 18216 37332 18222
rect 37280 18158 37332 18164
rect 37188 17876 37240 17882
rect 37188 17818 37240 17824
rect 37004 17536 37056 17542
rect 37004 17478 37056 17484
rect 37292 17338 37320 18158
rect 37280 17332 37332 17338
rect 37280 17274 37332 17280
rect 36912 17264 36964 17270
rect 36912 17206 36964 17212
rect 36820 16516 36872 16522
rect 36820 16458 36872 16464
rect 36924 16454 36952 17206
rect 37188 16992 37240 16998
rect 37188 16934 37240 16940
rect 37200 16794 37228 16934
rect 37188 16788 37240 16794
rect 37188 16730 37240 16736
rect 37094 16552 37150 16561
rect 37384 16538 37412 18226
rect 37462 18184 37518 18193
rect 37462 18119 37518 18128
rect 37476 18086 37504 18119
rect 37464 18080 37516 18086
rect 37464 18022 37516 18028
rect 37568 17678 37596 21286
rect 37752 19334 37780 21422
rect 37660 19306 37780 19334
rect 37556 17672 37608 17678
rect 37556 17614 37608 17620
rect 37660 17490 37688 19306
rect 37844 17814 37872 31726
rect 38016 30932 38068 30938
rect 38016 30874 38068 30880
rect 38028 28626 38056 30874
rect 38566 30152 38622 30161
rect 38566 30087 38622 30096
rect 38384 29776 38436 29782
rect 38384 29718 38436 29724
rect 38292 29028 38344 29034
rect 38292 28970 38344 28976
rect 38016 28620 38068 28626
rect 38016 28562 38068 28568
rect 38028 28218 38056 28562
rect 38200 28416 38252 28422
rect 38200 28358 38252 28364
rect 38016 28212 38068 28218
rect 38016 28154 38068 28160
rect 38016 28076 38068 28082
rect 38016 28018 38068 28024
rect 37922 26616 37978 26625
rect 37922 26551 37924 26560
rect 37976 26551 37978 26560
rect 37924 26522 37976 26528
rect 37924 25832 37976 25838
rect 37924 25774 37976 25780
rect 37936 22574 37964 25774
rect 38028 23322 38056 28018
rect 38016 23316 38068 23322
rect 38016 23258 38068 23264
rect 38108 23316 38160 23322
rect 38108 23258 38160 23264
rect 38120 22710 38148 23258
rect 38108 22704 38160 22710
rect 38108 22646 38160 22652
rect 38016 22636 38068 22642
rect 38016 22578 38068 22584
rect 37924 22568 37976 22574
rect 37924 22510 37976 22516
rect 38028 21486 38056 22578
rect 38108 21616 38160 21622
rect 38108 21558 38160 21564
rect 38016 21480 38068 21486
rect 38016 21422 38068 21428
rect 37924 20392 37976 20398
rect 37924 20334 37976 20340
rect 37832 17808 37884 17814
rect 37832 17750 37884 17756
rect 37568 17462 37688 17490
rect 37464 16788 37516 16794
rect 37464 16730 37516 16736
rect 37094 16487 37150 16496
rect 37292 16510 37412 16538
rect 36912 16448 36964 16454
rect 36912 16390 36964 16396
rect 36924 16114 36952 16390
rect 36912 16108 36964 16114
rect 36912 16050 36964 16056
rect 37004 16040 37056 16046
rect 37004 15982 37056 15988
rect 36728 15972 36780 15978
rect 36728 15914 36780 15920
rect 37016 15706 37044 15982
rect 37004 15700 37056 15706
rect 37004 15642 37056 15648
rect 37108 15366 37136 16487
rect 37188 15904 37240 15910
rect 37188 15846 37240 15852
rect 37200 15434 37228 15846
rect 37292 15706 37320 16510
rect 37372 16448 37424 16454
rect 37372 16390 37424 16396
rect 37280 15700 37332 15706
rect 37280 15642 37332 15648
rect 37188 15428 37240 15434
rect 37188 15370 37240 15376
rect 37096 15360 37148 15366
rect 37096 15302 37148 15308
rect 36176 15156 36228 15162
rect 36176 15098 36228 15104
rect 37384 15094 37412 16390
rect 37372 15088 37424 15094
rect 37372 15030 37424 15036
rect 37476 14521 37504 16730
rect 37462 14512 37518 14521
rect 37462 14447 37518 14456
rect 36084 13524 36136 13530
rect 36084 13466 36136 13472
rect 34426 13424 34482 13433
rect 31576 13388 31628 13394
rect 34426 13359 34482 13368
rect 31576 13330 31628 13336
rect 31668 13252 31720 13258
rect 31668 13194 31720 13200
rect 31484 12980 31536 12986
rect 31484 12922 31536 12928
rect 31116 12912 31168 12918
rect 31116 12854 31168 12860
rect 31680 12782 31708 13194
rect 37568 13190 37596 17462
rect 37648 17196 37700 17202
rect 37648 17138 37700 17144
rect 37660 16998 37688 17138
rect 37740 17060 37792 17066
rect 37740 17002 37792 17008
rect 37648 16992 37700 16998
rect 37648 16934 37700 16940
rect 37660 16538 37688 16934
rect 37752 16658 37780 17002
rect 37740 16652 37792 16658
rect 37740 16594 37792 16600
rect 37660 16510 37780 16538
rect 37844 16522 37872 17750
rect 37648 15496 37700 15502
rect 37648 15438 37700 15444
rect 37660 15026 37688 15438
rect 37752 15026 37780 16510
rect 37832 16516 37884 16522
rect 37832 16458 37884 16464
rect 37648 15020 37700 15026
rect 37648 14962 37700 14968
rect 37740 15020 37792 15026
rect 37740 14962 37792 14968
rect 37936 13394 37964 20334
rect 38028 17785 38056 21422
rect 38120 21350 38148 21558
rect 38108 21344 38160 21350
rect 38108 21286 38160 21292
rect 38212 20942 38240 28358
rect 38304 25514 38332 28970
rect 38396 28762 38424 29718
rect 38384 28756 38436 28762
rect 38384 28698 38436 28704
rect 38396 28506 38424 28698
rect 38580 28626 38608 30087
rect 38752 29164 38804 29170
rect 38752 29106 38804 29112
rect 38764 28762 38792 29106
rect 38752 28756 38804 28762
rect 38752 28698 38804 28704
rect 38568 28620 38620 28626
rect 38568 28562 38620 28568
rect 38396 28478 38608 28506
rect 38382 25936 38438 25945
rect 38580 25906 38608 28478
rect 38752 28484 38804 28490
rect 38752 28426 38804 28432
rect 38660 28416 38712 28422
rect 38660 28358 38712 28364
rect 38382 25871 38438 25880
rect 38568 25900 38620 25906
rect 38396 25702 38424 25871
rect 38568 25842 38620 25848
rect 38384 25696 38436 25702
rect 38384 25638 38436 25644
rect 38304 25486 38424 25514
rect 38292 24608 38344 24614
rect 38292 24550 38344 24556
rect 38304 24313 38332 24550
rect 38290 24304 38346 24313
rect 38290 24239 38346 24248
rect 38304 21554 38332 24239
rect 38396 22642 38424 25486
rect 38568 23112 38620 23118
rect 38568 23054 38620 23060
rect 38476 22976 38528 22982
rect 38476 22918 38528 22924
rect 38488 22778 38516 22918
rect 38476 22772 38528 22778
rect 38476 22714 38528 22720
rect 38384 22636 38436 22642
rect 38384 22578 38436 22584
rect 38384 22092 38436 22098
rect 38384 22034 38436 22040
rect 38292 21548 38344 21554
rect 38292 21490 38344 21496
rect 38396 21434 38424 22034
rect 38304 21406 38424 21434
rect 38304 21350 38332 21406
rect 38292 21344 38344 21350
rect 38292 21286 38344 21292
rect 38384 21344 38436 21350
rect 38384 21286 38436 21292
rect 38396 21146 38424 21286
rect 38384 21140 38436 21146
rect 38384 21082 38436 21088
rect 38200 20936 38252 20942
rect 38200 20878 38252 20884
rect 38292 20936 38344 20942
rect 38292 20878 38344 20884
rect 38304 20602 38332 20878
rect 38292 20596 38344 20602
rect 38292 20538 38344 20544
rect 38488 20534 38516 22714
rect 38476 20528 38528 20534
rect 38476 20470 38528 20476
rect 38580 19802 38608 23054
rect 38672 21962 38700 28358
rect 38764 27062 38792 28426
rect 38752 27056 38804 27062
rect 38752 26998 38804 27004
rect 38842 25256 38898 25265
rect 38842 25191 38898 25200
rect 38856 24818 38884 25191
rect 38844 24812 38896 24818
rect 38844 24754 38896 24760
rect 38752 24744 38804 24750
rect 38752 24686 38804 24692
rect 38660 21956 38712 21962
rect 38660 21898 38712 21904
rect 38764 21706 38792 24686
rect 38934 23760 38990 23769
rect 38934 23695 38936 23704
rect 38988 23695 38990 23704
rect 38936 23666 38988 23672
rect 38936 21956 38988 21962
rect 38936 21898 38988 21904
rect 38672 21678 38792 21706
rect 38948 21690 38976 21898
rect 38936 21684 38988 21690
rect 38672 20330 38700 21678
rect 38936 21626 38988 21632
rect 38752 21548 38804 21554
rect 38752 21490 38804 21496
rect 38844 21548 38896 21554
rect 38844 21490 38896 21496
rect 38660 20324 38712 20330
rect 38660 20266 38712 20272
rect 38764 19922 38792 21490
rect 38856 21146 38884 21490
rect 39040 21350 39068 32263
rect 40222 30288 40278 30297
rect 40222 30223 40278 30232
rect 39948 28960 40000 28966
rect 39948 28902 40000 28908
rect 39960 28558 39988 28902
rect 40040 28620 40092 28626
rect 40040 28562 40092 28568
rect 39948 28552 40000 28558
rect 39948 28494 40000 28500
rect 40052 27878 40080 28562
rect 40040 27872 40092 27878
rect 40040 27814 40092 27820
rect 39580 27396 39632 27402
rect 39580 27338 39632 27344
rect 39592 27130 39620 27338
rect 39580 27124 39632 27130
rect 39580 27066 39632 27072
rect 39854 27024 39910 27033
rect 39764 26988 39816 26994
rect 40052 26994 40080 27814
rect 39854 26959 39856 26968
rect 39764 26930 39816 26936
rect 39908 26959 39910 26968
rect 40040 26988 40092 26994
rect 39856 26930 39908 26936
rect 40040 26930 40092 26936
rect 39120 26512 39172 26518
rect 39120 26454 39172 26460
rect 39132 25974 39160 26454
rect 39120 25968 39172 25974
rect 39120 25910 39172 25916
rect 39776 25294 39804 26930
rect 39948 26920 40000 26926
rect 39948 26862 40000 26868
rect 40132 26920 40184 26926
rect 40132 26862 40184 26868
rect 39960 26450 39988 26862
rect 39948 26444 40000 26450
rect 39948 26386 40000 26392
rect 40144 26314 40172 26862
rect 40132 26308 40184 26314
rect 40132 26250 40184 26256
rect 39856 25900 39908 25906
rect 39856 25842 39908 25848
rect 39304 25288 39356 25294
rect 39304 25230 39356 25236
rect 39764 25288 39816 25294
rect 39764 25230 39816 25236
rect 39120 24608 39172 24614
rect 39120 24550 39172 24556
rect 39132 23526 39160 24550
rect 39212 23656 39264 23662
rect 39212 23598 39264 23604
rect 39120 23520 39172 23526
rect 39120 23462 39172 23468
rect 39224 23322 39252 23598
rect 39212 23316 39264 23322
rect 39212 23258 39264 23264
rect 39120 21480 39172 21486
rect 39120 21422 39172 21428
rect 39028 21344 39080 21350
rect 39028 21286 39080 21292
rect 38844 21140 38896 21146
rect 38844 21082 38896 21088
rect 39132 20602 39160 21422
rect 39120 20596 39172 20602
rect 39120 20538 39172 20544
rect 38752 19916 38804 19922
rect 38752 19858 38804 19864
rect 38488 19774 38608 19802
rect 38292 19304 38344 19310
rect 38292 19246 38344 19252
rect 38304 18766 38332 19246
rect 38488 19242 38516 19774
rect 38568 19712 38620 19718
rect 38568 19654 38620 19660
rect 38580 19378 38608 19654
rect 38568 19372 38620 19378
rect 38568 19314 38620 19320
rect 38660 19372 38712 19378
rect 38660 19314 38712 19320
rect 38476 19236 38528 19242
rect 38476 19178 38528 19184
rect 38672 18970 38700 19314
rect 38844 19168 38896 19174
rect 38844 19110 38896 19116
rect 38660 18964 38712 18970
rect 38660 18906 38712 18912
rect 38108 18760 38160 18766
rect 38108 18702 38160 18708
rect 38292 18760 38344 18766
rect 38292 18702 38344 18708
rect 38120 18086 38148 18702
rect 38200 18148 38252 18154
rect 38200 18090 38252 18096
rect 38108 18080 38160 18086
rect 38108 18022 38160 18028
rect 38014 17776 38070 17785
rect 38014 17711 38070 17720
rect 38212 17678 38240 18090
rect 38200 17672 38252 17678
rect 38200 17614 38252 17620
rect 38304 16998 38332 18702
rect 38752 18692 38804 18698
rect 38752 18634 38804 18640
rect 38660 18080 38712 18086
rect 38660 18022 38712 18028
rect 38476 17808 38528 17814
rect 38476 17750 38528 17756
rect 38488 17338 38516 17750
rect 38476 17332 38528 17338
rect 38476 17274 38528 17280
rect 38672 17202 38700 18022
rect 38764 17882 38792 18634
rect 38752 17876 38804 17882
rect 38752 17818 38804 17824
rect 38856 17678 38884 19110
rect 38936 18760 38988 18766
rect 38936 18702 38988 18708
rect 38948 17746 38976 18702
rect 38936 17740 38988 17746
rect 38936 17682 38988 17688
rect 38844 17672 38896 17678
rect 38750 17640 38806 17649
rect 38844 17614 38896 17620
rect 38750 17575 38752 17584
rect 38804 17575 38806 17584
rect 38752 17546 38804 17552
rect 38844 17264 38896 17270
rect 38844 17206 38896 17212
rect 38384 17196 38436 17202
rect 38384 17138 38436 17144
rect 38660 17196 38712 17202
rect 38660 17138 38712 17144
rect 38292 16992 38344 16998
rect 38292 16934 38344 16940
rect 38396 16726 38424 17138
rect 38856 17082 38884 17206
rect 38948 17202 38976 17682
rect 39028 17604 39080 17610
rect 39028 17546 39080 17552
rect 38936 17196 38988 17202
rect 38936 17138 38988 17144
rect 38580 17054 38884 17082
rect 38476 16992 38528 16998
rect 38476 16934 38528 16940
rect 38488 16794 38516 16934
rect 38476 16788 38528 16794
rect 38476 16730 38528 16736
rect 38384 16720 38436 16726
rect 38384 16662 38436 16668
rect 38580 16522 38608 17054
rect 39040 16697 39068 17546
rect 39316 16726 39344 25230
rect 39396 23724 39448 23730
rect 39396 23666 39448 23672
rect 39672 23724 39724 23730
rect 39672 23666 39724 23672
rect 39408 23254 39436 23666
rect 39396 23248 39448 23254
rect 39396 23190 39448 23196
rect 39396 21344 39448 21350
rect 39396 21286 39448 21292
rect 39408 21146 39436 21286
rect 39396 21140 39448 21146
rect 39396 21082 39448 21088
rect 39684 19854 39712 23666
rect 39868 23594 39896 25842
rect 39856 23588 39908 23594
rect 39856 23530 39908 23536
rect 39764 23316 39816 23322
rect 39764 23258 39816 23264
rect 39776 22438 39804 23258
rect 39868 23118 39896 23530
rect 39948 23316 40000 23322
rect 39948 23258 40000 23264
rect 39856 23112 39908 23118
rect 39856 23054 39908 23060
rect 39764 22432 39816 22438
rect 39764 22374 39816 22380
rect 39960 21894 39988 23258
rect 40040 22024 40092 22030
rect 40040 21966 40092 21972
rect 39948 21888 40000 21894
rect 39948 21830 40000 21836
rect 39672 19848 39724 19854
rect 39672 19790 39724 19796
rect 40052 19258 40080 21966
rect 40132 21888 40184 21894
rect 40132 21830 40184 21836
rect 40144 21622 40172 21830
rect 40132 21616 40184 21622
rect 40132 21558 40184 21564
rect 40236 20505 40264 30223
rect 44548 29640 44600 29646
rect 44548 29582 44600 29588
rect 42800 29504 42852 29510
rect 42800 29446 42852 29452
rect 41144 28688 41196 28694
rect 41144 28630 41196 28636
rect 40776 27872 40828 27878
rect 40776 27814 40828 27820
rect 40592 27668 40644 27674
rect 40592 27610 40644 27616
rect 40408 27464 40460 27470
rect 40408 27406 40460 27412
rect 40420 26994 40448 27406
rect 40408 26988 40460 26994
rect 40408 26930 40460 26936
rect 40500 26988 40552 26994
rect 40500 26930 40552 26936
rect 40512 26790 40540 26930
rect 40316 26784 40368 26790
rect 40316 26726 40368 26732
rect 40500 26784 40552 26790
rect 40500 26726 40552 26732
rect 40328 26382 40356 26726
rect 40604 26450 40632 27610
rect 40788 26994 40816 27814
rect 41052 27124 41104 27130
rect 41052 27066 41104 27072
rect 40958 27024 41014 27033
rect 40776 26988 40828 26994
rect 41064 26994 41092 27066
rect 40958 26959 40960 26968
rect 40776 26930 40828 26936
rect 41012 26959 41014 26968
rect 41052 26988 41104 26994
rect 40960 26930 41012 26936
rect 41052 26930 41104 26936
rect 40684 26920 40736 26926
rect 40684 26862 40736 26868
rect 40696 26586 40724 26862
rect 40684 26580 40736 26586
rect 40788 26568 40816 26930
rect 40788 26540 40908 26568
rect 40684 26522 40736 26528
rect 40592 26444 40644 26450
rect 40592 26386 40644 26392
rect 40316 26376 40368 26382
rect 40316 26318 40368 26324
rect 40592 25900 40644 25906
rect 40592 25842 40644 25848
rect 40604 25498 40632 25842
rect 40684 25696 40736 25702
rect 40684 25638 40736 25644
rect 40592 25492 40644 25498
rect 40592 25434 40644 25440
rect 40696 25430 40724 25638
rect 40684 25424 40736 25430
rect 40684 25366 40736 25372
rect 40880 25362 40908 26540
rect 40868 25356 40920 25362
rect 40868 25298 40920 25304
rect 40880 25158 40908 25298
rect 40868 25152 40920 25158
rect 40868 25094 40920 25100
rect 40316 24200 40368 24206
rect 40316 24142 40368 24148
rect 40328 23798 40356 24142
rect 41052 24132 41104 24138
rect 41052 24074 41104 24080
rect 40316 23792 40368 23798
rect 40316 23734 40368 23740
rect 40328 22642 40356 23734
rect 40684 23520 40736 23526
rect 40684 23462 40736 23468
rect 40696 23186 40724 23462
rect 41064 23254 41092 24074
rect 41052 23248 41104 23254
rect 41052 23190 41104 23196
rect 41156 23186 41184 28630
rect 41236 28552 41288 28558
rect 41236 28494 41288 28500
rect 41248 27674 41276 28494
rect 42064 28484 42116 28490
rect 42064 28426 42116 28432
rect 42076 27674 42104 28426
rect 42812 28150 42840 29446
rect 44560 29345 44588 29582
rect 44546 29336 44602 29345
rect 44546 29271 44602 29280
rect 44088 29028 44140 29034
rect 44088 28970 44140 28976
rect 44100 28665 44128 28970
rect 44086 28656 44142 28665
rect 44086 28591 44142 28600
rect 42984 28416 43036 28422
rect 42984 28358 43036 28364
rect 42800 28144 42852 28150
rect 42338 28112 42394 28121
rect 42800 28086 42852 28092
rect 42996 28082 43024 28358
rect 42338 28047 42394 28056
rect 42984 28076 43036 28082
rect 41236 27668 41288 27674
rect 41236 27610 41288 27616
rect 42064 27668 42116 27674
rect 42064 27610 42116 27616
rect 42352 27470 42380 28047
rect 42984 28018 43036 28024
rect 44454 27976 44510 27985
rect 44454 27911 44456 27920
rect 44508 27911 44510 27920
rect 44456 27882 44508 27888
rect 42432 27872 42484 27878
rect 42432 27814 42484 27820
rect 42616 27872 42668 27878
rect 42616 27814 42668 27820
rect 42444 27674 42472 27814
rect 42432 27668 42484 27674
rect 42432 27610 42484 27616
rect 42628 27470 42656 27814
rect 42248 27464 42300 27470
rect 42248 27406 42300 27412
rect 42340 27464 42392 27470
rect 42340 27406 42392 27412
rect 42616 27464 42668 27470
rect 42616 27406 42668 27412
rect 41328 27328 41380 27334
rect 41248 27276 41328 27282
rect 41248 27270 41380 27276
rect 41248 27254 41368 27270
rect 41248 26926 41276 27254
rect 42260 26994 42288 27406
rect 44456 27328 44508 27334
rect 44454 27296 44456 27305
rect 44508 27296 44510 27305
rect 44454 27231 44510 27240
rect 42432 27056 42484 27062
rect 42430 27024 42432 27033
rect 42484 27024 42486 27033
rect 42248 26988 42300 26994
rect 42430 26959 42486 26968
rect 42248 26930 42300 26936
rect 41236 26920 41288 26926
rect 41236 26862 41288 26868
rect 41328 26920 41380 26926
rect 41328 26862 41380 26868
rect 42064 26920 42116 26926
rect 42064 26862 42116 26868
rect 41340 26489 41368 26862
rect 42076 26586 42104 26862
rect 44272 26852 44324 26858
rect 44272 26794 44324 26800
rect 42248 26784 42300 26790
rect 42248 26726 42300 26732
rect 42064 26580 42116 26586
rect 42064 26522 42116 26528
rect 41326 26480 41382 26489
rect 41326 26415 41382 26424
rect 42260 26382 42288 26726
rect 44284 26586 44312 26794
rect 44456 26784 44508 26790
rect 44456 26726 44508 26732
rect 44468 26625 44496 26726
rect 44454 26616 44510 26625
rect 44272 26580 44324 26586
rect 44454 26551 44510 26560
rect 44272 26522 44324 26528
rect 44088 26512 44140 26518
rect 44088 26454 44140 26460
rect 41696 26376 41748 26382
rect 41696 26318 41748 26324
rect 42248 26376 42300 26382
rect 42248 26318 42300 26324
rect 43720 26376 43772 26382
rect 43720 26318 43772 26324
rect 41708 25974 41736 26318
rect 41696 25968 41748 25974
rect 41696 25910 41748 25916
rect 41512 25764 41564 25770
rect 41512 25706 41564 25712
rect 41524 25294 41552 25706
rect 41708 25294 41736 25910
rect 43732 25362 43760 26318
rect 44100 25945 44128 26454
rect 44086 25936 44142 25945
rect 44086 25871 44142 25880
rect 44180 25832 44232 25838
rect 44180 25774 44232 25780
rect 43720 25356 43772 25362
rect 43720 25298 43772 25304
rect 41512 25288 41564 25294
rect 41512 25230 41564 25236
rect 41696 25288 41748 25294
rect 41696 25230 41748 25236
rect 42800 25288 42852 25294
rect 42800 25230 42852 25236
rect 41602 24848 41658 24857
rect 41524 24792 41602 24800
rect 41524 24772 41604 24792
rect 41236 24744 41288 24750
rect 41236 24686 41288 24692
rect 41248 23662 41276 24686
rect 41236 23656 41288 23662
rect 41236 23598 41288 23604
rect 40684 23180 40736 23186
rect 40684 23122 40736 23128
rect 40776 23180 40828 23186
rect 40776 23122 40828 23128
rect 41144 23180 41196 23186
rect 41144 23122 41196 23128
rect 40408 22976 40460 22982
rect 40408 22918 40460 22924
rect 40420 22642 40448 22918
rect 40316 22636 40368 22642
rect 40316 22578 40368 22584
rect 40408 22636 40460 22642
rect 40408 22578 40460 22584
rect 40328 22166 40356 22578
rect 40316 22160 40368 22166
rect 40316 22102 40368 22108
rect 40328 21486 40356 22102
rect 40408 22024 40460 22030
rect 40408 21966 40460 21972
rect 40684 22024 40736 22030
rect 40788 22012 40816 23122
rect 41248 23118 41276 23598
rect 41524 23186 41552 24772
rect 41656 24783 41658 24792
rect 41604 24754 41656 24760
rect 41708 24732 41736 25230
rect 41972 24948 42024 24954
rect 41972 24890 42024 24896
rect 41880 24744 41932 24750
rect 41708 24704 41880 24732
rect 41604 24676 41656 24682
rect 41604 24618 41656 24624
rect 41616 23866 41644 24618
rect 41800 24206 41828 24704
rect 41880 24686 41932 24692
rect 41788 24200 41840 24206
rect 41788 24142 41840 24148
rect 41800 23866 41828 24142
rect 41880 24064 41932 24070
rect 41880 24006 41932 24012
rect 41604 23860 41656 23866
rect 41604 23802 41656 23808
rect 41788 23860 41840 23866
rect 41788 23802 41840 23808
rect 41892 23798 41920 24006
rect 41880 23792 41932 23798
rect 41880 23734 41932 23740
rect 41696 23520 41748 23526
rect 41696 23462 41748 23468
rect 41512 23180 41564 23186
rect 41512 23122 41564 23128
rect 41708 23118 41736 23462
rect 40868 23112 40920 23118
rect 40868 23054 40920 23060
rect 41236 23112 41288 23118
rect 41236 23054 41288 23060
rect 41696 23112 41748 23118
rect 41696 23054 41748 23060
rect 40880 22710 40908 23054
rect 40868 22704 40920 22710
rect 40868 22646 40920 22652
rect 41248 22234 41276 23054
rect 41788 22704 41840 22710
rect 41788 22646 41840 22652
rect 41878 22672 41934 22681
rect 41236 22228 41288 22234
rect 41236 22170 41288 22176
rect 40736 21984 40816 22012
rect 40684 21966 40736 21972
rect 40420 21554 40448 21966
rect 40408 21548 40460 21554
rect 40408 21490 40460 21496
rect 40316 21480 40368 21486
rect 40316 21422 40368 21428
rect 40328 21010 40356 21422
rect 40316 21004 40368 21010
rect 40316 20946 40368 20952
rect 40788 20534 40816 21984
rect 41328 21412 41380 21418
rect 41328 21354 41380 21360
rect 40776 20528 40828 20534
rect 40222 20496 40278 20505
rect 40776 20470 40828 20476
rect 40222 20431 40278 20440
rect 40776 19848 40828 19854
rect 40776 19790 40828 19796
rect 40408 19712 40460 19718
rect 40408 19654 40460 19660
rect 40420 19378 40448 19654
rect 40788 19514 40816 19790
rect 40776 19508 40828 19514
rect 40776 19450 40828 19456
rect 41052 19440 41104 19446
rect 41052 19382 41104 19388
rect 40316 19372 40368 19378
rect 40316 19314 40368 19320
rect 40408 19372 40460 19378
rect 40408 19314 40460 19320
rect 40052 19230 40172 19258
rect 40040 19168 40092 19174
rect 40040 19110 40092 19116
rect 40052 18902 40080 19110
rect 40040 18896 40092 18902
rect 40040 18838 40092 18844
rect 40144 18714 40172 19230
rect 40328 18766 40356 19314
rect 41064 18834 41092 19382
rect 41052 18828 41104 18834
rect 41052 18770 41104 18776
rect 40316 18760 40368 18766
rect 40052 18686 40172 18714
rect 40236 18720 40316 18748
rect 39580 18624 39632 18630
rect 39580 18566 39632 18572
rect 39592 17610 39620 18566
rect 40052 17882 40080 18686
rect 40132 18624 40184 18630
rect 40132 18566 40184 18572
rect 40040 17876 40092 17882
rect 40040 17818 40092 17824
rect 40144 17678 40172 18566
rect 39856 17672 39908 17678
rect 39856 17614 39908 17620
rect 40132 17672 40184 17678
rect 40132 17614 40184 17620
rect 39580 17604 39632 17610
rect 39580 17546 39632 17552
rect 39868 17270 39896 17614
rect 40236 17338 40264 18720
rect 40316 18702 40368 18708
rect 40868 18760 40920 18766
rect 40868 18702 40920 18708
rect 40880 18426 40908 18702
rect 41144 18692 41196 18698
rect 41340 18680 41368 21354
rect 41800 20874 41828 22646
rect 41878 22607 41934 22616
rect 41604 20868 41656 20874
rect 41604 20810 41656 20816
rect 41788 20868 41840 20874
rect 41788 20810 41840 20816
rect 41616 20602 41644 20810
rect 41604 20596 41656 20602
rect 41604 20538 41656 20544
rect 41800 20466 41828 20810
rect 41788 20460 41840 20466
rect 41788 20402 41840 20408
rect 41800 18970 41828 20402
rect 41788 18964 41840 18970
rect 41788 18906 41840 18912
rect 41196 18652 41368 18680
rect 41144 18634 41196 18640
rect 40868 18420 40920 18426
rect 40868 18362 40920 18368
rect 41340 18358 41368 18652
rect 41604 18692 41656 18698
rect 41604 18634 41656 18640
rect 41696 18692 41748 18698
rect 41696 18634 41748 18640
rect 41616 18426 41644 18634
rect 41604 18420 41656 18426
rect 41604 18362 41656 18368
rect 41328 18352 41380 18358
rect 41328 18294 41380 18300
rect 40316 18216 40368 18222
rect 40316 18158 40368 18164
rect 40328 17338 40356 18158
rect 41340 17678 41368 18294
rect 41708 18290 41736 18634
rect 41800 18290 41828 18906
rect 41892 18290 41920 22607
rect 41984 20466 42012 24890
rect 42432 23112 42484 23118
rect 42432 23054 42484 23060
rect 42444 22778 42472 23054
rect 42432 22772 42484 22778
rect 42432 22714 42484 22720
rect 42444 22642 42472 22714
rect 42432 22636 42484 22642
rect 42432 22578 42484 22584
rect 42812 21554 42840 25230
rect 43168 25220 43220 25226
rect 43168 25162 43220 25168
rect 42984 25152 43036 25158
rect 42984 25094 43036 25100
rect 43076 25152 43128 25158
rect 43076 25094 43128 25100
rect 42996 24818 43024 25094
rect 42984 24812 43036 24818
rect 42984 24754 43036 24760
rect 42996 24274 43024 24754
rect 43088 24614 43116 25094
rect 43076 24608 43128 24614
rect 43076 24550 43128 24556
rect 42984 24268 43036 24274
rect 42984 24210 43036 24216
rect 42984 24064 43036 24070
rect 42984 24006 43036 24012
rect 42996 23662 43024 24006
rect 43180 23866 43208 25162
rect 43732 24954 43760 25298
rect 43812 25220 43864 25226
rect 43812 25162 43864 25168
rect 43720 24948 43772 24954
rect 43720 24890 43772 24896
rect 43824 24857 43852 25162
rect 43810 24848 43866 24857
rect 43810 24783 43866 24792
rect 43628 24064 43680 24070
rect 43628 24006 43680 24012
rect 43168 23860 43220 23866
rect 43168 23802 43220 23808
rect 43640 23662 43668 24006
rect 43824 23730 43852 24783
rect 43812 23724 43864 23730
rect 43812 23666 43864 23672
rect 42984 23656 43036 23662
rect 42984 23598 43036 23604
rect 43628 23656 43680 23662
rect 43628 23598 43680 23604
rect 43536 23588 43588 23594
rect 43536 23530 43588 23536
rect 43548 22030 43576 23530
rect 44088 23520 44140 23526
rect 44088 23462 44140 23468
rect 44100 23225 44128 23462
rect 44086 23216 44142 23225
rect 44086 23151 44142 23160
rect 44192 22094 44220 25774
rect 44284 25294 44312 26522
rect 44272 25288 44324 25294
rect 44272 25230 44324 25236
rect 44454 25256 44510 25265
rect 44454 25191 44510 25200
rect 44468 25158 44496 25191
rect 44456 25152 44508 25158
rect 44456 25094 44508 25100
rect 44456 24608 44508 24614
rect 44454 24576 44456 24585
rect 44508 24576 44510 24585
rect 44454 24511 44510 24520
rect 44456 24064 44508 24070
rect 44456 24006 44508 24012
rect 44468 23905 44496 24006
rect 44454 23896 44510 23905
rect 44454 23831 44510 23840
rect 44454 22536 44510 22545
rect 44454 22471 44456 22480
rect 44508 22471 44510 22480
rect 44456 22442 44508 22448
rect 44192 22066 44312 22094
rect 43536 22024 43588 22030
rect 43536 21966 43588 21972
rect 43352 21956 43404 21962
rect 43352 21898 43404 21904
rect 43076 21888 43128 21894
rect 43076 21830 43128 21836
rect 43088 21554 43116 21830
rect 42800 21548 42852 21554
rect 42800 21490 42852 21496
rect 43076 21548 43128 21554
rect 43076 21490 43128 21496
rect 42616 20800 42668 20806
rect 42616 20742 42668 20748
rect 41972 20460 42024 20466
rect 41972 20402 42024 20408
rect 42628 20398 42656 20742
rect 42616 20392 42668 20398
rect 42616 20334 42668 20340
rect 42432 19372 42484 19378
rect 42432 19314 42484 19320
rect 42708 19372 42760 19378
rect 42708 19314 42760 19320
rect 41696 18284 41748 18290
rect 41696 18226 41748 18232
rect 41788 18284 41840 18290
rect 41788 18226 41840 18232
rect 41880 18284 41932 18290
rect 41880 18226 41932 18232
rect 41708 17814 41736 18226
rect 41800 18086 41828 18226
rect 41788 18080 41840 18086
rect 41788 18022 41840 18028
rect 41696 17808 41748 17814
rect 41696 17750 41748 17756
rect 41800 17678 41828 18022
rect 41328 17672 41380 17678
rect 41328 17614 41380 17620
rect 41788 17672 41840 17678
rect 41788 17614 41840 17620
rect 41800 17338 41828 17614
rect 40224 17332 40276 17338
rect 40224 17274 40276 17280
rect 40316 17332 40368 17338
rect 40316 17274 40368 17280
rect 41236 17332 41288 17338
rect 41236 17274 41288 17280
rect 41788 17332 41840 17338
rect 41788 17274 41840 17280
rect 39856 17264 39908 17270
rect 39856 17206 39908 17212
rect 39304 16720 39356 16726
rect 39026 16688 39082 16697
rect 38752 16652 38804 16658
rect 39304 16662 39356 16668
rect 39026 16623 39082 16632
rect 38752 16594 38804 16600
rect 38568 16516 38620 16522
rect 38568 16458 38620 16464
rect 38580 15502 38608 16458
rect 38764 16250 38792 16594
rect 40236 16590 40264 17274
rect 40328 16590 40356 17274
rect 41248 16998 41276 17274
rect 42444 17202 42472 19314
rect 42524 18624 42576 18630
rect 42524 18566 42576 18572
rect 42536 18222 42564 18566
rect 42524 18216 42576 18222
rect 42524 18158 42576 18164
rect 42524 18080 42576 18086
rect 42524 18022 42576 18028
rect 42536 17678 42564 18022
rect 42720 17814 42748 19314
rect 42708 17808 42760 17814
rect 42708 17750 42760 17756
rect 42524 17672 42576 17678
rect 42524 17614 42576 17620
rect 42708 17536 42760 17542
rect 42708 17478 42760 17484
rect 42720 17202 42748 17478
rect 42432 17196 42484 17202
rect 42432 17138 42484 17144
rect 42708 17196 42760 17202
rect 42708 17138 42760 17144
rect 41236 16992 41288 16998
rect 41236 16934 41288 16940
rect 40224 16584 40276 16590
rect 40224 16526 40276 16532
rect 40316 16584 40368 16590
rect 40316 16526 40368 16532
rect 38752 16244 38804 16250
rect 38752 16186 38804 16192
rect 39028 16108 39080 16114
rect 39028 16050 39080 16056
rect 38660 16040 38712 16046
rect 38660 15982 38712 15988
rect 38568 15496 38620 15502
rect 38568 15438 38620 15444
rect 38672 15366 38700 15982
rect 38660 15360 38712 15366
rect 38660 15302 38712 15308
rect 39040 15162 39068 16050
rect 40236 15502 40264 16526
rect 41248 15502 41276 16934
rect 42444 16522 42472 17138
rect 42432 16516 42484 16522
rect 42432 16458 42484 16464
rect 42444 15586 42472 16458
rect 42812 16182 42840 21490
rect 43364 21078 43392 21898
rect 43548 21690 43576 21966
rect 43536 21684 43588 21690
rect 43536 21626 43588 21632
rect 44180 21548 44232 21554
rect 44180 21490 44232 21496
rect 43904 21412 43956 21418
rect 43904 21354 43956 21360
rect 43812 21344 43864 21350
rect 43812 21286 43864 21292
rect 43824 21146 43852 21286
rect 43812 21140 43864 21146
rect 43812 21082 43864 21088
rect 43352 21072 43404 21078
rect 43352 21014 43404 21020
rect 43916 20942 43944 21354
rect 43260 20936 43312 20942
rect 43260 20878 43312 20884
rect 43904 20936 43956 20942
rect 43904 20878 43956 20884
rect 43272 19854 43300 20878
rect 44088 20800 44140 20806
rect 44088 20742 44140 20748
rect 44100 20505 44128 20742
rect 44086 20496 44142 20505
rect 44086 20431 44142 20440
rect 44192 19922 44220 21490
rect 44284 20942 44312 22066
rect 44456 21888 44508 21894
rect 44454 21856 44456 21865
rect 44508 21856 44510 21865
rect 44454 21791 44510 21800
rect 44456 21344 44508 21350
rect 44456 21286 44508 21292
rect 44468 21185 44496 21286
rect 44454 21176 44510 21185
rect 44454 21111 44510 21120
rect 44272 20936 44324 20942
rect 44272 20878 44324 20884
rect 44180 19916 44232 19922
rect 44180 19858 44232 19864
rect 43260 19848 43312 19854
rect 43260 19790 43312 19796
rect 44454 19816 44510 19825
rect 44454 19751 44510 19760
rect 44468 19718 44496 19751
rect 44456 19712 44508 19718
rect 44456 19654 44508 19660
rect 44088 19508 44140 19514
rect 44088 19450 44140 19456
rect 43812 19236 43864 19242
rect 43812 19178 43864 19184
rect 43824 18834 43852 19178
rect 44100 19145 44128 19450
rect 44086 19136 44142 19145
rect 44086 19071 44142 19080
rect 43812 18828 43864 18834
rect 43812 18770 43864 18776
rect 43168 18760 43220 18766
rect 43168 18702 43220 18708
rect 43180 18290 43208 18702
rect 43260 18624 43312 18630
rect 43260 18566 43312 18572
rect 44456 18624 44508 18630
rect 44456 18566 44508 18572
rect 43168 18284 43220 18290
rect 43168 18226 43220 18232
rect 43272 17882 43300 18566
rect 44468 18465 44496 18566
rect 44454 18456 44510 18465
rect 44454 18391 44510 18400
rect 44088 18080 44140 18086
rect 44088 18022 44140 18028
rect 43260 17876 43312 17882
rect 43260 17818 43312 17824
rect 44100 17785 44128 18022
rect 44086 17776 44142 17785
rect 44086 17711 44142 17720
rect 43812 17672 43864 17678
rect 43812 17614 43864 17620
rect 43824 17338 43852 17614
rect 43812 17332 43864 17338
rect 43812 17274 43864 17280
rect 44454 17096 44510 17105
rect 44454 17031 44456 17040
rect 44508 17031 44510 17040
rect 44456 17002 44508 17008
rect 44456 16448 44508 16454
rect 44454 16416 44456 16425
rect 44508 16416 44510 16425
rect 44454 16351 44510 16360
rect 42800 16176 42852 16182
rect 42800 16118 42852 16124
rect 44272 15972 44324 15978
rect 44272 15914 44324 15920
rect 41420 15564 41472 15570
rect 41420 15506 41472 15512
rect 42352 15558 42472 15586
rect 40224 15496 40276 15502
rect 40224 15438 40276 15444
rect 41236 15496 41288 15502
rect 41236 15438 41288 15444
rect 41432 15162 41460 15506
rect 42352 15502 42380 15558
rect 42340 15496 42392 15502
rect 42340 15438 42392 15444
rect 43076 15360 43128 15366
rect 43076 15302 43128 15308
rect 44088 15360 44140 15366
rect 44088 15302 44140 15308
rect 39028 15156 39080 15162
rect 39028 15098 39080 15104
rect 41420 15156 41472 15162
rect 41420 15098 41472 15104
rect 43088 14958 43116 15302
rect 44100 15065 44128 15302
rect 44086 15056 44142 15065
rect 44086 14991 44142 15000
rect 43076 14952 43128 14958
rect 43076 14894 43128 14900
rect 43088 13938 43116 14894
rect 44284 14414 44312 15914
rect 44456 15904 44508 15910
rect 44456 15846 44508 15852
rect 44468 15745 44496 15846
rect 44454 15736 44510 15745
rect 44454 15671 44510 15680
rect 44272 14408 44324 14414
rect 44272 14350 44324 14356
rect 44454 14376 44510 14385
rect 44454 14311 44510 14320
rect 44468 14278 44496 14311
rect 44456 14272 44508 14278
rect 44456 14214 44508 14220
rect 44088 14068 44140 14074
rect 44088 14010 44140 14016
rect 43076 13932 43128 13938
rect 43076 13874 43128 13880
rect 44100 13705 44128 14010
rect 44086 13696 44142 13705
rect 44086 13631 44142 13640
rect 37924 13388 37976 13394
rect 37924 13330 37976 13336
rect 37556 13184 37608 13190
rect 37556 13126 37608 13132
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 31668 12776 31720 12782
rect 31668 12718 31720 12724
rect 31024 12640 31076 12646
rect 31024 12582 31076 12588
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 30288 12436 30340 12442
rect 30288 12378 30340 12384
rect 29090 12200 29146 12209
rect 29090 12135 29146 12144
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 27618 10976 27674 10985
rect 4874 10908 5182 10917
rect 27618 10911 27674 10920
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 2502 19352 2558 19408
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4342 22616 4398 22672
rect 846 16532 848 16552
rect 848 16532 900 16552
rect 900 16532 902 16552
rect 846 16496 902 16532
rect 846 15816 902 15872
rect 1398 15000 1454 15056
rect 846 14456 902 14512
rect 1398 13640 1454 13696
rect 1398 12960 1454 13016
rect 846 12164 902 12200
rect 846 12144 848 12164
rect 848 12144 900 12164
rect 900 12144 902 12164
rect 3146 13232 3202 13288
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 5446 25900 5502 25936
rect 5446 25880 5448 25900
rect 5448 25880 5500 25900
rect 5500 25880 5502 25900
rect 6090 25336 6146 25392
rect 5538 23704 5594 23760
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 5170 22636 5226 22672
rect 5170 22616 5172 22636
rect 5172 22616 5224 22636
rect 5224 22616 5226 22636
rect 5078 22380 5080 22400
rect 5080 22380 5132 22400
rect 5132 22380 5134 22400
rect 5078 22344 5134 22380
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 5262 21528 5318 21584
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 5814 22636 5870 22672
rect 5814 22616 5816 22636
rect 5816 22616 5868 22636
rect 5868 22616 5870 22636
rect 5446 21528 5502 21584
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 5446 19080 5502 19136
rect 3698 16632 3754 16688
rect 4618 18400 4674 18456
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4894 18264 4950 18320
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4986 17212 4988 17232
rect 4988 17212 5040 17232
rect 5040 17212 5042 17232
rect 4986 17176 5042 17212
rect 4894 16632 4950 16688
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 5998 20204 6000 20224
rect 6000 20204 6052 20224
rect 6052 20204 6054 20224
rect 5998 20168 6054 20204
rect 5722 19624 5778 19680
rect 7654 29416 7710 29472
rect 6826 27940 6882 27976
rect 6826 27920 6828 27940
rect 6828 27920 6880 27940
rect 6880 27920 6882 27940
rect 6734 27668 6790 27704
rect 6734 27648 6736 27668
rect 6736 27648 6788 27668
rect 6788 27648 6790 27668
rect 6918 26424 6974 26480
rect 7010 21120 7066 21176
rect 5538 15544 5594 15600
rect 5078 13404 5080 13424
rect 5080 13404 5132 13424
rect 5132 13404 5134 13424
rect 5078 13368 5134 13404
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 6182 14592 6238 14648
rect 10046 30096 10102 30152
rect 8114 27376 8170 27432
rect 7930 24928 7986 24984
rect 8206 25644 8208 25664
rect 8208 25644 8260 25664
rect 8260 25644 8262 25664
rect 8206 25608 8262 25644
rect 8390 26868 8392 26888
rect 8392 26868 8444 26888
rect 8444 26868 8446 26888
rect 8390 26832 8446 26868
rect 8022 23840 8078 23896
rect 7930 23568 7986 23624
rect 7838 23468 7840 23488
rect 7840 23468 7892 23488
rect 7892 23468 7894 23488
rect 7838 23432 7894 23468
rect 7470 21936 7526 21992
rect 7102 18672 7158 18728
rect 7010 18536 7066 18592
rect 6918 17756 6920 17776
rect 6920 17756 6972 17776
rect 6972 17756 6974 17776
rect 6918 17720 6974 17756
rect 6642 17448 6698 17504
rect 6642 15952 6698 16008
rect 6734 15444 6736 15464
rect 6736 15444 6788 15464
rect 6788 15444 6790 15464
rect 6734 15408 6790 15444
rect 7286 16632 7342 16688
rect 7470 21392 7526 21448
rect 7930 23024 7986 23080
rect 7654 18672 7710 18728
rect 8206 20748 8208 20768
rect 8208 20748 8260 20768
rect 8260 20748 8262 20768
rect 8206 20712 8262 20748
rect 7930 18400 7986 18456
rect 7930 17720 7986 17776
rect 8298 19760 8354 19816
rect 8758 24692 8760 24712
rect 8760 24692 8812 24712
rect 8812 24692 8814 24712
rect 8758 24656 8814 24692
rect 8298 19216 8354 19272
rect 8482 18148 8538 18184
rect 8482 18128 8484 18148
rect 8484 18128 8536 18148
rect 8536 18128 8538 18148
rect 8114 17312 8170 17368
rect 7378 15444 7380 15464
rect 7380 15444 7432 15464
rect 7432 15444 7434 15464
rect 7378 15408 7434 15444
rect 7562 16516 7618 16552
rect 7562 16496 7564 16516
rect 7564 16496 7616 16516
rect 7616 16496 7618 16516
rect 7470 13368 7526 13424
rect 8666 18808 8722 18864
rect 9126 22516 9128 22536
rect 9128 22516 9180 22536
rect 9180 22516 9182 22536
rect 9586 27104 9642 27160
rect 10046 28056 10102 28112
rect 9586 24384 9642 24440
rect 9770 24248 9826 24304
rect 10506 30232 10562 30288
rect 10782 28872 10838 28928
rect 10414 28328 10470 28384
rect 10322 28056 10378 28112
rect 10598 28192 10654 28248
rect 10322 26560 10378 26616
rect 10322 26324 10324 26344
rect 10324 26324 10376 26344
rect 10376 26324 10378 26344
rect 10322 26288 10378 26324
rect 9954 24556 9956 24576
rect 9956 24556 10008 24576
rect 10008 24556 10010 24576
rect 9954 24520 10010 24556
rect 9678 23976 9734 24032
rect 9126 22480 9182 22516
rect 8850 21392 8906 21448
rect 9034 20848 9090 20904
rect 8850 20576 8906 20632
rect 8850 19352 8906 19408
rect 9034 18808 9090 18864
rect 8942 18400 8998 18456
rect 8850 17992 8906 18048
rect 8574 16668 8576 16688
rect 8576 16668 8628 16688
rect 8628 16668 8630 16688
rect 8574 16632 8630 16668
rect 8942 17720 8998 17776
rect 7930 14048 7986 14104
rect 7930 13640 7986 13696
rect 8758 16108 8814 16144
rect 8758 16088 8760 16108
rect 8760 16088 8812 16108
rect 8812 16088 8814 16108
rect 8850 13912 8906 13968
rect 9402 20304 9458 20360
rect 9402 20052 9458 20088
rect 9402 20032 9404 20052
rect 9404 20032 9456 20052
rect 9456 20032 9458 20052
rect 9678 21800 9734 21856
rect 10598 24928 10654 24984
rect 11150 31048 11206 31104
rect 11058 29588 11060 29608
rect 11060 29588 11112 29608
rect 11112 29588 11114 29608
rect 11058 29552 11114 29588
rect 11334 28464 11390 28520
rect 11150 26152 11206 26208
rect 10782 24792 10838 24848
rect 10414 24112 10470 24168
rect 10690 24268 10746 24304
rect 10690 24248 10692 24268
rect 10692 24248 10744 24268
rect 10744 24248 10746 24268
rect 10230 22616 10286 22672
rect 9678 20984 9734 21040
rect 9586 20576 9642 20632
rect 10046 20304 10102 20360
rect 9586 19896 9642 19952
rect 9770 19916 9826 19952
rect 9770 19896 9772 19916
rect 9772 19896 9824 19916
rect 9824 19896 9826 19916
rect 9218 18400 9274 18456
rect 9034 15680 9090 15736
rect 9402 16360 9458 16416
rect 9862 18964 9918 19000
rect 9862 18944 9864 18964
rect 9864 18944 9916 18964
rect 9916 18944 9918 18964
rect 9954 18264 10010 18320
rect 9954 17876 10010 17912
rect 9954 17856 9956 17876
rect 9956 17856 10008 17876
rect 10008 17856 10010 17876
rect 9678 16360 9734 16416
rect 9126 14728 9182 14784
rect 10230 21292 10232 21312
rect 10232 21292 10284 21312
rect 10284 21292 10286 21312
rect 10230 21256 10286 21292
rect 10506 20440 10562 20496
rect 10506 20324 10562 20360
rect 10506 20304 10508 20324
rect 10508 20304 10560 20324
rect 10560 20304 10562 20324
rect 10506 19896 10562 19952
rect 9954 15952 10010 16008
rect 10046 15816 10102 15872
rect 10414 17720 10470 17776
rect 10506 17584 10562 17640
rect 10874 23840 10930 23896
rect 10782 22888 10838 22944
rect 11058 22344 11114 22400
rect 11058 21936 11114 21992
rect 10690 18300 10692 18320
rect 10692 18300 10744 18320
rect 10744 18300 10746 18320
rect 10690 18264 10746 18300
rect 10414 17040 10470 17096
rect 10230 15972 10286 16008
rect 10230 15952 10232 15972
rect 10232 15952 10284 15972
rect 10284 15952 10286 15972
rect 10598 16360 10654 16416
rect 10690 16224 10746 16280
rect 10138 15408 10194 15464
rect 9126 14184 9182 14240
rect 8666 13504 8722 13560
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 846 11756 902 11792
rect 846 11736 848 11756
rect 848 11736 900 11756
rect 900 11736 902 11756
rect 8666 12824 8722 12880
rect 9126 13504 9182 13560
rect 9678 14048 9734 14104
rect 10966 17720 11022 17776
rect 11058 17176 11114 17232
rect 10966 16904 11022 16960
rect 11058 16768 11114 16824
rect 11702 26016 11758 26072
rect 11978 29144 12034 29200
rect 11978 26560 12034 26616
rect 12622 27512 12678 27568
rect 11794 24556 11796 24576
rect 11796 24556 11848 24576
rect 11848 24556 11850 24576
rect 11794 24520 11850 24556
rect 11518 22072 11574 22128
rect 11610 21936 11666 21992
rect 11610 21664 11666 21720
rect 11610 20984 11666 21040
rect 11518 20168 11574 20224
rect 11334 17176 11390 17232
rect 10782 15680 10838 15736
rect 10966 15680 11022 15736
rect 10782 15308 10784 15328
rect 10784 15308 10836 15328
rect 10836 15308 10838 15328
rect 10782 15272 10838 15308
rect 11058 15156 11114 15192
rect 11058 15136 11060 15156
rect 11060 15136 11112 15156
rect 11112 15136 11114 15156
rect 11150 15000 11206 15056
rect 10690 13096 10746 13152
rect 10782 12588 10784 12608
rect 10784 12588 10836 12608
rect 10836 12588 10838 12608
rect 10782 12552 10838 12588
rect 11150 12688 11206 12744
rect 11702 20712 11758 20768
rect 11702 18808 11758 18864
rect 11702 18264 11758 18320
rect 11518 16360 11574 16416
rect 11978 23432 12034 23488
rect 11886 23296 11942 23352
rect 13634 32272 13690 32328
rect 13450 31456 13506 31512
rect 13266 29044 13268 29064
rect 13268 29044 13320 29064
rect 13320 29044 13322 29064
rect 13266 29008 13322 29044
rect 13082 28908 13084 28928
rect 13084 28908 13136 28928
rect 13136 28908 13138 28928
rect 13082 28872 13138 28908
rect 12898 24148 12900 24168
rect 12900 24148 12952 24168
rect 12952 24148 12954 24168
rect 12898 24112 12954 24148
rect 13266 26988 13322 27024
rect 13266 26968 13268 26988
rect 13268 26968 13320 26988
rect 13320 26968 13322 26988
rect 13266 25644 13268 25664
rect 13268 25644 13320 25664
rect 13320 25644 13322 25664
rect 13266 25608 13322 25644
rect 13726 29960 13782 30016
rect 13542 29008 13598 29064
rect 13174 24520 13230 24576
rect 13174 24248 13230 24304
rect 11978 21256 12034 21312
rect 11978 20748 11980 20768
rect 11980 20748 12032 20768
rect 12032 20748 12034 20768
rect 11978 20712 12034 20748
rect 12438 22636 12494 22672
rect 13174 23160 13230 23216
rect 12438 22616 12440 22636
rect 12440 22616 12492 22636
rect 12492 22616 12494 22636
rect 12530 21392 12586 21448
rect 12346 21256 12402 21312
rect 12254 21020 12256 21040
rect 12256 21020 12308 21040
rect 12308 21020 12310 21040
rect 12254 20984 12310 21020
rect 12530 20984 12586 21040
rect 11978 19216 12034 19272
rect 11978 16360 12034 16416
rect 11794 13640 11850 13696
rect 12162 15000 12218 15056
rect 11978 13932 12034 13968
rect 11978 13912 11980 13932
rect 11980 13912 12032 13932
rect 12032 13912 12034 13932
rect 12070 13776 12126 13832
rect 13082 21256 13138 21312
rect 13358 22772 13414 22808
rect 13358 22752 13360 22772
rect 13360 22752 13412 22772
rect 13412 22752 13414 22772
rect 13266 21392 13322 21448
rect 13358 21256 13414 21312
rect 13818 28600 13874 28656
rect 13726 28192 13782 28248
rect 13634 27820 13636 27840
rect 13636 27820 13688 27840
rect 13688 27820 13690 27840
rect 13634 27784 13690 27820
rect 13634 27104 13690 27160
rect 13634 24248 13690 24304
rect 12990 20984 13046 21040
rect 12622 20748 12624 20768
rect 12624 20748 12676 20768
rect 12676 20748 12678 20768
rect 12622 20712 12678 20748
rect 12806 20712 12862 20768
rect 12898 19488 12954 19544
rect 12714 19216 12770 19272
rect 12898 18944 12954 19000
rect 13174 20576 13230 20632
rect 13358 20984 13414 21040
rect 13450 20712 13506 20768
rect 13082 20460 13138 20496
rect 13082 20440 13084 20460
rect 13084 20440 13136 20460
rect 13136 20440 13138 20460
rect 12990 17720 13046 17776
rect 12806 17584 12862 17640
rect 12530 17176 12586 17232
rect 12438 14048 12494 14104
rect 12254 13368 12310 13424
rect 11610 12980 11666 13016
rect 11610 12960 11612 12980
rect 11612 12960 11664 12980
rect 11664 12960 11666 12980
rect 11610 12416 11666 12472
rect 12990 17196 13046 17232
rect 12990 17176 12992 17196
rect 12992 17176 13044 17196
rect 13044 17176 13046 17196
rect 12898 15816 12954 15872
rect 12714 15444 12716 15464
rect 12716 15444 12768 15464
rect 12768 15444 12770 15464
rect 12714 15408 12770 15444
rect 12806 15136 12862 15192
rect 12990 15408 13046 15464
rect 13266 19488 13322 19544
rect 13910 23840 13966 23896
rect 13818 23568 13874 23624
rect 13818 22344 13874 22400
rect 14278 28872 14334 28928
rect 14554 31340 14610 31376
rect 14554 31320 14556 31340
rect 14556 31320 14608 31340
rect 14608 31320 14610 31340
rect 14462 30504 14518 30560
rect 14370 24656 14426 24712
rect 14278 24132 14334 24168
rect 14278 24112 14280 24132
rect 14280 24112 14332 24132
rect 14332 24112 14334 24132
rect 13818 22072 13874 22128
rect 13726 21936 13782 21992
rect 14186 23296 14242 23352
rect 14186 22752 14242 22808
rect 13266 17312 13322 17368
rect 13082 13912 13138 13968
rect 12530 12688 12586 12744
rect 12990 12688 13046 12744
rect 13266 15852 13268 15872
rect 13268 15852 13320 15872
rect 13320 15852 13322 15872
rect 13266 15816 13322 15852
rect 13266 14456 13322 14512
rect 13542 17312 13598 17368
rect 14094 19488 14150 19544
rect 13726 17756 13728 17776
rect 13728 17756 13780 17776
rect 13780 17756 13782 17776
rect 13726 17720 13782 17756
rect 13818 16768 13874 16824
rect 13910 16360 13966 16416
rect 13266 13232 13322 13288
rect 13634 13096 13690 13152
rect 13450 12708 13506 12744
rect 13450 12688 13452 12708
rect 13452 12688 13504 12708
rect 13504 12688 13506 12708
rect 15842 32136 15898 32192
rect 15474 31184 15530 31240
rect 15198 30912 15254 30968
rect 15014 28076 15070 28112
rect 15014 28056 15016 28076
rect 15016 28056 15068 28076
rect 15068 28056 15070 28076
rect 15198 26560 15254 26616
rect 15474 30368 15530 30424
rect 15474 30232 15530 30288
rect 15474 28076 15530 28112
rect 15474 28056 15476 28076
rect 15476 28056 15528 28076
rect 15528 28056 15530 28076
rect 14830 26152 14886 26208
rect 14646 22616 14702 22672
rect 14462 21392 14518 21448
rect 15106 25764 15162 25800
rect 15106 25744 15108 25764
rect 15108 25744 15160 25764
rect 15160 25744 15162 25764
rect 15474 26324 15476 26344
rect 15476 26324 15528 26344
rect 15528 26324 15530 26344
rect 15474 26288 15530 26324
rect 15106 24148 15108 24168
rect 15108 24148 15160 24168
rect 15160 24148 15162 24168
rect 15106 24112 15162 24148
rect 15198 23060 15200 23080
rect 15200 23060 15252 23080
rect 15252 23060 15254 23080
rect 15198 23024 15254 23060
rect 14922 21972 14924 21992
rect 14924 21972 14976 21992
rect 14976 21972 14978 21992
rect 14922 21936 14978 21972
rect 14738 21800 14794 21856
rect 14922 21664 14978 21720
rect 14370 19488 14426 19544
rect 15750 30252 15806 30288
rect 15750 30232 15752 30252
rect 15752 30232 15804 30252
rect 15804 30232 15806 30252
rect 15842 27376 15898 27432
rect 15658 23860 15714 23896
rect 15658 23840 15660 23860
rect 15660 23840 15712 23860
rect 15712 23840 15714 23860
rect 15934 26968 15990 27024
rect 17682 32020 17738 32056
rect 17682 32000 17684 32020
rect 17684 32000 17736 32020
rect 17736 32000 17738 32020
rect 16762 30368 16818 30424
rect 16762 29572 16818 29608
rect 16762 29552 16764 29572
rect 16764 29552 16816 29572
rect 16816 29552 16818 29572
rect 16210 26016 16266 26072
rect 16118 25472 16174 25528
rect 15934 24928 15990 24984
rect 14922 18284 14978 18320
rect 14922 18264 14924 18284
rect 14924 18264 14976 18284
rect 14976 18264 14978 18284
rect 14646 16768 14702 16824
rect 14738 15952 14794 16008
rect 15106 19352 15162 19408
rect 15106 17992 15162 18048
rect 15750 21392 15806 21448
rect 15198 17584 15254 17640
rect 15106 17448 15162 17504
rect 15014 16632 15070 16688
rect 16302 25220 16358 25256
rect 16302 25200 16304 25220
rect 16304 25200 16356 25220
rect 16356 25200 16358 25220
rect 16578 23976 16634 24032
rect 15198 16224 15254 16280
rect 15198 14592 15254 14648
rect 15198 13096 15254 13152
rect 14738 12688 14794 12744
rect 16486 22092 16542 22128
rect 16486 22072 16488 22092
rect 16488 22072 16540 22092
rect 16540 22072 16542 22092
rect 16486 20304 16542 20360
rect 16026 16360 16082 16416
rect 16210 15972 16266 16008
rect 16210 15952 16212 15972
rect 16212 15952 16264 15972
rect 16264 15952 16266 15972
rect 16394 16496 16450 16552
rect 16210 14728 16266 14784
rect 16394 13096 16450 13152
rect 17130 31456 17186 31512
rect 16854 22208 16910 22264
rect 16946 21664 17002 21720
rect 16854 20576 16910 20632
rect 17406 29824 17462 29880
rect 17314 29008 17370 29064
rect 17222 28056 17278 28112
rect 17222 27648 17278 27704
rect 17590 30096 17646 30152
rect 17590 29552 17646 29608
rect 17314 26560 17370 26616
rect 17406 26288 17462 26344
rect 17222 20884 17224 20904
rect 17224 20884 17276 20904
rect 17276 20884 17278 20904
rect 17222 20848 17278 20884
rect 17130 18808 17186 18864
rect 17038 18536 17094 18592
rect 17682 24812 17738 24848
rect 17682 24792 17684 24812
rect 17684 24792 17736 24812
rect 17736 24792 17738 24812
rect 18050 30096 18106 30152
rect 17866 27648 17922 27704
rect 17866 27104 17922 27160
rect 17590 21936 17646 21992
rect 17590 20884 17592 20904
rect 17592 20884 17644 20904
rect 17644 20884 17646 20904
rect 17590 20848 17646 20884
rect 17498 18808 17554 18864
rect 18050 24520 18106 24576
rect 18234 24676 18290 24712
rect 18234 24656 18236 24676
rect 18236 24656 18288 24676
rect 18288 24656 18290 24676
rect 17958 22888 18014 22944
rect 18786 30504 18842 30560
rect 18694 30096 18750 30152
rect 18878 29824 18934 29880
rect 18694 29688 18750 29744
rect 19430 31864 19486 31920
rect 19246 30912 19302 30968
rect 19982 31864 20038 31920
rect 19614 31628 19616 31648
rect 19616 31628 19668 31648
rect 19668 31628 19670 31648
rect 19614 31592 19670 31628
rect 19062 29688 19118 29744
rect 18970 29008 19026 29064
rect 18418 26288 18474 26344
rect 19062 28328 19118 28384
rect 19246 29008 19302 29064
rect 18786 27240 18842 27296
rect 19062 26560 19118 26616
rect 18142 20712 18198 20768
rect 18326 21528 18382 21584
rect 18510 24520 18566 24576
rect 18602 23432 18658 23488
rect 18234 20304 18290 20360
rect 18234 19624 18290 19680
rect 17498 18264 17554 18320
rect 16762 15136 16818 15192
rect 16670 14592 16726 14648
rect 17406 16768 17462 16824
rect 17314 16108 17370 16144
rect 17314 16088 17316 16108
rect 17316 16088 17368 16108
rect 17368 16088 17370 16108
rect 18050 17992 18106 18048
rect 18142 15680 18198 15736
rect 18050 15136 18106 15192
rect 17406 14048 17462 14104
rect 17222 13232 17278 13288
rect 16486 12552 16542 12608
rect 17682 13368 17738 13424
rect 18510 20304 18566 20360
rect 18510 19488 18566 19544
rect 18878 23160 18934 23216
rect 18878 22752 18934 22808
rect 18786 20032 18842 20088
rect 18970 20052 19026 20088
rect 18970 20032 18972 20052
rect 18972 20032 19024 20052
rect 19024 20032 19026 20052
rect 18878 19372 18934 19408
rect 18878 19352 18880 19372
rect 18880 19352 18932 19372
rect 18932 19352 18934 19372
rect 18326 16496 18382 16552
rect 18418 15816 18474 15872
rect 18602 18128 18658 18184
rect 18878 17176 18934 17232
rect 18878 16904 18934 16960
rect 18694 16360 18750 16416
rect 18510 15544 18566 15600
rect 18878 15544 18934 15600
rect 18786 15408 18842 15464
rect 18878 15136 18934 15192
rect 18510 13368 18566 13424
rect 18234 12960 18290 13016
rect 17682 12708 17738 12744
rect 17682 12688 17684 12708
rect 17684 12688 17736 12708
rect 17736 12688 17738 12708
rect 19338 27668 19394 27704
rect 19338 27648 19340 27668
rect 19340 27648 19392 27668
rect 19392 27648 19394 27668
rect 19982 30776 20038 30832
rect 19706 29280 19762 29336
rect 19798 28736 19854 28792
rect 19706 27124 19762 27160
rect 19706 27104 19708 27124
rect 19708 27104 19760 27124
rect 19760 27104 19762 27124
rect 19522 25492 19578 25528
rect 19522 25472 19524 25492
rect 19524 25472 19576 25492
rect 19576 25472 19578 25492
rect 19338 25336 19394 25392
rect 19338 25064 19394 25120
rect 19338 23024 19394 23080
rect 19338 22480 19394 22536
rect 20442 30540 20444 30560
rect 20444 30540 20496 30560
rect 20496 30540 20498 30560
rect 20442 30504 20498 30540
rect 19982 27396 20038 27432
rect 19982 27376 19984 27396
rect 19984 27376 20036 27396
rect 20036 27376 20038 27396
rect 19614 24928 19670 24984
rect 19890 25064 19946 25120
rect 19522 23432 19578 23488
rect 19706 23432 19762 23488
rect 19798 22752 19854 22808
rect 19154 17196 19210 17232
rect 19154 17176 19156 17196
rect 19156 17176 19208 17196
rect 19208 17176 19210 17196
rect 19338 17040 19394 17096
rect 20166 25336 20222 25392
rect 20626 29572 20682 29608
rect 20626 29552 20628 29572
rect 20628 29552 20680 29572
rect 20680 29552 20682 29572
rect 20626 26696 20682 26752
rect 19522 19236 19578 19272
rect 19522 19216 19524 19236
rect 19524 19216 19576 19236
rect 19576 19216 19578 19236
rect 19614 18284 19670 18320
rect 19614 18264 19616 18284
rect 19616 18264 19668 18284
rect 19668 18264 19670 18284
rect 19246 15680 19302 15736
rect 19798 18400 19854 18456
rect 19798 17992 19854 18048
rect 20166 19508 20222 19544
rect 20166 19488 20168 19508
rect 20168 19488 20220 19508
rect 20220 19488 20222 19508
rect 20166 19252 20168 19272
rect 20168 19252 20220 19272
rect 20220 19252 20222 19272
rect 20166 19216 20222 19252
rect 20166 18944 20222 19000
rect 22558 32136 22614 32192
rect 22558 31728 22614 31784
rect 21730 31048 21786 31104
rect 21086 29588 21088 29608
rect 21088 29588 21140 29608
rect 21140 29588 21142 29608
rect 21086 29552 21142 29588
rect 20902 26696 20958 26752
rect 20718 25744 20774 25800
rect 20534 23044 20590 23080
rect 20534 23024 20536 23044
rect 20536 23024 20588 23044
rect 20588 23024 20590 23044
rect 20626 22072 20682 22128
rect 20902 22888 20958 22944
rect 20810 22752 20866 22808
rect 20810 22072 20866 22128
rect 21178 23704 21234 23760
rect 21086 22208 21142 22264
rect 21086 21936 21142 21992
rect 20350 16108 20406 16144
rect 20350 16088 20352 16108
rect 20352 16088 20404 16108
rect 20404 16088 20406 16108
rect 19982 15272 20038 15328
rect 20350 14592 20406 14648
rect 20718 18400 20774 18456
rect 20534 14356 20536 14376
rect 20536 14356 20588 14376
rect 20588 14356 20590 14376
rect 20534 14320 20590 14356
rect 20166 13776 20222 13832
rect 20350 13640 20406 13696
rect 21086 21256 21142 21312
rect 20994 19896 21050 19952
rect 21914 29144 21970 29200
rect 21822 27648 21878 27704
rect 21270 19896 21326 19952
rect 21178 19216 21234 19272
rect 21086 18264 21142 18320
rect 20994 15816 21050 15872
rect 20994 15408 21050 15464
rect 22190 28328 22246 28384
rect 22190 26968 22246 27024
rect 22466 30776 22522 30832
rect 22374 29824 22430 29880
rect 22650 29960 22706 30016
rect 22098 24520 22154 24576
rect 22098 24248 22154 24304
rect 22282 23976 22338 24032
rect 22282 23588 22338 23624
rect 22282 23568 22284 23588
rect 22284 23568 22336 23588
rect 22336 23568 22338 23588
rect 22282 23432 22338 23488
rect 23294 32000 23350 32056
rect 24766 33224 24822 33280
rect 23938 31764 23940 31784
rect 23940 31764 23992 31784
rect 23992 31764 23994 31784
rect 23938 31728 23994 31764
rect 23386 30096 23442 30152
rect 22834 25880 22890 25936
rect 22558 24384 22614 24440
rect 22466 23432 22522 23488
rect 22374 22208 22430 22264
rect 22098 19624 22154 19680
rect 22650 23704 22706 23760
rect 22650 20204 22652 20224
rect 22652 20204 22704 20224
rect 22704 20204 22706 20224
rect 22650 20168 22706 20204
rect 22650 19488 22706 19544
rect 22282 18944 22338 19000
rect 22190 18672 22246 18728
rect 22466 18944 22522 19000
rect 22190 17856 22246 17912
rect 22466 18400 22522 18456
rect 22374 17448 22430 17504
rect 21362 15816 21418 15872
rect 22098 15952 22154 16008
rect 22098 15544 22154 15600
rect 22098 15272 22154 15328
rect 22006 14320 22062 14376
rect 22650 18148 22706 18184
rect 22650 18128 22652 18148
rect 22652 18128 22704 18148
rect 22704 18128 22706 18148
rect 22926 24520 22982 24576
rect 23386 28620 23442 28656
rect 23386 28600 23388 28620
rect 23388 28600 23440 28620
rect 23440 28600 23442 28620
rect 23386 27920 23442 27976
rect 23478 26560 23534 26616
rect 22834 24248 22890 24304
rect 23018 24248 23074 24304
rect 22926 23160 22982 23216
rect 22834 20848 22890 20904
rect 22834 18400 22890 18456
rect 22282 15952 22338 16008
rect 22466 15816 22522 15872
rect 22650 15816 22706 15872
rect 22282 15428 22338 15464
rect 22282 15408 22284 15428
rect 22284 15408 22336 15428
rect 22336 15408 22338 15428
rect 22466 14456 22522 14512
rect 23110 19624 23166 19680
rect 23018 17604 23074 17640
rect 23018 17584 23020 17604
rect 23020 17584 23072 17604
rect 23072 17584 23074 17604
rect 24122 32136 24178 32192
rect 24766 30504 24822 30560
rect 24030 29280 24086 29336
rect 24122 29008 24178 29064
rect 23386 24928 23442 24984
rect 23662 25608 23718 25664
rect 23570 25064 23626 25120
rect 23846 24520 23902 24576
rect 23754 24384 23810 24440
rect 23294 22616 23350 22672
rect 23478 22616 23534 22672
rect 23570 22344 23626 22400
rect 23294 20712 23350 20768
rect 23386 20168 23442 20224
rect 23846 22752 23902 22808
rect 23938 22616 23994 22672
rect 23754 21392 23810 21448
rect 24214 26560 24270 26616
rect 23938 20576 23994 20632
rect 23386 17992 23442 18048
rect 23018 16360 23074 16416
rect 23386 15272 23442 15328
rect 24582 29280 24638 29336
rect 24766 29144 24822 29200
rect 25042 29008 25098 29064
rect 24398 25780 24400 25800
rect 24400 25780 24452 25800
rect 24452 25780 24454 25800
rect 24398 25744 24454 25780
rect 24398 24520 24454 24576
rect 24398 24112 24454 24168
rect 24214 20712 24270 20768
rect 24214 20440 24270 20496
rect 24398 21956 24454 21992
rect 24398 21936 24400 21956
rect 24400 21936 24452 21956
rect 24452 21936 24454 21956
rect 24674 25744 24730 25800
rect 25042 25644 25044 25664
rect 25044 25644 25096 25664
rect 25096 25644 25098 25664
rect 25042 25608 25098 25644
rect 24674 25064 24730 25120
rect 24766 24112 24822 24168
rect 24950 23568 25006 23624
rect 24950 22888 25006 22944
rect 25318 26324 25320 26344
rect 25320 26324 25372 26344
rect 25372 26324 25374 26344
rect 25318 26288 25374 26324
rect 25318 25608 25374 25664
rect 25410 25472 25466 25528
rect 25226 23704 25282 23760
rect 25134 23160 25190 23216
rect 24490 21664 24546 21720
rect 25134 21972 25136 21992
rect 25136 21972 25188 21992
rect 25188 21972 25190 21992
rect 24858 21800 24914 21856
rect 24674 21392 24730 21448
rect 24490 20984 24546 21040
rect 24490 20712 24546 20768
rect 24030 17876 24086 17912
rect 24030 17856 24032 17876
rect 24032 17856 24084 17876
rect 24084 17856 24086 17876
rect 24030 16768 24086 16824
rect 22282 13524 22338 13560
rect 22282 13504 22284 13524
rect 22284 13504 22336 13524
rect 22336 13504 22338 13524
rect 23110 14068 23166 14104
rect 23110 14048 23112 14068
rect 23112 14048 23164 14068
rect 23164 14048 23166 14068
rect 23202 13232 23258 13288
rect 24214 14456 24270 14512
rect 23846 13640 23902 13696
rect 24398 13504 24454 13560
rect 23938 12960 23994 13016
rect 24858 20984 24914 21040
rect 25134 21936 25190 21972
rect 25134 21120 25190 21176
rect 24858 19216 24914 19272
rect 24766 16904 24822 16960
rect 25594 24284 25596 24304
rect 25596 24284 25648 24304
rect 25648 24284 25650 24304
rect 25594 24248 25650 24284
rect 25778 31592 25834 31648
rect 26422 32136 26478 32192
rect 26698 30776 26754 30832
rect 25962 29688 26018 29744
rect 26330 28736 26386 28792
rect 26330 27820 26332 27840
rect 26332 27820 26384 27840
rect 26384 27820 26386 27840
rect 25778 26288 25834 26344
rect 26330 27784 26386 27820
rect 25870 24928 25926 24984
rect 25778 24248 25834 24304
rect 26238 26288 26294 26344
rect 26054 24792 26110 24848
rect 26238 25100 26240 25120
rect 26240 25100 26292 25120
rect 26292 25100 26294 25120
rect 26238 25064 26294 25100
rect 26790 30232 26846 30288
rect 26698 29416 26754 29472
rect 26606 27376 26662 27432
rect 26606 26580 26662 26616
rect 26606 26560 26608 26580
rect 26608 26560 26660 26580
rect 26660 26560 26662 26580
rect 26882 27376 26938 27432
rect 26882 27104 26938 27160
rect 25686 21936 25742 21992
rect 25870 23724 25926 23760
rect 25870 23704 25872 23724
rect 25872 23704 25924 23724
rect 25924 23704 25926 23724
rect 25870 23432 25926 23488
rect 25410 18672 25466 18728
rect 25410 18400 25466 18456
rect 25410 18028 25412 18048
rect 25412 18028 25464 18048
rect 25464 18028 25466 18048
rect 25410 17992 25466 18028
rect 25686 19916 25742 19952
rect 25686 19896 25688 19916
rect 25688 19896 25740 19916
rect 25740 19896 25742 19916
rect 26422 24792 26478 24848
rect 26698 25064 26754 25120
rect 26606 24792 26662 24848
rect 26330 24248 26386 24304
rect 26790 24928 26846 24984
rect 26698 23840 26754 23896
rect 26238 23432 26294 23488
rect 26146 22480 26202 22536
rect 26514 23704 26570 23760
rect 27066 30504 27122 30560
rect 27158 28736 27214 28792
rect 27158 27920 27214 27976
rect 26882 23704 26938 23760
rect 27250 26560 27306 26616
rect 27066 22752 27122 22808
rect 26882 22480 26938 22536
rect 26238 22344 26294 22400
rect 25962 21528 26018 21584
rect 26146 21528 26202 21584
rect 26146 21256 26202 21312
rect 26422 21120 26478 21176
rect 26054 20576 26110 20632
rect 25410 14728 25466 14784
rect 24398 12824 24454 12880
rect 23202 12588 23204 12608
rect 23204 12588 23256 12608
rect 23256 12588 23258 12608
rect 23202 12552 23258 12588
rect 25594 15408 25650 15464
rect 26790 22344 26846 22400
rect 26790 20712 26846 20768
rect 26146 17856 26202 17912
rect 27618 27648 27674 27704
rect 27894 31592 27950 31648
rect 27894 31048 27950 31104
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 28078 32000 28134 32056
rect 28170 31864 28226 31920
rect 28078 29416 28134 29472
rect 27986 28056 28042 28112
rect 27986 27648 28042 27704
rect 27434 26288 27490 26344
rect 27526 26016 27582 26072
rect 27434 25472 27490 25528
rect 27434 25200 27490 25256
rect 27618 25200 27674 25256
rect 27526 24284 27528 24304
rect 27528 24284 27580 24304
rect 27580 24284 27582 24304
rect 27526 24248 27582 24284
rect 26974 20712 27030 20768
rect 26514 19660 26516 19680
rect 26516 19660 26568 19680
rect 26568 19660 26570 19680
rect 26514 19624 26570 19660
rect 26974 19080 27030 19136
rect 27066 18400 27122 18456
rect 26422 15952 26478 16008
rect 26790 17720 26846 17776
rect 26974 17312 27030 17368
rect 27250 20576 27306 20632
rect 27986 26832 28042 26888
rect 28078 24284 28080 24304
rect 28080 24284 28132 24304
rect 28132 24284 28134 24304
rect 28078 24248 28134 24284
rect 27802 23724 27858 23760
rect 27802 23704 27804 23724
rect 27804 23704 27856 23724
rect 27856 23704 27858 23724
rect 27802 23432 27858 23488
rect 27802 22888 27858 22944
rect 28354 32000 28410 32056
rect 28538 31456 28594 31512
rect 28262 31048 28318 31104
rect 28722 30932 28778 30968
rect 28722 30912 28724 30932
rect 28724 30912 28776 30932
rect 28776 30912 28778 30932
rect 28262 28328 28318 28384
rect 28630 30096 28686 30152
rect 28354 28192 28410 28248
rect 29550 29824 29606 29880
rect 29550 29688 29606 29744
rect 28906 28736 28962 28792
rect 28630 28328 28686 28384
rect 29090 28192 29146 28248
rect 29366 29008 29422 29064
rect 28538 26832 28594 26888
rect 28630 25880 28686 25936
rect 28170 23432 28226 23488
rect 27986 22092 28042 22128
rect 28262 22616 28318 22672
rect 27986 22072 27988 22092
rect 27988 22072 28040 22092
rect 28040 22072 28042 22092
rect 28078 21972 28080 21992
rect 28080 21972 28132 21992
rect 28132 21972 28134 21992
rect 28078 21936 28134 21972
rect 27894 20984 27950 21040
rect 27710 20712 27766 20768
rect 27434 19624 27490 19680
rect 27342 19352 27398 19408
rect 26422 15544 26478 15600
rect 26054 12960 26110 13016
rect 26330 14864 26386 14920
rect 26698 15816 26754 15872
rect 26698 15272 26754 15328
rect 26514 13932 26570 13968
rect 26514 13912 26516 13932
rect 26516 13912 26568 13932
rect 26568 13912 26570 13932
rect 26882 16224 26938 16280
rect 26882 15816 26938 15872
rect 25686 12416 25742 12472
rect 27342 16496 27398 16552
rect 27342 16224 27398 16280
rect 27342 15156 27398 15192
rect 27342 15136 27344 15156
rect 27344 15136 27396 15156
rect 27396 15136 27398 15156
rect 27894 20712 27950 20768
rect 27986 20596 28042 20632
rect 27986 20576 27988 20596
rect 27988 20576 28040 20596
rect 28040 20576 28042 20596
rect 28170 21528 28226 21584
rect 28446 22228 28502 22264
rect 28446 22208 28448 22228
rect 28448 22208 28500 22228
rect 28500 22208 28502 22228
rect 28354 21936 28410 21992
rect 27802 19216 27858 19272
rect 27802 17992 27858 18048
rect 27526 17176 27582 17232
rect 27158 12280 27214 12336
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 27986 17856 28042 17912
rect 28078 17196 28134 17232
rect 28078 17176 28080 17196
rect 28080 17176 28132 17196
rect 28132 17176 28134 17196
rect 27894 16768 27950 16824
rect 28446 20984 28502 21040
rect 28630 22208 28686 22264
rect 28814 27784 28870 27840
rect 28998 27104 29054 27160
rect 28906 26560 28962 26616
rect 28814 25472 28870 25528
rect 29366 27784 29422 27840
rect 30378 32136 30434 32192
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 30378 31728 30434 31784
rect 30562 31048 30618 31104
rect 30286 30504 30342 30560
rect 30102 30132 30104 30152
rect 30104 30132 30156 30152
rect 30156 30132 30158 30152
rect 30102 30096 30158 30132
rect 30286 29960 30342 30016
rect 30010 29280 30066 29336
rect 29090 25472 29146 25528
rect 28906 24928 28962 24984
rect 29090 23840 29146 23896
rect 28998 22380 29000 22400
rect 29000 22380 29052 22400
rect 29052 22380 29054 22400
rect 28998 22344 29054 22380
rect 29366 22480 29422 22536
rect 29090 22208 29146 22264
rect 29182 21664 29238 21720
rect 29090 20340 29092 20360
rect 29092 20340 29144 20360
rect 29144 20340 29146 20360
rect 29090 20304 29146 20340
rect 28998 20032 29054 20088
rect 28538 17992 28594 18048
rect 28354 17176 28410 17232
rect 28814 18944 28870 19000
rect 29090 19080 29146 19136
rect 29366 21392 29422 21448
rect 29274 20984 29330 21040
rect 29274 20032 29330 20088
rect 29274 19624 29330 19680
rect 29274 18536 29330 18592
rect 29366 17856 29422 17912
rect 29826 28328 29882 28384
rect 30010 27920 30066 27976
rect 30102 26016 30158 26072
rect 29826 24928 29882 24984
rect 29734 24248 29790 24304
rect 29734 23840 29790 23896
rect 29826 23468 29828 23488
rect 29828 23468 29880 23488
rect 29880 23468 29882 23488
rect 29826 23432 29882 23468
rect 29734 21412 29790 21448
rect 29734 21392 29736 21412
rect 29736 21392 29788 21412
rect 29788 21392 29790 21412
rect 30010 20576 30066 20632
rect 29734 19488 29790 19544
rect 29734 17992 29790 18048
rect 29550 17604 29606 17640
rect 29550 17584 29552 17604
rect 29552 17584 29604 17604
rect 29604 17584 29606 17604
rect 27802 14764 27804 14784
rect 27804 14764 27856 14784
rect 27856 14764 27858 14784
rect 27802 14728 27858 14764
rect 27710 14592 27766 14648
rect 28906 16496 28962 16552
rect 28078 14068 28134 14104
rect 28078 14048 28080 14068
rect 28080 14048 28132 14068
rect 28132 14048 28134 14068
rect 28354 13096 28410 13152
rect 29642 16360 29698 16416
rect 29550 15952 29606 16008
rect 29734 15952 29790 16008
rect 29550 15544 29606 15600
rect 29826 13504 29882 13560
rect 30746 29552 30802 29608
rect 30378 25608 30434 25664
rect 30378 24928 30434 24984
rect 30194 17312 30250 17368
rect 30562 19624 30618 19680
rect 30746 29008 30802 29064
rect 30746 25608 30802 25664
rect 30746 24112 30802 24168
rect 30930 29688 30986 29744
rect 31482 31592 31538 31648
rect 31666 30268 31668 30288
rect 31668 30268 31720 30288
rect 31720 30268 31722 30288
rect 31666 30232 31722 30268
rect 31390 29708 31446 29744
rect 31390 29688 31392 29708
rect 31392 29688 31444 29708
rect 31444 29688 31446 29708
rect 31114 29588 31116 29608
rect 31116 29588 31168 29608
rect 31168 29588 31170 29608
rect 31114 29552 31170 29588
rect 31206 29144 31262 29200
rect 31574 30096 31630 30152
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 31666 29280 31722 29336
rect 31482 29008 31538 29064
rect 31022 26424 31078 26480
rect 30930 26288 30986 26344
rect 30838 23704 30894 23760
rect 31482 25064 31538 25120
rect 31758 29008 31814 29064
rect 32126 29144 32182 29200
rect 32126 27276 32128 27296
rect 32128 27276 32180 27296
rect 32180 27276 32182 27296
rect 32126 27240 32182 27276
rect 31666 26288 31722 26344
rect 31850 25064 31906 25120
rect 31666 24520 31722 24576
rect 31666 24112 31722 24168
rect 31666 23840 31722 23896
rect 30930 20576 30986 20632
rect 30930 19352 30986 19408
rect 30654 14900 30656 14920
rect 30656 14900 30708 14920
rect 30708 14900 30710 14920
rect 30654 14864 30710 14900
rect 30838 15136 30894 15192
rect 31022 18400 31078 18456
rect 31390 20576 31446 20632
rect 31390 19488 31446 19544
rect 31574 20576 31630 20632
rect 31574 20304 31630 20360
rect 31942 24792 31998 24848
rect 31942 24112 31998 24168
rect 31942 23568 31998 23624
rect 31758 22752 31814 22808
rect 31942 22616 31998 22672
rect 32862 31184 32918 31240
rect 32402 29552 32458 29608
rect 32586 29960 32642 30016
rect 32310 26560 32366 26616
rect 32310 26152 32366 26208
rect 32218 24656 32274 24712
rect 32310 24520 32366 24576
rect 32310 24248 32366 24304
rect 32218 24112 32274 24168
rect 31482 19116 31484 19136
rect 31484 19116 31536 19136
rect 31536 19116 31538 19136
rect 31206 18808 31262 18864
rect 31482 19080 31538 19116
rect 31390 16360 31446 16416
rect 31022 15000 31078 15056
rect 30930 14612 30986 14648
rect 30930 14592 30932 14612
rect 30932 14592 30984 14612
rect 30984 14592 30986 14612
rect 30930 13640 30986 13696
rect 31022 13504 31078 13560
rect 31666 18536 31722 18592
rect 31942 18536 31998 18592
rect 31942 17856 31998 17912
rect 32218 21800 32274 21856
rect 32862 29416 32918 29472
rect 32678 28364 32680 28384
rect 32680 28364 32732 28384
rect 32732 28364 32734 28384
rect 32678 28328 32734 28364
rect 32770 27648 32826 27704
rect 32770 26832 32826 26888
rect 32586 22480 32642 22536
rect 33138 28736 33194 28792
rect 33414 30640 33470 30696
rect 33414 27920 33470 27976
rect 32770 23432 32826 23488
rect 32954 23432 33010 23488
rect 32678 22208 32734 22264
rect 32310 21392 32366 21448
rect 32218 20712 32274 20768
rect 32310 19488 32366 19544
rect 32218 19252 32220 19272
rect 32220 19252 32272 19272
rect 32272 19252 32274 19272
rect 32218 19216 32274 19252
rect 32126 19116 32128 19136
rect 32128 19116 32180 19136
rect 32180 19116 32182 19136
rect 32126 19080 32182 19116
rect 32218 17992 32274 18048
rect 32402 16768 32458 16824
rect 32586 21664 32642 21720
rect 33046 22480 33102 22536
rect 32862 21936 32918 21992
rect 32586 17856 32642 17912
rect 32586 17448 32642 17504
rect 32402 16244 32458 16280
rect 32402 16224 32404 16244
rect 32404 16224 32456 16244
rect 32456 16224 32458 16244
rect 32586 16108 32642 16144
rect 32586 16088 32588 16108
rect 32588 16088 32640 16108
rect 32640 16088 32642 16108
rect 31574 15020 31630 15056
rect 31574 15000 31576 15020
rect 31576 15000 31628 15020
rect 31628 15000 31630 15020
rect 31574 14764 31576 14784
rect 31576 14764 31628 14784
rect 31628 14764 31630 14784
rect 31574 14728 31630 14764
rect 33414 27240 33470 27296
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 33598 24384 33654 24440
rect 33230 21936 33286 21992
rect 33230 21684 33286 21720
rect 33230 21664 33232 21684
rect 33232 21664 33284 21684
rect 33284 21664 33286 21684
rect 33230 21256 33286 21312
rect 33874 29008 33930 29064
rect 34150 28600 34206 28656
rect 33874 24520 33930 24576
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34702 30368 34758 30424
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35070 29280 35126 29336
rect 34702 29008 34758 29064
rect 34702 28872 34758 28928
rect 34518 28192 34574 28248
rect 34242 25608 34298 25664
rect 34242 25472 34298 25528
rect 33598 21936 33654 21992
rect 33506 21664 33562 21720
rect 32954 16088 33010 16144
rect 32862 15700 32918 15736
rect 32862 15680 32864 15700
rect 32864 15680 32916 15700
rect 32916 15680 32918 15700
rect 32862 15428 32918 15464
rect 32862 15408 32864 15428
rect 32864 15408 32916 15428
rect 32916 15408 32918 15428
rect 33322 17040 33378 17096
rect 33230 16224 33286 16280
rect 33414 16360 33470 16416
rect 34426 24928 34482 24984
rect 34426 23976 34482 24032
rect 34702 27668 34758 27704
rect 34702 27648 34704 27668
rect 34704 27648 34756 27668
rect 34756 27648 34758 27668
rect 34886 29008 34942 29064
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 36174 31320 36230 31376
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35622 28484 35678 28520
rect 35622 28464 35624 28484
rect 35624 28464 35676 28484
rect 35676 28464 35678 28484
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 35530 27668 35586 27704
rect 35530 27648 35532 27668
rect 35532 27648 35584 27668
rect 35584 27648 35586 27668
rect 35254 27240 35310 27296
rect 34610 24112 34666 24168
rect 34518 23840 34574 23896
rect 34242 22208 34298 22264
rect 34058 21256 34114 21312
rect 33966 21120 34022 21176
rect 33966 20032 34022 20088
rect 33966 19780 34022 19816
rect 33966 19760 33968 19780
rect 33968 19760 34020 19780
rect 34020 19760 34022 19780
rect 34242 21936 34298 21992
rect 34242 21800 34298 21856
rect 34426 23296 34482 23352
rect 34518 23160 34574 23216
rect 34518 22344 34574 22400
rect 34334 20984 34390 21040
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35162 26016 35218 26072
rect 34794 25608 34850 25664
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34886 24792 34942 24848
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34978 23976 35034 24032
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34886 23196 34888 23216
rect 34888 23196 34940 23216
rect 34940 23196 34942 23216
rect 34886 23160 34942 23196
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34610 20340 34612 20360
rect 34612 20340 34664 20360
rect 34664 20340 34666 20360
rect 34610 20304 34666 20340
rect 33874 19352 33930 19408
rect 33782 17720 33838 17776
rect 34242 18400 34298 18456
rect 34150 17040 34206 17096
rect 32678 14592 32734 14648
rect 33598 15444 33600 15464
rect 33600 15444 33652 15464
rect 33652 15444 33654 15464
rect 33598 15408 33654 15444
rect 33690 15020 33746 15056
rect 33690 15000 33692 15020
rect 33692 15000 33744 15020
rect 33744 15000 33746 15020
rect 33506 14864 33562 14920
rect 34518 19760 34574 19816
rect 35070 21664 35126 21720
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 35438 27104 35494 27160
rect 35530 26580 35586 26616
rect 35530 26560 35532 26580
rect 35532 26560 35584 26580
rect 35584 26560 35586 26580
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 36082 26016 36138 26072
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35530 21956 35586 21992
rect 35530 21936 35532 21956
rect 35532 21936 35584 21956
rect 35584 21936 35586 21956
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 36450 25336 36506 25392
rect 36634 27376 36690 27432
rect 36450 22480 36506 22536
rect 35438 20848 35494 20904
rect 34702 18284 34758 18320
rect 34702 18264 34704 18284
rect 34704 18264 34756 18284
rect 34756 18264 34758 18284
rect 34518 18028 34520 18048
rect 34520 18028 34572 18048
rect 34572 18028 34574 18048
rect 34518 17992 34574 18028
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 35346 18264 35402 18320
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35346 17720 35402 17776
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 35070 17312 35126 17368
rect 35346 17176 35402 17232
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34794 14320 34850 14376
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 36542 20984 36598 21040
rect 39026 32272 39082 32328
rect 37738 29960 37794 30016
rect 37370 29688 37426 29744
rect 37186 26868 37188 26888
rect 37188 26868 37240 26888
rect 37240 26868 37242 26888
rect 37186 26832 37242 26868
rect 36726 23724 36782 23760
rect 36726 23704 36728 23724
rect 36728 23704 36780 23724
rect 36780 23704 36782 23724
rect 36818 21528 36874 21584
rect 37278 25764 37334 25800
rect 37278 25744 37280 25764
rect 37280 25744 37332 25764
rect 37332 25744 37334 25764
rect 37278 23160 37334 23216
rect 37646 26288 37702 26344
rect 37462 24928 37518 24984
rect 37462 23568 37518 23624
rect 37462 21548 37518 21584
rect 37462 21528 37464 21548
rect 37464 21528 37516 21548
rect 37516 21528 37518 21548
rect 37094 19896 37150 19952
rect 36634 17196 36690 17232
rect 36634 17176 36636 17196
rect 36636 17176 36688 17196
rect 36688 17176 36690 17196
rect 36542 17076 36544 17096
rect 36544 17076 36596 17096
rect 36596 17076 36598 17096
rect 36542 17040 36598 17076
rect 36634 16088 36690 16144
rect 36910 18672 36966 18728
rect 37094 16496 37150 16552
rect 37462 18128 37518 18184
rect 38566 30096 38622 30152
rect 37922 26580 37978 26616
rect 37922 26560 37924 26580
rect 37924 26560 37976 26580
rect 37976 26560 37978 26580
rect 37462 14456 37518 14512
rect 34426 13368 34482 13424
rect 38382 25880 38438 25936
rect 38290 24248 38346 24304
rect 38842 25200 38898 25256
rect 38934 23724 38990 23760
rect 38934 23704 38936 23724
rect 38936 23704 38988 23724
rect 38988 23704 38990 23724
rect 40222 30232 40278 30288
rect 39854 26988 39910 27024
rect 39854 26968 39856 26988
rect 39856 26968 39908 26988
rect 39908 26968 39910 26988
rect 38014 17720 38070 17776
rect 38750 17604 38806 17640
rect 38750 17584 38752 17604
rect 38752 17584 38804 17604
rect 38804 17584 38806 17604
rect 40958 26988 41014 27024
rect 40958 26968 40960 26988
rect 40960 26968 41012 26988
rect 41012 26968 41014 26988
rect 44546 29280 44602 29336
rect 44086 28600 44142 28656
rect 42338 28056 42394 28112
rect 44454 27940 44510 27976
rect 44454 27920 44456 27940
rect 44456 27920 44508 27940
rect 44508 27920 44510 27940
rect 44454 27276 44456 27296
rect 44456 27276 44508 27296
rect 44508 27276 44510 27296
rect 44454 27240 44510 27276
rect 42430 27004 42432 27024
rect 42432 27004 42484 27024
rect 42484 27004 42486 27024
rect 42430 26968 42486 27004
rect 41326 26424 41382 26480
rect 44454 26560 44510 26616
rect 44086 25880 44142 25936
rect 41602 24812 41658 24848
rect 41602 24792 41604 24812
rect 41604 24792 41656 24812
rect 41656 24792 41658 24812
rect 40222 20440 40278 20496
rect 41878 22616 41934 22672
rect 43810 24792 43866 24848
rect 44086 23160 44142 23216
rect 44454 25200 44510 25256
rect 44454 24556 44456 24576
rect 44456 24556 44508 24576
rect 44508 24556 44510 24576
rect 44454 24520 44510 24556
rect 44454 23840 44510 23896
rect 44454 22500 44510 22536
rect 44454 22480 44456 22500
rect 44456 22480 44508 22500
rect 44508 22480 44510 22500
rect 39026 16632 39082 16688
rect 44086 20440 44142 20496
rect 44454 21836 44456 21856
rect 44456 21836 44508 21856
rect 44508 21836 44510 21856
rect 44454 21800 44510 21836
rect 44454 21120 44510 21176
rect 44454 19760 44510 19816
rect 44086 19080 44142 19136
rect 44454 18400 44510 18456
rect 44086 17720 44142 17776
rect 44454 17060 44510 17096
rect 44454 17040 44456 17060
rect 44456 17040 44508 17060
rect 44508 17040 44510 17060
rect 44454 16396 44456 16416
rect 44456 16396 44508 16416
rect 44508 16396 44510 16416
rect 44454 16360 44510 16396
rect 44086 15000 44142 15056
rect 44454 15680 44510 15736
rect 44454 14320 44510 14376
rect 44086 13640 44142 13696
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 29090 12144 29146 12200
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 27618 10920 27674 10976
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 24761 33282 24827 33285
rect 25078 33282 25084 33284
rect 24761 33280 25084 33282
rect 24761 33224 24766 33280
rect 24822 33224 25084 33280
rect 24761 33222 25084 33224
rect 24761 33219 24827 33222
rect 25078 33220 25084 33222
rect 25148 33220 25154 33284
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 13629 32330 13695 32333
rect 39021 32330 39087 32333
rect 13629 32328 39087 32330
rect 13629 32272 13634 32328
rect 13690 32272 39026 32328
rect 39082 32272 39087 32328
rect 13629 32270 39087 32272
rect 13629 32267 13695 32270
rect 39021 32267 39087 32270
rect 15837 32194 15903 32197
rect 22553 32194 22619 32197
rect 24117 32194 24183 32197
rect 26417 32194 26483 32197
rect 15837 32192 22619 32194
rect 15837 32136 15842 32192
rect 15898 32136 22558 32192
rect 22614 32136 22619 32192
rect 15837 32134 22619 32136
rect 15837 32131 15903 32134
rect 22553 32131 22619 32134
rect 23062 32134 24042 32194
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 17677 32058 17743 32061
rect 23062 32058 23122 32134
rect 23289 32060 23355 32061
rect 23238 32058 23244 32060
rect 17677 32056 23122 32058
rect 17677 32000 17682 32056
rect 17738 32000 23122 32056
rect 17677 31998 23122 32000
rect 23198 31998 23244 32058
rect 23308 32056 23355 32060
rect 23350 32000 23355 32056
rect 17677 31995 17743 31998
rect 23238 31996 23244 31998
rect 23308 31996 23355 32000
rect 23982 32058 24042 32134
rect 24117 32192 26483 32194
rect 24117 32136 24122 32192
rect 24178 32136 26422 32192
rect 26478 32136 26483 32192
rect 24117 32134 26483 32136
rect 24117 32131 24183 32134
rect 26417 32131 26483 32134
rect 28022 32132 28028 32196
rect 28092 32194 28098 32196
rect 30373 32194 30439 32197
rect 28092 32192 30439 32194
rect 28092 32136 30378 32192
rect 30434 32136 30439 32192
rect 28092 32134 30439 32136
rect 28092 32132 28098 32134
rect 30373 32131 30439 32134
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 28073 32058 28139 32061
rect 23982 32056 28139 32058
rect 23982 32000 28078 32056
rect 28134 32000 28139 32056
rect 23982 31998 28139 32000
rect 23289 31995 23355 31996
rect 28073 31995 28139 31998
rect 28206 31996 28212 32060
rect 28276 32058 28282 32060
rect 28349 32058 28415 32061
rect 28276 32056 28415 32058
rect 28276 32000 28354 32056
rect 28410 32000 28415 32056
rect 28276 31998 28415 32000
rect 28276 31996 28282 31998
rect 28349 31995 28415 31998
rect 19425 31922 19491 31925
rect 19977 31922 20043 31925
rect 28165 31922 28231 31925
rect 19425 31920 28231 31922
rect 19425 31864 19430 31920
rect 19486 31864 19982 31920
rect 20038 31864 28170 31920
rect 28226 31864 28231 31920
rect 19425 31862 28231 31864
rect 19425 31859 19491 31862
rect 19977 31859 20043 31862
rect 28165 31859 28231 31862
rect 22553 31786 22619 31789
rect 23933 31786 23999 31789
rect 30373 31786 30439 31789
rect 22553 31784 30439 31786
rect 22553 31728 22558 31784
rect 22614 31728 23938 31784
rect 23994 31728 30378 31784
rect 30434 31728 30439 31784
rect 22553 31726 30439 31728
rect 22553 31723 22619 31726
rect 23933 31723 23999 31726
rect 30373 31723 30439 31726
rect 19609 31650 19675 31653
rect 25773 31650 25839 31653
rect 19609 31648 25839 31650
rect 19609 31592 19614 31648
rect 19670 31592 25778 31648
rect 25834 31592 25839 31648
rect 19609 31590 25839 31592
rect 19609 31587 19675 31590
rect 25773 31587 25839 31590
rect 27889 31650 27955 31653
rect 31477 31650 31543 31653
rect 27889 31648 31543 31650
rect 27889 31592 27894 31648
rect 27950 31592 31482 31648
rect 31538 31592 31543 31648
rect 27889 31590 31543 31592
rect 27889 31587 27955 31590
rect 31477 31587 31543 31590
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 13445 31514 13511 31517
rect 17125 31514 17191 31517
rect 28533 31514 28599 31517
rect 13445 31512 28599 31514
rect 13445 31456 13450 31512
rect 13506 31456 17130 31512
rect 17186 31456 28538 31512
rect 28594 31456 28599 31512
rect 13445 31454 28599 31456
rect 13445 31451 13511 31454
rect 17125 31451 17191 31454
rect 28533 31451 28599 31454
rect 14549 31378 14615 31381
rect 36169 31378 36235 31381
rect 14549 31376 36235 31378
rect 14549 31320 14554 31376
rect 14610 31320 36174 31376
rect 36230 31320 36235 31376
rect 14549 31318 36235 31320
rect 14549 31315 14615 31318
rect 36169 31315 36235 31318
rect 15469 31242 15535 31245
rect 19190 31242 19196 31244
rect 15469 31240 19196 31242
rect 15469 31184 15474 31240
rect 15530 31184 19196 31240
rect 15469 31182 19196 31184
rect 15469 31179 15535 31182
rect 19190 31180 19196 31182
rect 19260 31242 19266 31244
rect 32857 31242 32923 31245
rect 19260 31240 32923 31242
rect 19260 31184 32862 31240
rect 32918 31184 32923 31240
rect 19260 31182 32923 31184
rect 19260 31180 19266 31182
rect 32857 31179 32923 31182
rect 11145 31106 11211 31109
rect 19926 31106 19932 31108
rect 11145 31104 19932 31106
rect 11145 31048 11150 31104
rect 11206 31048 19932 31104
rect 11145 31046 19932 31048
rect 11145 31043 11211 31046
rect 19926 31044 19932 31046
rect 19996 31044 20002 31108
rect 21725 31106 21791 31109
rect 27889 31106 27955 31109
rect 21725 31104 27955 31106
rect 21725 31048 21730 31104
rect 21786 31048 27894 31104
rect 27950 31048 27955 31104
rect 21725 31046 27955 31048
rect 21725 31043 21791 31046
rect 27889 31043 27955 31046
rect 28257 31106 28323 31109
rect 30557 31106 30623 31109
rect 28257 31104 30623 31106
rect 28257 31048 28262 31104
rect 28318 31048 30562 31104
rect 30618 31048 30623 31104
rect 28257 31046 30623 31048
rect 28257 31043 28323 31046
rect 30557 31043 30623 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 15193 30970 15259 30973
rect 19241 30970 19307 30973
rect 28717 30970 28783 30973
rect 15193 30968 28783 30970
rect 15193 30912 15198 30968
rect 15254 30912 19246 30968
rect 19302 30912 28722 30968
rect 28778 30912 28783 30968
rect 15193 30910 28783 30912
rect 15193 30907 15259 30910
rect 19241 30907 19307 30910
rect 28717 30907 28783 30910
rect 19977 30834 20043 30837
rect 22461 30834 22527 30837
rect 26693 30834 26759 30837
rect 19977 30832 26759 30834
rect 19977 30776 19982 30832
rect 20038 30776 22466 30832
rect 22522 30776 26698 30832
rect 26754 30776 26759 30832
rect 19977 30774 26759 30776
rect 19977 30771 20043 30774
rect 22461 30771 22527 30774
rect 26693 30771 26759 30774
rect 33409 30700 33475 30701
rect 33358 30698 33364 30700
rect 22050 30638 33364 30698
rect 33428 30698 33475 30700
rect 33428 30696 33556 30698
rect 33470 30640 33556 30696
rect 14457 30562 14523 30565
rect 18781 30562 18847 30565
rect 14457 30560 18847 30562
rect 14457 30504 14462 30560
rect 14518 30504 18786 30560
rect 18842 30504 18847 30560
rect 14457 30502 18847 30504
rect 14457 30499 14523 30502
rect 18781 30499 18847 30502
rect 19742 30500 19748 30564
rect 19812 30562 19818 30564
rect 20437 30562 20503 30565
rect 22050 30562 22110 30638
rect 33358 30636 33364 30638
rect 33428 30638 33556 30640
rect 33428 30636 33475 30638
rect 33409 30635 33475 30636
rect 19812 30560 22110 30562
rect 19812 30504 20442 30560
rect 20498 30504 22110 30560
rect 19812 30502 22110 30504
rect 24761 30562 24827 30565
rect 27061 30562 27127 30565
rect 24761 30560 27127 30562
rect 24761 30504 24766 30560
rect 24822 30504 27066 30560
rect 27122 30504 27127 30560
rect 24761 30502 27127 30504
rect 19812 30500 19818 30502
rect 20437 30499 20503 30502
rect 24761 30499 24827 30502
rect 27061 30499 27127 30502
rect 29678 30500 29684 30564
rect 29748 30562 29754 30564
rect 30281 30562 30347 30565
rect 29748 30560 30347 30562
rect 29748 30504 30286 30560
rect 30342 30504 30347 30560
rect 29748 30502 30347 30504
rect 29748 30500 29754 30502
rect 30281 30499 30347 30502
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 15469 30426 15535 30429
rect 15150 30424 15535 30426
rect 15150 30368 15474 30424
rect 15530 30368 15535 30424
rect 15150 30366 15535 30368
rect 10501 30290 10567 30293
rect 15150 30290 15210 30366
rect 15469 30363 15535 30366
rect 16757 30426 16823 30429
rect 34697 30426 34763 30429
rect 16757 30424 34763 30426
rect 16757 30368 16762 30424
rect 16818 30368 34702 30424
rect 34758 30368 34763 30424
rect 16757 30366 34763 30368
rect 16757 30363 16823 30366
rect 34697 30363 34763 30366
rect 15469 30290 15535 30293
rect 15745 30290 15811 30293
rect 26785 30290 26851 30293
rect 10501 30288 15210 30290
rect 10501 30232 10506 30288
rect 10562 30232 15210 30288
rect 10501 30230 15210 30232
rect 15334 30288 16314 30290
rect 15334 30232 15474 30288
rect 15530 30232 15750 30288
rect 15806 30232 16314 30288
rect 15334 30230 16314 30232
rect 10501 30227 10567 30230
rect 10041 30154 10107 30157
rect 15334 30154 15394 30230
rect 15469 30227 15535 30230
rect 15745 30227 15811 30230
rect 10041 30152 15394 30154
rect 10041 30096 10046 30152
rect 10102 30096 15394 30152
rect 10041 30094 15394 30096
rect 10041 30091 10107 30094
rect 13721 30018 13787 30021
rect 15326 30018 15332 30020
rect 13721 30016 15332 30018
rect 13721 29960 13726 30016
rect 13782 29960 15332 30016
rect 13721 29958 15332 29960
rect 13721 29955 13787 29958
rect 15326 29956 15332 29958
rect 15396 29956 15402 30020
rect 16254 30018 16314 30230
rect 17588 30288 26851 30290
rect 17588 30232 26790 30288
rect 26846 30232 26851 30288
rect 17588 30230 26851 30232
rect 17588 30157 17648 30230
rect 26785 30227 26851 30230
rect 31661 30290 31727 30293
rect 40217 30290 40283 30293
rect 31661 30288 40283 30290
rect 31661 30232 31666 30288
rect 31722 30232 40222 30288
rect 40278 30232 40283 30288
rect 31661 30230 40283 30232
rect 31661 30227 31727 30230
rect 40217 30227 40283 30230
rect 17585 30156 17651 30157
rect 17534 30092 17540 30156
rect 17604 30154 17651 30156
rect 18045 30154 18111 30157
rect 18689 30154 18755 30157
rect 23381 30154 23447 30157
rect 28625 30154 28691 30157
rect 17604 30152 17696 30154
rect 17646 30096 17696 30152
rect 17604 30094 17696 30096
rect 18045 30152 18755 30154
rect 18045 30096 18050 30152
rect 18106 30096 18694 30152
rect 18750 30096 18755 30152
rect 18045 30094 18755 30096
rect 17604 30092 17651 30094
rect 17585 30091 17651 30092
rect 18045 30091 18111 30094
rect 18689 30091 18755 30094
rect 22878 30152 28691 30154
rect 22878 30096 23386 30152
rect 23442 30096 28630 30152
rect 28686 30096 28691 30152
rect 22878 30094 28691 30096
rect 22645 30018 22711 30021
rect 16254 30016 22711 30018
rect 16254 29960 22650 30016
rect 22706 29960 22711 30016
rect 16254 29958 22711 29960
rect 22645 29955 22711 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 17401 29882 17467 29885
rect 18873 29882 18939 29885
rect 17401 29880 18939 29882
rect 17401 29824 17406 29880
rect 17462 29824 18878 29880
rect 18934 29824 18939 29880
rect 17401 29822 18939 29824
rect 17401 29819 17467 29822
rect 18873 29819 18939 29822
rect 22369 29882 22435 29885
rect 22878 29882 22938 30094
rect 23381 30091 23447 30094
rect 28625 30091 28691 30094
rect 30097 30154 30163 30157
rect 31569 30154 31635 30157
rect 38561 30154 38627 30157
rect 30097 30152 31635 30154
rect 30097 30096 30102 30152
rect 30158 30096 31574 30152
rect 31630 30096 31635 30152
rect 30097 30094 31635 30096
rect 30097 30091 30163 30094
rect 31569 30091 31635 30094
rect 34700 30152 38627 30154
rect 34700 30096 38566 30152
rect 38622 30096 38627 30152
rect 34700 30094 38627 30096
rect 30281 30018 30347 30021
rect 32581 30018 32647 30021
rect 30281 30016 32647 30018
rect 30281 29960 30286 30016
rect 30342 29960 32586 30016
rect 32642 29960 32647 30016
rect 30281 29958 32647 29960
rect 30281 29955 30347 29958
rect 32581 29955 32647 29958
rect 22369 29880 22938 29882
rect 22369 29824 22374 29880
rect 22430 29824 22938 29880
rect 22369 29822 22938 29824
rect 29545 29882 29611 29885
rect 34700 29882 34760 30094
rect 38561 30091 38627 30094
rect 37733 30018 37799 30021
rect 45200 30018 46000 30048
rect 37733 30016 46000 30018
rect 37733 29960 37738 30016
rect 37794 29960 46000 30016
rect 37733 29958 46000 29960
rect 37733 29955 37799 29958
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 45200 29928 46000 29958
rect 34930 29887 35246 29888
rect 29545 29880 34760 29882
rect 29545 29824 29550 29880
rect 29606 29824 34760 29880
rect 29545 29822 34760 29824
rect 22369 29819 22435 29822
rect 29545 29819 29611 29822
rect 18689 29746 18755 29749
rect 19057 29746 19123 29749
rect 25957 29746 26023 29749
rect 18689 29744 19123 29746
rect 18689 29688 18694 29744
rect 18750 29688 19062 29744
rect 19118 29688 19123 29744
rect 18689 29686 19123 29688
rect 18689 29683 18755 29686
rect 19057 29683 19123 29686
rect 20670 29744 26023 29746
rect 20670 29688 25962 29744
rect 26018 29688 26023 29744
rect 20670 29686 26023 29688
rect 20670 29613 20730 29686
rect 25957 29683 26023 29686
rect 29545 29746 29611 29749
rect 30925 29746 30991 29749
rect 29545 29744 30991 29746
rect 29545 29688 29550 29744
rect 29606 29688 30930 29744
rect 30986 29688 30991 29744
rect 29545 29686 30991 29688
rect 29545 29683 29611 29686
rect 30925 29683 30991 29686
rect 31385 29746 31451 29749
rect 37365 29746 37431 29749
rect 31385 29744 37431 29746
rect 31385 29688 31390 29744
rect 31446 29688 37370 29744
rect 37426 29688 37431 29744
rect 31385 29686 37431 29688
rect 31385 29683 31451 29686
rect 37365 29683 37431 29686
rect 11053 29610 11119 29613
rect 16757 29610 16823 29613
rect 11053 29608 16823 29610
rect 11053 29552 11058 29608
rect 11114 29552 16762 29608
rect 16818 29552 16823 29608
rect 11053 29550 16823 29552
rect 11053 29547 11119 29550
rect 16757 29547 16823 29550
rect 17585 29610 17651 29613
rect 20621 29610 20730 29613
rect 17585 29608 20730 29610
rect 17585 29552 17590 29608
rect 17646 29552 20626 29608
rect 20682 29552 20730 29608
rect 17585 29550 20730 29552
rect 21081 29610 21147 29613
rect 21582 29610 21588 29612
rect 21081 29608 21588 29610
rect 21081 29552 21086 29608
rect 21142 29552 21588 29608
rect 21081 29550 21588 29552
rect 17585 29547 17651 29550
rect 20621 29547 20687 29550
rect 21081 29547 21147 29550
rect 21582 29548 21588 29550
rect 21652 29610 21658 29612
rect 30741 29610 30807 29613
rect 21652 29608 30807 29610
rect 21652 29552 30746 29608
rect 30802 29552 30807 29608
rect 21652 29550 30807 29552
rect 21652 29548 21658 29550
rect 30741 29547 30807 29550
rect 31109 29610 31175 29613
rect 32397 29610 32463 29613
rect 31109 29608 32463 29610
rect 31109 29552 31114 29608
rect 31170 29552 32402 29608
rect 32458 29552 32463 29608
rect 31109 29550 32463 29552
rect 31109 29547 31175 29550
rect 32397 29547 32463 29550
rect 7649 29474 7715 29477
rect 26693 29474 26759 29477
rect 7649 29472 26759 29474
rect 7649 29416 7654 29472
rect 7710 29416 26698 29472
rect 26754 29416 26759 29472
rect 7649 29414 26759 29416
rect 7649 29411 7715 29414
rect 26693 29411 26759 29414
rect 28073 29474 28139 29477
rect 32857 29474 32923 29477
rect 28073 29472 32923 29474
rect 28073 29416 28078 29472
rect 28134 29416 32862 29472
rect 32918 29416 32923 29472
rect 28073 29414 32923 29416
rect 28073 29411 28139 29414
rect 32857 29411 32923 29414
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 19701 29338 19767 29341
rect 24025 29338 24091 29341
rect 24577 29338 24643 29341
rect 30005 29338 30071 29341
rect 19701 29336 24410 29338
rect 19701 29280 19706 29336
rect 19762 29280 24030 29336
rect 24086 29280 24410 29336
rect 19701 29278 24410 29280
rect 19701 29275 19767 29278
rect 24025 29275 24091 29278
rect 11973 29202 12039 29205
rect 15694 29202 15700 29204
rect 11973 29200 15700 29202
rect 11973 29144 11978 29200
rect 12034 29144 15700 29200
rect 11973 29142 15700 29144
rect 11973 29139 12039 29142
rect 15694 29140 15700 29142
rect 15764 29140 15770 29204
rect 21909 29202 21975 29205
rect 15840 29200 21975 29202
rect 15840 29144 21914 29200
rect 21970 29144 21975 29200
rect 15840 29142 21975 29144
rect 24350 29202 24410 29278
rect 24577 29336 30071 29338
rect 24577 29280 24582 29336
rect 24638 29280 30010 29336
rect 30066 29280 30071 29336
rect 24577 29278 30071 29280
rect 24577 29275 24643 29278
rect 30005 29275 30071 29278
rect 31661 29338 31727 29341
rect 35065 29338 35131 29341
rect 31661 29336 35131 29338
rect 31661 29280 31666 29336
rect 31722 29280 35070 29336
rect 35126 29280 35131 29336
rect 31661 29278 35131 29280
rect 31661 29275 31727 29278
rect 35065 29275 35131 29278
rect 44541 29338 44607 29341
rect 45200 29338 46000 29368
rect 44541 29336 46000 29338
rect 44541 29280 44546 29336
rect 44602 29280 46000 29336
rect 44541 29278 46000 29280
rect 44541 29275 44607 29278
rect 45200 29248 46000 29278
rect 24761 29202 24827 29205
rect 31201 29202 31267 29205
rect 24350 29200 24827 29202
rect 24350 29144 24766 29200
rect 24822 29144 24827 29200
rect 24350 29142 24827 29144
rect 13261 29068 13327 29069
rect 13537 29068 13603 29069
rect 13261 29064 13308 29068
rect 13372 29066 13378 29068
rect 13261 29008 13266 29064
rect 13261 29004 13308 29008
rect 13372 29006 13418 29066
rect 13372 29004 13378 29006
rect 13486 29004 13492 29068
rect 13556 29066 13603 29068
rect 15840 29066 15900 29142
rect 21909 29139 21975 29142
rect 24761 29139 24827 29142
rect 24902 29200 31267 29202
rect 24902 29144 31206 29200
rect 31262 29144 31267 29200
rect 24902 29142 31267 29144
rect 13556 29064 15900 29066
rect 13598 29008 15900 29064
rect 13556 29006 15900 29008
rect 17309 29068 17375 29069
rect 17309 29064 17356 29068
rect 17420 29066 17426 29068
rect 18965 29066 19031 29069
rect 19241 29066 19307 29069
rect 17309 29008 17314 29064
rect 13556 29004 13603 29006
rect 13261 29003 13327 29004
rect 13537 29003 13603 29004
rect 17309 29004 17356 29008
rect 17420 29006 17466 29066
rect 18965 29064 19307 29066
rect 18965 29008 18970 29064
rect 19026 29008 19246 29064
rect 19302 29008 19307 29064
rect 18965 29006 19307 29008
rect 17420 29004 17426 29006
rect 17309 29003 17375 29004
rect 18965 29003 19031 29006
rect 19241 29003 19307 29006
rect 23974 29004 23980 29068
rect 24044 29066 24050 29068
rect 24117 29066 24183 29069
rect 24902 29066 24962 29142
rect 31201 29139 31267 29142
rect 32121 29202 32187 29205
rect 36118 29202 36124 29204
rect 32121 29200 36124 29202
rect 32121 29144 32126 29200
rect 32182 29144 36124 29200
rect 32121 29142 36124 29144
rect 32121 29139 32187 29142
rect 36118 29140 36124 29142
rect 36188 29140 36194 29204
rect 24044 29064 24962 29066
rect 24044 29008 24122 29064
rect 24178 29008 24962 29064
rect 24044 29006 24962 29008
rect 25037 29066 25103 29069
rect 28574 29066 28580 29068
rect 25037 29064 28580 29066
rect 25037 29008 25042 29064
rect 25098 29008 28580 29064
rect 25037 29006 28580 29008
rect 24044 29004 24050 29006
rect 24117 29003 24183 29006
rect 25037 29003 25103 29006
rect 28574 29004 28580 29006
rect 28644 29004 28650 29068
rect 29361 29066 29427 29069
rect 30741 29066 30807 29069
rect 29361 29064 30807 29066
rect 29361 29008 29366 29064
rect 29422 29008 30746 29064
rect 30802 29008 30807 29064
rect 29361 29006 30807 29008
rect 29361 29003 29427 29006
rect 30741 29003 30807 29006
rect 31477 29068 31543 29069
rect 31477 29064 31524 29068
rect 31588 29066 31594 29068
rect 31753 29066 31819 29069
rect 33869 29066 33935 29069
rect 31477 29008 31482 29064
rect 31477 29004 31524 29008
rect 31588 29006 31634 29066
rect 31753 29064 33935 29066
rect 31753 29008 31758 29064
rect 31814 29008 33874 29064
rect 33930 29008 33935 29064
rect 31753 29006 33935 29008
rect 31588 29004 31594 29006
rect 31477 29003 31543 29004
rect 31753 29003 31819 29006
rect 33869 29003 33935 29006
rect 34697 29066 34763 29069
rect 34881 29066 34947 29069
rect 34697 29064 34947 29066
rect 34697 29008 34702 29064
rect 34758 29008 34886 29064
rect 34942 29008 34947 29064
rect 34697 29006 34947 29008
rect 34697 29003 34763 29006
rect 34881 29003 34947 29006
rect 10777 28930 10843 28933
rect 13077 28930 13143 28933
rect 10777 28928 13143 28930
rect 10777 28872 10782 28928
rect 10838 28872 13082 28928
rect 13138 28872 13143 28928
rect 10777 28870 13143 28872
rect 10777 28867 10843 28870
rect 13077 28867 13143 28870
rect 14273 28930 14339 28933
rect 34697 28930 34763 28933
rect 14273 28928 34763 28930
rect 14273 28872 14278 28928
rect 14334 28872 34702 28928
rect 34758 28872 34763 28928
rect 14273 28870 34763 28872
rect 14273 28867 14339 28870
rect 34697 28867 34763 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19558 28732 19564 28796
rect 19628 28794 19634 28796
rect 19793 28794 19859 28797
rect 26325 28794 26391 28797
rect 27153 28794 27219 28797
rect 19628 28792 19859 28794
rect 19628 28736 19798 28792
rect 19854 28736 19859 28792
rect 19628 28734 19859 28736
rect 19628 28732 19634 28734
rect 19793 28731 19859 28734
rect 22050 28792 27219 28794
rect 22050 28736 26330 28792
rect 26386 28736 27158 28792
rect 27214 28736 27219 28792
rect 22050 28734 27219 28736
rect 13813 28658 13879 28661
rect 22050 28658 22110 28734
rect 26325 28731 26391 28734
rect 27153 28731 27219 28734
rect 28901 28794 28967 28797
rect 33133 28794 33199 28797
rect 28901 28792 33199 28794
rect 28901 28736 28906 28792
rect 28962 28736 33138 28792
rect 33194 28736 33199 28792
rect 28901 28734 33199 28736
rect 28901 28731 28967 28734
rect 33133 28731 33199 28734
rect 13813 28656 22110 28658
rect 13813 28600 13818 28656
rect 13874 28600 22110 28656
rect 13813 28598 22110 28600
rect 23381 28658 23447 28661
rect 34145 28658 34211 28661
rect 23381 28656 34211 28658
rect 23381 28600 23386 28656
rect 23442 28600 34150 28656
rect 34206 28600 34211 28656
rect 23381 28598 34211 28600
rect 13813 28595 13879 28598
rect 23381 28595 23447 28598
rect 34145 28595 34211 28598
rect 44081 28658 44147 28661
rect 45200 28658 46000 28688
rect 44081 28656 46000 28658
rect 44081 28600 44086 28656
rect 44142 28600 46000 28656
rect 44081 28598 46000 28600
rect 44081 28595 44147 28598
rect 45200 28568 46000 28598
rect 11329 28522 11395 28525
rect 35617 28522 35683 28525
rect 11329 28520 35683 28522
rect 11329 28464 11334 28520
rect 11390 28464 35622 28520
rect 35678 28464 35683 28520
rect 11329 28462 35683 28464
rect 11329 28459 11395 28462
rect 35617 28459 35683 28462
rect 10409 28386 10475 28389
rect 19057 28386 19123 28389
rect 10409 28384 19123 28386
rect 10409 28328 10414 28384
rect 10470 28328 19062 28384
rect 19118 28328 19123 28384
rect 10409 28326 19123 28328
rect 10409 28323 10475 28326
rect 19057 28323 19123 28326
rect 22185 28386 22251 28389
rect 28257 28386 28323 28389
rect 22185 28384 28323 28386
rect 22185 28328 22190 28384
rect 22246 28328 28262 28384
rect 28318 28328 28323 28384
rect 22185 28326 28323 28328
rect 22185 28323 22251 28326
rect 28257 28323 28323 28326
rect 28625 28386 28691 28389
rect 29821 28386 29887 28389
rect 28625 28384 29887 28386
rect 28625 28328 28630 28384
rect 28686 28328 29826 28384
rect 29882 28328 29887 28384
rect 28625 28326 29887 28328
rect 28625 28323 28691 28326
rect 29821 28323 29887 28326
rect 32254 28324 32260 28388
rect 32324 28386 32330 28388
rect 32673 28386 32739 28389
rect 32324 28384 32739 28386
rect 32324 28328 32678 28384
rect 32734 28328 32739 28384
rect 32324 28326 32739 28328
rect 32324 28324 32330 28326
rect 32673 28323 32739 28326
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 10593 28250 10659 28253
rect 10726 28250 10732 28252
rect 10593 28248 10732 28250
rect 10593 28192 10598 28248
rect 10654 28192 10732 28248
rect 10593 28190 10732 28192
rect 10593 28187 10659 28190
rect 10726 28188 10732 28190
rect 10796 28188 10802 28252
rect 13721 28250 13787 28253
rect 28349 28250 28415 28253
rect 28942 28250 28948 28252
rect 13721 28248 28948 28250
rect 13721 28192 13726 28248
rect 13782 28192 28354 28248
rect 28410 28192 28948 28248
rect 13721 28190 28948 28192
rect 13721 28187 13787 28190
rect 28349 28187 28415 28190
rect 28942 28188 28948 28190
rect 29012 28188 29018 28252
rect 29085 28250 29151 28253
rect 34513 28250 34579 28253
rect 29085 28248 34579 28250
rect 29085 28192 29090 28248
rect 29146 28192 34518 28248
rect 34574 28192 34579 28248
rect 29085 28190 34579 28192
rect 29085 28187 29151 28190
rect 34513 28187 34579 28190
rect 10041 28114 10107 28117
rect 10317 28114 10383 28117
rect 15009 28114 15075 28117
rect 10041 28112 15075 28114
rect 10041 28056 10046 28112
rect 10102 28056 10322 28112
rect 10378 28056 15014 28112
rect 15070 28056 15075 28112
rect 10041 28054 15075 28056
rect 10041 28051 10107 28054
rect 10317 28051 10383 28054
rect 15009 28051 15075 28054
rect 15469 28116 15535 28117
rect 15469 28112 15516 28116
rect 15580 28114 15586 28116
rect 17217 28114 17283 28117
rect 27981 28114 28047 28117
rect 42333 28114 42399 28117
rect 15469 28056 15474 28112
rect 15469 28052 15516 28056
rect 15580 28054 15626 28114
rect 17217 28112 26618 28114
rect 17217 28056 17222 28112
rect 17278 28056 26618 28112
rect 17217 28054 26618 28056
rect 15580 28052 15586 28054
rect 15469 28051 15535 28052
rect 17217 28051 17283 28054
rect 6821 27978 6887 27981
rect 23381 27978 23447 27981
rect 6821 27976 23447 27978
rect 6821 27920 6826 27976
rect 6882 27920 23386 27976
rect 23442 27920 23447 27976
rect 6821 27918 23447 27920
rect 6821 27915 6887 27918
rect 23381 27915 23447 27918
rect 13629 27842 13695 27845
rect 26325 27842 26391 27845
rect 13629 27840 26391 27842
rect 13629 27784 13634 27840
rect 13690 27784 26330 27840
rect 26386 27784 26391 27840
rect 13629 27782 26391 27784
rect 26558 27842 26618 28054
rect 27981 28112 42399 28114
rect 27981 28056 27986 28112
rect 28042 28056 42338 28112
rect 42394 28056 42399 28112
rect 27981 28054 42399 28056
rect 27981 28051 28047 28054
rect 42333 28051 42399 28054
rect 27153 27978 27219 27981
rect 30005 27978 30071 27981
rect 33409 27978 33475 27981
rect 27153 27976 33475 27978
rect 27153 27920 27158 27976
rect 27214 27920 30010 27976
rect 30066 27920 33414 27976
rect 33470 27920 33475 27976
rect 27153 27918 33475 27920
rect 27153 27915 27219 27918
rect 30005 27915 30071 27918
rect 33409 27915 33475 27918
rect 44449 27978 44515 27981
rect 45200 27978 46000 28008
rect 44449 27976 46000 27978
rect 44449 27920 44454 27976
rect 44510 27920 46000 27976
rect 44449 27918 46000 27920
rect 44449 27915 44515 27918
rect 45200 27888 46000 27918
rect 28809 27842 28875 27845
rect 26558 27840 28875 27842
rect 26558 27784 28814 27840
rect 28870 27784 28875 27840
rect 26558 27782 28875 27784
rect 13629 27779 13695 27782
rect 26325 27779 26391 27782
rect 28809 27779 28875 27782
rect 29361 27840 29427 27845
rect 29361 27784 29366 27840
rect 29422 27784 29427 27840
rect 29361 27779 29427 27784
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 6729 27706 6795 27709
rect 17217 27706 17283 27709
rect 6729 27704 17283 27706
rect 6729 27648 6734 27704
rect 6790 27648 17222 27704
rect 17278 27648 17283 27704
rect 6729 27646 17283 27648
rect 6729 27643 6795 27646
rect 17217 27643 17283 27646
rect 17861 27706 17927 27709
rect 19333 27706 19399 27709
rect 17861 27704 19399 27706
rect 17861 27648 17866 27704
rect 17922 27648 19338 27704
rect 19394 27648 19399 27704
rect 17861 27646 19399 27648
rect 17861 27643 17927 27646
rect 19333 27643 19399 27646
rect 21817 27706 21883 27709
rect 27613 27706 27679 27709
rect 21817 27704 27679 27706
rect 21817 27648 21822 27704
rect 21878 27648 27618 27704
rect 27674 27648 27679 27704
rect 21817 27646 27679 27648
rect 21817 27643 21883 27646
rect 27613 27643 27679 27646
rect 27981 27706 28047 27709
rect 29364 27706 29424 27779
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 27981 27704 29424 27706
rect 27981 27648 27986 27704
rect 28042 27648 29424 27704
rect 27981 27646 29424 27648
rect 32765 27708 32831 27709
rect 32765 27704 32812 27708
rect 32876 27706 32882 27708
rect 32765 27648 32770 27704
rect 27981 27643 28047 27646
rect 32765 27644 32812 27648
rect 32876 27646 32922 27706
rect 32876 27644 32882 27646
rect 34462 27644 34468 27708
rect 34532 27706 34538 27708
rect 34697 27706 34763 27709
rect 34532 27704 34763 27706
rect 34532 27648 34702 27704
rect 34758 27648 34763 27704
rect 34532 27646 34763 27648
rect 34532 27644 34538 27646
rect 32765 27643 32831 27644
rect 34697 27643 34763 27646
rect 35382 27644 35388 27708
rect 35452 27706 35458 27708
rect 35525 27706 35591 27709
rect 35452 27704 35591 27706
rect 35452 27648 35530 27704
rect 35586 27648 35591 27704
rect 35452 27646 35591 27648
rect 35452 27644 35458 27646
rect 35525 27643 35591 27646
rect 12617 27570 12683 27573
rect 37222 27570 37228 27572
rect 12617 27568 37228 27570
rect 12617 27512 12622 27568
rect 12678 27512 37228 27568
rect 12617 27510 37228 27512
rect 12617 27507 12683 27510
rect 37222 27508 37228 27510
rect 37292 27508 37298 27572
rect 8109 27434 8175 27437
rect 15837 27434 15903 27437
rect 8109 27432 15903 27434
rect 8109 27376 8114 27432
rect 8170 27376 15842 27432
rect 15898 27376 15903 27432
rect 8109 27374 15903 27376
rect 8109 27371 8175 27374
rect 15837 27371 15903 27374
rect 19977 27434 20043 27437
rect 26601 27434 26667 27437
rect 19977 27432 26667 27434
rect 19977 27376 19982 27432
rect 20038 27376 26606 27432
rect 26662 27376 26667 27432
rect 19977 27374 26667 27376
rect 19977 27371 20043 27374
rect 26601 27371 26667 27374
rect 26877 27434 26943 27437
rect 36629 27434 36695 27437
rect 26877 27432 36695 27434
rect 26877 27376 26882 27432
rect 26938 27376 36634 27432
rect 36690 27376 36695 27432
rect 26877 27374 36695 27376
rect 26877 27371 26943 27374
rect 36629 27371 36695 27374
rect 18781 27298 18847 27301
rect 32121 27298 32187 27301
rect 18781 27296 32187 27298
rect 18781 27240 18786 27296
rect 18842 27240 32126 27296
rect 32182 27240 32187 27296
rect 18781 27238 32187 27240
rect 18781 27235 18847 27238
rect 32121 27235 32187 27238
rect 33409 27298 33475 27301
rect 35249 27298 35315 27301
rect 33409 27296 35315 27298
rect 33409 27240 33414 27296
rect 33470 27240 35254 27296
rect 35310 27240 35315 27296
rect 33409 27238 35315 27240
rect 33409 27235 33475 27238
rect 35249 27235 35315 27238
rect 44449 27298 44515 27301
rect 45200 27298 46000 27328
rect 44449 27296 46000 27298
rect 44449 27240 44454 27296
rect 44510 27240 46000 27296
rect 44449 27238 46000 27240
rect 44449 27235 44515 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 45200 27208 46000 27238
rect 35590 27167 35906 27168
rect 9254 27100 9260 27164
rect 9324 27162 9330 27164
rect 9581 27162 9647 27165
rect 9324 27160 9647 27162
rect 9324 27104 9586 27160
rect 9642 27104 9647 27160
rect 9324 27102 9647 27104
rect 9324 27100 9330 27102
rect 9581 27099 9647 27102
rect 13629 27162 13695 27165
rect 17861 27162 17927 27165
rect 13629 27160 17927 27162
rect 13629 27104 13634 27160
rect 13690 27104 17866 27160
rect 17922 27104 17927 27160
rect 13629 27102 17927 27104
rect 13629 27099 13695 27102
rect 17861 27099 17927 27102
rect 19701 27162 19767 27165
rect 26877 27162 26943 27165
rect 19701 27160 26943 27162
rect 19701 27104 19706 27160
rect 19762 27104 26882 27160
rect 26938 27104 26943 27160
rect 19701 27102 26943 27104
rect 19701 27099 19767 27102
rect 26877 27099 26943 27102
rect 28993 27162 29059 27165
rect 34646 27162 34652 27164
rect 28993 27160 34652 27162
rect 28993 27104 28998 27160
rect 29054 27104 34652 27160
rect 28993 27102 34652 27104
rect 28993 27099 29059 27102
rect 34646 27100 34652 27102
rect 34716 27162 34722 27164
rect 35433 27162 35499 27165
rect 34716 27160 35499 27162
rect 34716 27104 35438 27160
rect 35494 27104 35499 27160
rect 34716 27102 35499 27104
rect 34716 27100 34722 27102
rect 35433 27099 35499 27102
rect 13261 27026 13327 27029
rect 15929 27026 15995 27029
rect 13261 27024 15995 27026
rect 13261 26968 13266 27024
rect 13322 26968 15934 27024
rect 15990 26968 15995 27024
rect 13261 26966 15995 26968
rect 13261 26963 13327 26966
rect 15929 26963 15995 26966
rect 22185 27026 22251 27029
rect 39849 27026 39915 27029
rect 22185 27024 39915 27026
rect 22185 26968 22190 27024
rect 22246 26968 39854 27024
rect 39910 26968 39915 27024
rect 22185 26966 39915 26968
rect 22185 26963 22251 26966
rect 39849 26963 39915 26966
rect 40953 27026 41019 27029
rect 42425 27026 42491 27029
rect 40953 27024 42491 27026
rect 40953 26968 40958 27024
rect 41014 26968 42430 27024
rect 42486 26968 42491 27024
rect 40953 26966 42491 26968
rect 40953 26963 41019 26966
rect 42425 26963 42491 26966
rect 8385 26890 8451 26893
rect 27102 26890 27108 26892
rect 8385 26888 27108 26890
rect 8385 26832 8390 26888
rect 8446 26832 27108 26888
rect 8385 26830 27108 26832
rect 8385 26827 8451 26830
rect 27102 26828 27108 26830
rect 27172 26890 27178 26892
rect 27981 26890 28047 26893
rect 27172 26888 28047 26890
rect 27172 26832 27986 26888
rect 28042 26832 28047 26888
rect 27172 26830 28047 26832
rect 27172 26828 27178 26830
rect 27981 26827 28047 26830
rect 28533 26890 28599 26893
rect 32765 26890 32831 26893
rect 37181 26890 37247 26893
rect 28533 26888 31770 26890
rect 28533 26832 28538 26888
rect 28594 26832 31770 26888
rect 28533 26830 31770 26832
rect 28533 26827 28599 26830
rect 20621 26756 20687 26757
rect 20621 26754 20668 26756
rect 20576 26752 20668 26754
rect 20576 26696 20626 26752
rect 20576 26694 20668 26696
rect 20621 26692 20668 26694
rect 20732 26692 20738 26756
rect 20897 26754 20963 26757
rect 31710 26754 31770 26830
rect 32765 26888 37247 26890
rect 32765 26832 32770 26888
rect 32826 26832 37186 26888
rect 37242 26832 37247 26888
rect 32765 26830 37247 26832
rect 32765 26827 32831 26830
rect 37181 26827 37247 26830
rect 34278 26754 34284 26756
rect 20897 26752 31402 26754
rect 20897 26696 20902 26752
rect 20958 26696 31402 26752
rect 20897 26694 31402 26696
rect 31710 26694 34284 26754
rect 20621 26691 20687 26692
rect 20897 26691 20963 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 10317 26618 10383 26621
rect 11973 26618 12039 26621
rect 15193 26618 15259 26621
rect 10317 26616 15259 26618
rect 10317 26560 10322 26616
rect 10378 26560 11978 26616
rect 12034 26560 15198 26616
rect 15254 26560 15259 26616
rect 10317 26558 15259 26560
rect 10317 26555 10383 26558
rect 11973 26555 12039 26558
rect 15193 26555 15259 26558
rect 17309 26618 17375 26621
rect 19057 26618 19123 26621
rect 17309 26616 19123 26618
rect 17309 26560 17314 26616
rect 17370 26560 19062 26616
rect 19118 26560 19123 26616
rect 17309 26558 19123 26560
rect 17309 26555 17375 26558
rect 19057 26555 19123 26558
rect 22686 26556 22692 26620
rect 22756 26618 22762 26620
rect 23473 26618 23539 26621
rect 22756 26616 23539 26618
rect 22756 26560 23478 26616
rect 23534 26560 23539 26616
rect 22756 26558 23539 26560
rect 22756 26556 22762 26558
rect 23473 26555 23539 26558
rect 24209 26618 24275 26621
rect 26601 26618 26667 26621
rect 24209 26616 26667 26618
rect 24209 26560 24214 26616
rect 24270 26560 26606 26616
rect 26662 26560 26667 26616
rect 24209 26558 26667 26560
rect 24209 26555 24275 26558
rect 26601 26555 26667 26558
rect 27245 26618 27311 26621
rect 28901 26618 28967 26621
rect 27245 26616 28967 26618
rect 27245 26560 27250 26616
rect 27306 26560 28906 26616
rect 28962 26560 28967 26616
rect 27245 26558 28967 26560
rect 27245 26555 27311 26558
rect 28901 26555 28967 26558
rect 6913 26482 6979 26485
rect 31017 26482 31083 26485
rect 6913 26480 31083 26482
rect 6913 26424 6918 26480
rect 6974 26424 31022 26480
rect 31078 26424 31083 26480
rect 6913 26422 31083 26424
rect 31342 26482 31402 26694
rect 34278 26692 34284 26694
rect 34348 26692 34354 26756
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 32305 26618 32371 26621
rect 32438 26618 32444 26620
rect 32305 26616 32444 26618
rect 32305 26560 32310 26616
rect 32366 26560 32444 26616
rect 32305 26558 32444 26560
rect 32305 26555 32371 26558
rect 32438 26556 32444 26558
rect 32508 26556 32514 26620
rect 35525 26618 35591 26621
rect 37917 26618 37983 26621
rect 35525 26616 37983 26618
rect 35525 26560 35530 26616
rect 35586 26560 37922 26616
rect 37978 26560 37983 26616
rect 35525 26558 37983 26560
rect 35525 26555 35591 26558
rect 37917 26555 37983 26558
rect 44449 26618 44515 26621
rect 45200 26618 46000 26648
rect 44449 26616 46000 26618
rect 44449 26560 44454 26616
rect 44510 26560 46000 26616
rect 44449 26558 46000 26560
rect 44449 26555 44515 26558
rect 45200 26528 46000 26558
rect 41321 26482 41387 26485
rect 31342 26480 41387 26482
rect 31342 26424 41326 26480
rect 41382 26424 41387 26480
rect 31342 26422 41387 26424
rect 6913 26419 6979 26422
rect 31017 26419 31083 26422
rect 41321 26419 41387 26422
rect 10317 26346 10383 26349
rect 15469 26346 15535 26349
rect 17401 26346 17467 26349
rect 10317 26344 17467 26346
rect 10317 26288 10322 26344
rect 10378 26288 15474 26344
rect 15530 26288 17406 26344
rect 17462 26288 17467 26344
rect 10317 26286 17467 26288
rect 10317 26283 10383 26286
rect 15469 26283 15535 26286
rect 17401 26283 17467 26286
rect 18270 26284 18276 26348
rect 18340 26346 18346 26348
rect 18413 26346 18479 26349
rect 18340 26344 18479 26346
rect 18340 26288 18418 26344
rect 18474 26288 18479 26344
rect 18340 26286 18479 26288
rect 18340 26284 18346 26286
rect 18413 26283 18479 26286
rect 25313 26346 25379 26349
rect 25773 26348 25839 26349
rect 25630 26346 25636 26348
rect 25313 26344 25636 26346
rect 25313 26288 25318 26344
rect 25374 26288 25636 26344
rect 25313 26286 25636 26288
rect 25313 26283 25379 26286
rect 25630 26284 25636 26286
rect 25700 26284 25706 26348
rect 25773 26344 25820 26348
rect 25884 26346 25890 26348
rect 26233 26346 26299 26349
rect 27429 26346 27495 26349
rect 25773 26288 25778 26344
rect 25773 26284 25820 26288
rect 25884 26286 25930 26346
rect 26233 26344 27495 26346
rect 26233 26288 26238 26344
rect 26294 26288 27434 26344
rect 27490 26288 27495 26344
rect 26233 26286 27495 26288
rect 25884 26284 25890 26286
rect 25773 26283 25839 26284
rect 26233 26283 26299 26286
rect 27429 26283 27495 26286
rect 30782 26284 30788 26348
rect 30852 26346 30858 26348
rect 30925 26346 30991 26349
rect 30852 26344 30991 26346
rect 30852 26288 30930 26344
rect 30986 26288 30991 26344
rect 30852 26286 30991 26288
rect 30852 26284 30858 26286
rect 30925 26283 30991 26286
rect 31661 26346 31727 26349
rect 37641 26346 37707 26349
rect 31661 26344 37707 26346
rect 31661 26288 31666 26344
rect 31722 26288 37646 26344
rect 37702 26288 37707 26344
rect 31661 26286 37707 26288
rect 31661 26283 31727 26286
rect 37641 26283 37707 26286
rect 11145 26210 11211 26213
rect 14825 26210 14891 26213
rect 11145 26208 14891 26210
rect 11145 26152 11150 26208
rect 11206 26152 14830 26208
rect 14886 26152 14891 26208
rect 11145 26150 14891 26152
rect 11145 26147 11211 26150
rect 14825 26147 14891 26150
rect 21950 26148 21956 26212
rect 22020 26210 22026 26212
rect 32305 26210 32371 26213
rect 22020 26208 32371 26210
rect 22020 26152 32310 26208
rect 32366 26152 32371 26208
rect 22020 26150 32371 26152
rect 22020 26148 22026 26150
rect 32305 26147 32371 26150
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 11697 26074 11763 26077
rect 11830 26074 11836 26076
rect 11697 26072 11836 26074
rect 11697 26016 11702 26072
rect 11758 26016 11836 26072
rect 11697 26014 11836 26016
rect 11697 26011 11763 26014
rect 11830 26012 11836 26014
rect 11900 26012 11906 26076
rect 16205 26074 16271 26077
rect 27521 26074 27587 26077
rect 16205 26072 27587 26074
rect 16205 26016 16210 26072
rect 16266 26016 27526 26072
rect 27582 26016 27587 26072
rect 16205 26014 27587 26016
rect 16205 26011 16271 26014
rect 27521 26011 27587 26014
rect 30097 26074 30163 26077
rect 30097 26072 31954 26074
rect 30097 26016 30102 26072
rect 30158 26016 31954 26072
rect 30097 26014 31954 26016
rect 30097 26011 30163 26014
rect 5441 25938 5507 25941
rect 22829 25938 22895 25941
rect 28625 25938 28691 25941
rect 5441 25936 22754 25938
rect 5441 25880 5446 25936
rect 5502 25880 22754 25936
rect 5441 25878 22754 25880
rect 5441 25875 5507 25878
rect 15101 25802 15167 25805
rect 20713 25802 20779 25805
rect 15101 25800 20779 25802
rect 15101 25744 15106 25800
rect 15162 25744 20718 25800
rect 20774 25744 20779 25800
rect 15101 25742 20779 25744
rect 22694 25802 22754 25878
rect 22829 25936 28691 25938
rect 22829 25880 22834 25936
rect 22890 25880 28630 25936
rect 28686 25880 28691 25936
rect 22829 25878 28691 25880
rect 31894 25938 31954 26014
rect 33542 26012 33548 26076
rect 33612 26074 33618 26076
rect 35157 26074 35223 26077
rect 33612 26072 35223 26074
rect 33612 26016 35162 26072
rect 35218 26016 35223 26072
rect 33612 26014 35223 26016
rect 33612 26012 33618 26014
rect 35157 26011 35223 26014
rect 36077 26074 36143 26077
rect 36302 26074 36308 26076
rect 36077 26072 36308 26074
rect 36077 26016 36082 26072
rect 36138 26016 36308 26072
rect 36077 26014 36308 26016
rect 36077 26011 36143 26014
rect 36302 26012 36308 26014
rect 36372 26012 36378 26076
rect 38377 25938 38443 25941
rect 31894 25936 38443 25938
rect 31894 25880 38382 25936
rect 38438 25880 38443 25936
rect 31894 25878 38443 25880
rect 22829 25875 22895 25878
rect 28625 25875 28691 25878
rect 38377 25875 38443 25878
rect 44081 25938 44147 25941
rect 45200 25938 46000 25968
rect 44081 25936 46000 25938
rect 44081 25880 44086 25936
rect 44142 25880 46000 25936
rect 44081 25878 46000 25880
rect 44081 25875 44147 25878
rect 45200 25848 46000 25878
rect 24393 25802 24459 25805
rect 22694 25800 24459 25802
rect 22694 25744 24398 25800
rect 24454 25744 24459 25800
rect 22694 25742 24459 25744
rect 15101 25739 15167 25742
rect 20713 25739 20779 25742
rect 24393 25739 24459 25742
rect 24669 25802 24735 25805
rect 37273 25802 37339 25805
rect 24669 25800 37339 25802
rect 24669 25744 24674 25800
rect 24730 25744 37278 25800
rect 37334 25744 37339 25800
rect 24669 25742 37339 25744
rect 24669 25739 24735 25742
rect 37273 25739 37339 25742
rect 8201 25668 8267 25669
rect 8150 25604 8156 25668
rect 8220 25666 8267 25668
rect 13261 25666 13327 25669
rect 23657 25666 23723 25669
rect 8220 25664 12450 25666
rect 8262 25608 12450 25664
rect 8220 25606 12450 25608
rect 8220 25604 8267 25606
rect 8201 25603 8267 25604
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 12390 25530 12450 25606
rect 13261 25664 23723 25666
rect 13261 25608 13266 25664
rect 13322 25608 23662 25664
rect 23718 25608 23723 25664
rect 13261 25606 23723 25608
rect 24396 25666 24456 25739
rect 25037 25666 25103 25669
rect 24396 25664 25103 25666
rect 24396 25608 25042 25664
rect 25098 25608 25103 25664
rect 24396 25606 25103 25608
rect 13261 25603 13327 25606
rect 23657 25603 23723 25606
rect 25037 25603 25103 25606
rect 25313 25666 25379 25669
rect 25446 25666 25452 25668
rect 25313 25664 25452 25666
rect 25313 25608 25318 25664
rect 25374 25608 25452 25664
rect 25313 25606 25452 25608
rect 25313 25603 25379 25606
rect 25446 25604 25452 25606
rect 25516 25666 25522 25668
rect 30373 25666 30439 25669
rect 25516 25664 30439 25666
rect 25516 25608 30378 25664
rect 30434 25608 30439 25664
rect 25516 25606 30439 25608
rect 25516 25604 25522 25606
rect 30373 25603 30439 25606
rect 30741 25666 30807 25669
rect 33542 25666 33548 25668
rect 30741 25664 33548 25666
rect 30741 25608 30746 25664
rect 30802 25608 33548 25664
rect 30741 25606 33548 25608
rect 30741 25603 30807 25606
rect 33542 25604 33548 25606
rect 33612 25604 33618 25668
rect 34237 25666 34303 25669
rect 34789 25666 34855 25669
rect 34237 25664 34855 25666
rect 34237 25608 34242 25664
rect 34298 25608 34794 25664
rect 34850 25608 34855 25664
rect 34237 25606 34855 25608
rect 34237 25603 34303 25606
rect 34789 25603 34855 25606
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 16113 25530 16179 25533
rect 12390 25528 16179 25530
rect 12390 25472 16118 25528
rect 16174 25472 16179 25528
rect 12390 25470 16179 25472
rect 16113 25467 16179 25470
rect 19517 25530 19583 25533
rect 25405 25530 25471 25533
rect 19517 25528 25471 25530
rect 19517 25472 19522 25528
rect 19578 25472 25410 25528
rect 25466 25472 25471 25528
rect 19517 25470 25471 25472
rect 19517 25467 19583 25470
rect 25405 25467 25471 25470
rect 27429 25530 27495 25533
rect 28809 25530 28875 25533
rect 27429 25528 28875 25530
rect 27429 25472 27434 25528
rect 27490 25472 28814 25528
rect 28870 25472 28875 25528
rect 27429 25470 28875 25472
rect 27429 25467 27495 25470
rect 28809 25467 28875 25470
rect 29085 25530 29151 25533
rect 34237 25530 34303 25533
rect 29085 25528 34303 25530
rect 29085 25472 29090 25528
rect 29146 25472 34242 25528
rect 34298 25472 34303 25528
rect 29085 25470 34303 25472
rect 29085 25467 29151 25470
rect 34237 25467 34303 25470
rect 6085 25394 6151 25397
rect 19333 25394 19399 25397
rect 6085 25392 19399 25394
rect 6085 25336 6090 25392
rect 6146 25336 19338 25392
rect 19394 25336 19399 25392
rect 6085 25334 19399 25336
rect 6085 25331 6151 25334
rect 19333 25331 19399 25334
rect 20161 25394 20227 25397
rect 36445 25394 36511 25397
rect 20161 25392 36511 25394
rect 20161 25336 20166 25392
rect 20222 25336 36450 25392
rect 36506 25336 36511 25392
rect 20161 25334 36511 25336
rect 20161 25331 20227 25334
rect 36445 25331 36511 25334
rect 16297 25260 16363 25261
rect 16246 25258 16252 25260
rect 16170 25198 16252 25258
rect 16316 25258 16363 25260
rect 27429 25258 27495 25261
rect 16316 25256 27495 25258
rect 16358 25200 27434 25256
rect 27490 25200 27495 25256
rect 16246 25196 16252 25198
rect 16316 25198 27495 25200
rect 16316 25196 16363 25198
rect 16297 25195 16363 25196
rect 27429 25195 27495 25198
rect 27613 25258 27679 25261
rect 38837 25258 38903 25261
rect 27613 25256 38903 25258
rect 27613 25200 27618 25256
rect 27674 25200 38842 25256
rect 38898 25200 38903 25256
rect 27613 25198 38903 25200
rect 27613 25195 27679 25198
rect 38837 25195 38903 25198
rect 44449 25258 44515 25261
rect 45200 25258 46000 25288
rect 44449 25256 46000 25258
rect 44449 25200 44454 25256
rect 44510 25200 46000 25256
rect 44449 25198 46000 25200
rect 44449 25195 44515 25198
rect 45200 25168 46000 25198
rect 19333 25122 19399 25125
rect 19885 25122 19951 25125
rect 23565 25122 23631 25125
rect 19333 25120 23631 25122
rect 19333 25064 19338 25120
rect 19394 25064 19890 25120
rect 19946 25064 23570 25120
rect 23626 25064 23631 25120
rect 19333 25062 23631 25064
rect 19333 25059 19399 25062
rect 19885 25059 19951 25062
rect 23565 25059 23631 25062
rect 24669 25122 24735 25125
rect 26233 25122 26299 25125
rect 24669 25120 26299 25122
rect 24669 25064 24674 25120
rect 24730 25064 26238 25120
rect 26294 25064 26299 25120
rect 24669 25062 26299 25064
rect 24669 25059 24735 25062
rect 26233 25059 26299 25062
rect 26693 25122 26759 25125
rect 31477 25122 31543 25125
rect 31845 25122 31911 25125
rect 26693 25120 31543 25122
rect 26693 25064 26698 25120
rect 26754 25064 31482 25120
rect 31538 25064 31543 25120
rect 26693 25062 31543 25064
rect 26693 25059 26759 25062
rect 31477 25059 31543 25062
rect 31710 25120 35450 25122
rect 31710 25064 31850 25120
rect 31906 25064 35450 25120
rect 31710 25062 35450 25064
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 7925 24988 7991 24989
rect 10593 24988 10659 24989
rect 7925 24984 7972 24988
rect 8036 24986 8042 24988
rect 10542 24986 10548 24988
rect 7925 24928 7930 24984
rect 7925 24924 7972 24928
rect 8036 24926 8082 24986
rect 10502 24926 10548 24986
rect 10612 24984 10659 24988
rect 10654 24928 10659 24984
rect 8036 24924 8042 24926
rect 10542 24924 10548 24926
rect 10612 24924 10659 24928
rect 7925 24923 7991 24924
rect 10593 24923 10659 24924
rect 15929 24986 15995 24989
rect 15929 24984 17970 24986
rect 15929 24928 15934 24984
rect 15990 24928 17970 24984
rect 15929 24926 17970 24928
rect 15929 24923 15995 24926
rect 10777 24850 10843 24853
rect 17677 24850 17743 24853
rect 10777 24848 17743 24850
rect 10777 24792 10782 24848
rect 10838 24792 17682 24848
rect 17738 24792 17743 24848
rect 10777 24790 17743 24792
rect 17910 24850 17970 24926
rect 19374 24924 19380 24988
rect 19444 24986 19450 24988
rect 19609 24986 19675 24989
rect 19444 24984 19675 24986
rect 19444 24928 19614 24984
rect 19670 24928 19675 24984
rect 19444 24926 19675 24928
rect 19444 24924 19450 24926
rect 19609 24923 19675 24926
rect 23381 24986 23447 24989
rect 24710 24986 24716 24988
rect 23381 24984 24716 24986
rect 23381 24928 23386 24984
rect 23442 24928 24716 24984
rect 23381 24926 24716 24928
rect 23381 24923 23447 24926
rect 24710 24924 24716 24926
rect 24780 24924 24786 24988
rect 25865 24986 25931 24989
rect 26550 24986 26556 24988
rect 25865 24984 26556 24986
rect 25865 24928 25870 24984
rect 25926 24928 26556 24984
rect 25865 24926 26556 24928
rect 25865 24923 25931 24926
rect 26550 24924 26556 24926
rect 26620 24924 26626 24988
rect 26785 24986 26851 24989
rect 27286 24986 27292 24988
rect 26785 24984 27292 24986
rect 26785 24928 26790 24984
rect 26846 24928 27292 24984
rect 26785 24926 27292 24928
rect 26785 24923 26851 24926
rect 27286 24924 27292 24926
rect 27356 24924 27362 24988
rect 28758 24924 28764 24988
rect 28828 24986 28834 24988
rect 28901 24986 28967 24989
rect 28828 24984 28967 24986
rect 28828 24928 28906 24984
rect 28962 24928 28967 24984
rect 28828 24926 28967 24928
rect 28828 24924 28834 24926
rect 28901 24923 28967 24926
rect 29821 24986 29887 24989
rect 30046 24986 30052 24988
rect 29821 24984 30052 24986
rect 29821 24928 29826 24984
rect 29882 24928 30052 24984
rect 29821 24926 30052 24928
rect 29821 24923 29887 24926
rect 30046 24924 30052 24926
rect 30116 24924 30122 24988
rect 30373 24986 30439 24989
rect 31710 24986 31770 25062
rect 31845 25059 31911 25062
rect 30373 24984 31770 24986
rect 30373 24928 30378 24984
rect 30434 24928 31770 24984
rect 30373 24926 31770 24928
rect 30373 24923 30439 24926
rect 34094 24924 34100 24988
rect 34164 24986 34170 24988
rect 34421 24986 34487 24989
rect 34164 24984 34487 24986
rect 34164 24928 34426 24984
rect 34482 24928 34487 24984
rect 34164 24926 34487 24928
rect 34164 24924 34170 24926
rect 34421 24923 34487 24926
rect 26049 24850 26115 24853
rect 26417 24852 26483 24853
rect 26366 24850 26372 24852
rect 17910 24848 26115 24850
rect 17910 24792 26054 24848
rect 26110 24792 26115 24848
rect 17910 24790 26115 24792
rect 26326 24790 26372 24850
rect 26436 24848 26483 24852
rect 26478 24792 26483 24848
rect 10777 24787 10843 24790
rect 17677 24787 17743 24790
rect 26049 24787 26115 24790
rect 26366 24788 26372 24790
rect 26436 24788 26483 24792
rect 26417 24787 26483 24788
rect 26601 24850 26667 24853
rect 26918 24850 26924 24852
rect 26601 24848 26924 24850
rect 26601 24792 26606 24848
rect 26662 24792 26924 24848
rect 26601 24790 26924 24792
rect 26601 24787 26667 24790
rect 26918 24788 26924 24790
rect 26988 24788 26994 24852
rect 31937 24850 32003 24853
rect 34881 24850 34947 24853
rect 31937 24848 34947 24850
rect 31937 24792 31942 24848
rect 31998 24792 34886 24848
rect 34942 24792 34947 24848
rect 31937 24790 34947 24792
rect 35390 24850 35450 25062
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 37457 24986 37523 24989
rect 36126 24984 37523 24986
rect 36126 24928 37462 24984
rect 37518 24928 37523 24984
rect 36126 24926 37523 24928
rect 36126 24850 36186 24926
rect 37457 24923 37523 24926
rect 35390 24790 36186 24850
rect 41597 24850 41663 24853
rect 43805 24850 43871 24853
rect 41597 24848 43871 24850
rect 41597 24792 41602 24848
rect 41658 24792 43810 24848
rect 43866 24792 43871 24848
rect 41597 24790 43871 24792
rect 31937 24787 32003 24790
rect 34881 24787 34947 24790
rect 41597 24787 41663 24790
rect 43805 24787 43871 24790
rect 8753 24716 8819 24717
rect 8702 24652 8708 24716
rect 8772 24714 8819 24716
rect 14365 24716 14431 24717
rect 8772 24712 8864 24714
rect 8814 24656 8864 24712
rect 8772 24654 8864 24656
rect 14365 24712 14412 24716
rect 14476 24714 14482 24716
rect 18229 24714 18295 24717
rect 32213 24714 32279 24717
rect 14365 24656 14370 24712
rect 8772 24652 8819 24654
rect 8753 24651 8819 24652
rect 14365 24652 14412 24656
rect 14476 24654 14522 24714
rect 18229 24712 32279 24714
rect 18229 24656 18234 24712
rect 18290 24656 32218 24712
rect 32274 24656 32279 24712
rect 18229 24654 32279 24656
rect 14476 24652 14482 24654
rect 14365 24651 14431 24652
rect 18229 24651 18295 24654
rect 32213 24651 32279 24654
rect 9949 24580 10015 24581
rect 9949 24578 9996 24580
rect 9904 24576 9996 24578
rect 9904 24520 9954 24576
rect 9904 24518 9996 24520
rect 9949 24516 9996 24518
rect 10060 24516 10066 24580
rect 11094 24516 11100 24580
rect 11164 24578 11170 24580
rect 11789 24578 11855 24581
rect 11164 24576 11855 24578
rect 11164 24520 11794 24576
rect 11850 24520 11855 24576
rect 11164 24518 11855 24520
rect 11164 24516 11170 24518
rect 9949 24515 10015 24516
rect 11789 24515 11855 24518
rect 13169 24578 13235 24581
rect 18045 24578 18111 24581
rect 18505 24578 18571 24581
rect 13169 24576 18571 24578
rect 13169 24520 13174 24576
rect 13230 24520 18050 24576
rect 18106 24520 18510 24576
rect 18566 24520 18571 24576
rect 13169 24518 18571 24520
rect 13169 24515 13235 24518
rect 18045 24515 18111 24518
rect 18505 24515 18571 24518
rect 22093 24578 22159 24581
rect 22921 24580 22987 24581
rect 22093 24576 22754 24578
rect 22093 24520 22098 24576
rect 22154 24520 22754 24576
rect 22093 24518 22754 24520
rect 22093 24515 22159 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 9581 24442 9647 24445
rect 21766 24442 21772 24444
rect 9581 24440 21772 24442
rect 9581 24384 9586 24440
rect 9642 24384 21772 24440
rect 9581 24382 21772 24384
rect 9581 24379 9647 24382
rect 21766 24380 21772 24382
rect 21836 24442 21842 24444
rect 22553 24442 22619 24445
rect 21836 24440 22619 24442
rect 21836 24384 22558 24440
rect 22614 24384 22619 24440
rect 21836 24382 22619 24384
rect 22694 24442 22754 24518
rect 22870 24516 22876 24580
rect 22940 24578 22987 24580
rect 23841 24578 23907 24581
rect 22940 24576 23032 24578
rect 22982 24520 23032 24576
rect 22940 24518 23032 24520
rect 23108 24576 23907 24578
rect 23108 24520 23846 24576
rect 23902 24520 23907 24576
rect 23108 24518 23907 24520
rect 22940 24516 22987 24518
rect 22921 24515 22987 24516
rect 23108 24442 23168 24518
rect 23841 24515 23907 24518
rect 24393 24578 24459 24581
rect 31661 24578 31727 24581
rect 24393 24576 31727 24578
rect 24393 24520 24398 24576
rect 24454 24520 31666 24576
rect 31722 24520 31727 24576
rect 24393 24518 31727 24520
rect 24393 24515 24459 24518
rect 31661 24515 31727 24518
rect 32305 24578 32371 24581
rect 33869 24578 33935 24581
rect 32305 24576 33935 24578
rect 32305 24520 32310 24576
rect 32366 24520 33874 24576
rect 33930 24520 33935 24576
rect 32305 24518 33935 24520
rect 32305 24515 32371 24518
rect 33869 24515 33935 24518
rect 44449 24578 44515 24581
rect 45200 24578 46000 24608
rect 44449 24576 46000 24578
rect 44449 24520 44454 24576
rect 44510 24520 46000 24576
rect 44449 24518 46000 24520
rect 44449 24515 44515 24518
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 45200 24488 46000 24518
rect 34930 24447 35246 24448
rect 22694 24382 23168 24442
rect 23749 24442 23815 24445
rect 33593 24442 33659 24445
rect 23749 24440 33659 24442
rect 23749 24384 23754 24440
rect 23810 24384 33598 24440
rect 33654 24384 33659 24440
rect 23749 24382 33659 24384
rect 21836 24380 21842 24382
rect 22553 24379 22619 24382
rect 23749 24379 23815 24382
rect 33593 24379 33659 24382
rect 9765 24306 9831 24309
rect 10685 24306 10751 24309
rect 13169 24306 13235 24309
rect 13629 24308 13695 24309
rect 13629 24306 13676 24308
rect 9765 24304 13235 24306
rect 9765 24248 9770 24304
rect 9826 24248 10690 24304
rect 10746 24248 13174 24304
rect 13230 24248 13235 24304
rect 9765 24246 13235 24248
rect 13588 24304 13676 24306
rect 13740 24306 13746 24308
rect 22093 24306 22159 24309
rect 13740 24304 22159 24306
rect 13588 24248 13634 24304
rect 13740 24248 22098 24304
rect 22154 24248 22159 24304
rect 13588 24246 13676 24248
rect 9765 24243 9831 24246
rect 10685 24243 10751 24246
rect 13169 24243 13235 24246
rect 13629 24244 13676 24246
rect 13740 24246 22159 24248
rect 13740 24244 13746 24246
rect 13629 24243 13695 24244
rect 22093 24243 22159 24246
rect 22502 24244 22508 24308
rect 22572 24306 22578 24308
rect 22829 24306 22895 24309
rect 22572 24304 22895 24306
rect 22572 24248 22834 24304
rect 22890 24248 22895 24304
rect 22572 24246 22895 24248
rect 22572 24244 22578 24246
rect 22829 24243 22895 24246
rect 23013 24306 23079 24309
rect 25589 24306 25655 24309
rect 23013 24304 25655 24306
rect 23013 24248 23018 24304
rect 23074 24248 25594 24304
rect 25650 24248 25655 24304
rect 23013 24246 25655 24248
rect 23013 24243 23079 24246
rect 25589 24243 25655 24246
rect 25773 24306 25839 24309
rect 25998 24306 26004 24308
rect 25773 24304 26004 24306
rect 25773 24248 25778 24304
rect 25834 24248 26004 24304
rect 25773 24246 26004 24248
rect 25773 24243 25839 24246
rect 25998 24244 26004 24246
rect 26068 24244 26074 24308
rect 26182 24244 26188 24308
rect 26252 24306 26258 24308
rect 26325 24306 26391 24309
rect 26252 24304 26391 24306
rect 26252 24248 26330 24304
rect 26386 24248 26391 24304
rect 26252 24246 26391 24248
rect 26252 24244 26258 24246
rect 26325 24243 26391 24246
rect 27521 24306 27587 24309
rect 28073 24306 28139 24309
rect 27521 24304 28139 24306
rect 27521 24248 27526 24304
rect 27582 24248 28078 24304
rect 28134 24248 28139 24304
rect 27521 24246 28139 24248
rect 27521 24243 27587 24246
rect 28073 24243 28139 24246
rect 29729 24306 29795 24309
rect 32305 24306 32371 24309
rect 38285 24306 38351 24309
rect 29729 24304 38351 24306
rect 29729 24248 29734 24304
rect 29790 24248 32310 24304
rect 32366 24248 38290 24304
rect 38346 24248 38351 24304
rect 29729 24246 38351 24248
rect 29729 24243 29795 24246
rect 32305 24243 32371 24246
rect 38285 24243 38351 24246
rect 10409 24170 10475 24173
rect 12893 24170 12959 24173
rect 10409 24168 12959 24170
rect 10409 24112 10414 24168
rect 10470 24112 12898 24168
rect 12954 24112 12959 24168
rect 10409 24110 12959 24112
rect 10409 24107 10475 24110
rect 12893 24107 12959 24110
rect 14038 24108 14044 24172
rect 14108 24170 14114 24172
rect 14273 24170 14339 24173
rect 15101 24172 15167 24173
rect 15101 24170 15148 24172
rect 14108 24168 14339 24170
rect 14108 24112 14278 24168
rect 14334 24112 14339 24168
rect 14108 24110 14339 24112
rect 15056 24168 15148 24170
rect 15056 24112 15106 24168
rect 15056 24110 15148 24112
rect 14108 24108 14114 24110
rect 14273 24107 14339 24110
rect 15101 24108 15148 24110
rect 15212 24108 15218 24172
rect 22686 24108 22692 24172
rect 22756 24170 22762 24172
rect 24393 24170 24459 24173
rect 22756 24168 24459 24170
rect 22756 24112 24398 24168
rect 24454 24112 24459 24168
rect 22756 24110 24459 24112
rect 22756 24108 22762 24110
rect 15101 24107 15167 24108
rect 24393 24107 24459 24110
rect 24761 24170 24827 24173
rect 24894 24170 24900 24172
rect 24761 24168 24900 24170
rect 24761 24112 24766 24168
rect 24822 24112 24900 24168
rect 24761 24110 24900 24112
rect 24761 24107 24827 24110
rect 24894 24108 24900 24110
rect 24964 24108 24970 24172
rect 26550 24108 26556 24172
rect 26620 24170 26626 24172
rect 30741 24170 30807 24173
rect 26620 24168 30807 24170
rect 26620 24112 30746 24168
rect 30802 24112 30807 24168
rect 26620 24110 30807 24112
rect 26620 24108 26626 24110
rect 30741 24107 30807 24110
rect 31661 24170 31727 24173
rect 31937 24170 32003 24173
rect 31661 24168 32003 24170
rect 31661 24112 31666 24168
rect 31722 24112 31942 24168
rect 31998 24112 32003 24168
rect 31661 24110 32003 24112
rect 31661 24107 31727 24110
rect 31937 24107 32003 24110
rect 32213 24170 32279 24173
rect 34605 24170 34671 24173
rect 32213 24168 34671 24170
rect 32213 24112 32218 24168
rect 32274 24112 34610 24168
rect 34666 24112 34671 24168
rect 32213 24110 34671 24112
rect 32213 24107 32279 24110
rect 34605 24107 34671 24110
rect 9673 24034 9739 24037
rect 16573 24034 16639 24037
rect 9673 24032 16639 24034
rect 9673 23976 9678 24032
rect 9734 23976 16578 24032
rect 16634 23976 16639 24032
rect 9673 23974 16639 23976
rect 9673 23971 9739 23974
rect 16573 23971 16639 23974
rect 22277 24034 22343 24037
rect 34421 24036 34487 24037
rect 34421 24034 34468 24036
rect 22277 24032 34468 24034
rect 22277 23976 22282 24032
rect 22338 23976 34426 24032
rect 22277 23974 34468 23976
rect 22277 23971 22343 23974
rect 34421 23972 34468 23974
rect 34532 23972 34538 24036
rect 34646 23972 34652 24036
rect 34716 24034 34722 24036
rect 34973 24034 35039 24037
rect 34716 24032 35039 24034
rect 34716 23976 34978 24032
rect 35034 23976 35039 24032
rect 34716 23974 35039 23976
rect 34716 23972 34722 23974
rect 34421 23971 34487 23972
rect 34973 23971 35039 23974
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 8017 23898 8083 23901
rect 10869 23898 10935 23901
rect 13905 23898 13971 23901
rect 8017 23896 13971 23898
rect 8017 23840 8022 23896
rect 8078 23840 10874 23896
rect 10930 23840 13910 23896
rect 13966 23840 13971 23896
rect 8017 23838 13971 23840
rect 8017 23835 8083 23838
rect 10869 23835 10935 23838
rect 13905 23835 13971 23838
rect 15653 23898 15719 23901
rect 26693 23898 26759 23901
rect 15653 23896 26759 23898
rect 15653 23840 15658 23896
rect 15714 23840 26698 23896
rect 26754 23840 26759 23896
rect 15653 23838 26759 23840
rect 15653 23835 15719 23838
rect 26693 23835 26759 23838
rect 29085 23898 29151 23901
rect 29729 23898 29795 23901
rect 29085 23896 29795 23898
rect 29085 23840 29090 23896
rect 29146 23840 29734 23896
rect 29790 23840 29795 23896
rect 29085 23838 29795 23840
rect 29085 23835 29151 23838
rect 29729 23835 29795 23838
rect 31661 23898 31727 23901
rect 34513 23898 34579 23901
rect 31661 23896 34579 23898
rect 31661 23840 31666 23896
rect 31722 23840 34518 23896
rect 34574 23840 34579 23896
rect 31661 23838 34579 23840
rect 31661 23835 31727 23838
rect 34513 23835 34579 23838
rect 44449 23898 44515 23901
rect 45200 23898 46000 23928
rect 44449 23896 46000 23898
rect 44449 23840 44454 23896
rect 44510 23840 46000 23896
rect 44449 23838 46000 23840
rect 44449 23835 44515 23838
rect 45200 23808 46000 23838
rect 5533 23762 5599 23765
rect 21173 23762 21239 23765
rect 5533 23760 21239 23762
rect 5533 23704 5538 23760
rect 5594 23704 21178 23760
rect 21234 23704 21239 23760
rect 5533 23702 21239 23704
rect 5533 23699 5599 23702
rect 21173 23699 21239 23702
rect 22645 23762 22711 23765
rect 25221 23762 25287 23765
rect 22645 23760 25287 23762
rect 22645 23704 22650 23760
rect 22706 23704 25226 23760
rect 25282 23704 25287 23760
rect 22645 23702 25287 23704
rect 22645 23699 22711 23702
rect 25221 23699 25287 23702
rect 25865 23762 25931 23765
rect 26509 23762 26575 23765
rect 25865 23760 26575 23762
rect 25865 23704 25870 23760
rect 25926 23704 26514 23760
rect 26570 23704 26575 23760
rect 25865 23702 26575 23704
rect 25865 23699 25931 23702
rect 26509 23699 26575 23702
rect 26877 23762 26943 23765
rect 27797 23762 27863 23765
rect 26877 23760 27863 23762
rect 26877 23704 26882 23760
rect 26938 23704 27802 23760
rect 27858 23704 27863 23760
rect 26877 23702 27863 23704
rect 26877 23699 26943 23702
rect 27797 23699 27863 23702
rect 30833 23762 30899 23765
rect 30966 23762 30972 23764
rect 30833 23760 30972 23762
rect 30833 23704 30838 23760
rect 30894 23704 30972 23760
rect 30833 23702 30972 23704
rect 30833 23699 30899 23702
rect 30966 23700 30972 23702
rect 31036 23762 31042 23764
rect 36721 23762 36787 23765
rect 31036 23760 36787 23762
rect 31036 23704 36726 23760
rect 36782 23704 36787 23760
rect 31036 23702 36787 23704
rect 31036 23700 31042 23702
rect 36721 23699 36787 23702
rect 37222 23700 37228 23764
rect 37292 23762 37298 23764
rect 38929 23762 38995 23765
rect 37292 23760 38995 23762
rect 37292 23704 38934 23760
rect 38990 23704 38995 23760
rect 37292 23702 38995 23704
rect 37292 23700 37298 23702
rect 38929 23699 38995 23702
rect 7046 23564 7052 23628
rect 7116 23626 7122 23628
rect 7925 23626 7991 23629
rect 7116 23624 7991 23626
rect 7116 23568 7930 23624
rect 7986 23568 7991 23624
rect 7116 23566 7991 23568
rect 7116 23564 7122 23566
rect 7925 23563 7991 23566
rect 13813 23626 13879 23629
rect 19006 23626 19012 23628
rect 13813 23624 19012 23626
rect 13813 23568 13818 23624
rect 13874 23568 19012 23624
rect 13813 23566 19012 23568
rect 13813 23563 13879 23566
rect 19006 23564 19012 23566
rect 19076 23564 19082 23628
rect 22277 23626 22343 23629
rect 24945 23626 25011 23629
rect 31937 23626 32003 23629
rect 37457 23626 37523 23629
rect 22277 23624 29746 23626
rect 22277 23568 22282 23624
rect 22338 23568 24950 23624
rect 25006 23568 29746 23624
rect 22277 23566 29746 23568
rect 22277 23563 22343 23566
rect 24945 23563 25011 23566
rect 7833 23492 7899 23493
rect 7782 23490 7788 23492
rect 7742 23430 7788 23490
rect 7852 23488 7899 23492
rect 7894 23432 7899 23488
rect 7782 23428 7788 23430
rect 7852 23428 7899 23432
rect 7833 23427 7899 23428
rect 11973 23490 12039 23493
rect 12198 23490 12204 23492
rect 11973 23488 12204 23490
rect 11973 23432 11978 23488
rect 12034 23432 12204 23488
rect 11973 23430 12204 23432
rect 11973 23427 12039 23430
rect 12198 23428 12204 23430
rect 12268 23428 12274 23492
rect 18597 23490 18663 23493
rect 19517 23490 19583 23493
rect 18597 23488 19583 23490
rect 18597 23432 18602 23488
rect 18658 23432 19522 23488
rect 19578 23432 19583 23488
rect 18597 23430 19583 23432
rect 18597 23427 18663 23430
rect 19517 23427 19583 23430
rect 19701 23490 19767 23493
rect 22277 23490 22343 23493
rect 22461 23490 22527 23493
rect 25865 23490 25931 23493
rect 19701 23488 22110 23490
rect 19701 23432 19706 23488
rect 19762 23432 22110 23488
rect 19701 23430 22110 23432
rect 19701 23427 19767 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 11646 23292 11652 23356
rect 11716 23354 11722 23356
rect 11881 23354 11947 23357
rect 14181 23354 14247 23357
rect 11716 23352 11947 23354
rect 11716 23296 11886 23352
rect 11942 23296 11947 23352
rect 11716 23294 11947 23296
rect 11716 23292 11722 23294
rect 11881 23291 11947 23294
rect 12988 23352 14247 23354
rect 12988 23296 14186 23352
rect 14242 23296 14247 23352
rect 12988 23294 14247 23296
rect 22050 23354 22110 23430
rect 22277 23488 25931 23490
rect 22277 23432 22282 23488
rect 22338 23432 22466 23488
rect 22522 23432 25870 23488
rect 25926 23432 25931 23488
rect 22277 23430 25931 23432
rect 22277 23427 22343 23430
rect 22461 23427 22527 23430
rect 25865 23427 25931 23430
rect 26233 23490 26299 23493
rect 27797 23490 27863 23493
rect 26233 23488 27863 23490
rect 26233 23432 26238 23488
rect 26294 23432 27802 23488
rect 27858 23432 27863 23488
rect 26233 23430 27863 23432
rect 26233 23427 26299 23430
rect 27797 23427 27863 23430
rect 28165 23490 28231 23493
rect 29310 23490 29316 23492
rect 28165 23488 29316 23490
rect 28165 23432 28170 23488
rect 28226 23432 29316 23488
rect 28165 23430 29316 23432
rect 28165 23427 28231 23430
rect 29310 23428 29316 23430
rect 29380 23428 29386 23492
rect 29686 23490 29746 23566
rect 31937 23624 37523 23626
rect 31937 23568 31942 23624
rect 31998 23568 37462 23624
rect 37518 23568 37523 23624
rect 31937 23566 37523 23568
rect 31937 23563 32003 23566
rect 37457 23563 37523 23566
rect 29821 23490 29887 23493
rect 29686 23488 29887 23490
rect 29686 23432 29826 23488
rect 29882 23432 29887 23488
rect 29686 23430 29887 23432
rect 29821 23427 29887 23430
rect 31886 23428 31892 23492
rect 31956 23490 31962 23492
rect 32765 23490 32831 23493
rect 31956 23488 32831 23490
rect 31956 23432 32770 23488
rect 32826 23432 32831 23488
rect 31956 23430 32831 23432
rect 31956 23428 31962 23430
rect 32765 23427 32831 23430
rect 32949 23492 33015 23493
rect 32949 23488 32996 23492
rect 33060 23490 33066 23492
rect 32949 23432 32954 23488
rect 32949 23428 32996 23432
rect 33060 23430 33106 23490
rect 33060 23428 33066 23430
rect 32949 23427 33015 23428
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 34421 23354 34487 23357
rect 22050 23352 34487 23354
rect 22050 23296 34426 23352
rect 34482 23296 34487 23352
rect 22050 23294 34487 23296
rect 9990 23156 9996 23220
rect 10060 23218 10066 23220
rect 12988 23218 13048 23294
rect 14181 23291 14247 23294
rect 34421 23291 34487 23294
rect 10060 23158 13048 23218
rect 13169 23218 13235 23221
rect 18873 23218 18939 23221
rect 13169 23216 18939 23218
rect 13169 23160 13174 23216
rect 13230 23160 18878 23216
rect 18934 23160 18939 23216
rect 13169 23158 18939 23160
rect 10060 23156 10066 23158
rect 13169 23155 13235 23158
rect 18873 23155 18939 23158
rect 22686 23156 22692 23220
rect 22756 23218 22762 23220
rect 22921 23218 22987 23221
rect 22756 23216 22987 23218
rect 22756 23160 22926 23216
rect 22982 23160 22987 23216
rect 22756 23158 22987 23160
rect 22756 23156 22762 23158
rect 22921 23155 22987 23158
rect 25129 23218 25195 23221
rect 29678 23218 29684 23220
rect 25129 23216 29684 23218
rect 25129 23160 25134 23216
rect 25190 23160 29684 23216
rect 25129 23158 29684 23160
rect 25129 23155 25195 23158
rect 29678 23156 29684 23158
rect 29748 23156 29754 23220
rect 34278 23156 34284 23220
rect 34348 23218 34354 23220
rect 34513 23218 34579 23221
rect 34348 23216 34579 23218
rect 34348 23160 34518 23216
rect 34574 23160 34579 23216
rect 34348 23158 34579 23160
rect 34348 23156 34354 23158
rect 34513 23155 34579 23158
rect 34881 23218 34947 23221
rect 37273 23218 37339 23221
rect 34881 23216 37339 23218
rect 34881 23160 34886 23216
rect 34942 23160 37278 23216
rect 37334 23160 37339 23216
rect 34881 23158 37339 23160
rect 34881 23155 34947 23158
rect 37273 23155 37339 23158
rect 44081 23218 44147 23221
rect 45200 23218 46000 23248
rect 44081 23216 46000 23218
rect 44081 23160 44086 23216
rect 44142 23160 46000 23216
rect 44081 23158 46000 23160
rect 44081 23155 44147 23158
rect 45200 23128 46000 23158
rect 7925 23082 7991 23085
rect 15193 23082 15259 23085
rect 7925 23080 15259 23082
rect 7925 23024 7930 23080
rect 7986 23024 15198 23080
rect 15254 23024 15259 23080
rect 7925 23022 15259 23024
rect 7925 23019 7991 23022
rect 15193 23019 15259 23022
rect 19333 23082 19399 23085
rect 20529 23082 20595 23085
rect 35382 23082 35388 23084
rect 19333 23080 35388 23082
rect 19333 23024 19338 23080
rect 19394 23024 20534 23080
rect 20590 23024 35388 23080
rect 19333 23022 35388 23024
rect 19333 23019 19399 23022
rect 20529 23019 20595 23022
rect 35382 23020 35388 23022
rect 35452 23020 35458 23084
rect 10777 22948 10843 22949
rect 10726 22946 10732 22948
rect 10650 22886 10732 22946
rect 10796 22946 10843 22948
rect 17953 22946 18019 22949
rect 20897 22946 20963 22949
rect 24945 22946 25011 22949
rect 10796 22944 20963 22946
rect 10838 22888 17958 22944
rect 18014 22888 20902 22944
rect 20958 22888 20963 22944
rect 10726 22884 10732 22886
rect 10796 22886 20963 22888
rect 10796 22884 10843 22886
rect 10777 22883 10843 22884
rect 17953 22883 18019 22886
rect 20897 22883 20963 22886
rect 21038 22944 25011 22946
rect 21038 22888 24950 22944
rect 25006 22888 25011 22944
rect 21038 22886 25011 22888
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 13353 22812 13419 22813
rect 13302 22748 13308 22812
rect 13372 22810 13419 22812
rect 14181 22810 14247 22813
rect 18873 22810 18939 22813
rect 19374 22810 19380 22812
rect 13372 22808 13464 22810
rect 13414 22752 13464 22808
rect 13372 22750 13464 22752
rect 14181 22808 16590 22810
rect 14181 22752 14186 22808
rect 14242 22752 16590 22808
rect 14181 22750 16590 22752
rect 13372 22748 13419 22750
rect 13353 22747 13419 22748
rect 14181 22747 14247 22750
rect 4337 22674 4403 22677
rect 5165 22674 5231 22677
rect 5809 22674 5875 22677
rect 4337 22672 5875 22674
rect 4337 22616 4342 22672
rect 4398 22616 5170 22672
rect 5226 22616 5814 22672
rect 5870 22616 5875 22672
rect 4337 22614 5875 22616
rect 4337 22611 4403 22614
rect 5165 22611 5231 22614
rect 5809 22611 5875 22614
rect 10225 22674 10291 22677
rect 12433 22674 12499 22677
rect 14641 22674 14707 22677
rect 10225 22672 14707 22674
rect 10225 22616 10230 22672
rect 10286 22616 12438 22672
rect 12494 22616 14646 22672
rect 14702 22616 14707 22672
rect 10225 22614 14707 22616
rect 16530 22674 16590 22750
rect 18873 22808 19380 22810
rect 18873 22752 18878 22808
rect 18934 22752 19380 22808
rect 18873 22750 19380 22752
rect 18873 22747 18939 22750
rect 19374 22748 19380 22750
rect 19444 22810 19450 22812
rect 19793 22810 19859 22813
rect 19444 22808 19859 22810
rect 19444 22752 19798 22808
rect 19854 22752 19859 22808
rect 19444 22750 19859 22752
rect 19444 22748 19450 22750
rect 19793 22747 19859 22750
rect 20805 22810 20871 22813
rect 21038 22810 21098 22886
rect 24945 22883 25011 22886
rect 25630 22884 25636 22948
rect 25700 22946 25706 22948
rect 27797 22946 27863 22949
rect 31150 22946 31156 22948
rect 25700 22886 27722 22946
rect 25700 22884 25706 22886
rect 20805 22808 21098 22810
rect 20805 22752 20810 22808
rect 20866 22752 21098 22808
rect 20805 22750 21098 22752
rect 23841 22810 23907 22813
rect 27061 22810 27127 22813
rect 23841 22808 27127 22810
rect 23841 22752 23846 22808
rect 23902 22752 27066 22808
rect 27122 22752 27127 22808
rect 23841 22750 27127 22752
rect 27662 22810 27722 22886
rect 27797 22944 31156 22946
rect 27797 22888 27802 22944
rect 27858 22888 31156 22944
rect 27797 22886 31156 22888
rect 27797 22883 27863 22886
rect 31150 22884 31156 22886
rect 31220 22884 31226 22948
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 31753 22810 31819 22813
rect 27662 22808 31819 22810
rect 27662 22752 31758 22808
rect 31814 22752 31819 22808
rect 27662 22750 31819 22752
rect 20805 22747 20871 22750
rect 23841 22747 23907 22750
rect 27061 22747 27127 22750
rect 31753 22747 31819 22750
rect 23289 22674 23355 22677
rect 16530 22672 23355 22674
rect 16530 22616 23294 22672
rect 23350 22616 23355 22672
rect 16530 22614 23355 22616
rect 10225 22611 10291 22614
rect 12433 22611 12499 22614
rect 14641 22611 14707 22614
rect 23289 22611 23355 22614
rect 23473 22674 23539 22677
rect 23933 22674 23999 22677
rect 28257 22674 28323 22677
rect 23473 22672 28323 22674
rect 23473 22616 23478 22672
rect 23534 22616 23938 22672
rect 23994 22616 28262 22672
rect 28318 22616 28323 22672
rect 23473 22614 28323 22616
rect 23473 22611 23539 22614
rect 23933 22611 23999 22614
rect 28257 22611 28323 22614
rect 31937 22674 32003 22677
rect 41873 22674 41939 22677
rect 31937 22672 41939 22674
rect 31937 22616 31942 22672
rect 31998 22616 41878 22672
rect 41934 22616 41939 22672
rect 31937 22614 41939 22616
rect 31937 22611 32003 22614
rect 41873 22611 41939 22614
rect 8886 22476 8892 22540
rect 8956 22538 8962 22540
rect 9121 22538 9187 22541
rect 17902 22538 17908 22540
rect 8956 22536 9187 22538
rect 8956 22480 9126 22536
rect 9182 22480 9187 22536
rect 8956 22478 9187 22480
rect 8956 22476 8962 22478
rect 9121 22475 9187 22478
rect 9262 22478 17908 22538
rect 5073 22402 5139 22405
rect 9262 22402 9322 22478
rect 17902 22476 17908 22478
rect 17972 22476 17978 22540
rect 19333 22538 19399 22541
rect 26141 22538 26207 22541
rect 26877 22538 26943 22541
rect 19333 22536 26207 22538
rect 19333 22480 19338 22536
rect 19394 22480 26146 22536
rect 26202 22480 26207 22536
rect 19333 22478 26207 22480
rect 19333 22475 19399 22478
rect 26141 22475 26207 22478
rect 26374 22536 26943 22538
rect 26374 22480 26882 22536
rect 26938 22480 26943 22536
rect 26374 22478 26943 22480
rect 5073 22400 9322 22402
rect 5073 22344 5078 22400
rect 5134 22344 9322 22400
rect 5073 22342 9322 22344
rect 5073 22339 5139 22342
rect 10726 22340 10732 22404
rect 10796 22402 10802 22404
rect 11053 22402 11119 22405
rect 13813 22402 13879 22405
rect 18270 22402 18276 22404
rect 10796 22400 18276 22402
rect 10796 22344 11058 22400
rect 11114 22344 13818 22400
rect 13874 22344 18276 22400
rect 10796 22342 18276 22344
rect 10796 22340 10802 22342
rect 11053 22339 11119 22342
rect 13813 22339 13879 22342
rect 18270 22340 18276 22342
rect 18340 22402 18346 22404
rect 23565 22402 23631 22405
rect 18340 22400 23631 22402
rect 18340 22344 23570 22400
rect 23626 22344 23631 22400
rect 18340 22342 23631 22344
rect 18340 22340 18346 22342
rect 23565 22339 23631 22342
rect 26233 22402 26299 22405
rect 26374 22402 26434 22478
rect 26877 22475 26943 22478
rect 29361 22538 29427 22541
rect 32581 22538 32647 22541
rect 29361 22536 32647 22538
rect 29361 22480 29366 22536
rect 29422 22480 32586 22536
rect 32642 22480 32647 22536
rect 29361 22478 32647 22480
rect 29361 22475 29427 22478
rect 32581 22475 32647 22478
rect 33041 22538 33107 22541
rect 36445 22538 36511 22541
rect 33041 22536 36511 22538
rect 33041 22480 33046 22536
rect 33102 22480 36450 22536
rect 36506 22480 36511 22536
rect 33041 22478 36511 22480
rect 33041 22475 33107 22478
rect 36445 22475 36511 22478
rect 44449 22538 44515 22541
rect 45200 22538 46000 22568
rect 44449 22536 46000 22538
rect 44449 22480 44454 22536
rect 44510 22480 46000 22536
rect 44449 22478 46000 22480
rect 44449 22475 44515 22478
rect 45200 22448 46000 22478
rect 26233 22400 26434 22402
rect 26233 22344 26238 22400
rect 26294 22344 26434 22400
rect 26233 22342 26434 22344
rect 26233 22339 26299 22342
rect 26550 22340 26556 22404
rect 26620 22402 26626 22404
rect 26785 22402 26851 22405
rect 28993 22404 29059 22405
rect 26620 22400 26851 22402
rect 26620 22344 26790 22400
rect 26846 22344 26851 22400
rect 26620 22342 26851 22344
rect 26620 22340 26626 22342
rect 26785 22339 26851 22342
rect 28942 22340 28948 22404
rect 29012 22402 29059 22404
rect 34513 22402 34579 22405
rect 29012 22400 29104 22402
rect 29054 22344 29104 22400
rect 29012 22342 29104 22344
rect 32446 22400 34579 22402
rect 32446 22344 34518 22400
rect 34574 22344 34579 22400
rect 32446 22342 34579 22344
rect 29012 22340 29059 22342
rect 28993 22339 29059 22340
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 16849 22266 16915 22269
rect 13816 22264 16915 22266
rect 13816 22208 16854 22264
rect 16910 22208 16915 22264
rect 13816 22206 16915 22208
rect 13816 22133 13876 22206
rect 16849 22203 16915 22206
rect 21081 22264 21147 22269
rect 21081 22208 21086 22264
rect 21142 22208 21147 22264
rect 21081 22203 21147 22208
rect 22369 22266 22435 22269
rect 28441 22266 28507 22269
rect 22369 22264 28507 22266
rect 22369 22208 22374 22264
rect 22430 22208 28446 22264
rect 28502 22208 28507 22264
rect 22369 22206 28507 22208
rect 22369 22203 22435 22206
rect 28441 22203 28507 22206
rect 28625 22264 28691 22269
rect 28625 22208 28630 22264
rect 28686 22208 28691 22264
rect 28625 22203 28691 22208
rect 29085 22266 29151 22269
rect 32446 22266 32506 22342
rect 34513 22339 34579 22342
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 32673 22268 32739 22269
rect 32622 22266 32628 22268
rect 29085 22264 32506 22266
rect 29085 22208 29090 22264
rect 29146 22208 32506 22264
rect 29085 22206 32506 22208
rect 32582 22206 32628 22266
rect 32692 22264 32739 22268
rect 32734 22208 32739 22264
rect 29085 22203 29151 22206
rect 32622 22204 32628 22206
rect 32692 22204 32739 22208
rect 32673 22203 32739 22204
rect 34237 22264 34303 22269
rect 34237 22208 34242 22264
rect 34298 22208 34303 22264
rect 34237 22203 34303 22208
rect 11513 22130 11579 22133
rect 13813 22130 13879 22133
rect 11513 22128 13879 22130
rect 11513 22072 11518 22128
rect 11574 22072 13818 22128
rect 13874 22072 13879 22128
rect 11513 22070 13879 22072
rect 11513 22067 11579 22070
rect 13813 22067 13879 22070
rect 16481 22130 16547 22133
rect 20621 22130 20687 22133
rect 16481 22128 20687 22130
rect 16481 22072 16486 22128
rect 16542 22072 20626 22128
rect 20682 22072 20687 22128
rect 16481 22070 20687 22072
rect 16481 22067 16547 22070
rect 20621 22067 20687 22070
rect 20805 22130 20871 22133
rect 21084 22130 21144 22203
rect 20805 22128 21144 22130
rect 20805 22072 20810 22128
rect 20866 22072 21144 22128
rect 20805 22070 21144 22072
rect 20805 22067 20871 22070
rect 24710 22068 24716 22132
rect 24780 22130 24786 22132
rect 27981 22130 28047 22133
rect 24780 22128 28047 22130
rect 24780 22072 27986 22128
rect 28042 22072 28047 22128
rect 24780 22070 28047 22072
rect 24780 22068 24786 22070
rect 27981 22067 28047 22070
rect 7465 21994 7531 21997
rect 11053 21994 11119 21997
rect 11605 21994 11671 21997
rect 7465 21992 11671 21994
rect 7465 21936 7470 21992
rect 7526 21936 11058 21992
rect 11114 21936 11610 21992
rect 11666 21936 11671 21992
rect 7465 21934 11671 21936
rect 7465 21931 7531 21934
rect 11053 21931 11119 21934
rect 11605 21931 11671 21934
rect 12934 21932 12940 21996
rect 13004 21994 13010 21996
rect 13721 21994 13787 21997
rect 13004 21992 13787 21994
rect 13004 21936 13726 21992
rect 13782 21936 13787 21992
rect 13004 21934 13787 21936
rect 13004 21932 13010 21934
rect 13721 21931 13787 21934
rect 14917 21994 14983 21997
rect 17585 21994 17651 21997
rect 14917 21992 17651 21994
rect 14917 21936 14922 21992
rect 14978 21936 17590 21992
rect 17646 21936 17651 21992
rect 14917 21934 17651 21936
rect 14917 21931 14983 21934
rect 17585 21931 17651 21934
rect 21081 21994 21147 21997
rect 24393 21994 24459 21997
rect 21081 21992 24459 21994
rect 21081 21936 21086 21992
rect 21142 21936 24398 21992
rect 24454 21936 24459 21992
rect 21081 21934 24459 21936
rect 21081 21931 21147 21934
rect 24393 21931 24459 21934
rect 25129 21994 25195 21997
rect 25262 21994 25268 21996
rect 25129 21992 25268 21994
rect 25129 21936 25134 21992
rect 25190 21936 25268 21992
rect 25129 21934 25268 21936
rect 25129 21931 25195 21934
rect 25262 21932 25268 21934
rect 25332 21932 25338 21996
rect 25681 21994 25747 21997
rect 28073 21994 28139 21997
rect 25681 21992 28139 21994
rect 25681 21936 25686 21992
rect 25742 21936 28078 21992
rect 28134 21936 28139 21992
rect 25681 21934 28139 21936
rect 25681 21931 25747 21934
rect 28073 21931 28139 21934
rect 28349 21994 28415 21997
rect 28628 21994 28688 22203
rect 34240 21997 34300 22203
rect 28349 21992 28688 21994
rect 28349 21936 28354 21992
rect 28410 21936 28688 21992
rect 28349 21934 28688 21936
rect 28349 21931 28415 21934
rect 32438 21932 32444 21996
rect 32508 21994 32514 21996
rect 32857 21994 32923 21997
rect 33225 21994 33291 21997
rect 32508 21992 33291 21994
rect 32508 21936 32862 21992
rect 32918 21936 33230 21992
rect 33286 21936 33291 21992
rect 32508 21934 33291 21936
rect 32508 21932 32514 21934
rect 32857 21931 32923 21934
rect 33225 21931 33291 21934
rect 33593 21994 33659 21997
rect 33593 21992 34162 21994
rect 33593 21936 33598 21992
rect 33654 21936 34162 21992
rect 33593 21934 34162 21936
rect 33593 21931 33659 21934
rect 9673 21858 9739 21861
rect 14733 21858 14799 21861
rect 9673 21856 14799 21858
rect 9673 21800 9678 21856
rect 9734 21800 14738 21856
rect 14794 21800 14799 21856
rect 9673 21798 14799 21800
rect 9673 21795 9739 21798
rect 14733 21795 14799 21798
rect 17902 21796 17908 21860
rect 17972 21858 17978 21860
rect 24853 21858 24919 21861
rect 32213 21858 32279 21861
rect 34102 21858 34162 21934
rect 34237 21992 34303 21997
rect 34237 21936 34242 21992
rect 34298 21936 34303 21992
rect 34237 21931 34303 21936
rect 34646 21932 34652 21996
rect 34716 21994 34722 21996
rect 35525 21994 35591 21997
rect 36302 21994 36308 21996
rect 34716 21992 36308 21994
rect 34716 21936 35530 21992
rect 35586 21936 36308 21992
rect 34716 21934 36308 21936
rect 34716 21932 34722 21934
rect 35525 21931 35591 21934
rect 36302 21932 36308 21934
rect 36372 21932 36378 21996
rect 34237 21858 34303 21861
rect 17972 21856 34024 21858
rect 17972 21800 24858 21856
rect 24914 21800 32218 21856
rect 32274 21800 34024 21856
rect 17972 21798 34024 21800
rect 34102 21856 34303 21858
rect 34102 21800 34242 21856
rect 34298 21800 34303 21856
rect 34102 21798 34303 21800
rect 17972 21796 17978 21798
rect 24853 21795 24919 21798
rect 32213 21795 32279 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 11605 21722 11671 21725
rect 14917 21722 14983 21725
rect 11605 21720 14983 21722
rect 11605 21664 11610 21720
rect 11666 21664 14922 21720
rect 14978 21664 14983 21720
rect 11605 21662 14983 21664
rect 11605 21659 11671 21662
rect 14917 21659 14983 21662
rect 16941 21722 17007 21725
rect 21582 21722 21588 21724
rect 16941 21720 21588 21722
rect 16941 21664 16946 21720
rect 17002 21664 21588 21720
rect 16941 21662 21588 21664
rect 16941 21659 17007 21662
rect 21582 21660 21588 21662
rect 21652 21660 21658 21724
rect 24485 21722 24551 21725
rect 29177 21722 29243 21725
rect 32581 21722 32647 21725
rect 33225 21724 33291 21725
rect 24485 21720 32647 21722
rect 24485 21664 24490 21720
rect 24546 21664 29182 21720
rect 29238 21664 32586 21720
rect 32642 21664 32647 21720
rect 24485 21662 32647 21664
rect 24485 21659 24551 21662
rect 29177 21659 29243 21662
rect 32581 21659 32647 21662
rect 33174 21660 33180 21724
rect 33244 21722 33291 21724
rect 33501 21722 33567 21725
rect 33244 21720 33567 21722
rect 33286 21664 33506 21720
rect 33562 21664 33567 21720
rect 33244 21662 33567 21664
rect 33964 21722 34024 21798
rect 34237 21795 34303 21798
rect 44449 21858 44515 21861
rect 45200 21858 46000 21888
rect 44449 21856 46000 21858
rect 44449 21800 44454 21856
rect 44510 21800 46000 21856
rect 44449 21798 46000 21800
rect 44449 21795 44515 21798
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 45200 21768 46000 21798
rect 35590 21727 35906 21728
rect 35065 21722 35131 21725
rect 33964 21720 35131 21722
rect 33964 21664 35070 21720
rect 35126 21664 35131 21720
rect 33964 21662 35131 21664
rect 33244 21660 33291 21662
rect 33225 21659 33291 21660
rect 33501 21659 33567 21662
rect 35065 21659 35131 21662
rect 5257 21586 5323 21589
rect 5441 21586 5507 21589
rect 18321 21586 18387 21589
rect 25957 21588 26023 21589
rect 22318 21586 22324 21588
rect 5257 21584 22324 21586
rect 5257 21528 5262 21584
rect 5318 21528 5446 21584
rect 5502 21528 18326 21584
rect 18382 21528 22324 21584
rect 5257 21526 22324 21528
rect 5257 21523 5323 21526
rect 5441 21523 5507 21526
rect 18321 21523 18387 21526
rect 22318 21524 22324 21526
rect 22388 21586 22394 21588
rect 25957 21586 26004 21588
rect 22388 21526 24962 21586
rect 25912 21584 26004 21586
rect 25912 21528 25962 21584
rect 25912 21526 26004 21528
rect 22388 21524 22394 21526
rect 7465 21450 7531 21453
rect 8845 21450 8911 21453
rect 7465 21448 8911 21450
rect 7465 21392 7470 21448
rect 7526 21392 8850 21448
rect 8906 21392 8911 21448
rect 7465 21390 8911 21392
rect 7465 21387 7531 21390
rect 8845 21387 8911 21390
rect 12525 21450 12591 21453
rect 13261 21450 13327 21453
rect 12525 21448 13327 21450
rect 12525 21392 12530 21448
rect 12586 21392 13266 21448
rect 13322 21392 13327 21448
rect 12525 21390 13327 21392
rect 12525 21387 12591 21390
rect 13261 21387 13327 21390
rect 14457 21450 14523 21453
rect 15745 21450 15811 21453
rect 14457 21448 15811 21450
rect 14457 21392 14462 21448
rect 14518 21392 15750 21448
rect 15806 21392 15811 21448
rect 14457 21390 15811 21392
rect 14457 21387 14523 21390
rect 15745 21387 15811 21390
rect 23749 21450 23815 21453
rect 24669 21450 24735 21453
rect 23749 21448 24735 21450
rect 23749 21392 23754 21448
rect 23810 21392 24674 21448
rect 24730 21392 24735 21448
rect 23749 21390 24735 21392
rect 24902 21450 24962 21526
rect 25957 21524 26004 21526
rect 26068 21524 26074 21588
rect 26141 21586 26207 21589
rect 28165 21586 28231 21589
rect 36813 21586 36879 21589
rect 37457 21586 37523 21589
rect 26141 21584 37523 21586
rect 26141 21528 26146 21584
rect 26202 21528 28170 21584
rect 28226 21528 36818 21584
rect 36874 21528 37462 21584
rect 37518 21528 37523 21584
rect 26141 21526 37523 21528
rect 25957 21523 26023 21524
rect 26141 21523 26207 21526
rect 28165 21523 28231 21526
rect 36813 21523 36879 21526
rect 37457 21523 37523 21526
rect 29361 21450 29427 21453
rect 24902 21448 29427 21450
rect 24902 21392 29366 21448
rect 29422 21392 29427 21448
rect 24902 21390 29427 21392
rect 23749 21387 23815 21390
rect 24669 21387 24735 21390
rect 29361 21387 29427 21390
rect 29729 21450 29795 21453
rect 32305 21450 32371 21453
rect 29729 21448 32371 21450
rect 29729 21392 29734 21448
rect 29790 21392 32310 21448
rect 32366 21392 32371 21448
rect 29729 21390 32371 21392
rect 29729 21387 29795 21390
rect 32305 21387 32371 21390
rect 10225 21314 10291 21317
rect 11973 21314 12039 21317
rect 10225 21312 12039 21314
rect 10225 21256 10230 21312
rect 10286 21256 11978 21312
rect 12034 21256 12039 21312
rect 10225 21254 12039 21256
rect 10225 21251 10291 21254
rect 11973 21251 12039 21254
rect 12341 21314 12407 21317
rect 13077 21314 13143 21317
rect 12341 21312 13143 21314
rect 12341 21256 12346 21312
rect 12402 21256 13082 21312
rect 13138 21256 13143 21312
rect 12341 21254 13143 21256
rect 12341 21251 12407 21254
rect 13077 21251 13143 21254
rect 13353 21314 13419 21317
rect 21081 21314 21147 21317
rect 26141 21314 26207 21317
rect 13353 21312 21147 21314
rect 13353 21256 13358 21312
rect 13414 21256 21086 21312
rect 21142 21256 21147 21312
rect 13353 21254 21147 21256
rect 13353 21251 13419 21254
rect 21081 21251 21147 21254
rect 24902 21312 26207 21314
rect 24902 21256 26146 21312
rect 26202 21256 26207 21312
rect 24902 21254 26207 21256
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 7005 21178 7071 21181
rect 24902 21178 24962 21254
rect 26141 21251 26207 21254
rect 33225 21314 33291 21317
rect 34053 21314 34119 21317
rect 33225 21312 34119 21314
rect 33225 21256 33230 21312
rect 33286 21256 34058 21312
rect 34114 21256 34119 21312
rect 33225 21254 34119 21256
rect 33225 21251 33291 21254
rect 34053 21251 34119 21254
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 25129 21180 25195 21181
rect 26417 21180 26483 21181
rect 7005 21176 24962 21178
rect 7005 21120 7010 21176
rect 7066 21120 24962 21176
rect 7005 21118 24962 21120
rect 7005 21115 7071 21118
rect 25078 21116 25084 21180
rect 25148 21178 25195 21180
rect 25148 21176 25240 21178
rect 25190 21120 25240 21176
rect 25148 21118 25240 21120
rect 25148 21116 25195 21118
rect 26366 21116 26372 21180
rect 26436 21178 26483 21180
rect 26436 21176 26528 21178
rect 26478 21120 26528 21176
rect 26436 21118 26528 21120
rect 26436 21116 26483 21118
rect 27286 21116 27292 21180
rect 27356 21178 27362 21180
rect 33961 21178 34027 21181
rect 27356 21176 34027 21178
rect 27356 21120 33966 21176
rect 34022 21120 34027 21176
rect 27356 21118 34027 21120
rect 27356 21116 27362 21118
rect 25129 21115 25195 21116
rect 26417 21115 26483 21116
rect 33961 21115 34027 21118
rect 44449 21178 44515 21181
rect 45200 21178 46000 21208
rect 44449 21176 46000 21178
rect 44449 21120 44454 21176
rect 44510 21120 46000 21176
rect 44449 21118 46000 21120
rect 44449 21115 44515 21118
rect 45200 21088 46000 21118
rect 9673 21042 9739 21045
rect 11605 21042 11671 21045
rect 9673 21040 11671 21042
rect 9673 20984 9678 21040
rect 9734 20984 11610 21040
rect 11666 20984 11671 21040
rect 9673 20982 11671 20984
rect 9673 20979 9739 20982
rect 11605 20979 11671 20982
rect 12249 21042 12315 21045
rect 12525 21042 12591 21045
rect 12249 21040 12591 21042
rect 12249 20984 12254 21040
rect 12310 20984 12530 21040
rect 12586 20984 12591 21040
rect 12249 20982 12591 20984
rect 12249 20979 12315 20982
rect 12525 20979 12591 20982
rect 12985 21042 13051 21045
rect 13353 21042 13419 21045
rect 24485 21042 24551 21045
rect 12985 21040 13419 21042
rect 12985 20984 12990 21040
rect 13046 20984 13358 21040
rect 13414 20984 13419 21040
rect 12985 20982 13419 20984
rect 12985 20979 13051 20982
rect 13353 20979 13419 20982
rect 18094 21040 24551 21042
rect 18094 20984 24490 21040
rect 24546 20984 24551 21040
rect 18094 20982 24551 20984
rect 9029 20906 9095 20909
rect 17217 20906 17283 20909
rect 9029 20904 17283 20906
rect 9029 20848 9034 20904
rect 9090 20848 17222 20904
rect 17278 20848 17283 20904
rect 9029 20846 17283 20848
rect 9029 20843 9095 20846
rect 17217 20843 17283 20846
rect 17585 20906 17651 20909
rect 18094 20906 18154 20982
rect 24485 20979 24551 20982
rect 24853 21042 24919 21045
rect 27889 21042 27955 21045
rect 24853 21040 27955 21042
rect 24853 20984 24858 21040
rect 24914 20984 27894 21040
rect 27950 20984 27955 21040
rect 24853 20982 27955 20984
rect 24853 20979 24919 20982
rect 27889 20979 27955 20982
rect 28441 21042 28507 21045
rect 29269 21042 29335 21045
rect 28441 21040 29335 21042
rect 28441 20984 28446 21040
rect 28502 20984 29274 21040
rect 29330 20984 29335 21040
rect 28441 20982 29335 20984
rect 28441 20979 28507 20982
rect 29269 20979 29335 20982
rect 34329 21042 34395 21045
rect 36537 21042 36603 21045
rect 34329 21040 36603 21042
rect 34329 20984 34334 21040
rect 34390 20984 36542 21040
rect 36598 20984 36603 21040
rect 34329 20982 36603 20984
rect 34329 20979 34395 20982
rect 36537 20979 36603 20982
rect 17585 20904 18154 20906
rect 17585 20848 17590 20904
rect 17646 20848 18154 20904
rect 17585 20846 18154 20848
rect 17585 20843 17651 20846
rect 20662 20844 20668 20908
rect 20732 20906 20738 20908
rect 22829 20906 22895 20909
rect 35433 20906 35499 20909
rect 20732 20904 22895 20906
rect 20732 20848 22834 20904
rect 22890 20848 22895 20904
rect 20732 20846 22895 20848
rect 20732 20844 20738 20846
rect 22829 20843 22895 20846
rect 23062 20904 35499 20906
rect 23062 20848 35438 20904
rect 35494 20848 35499 20904
rect 23062 20846 35499 20848
rect 8201 20770 8267 20773
rect 11697 20770 11763 20773
rect 8201 20768 11763 20770
rect 8201 20712 8206 20768
rect 8262 20712 11702 20768
rect 11758 20712 11763 20768
rect 8201 20710 11763 20712
rect 8201 20707 8267 20710
rect 11697 20707 11763 20710
rect 11973 20770 12039 20773
rect 12617 20770 12683 20773
rect 11973 20768 12683 20770
rect 11973 20712 11978 20768
rect 12034 20712 12622 20768
rect 12678 20712 12683 20768
rect 11973 20710 12683 20712
rect 11973 20707 12039 20710
rect 12617 20707 12683 20710
rect 12801 20770 12867 20773
rect 12934 20770 12940 20772
rect 12801 20768 12940 20770
rect 12801 20712 12806 20768
rect 12862 20712 12940 20768
rect 12801 20710 12940 20712
rect 12801 20707 12867 20710
rect 12934 20708 12940 20710
rect 13004 20708 13010 20772
rect 13445 20770 13511 20773
rect 13445 20768 13554 20770
rect 13445 20712 13450 20768
rect 13506 20712 13554 20768
rect 13445 20707 13554 20712
rect 17902 20708 17908 20772
rect 17972 20770 17978 20772
rect 18137 20770 18203 20773
rect 17972 20768 18203 20770
rect 17972 20712 18142 20768
rect 18198 20712 18203 20768
rect 17972 20710 18203 20712
rect 17972 20708 17978 20710
rect 18137 20707 18203 20710
rect 21582 20708 21588 20772
rect 21652 20770 21658 20772
rect 23062 20770 23122 20846
rect 35433 20843 35499 20846
rect 23289 20772 23355 20773
rect 21652 20710 23122 20770
rect 21652 20708 21658 20710
rect 23238 20708 23244 20772
rect 23308 20770 23355 20772
rect 24209 20770 24275 20773
rect 24485 20770 24551 20773
rect 26785 20770 26851 20773
rect 23308 20768 23400 20770
rect 23350 20712 23400 20768
rect 23308 20710 23400 20712
rect 24209 20768 24551 20770
rect 24209 20712 24214 20768
rect 24270 20712 24490 20768
rect 24546 20712 24551 20768
rect 24209 20710 24551 20712
rect 23308 20708 23355 20710
rect 23289 20707 23355 20708
rect 24209 20707 24275 20710
rect 24485 20707 24551 20710
rect 24902 20768 26851 20770
rect 24902 20712 26790 20768
rect 26846 20712 26851 20768
rect 24902 20710 26851 20712
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 8845 20634 8911 20637
rect 9438 20634 9444 20636
rect 8845 20632 9444 20634
rect 8845 20576 8850 20632
rect 8906 20576 9444 20632
rect 8845 20574 9444 20576
rect 8845 20571 8911 20574
rect 9438 20572 9444 20574
rect 9508 20634 9514 20636
rect 9581 20634 9647 20637
rect 9508 20632 9647 20634
rect 9508 20576 9586 20632
rect 9642 20576 9647 20632
rect 9508 20574 9647 20576
rect 9508 20572 9514 20574
rect 9581 20571 9647 20574
rect 13169 20634 13235 20637
rect 13302 20634 13308 20636
rect 13169 20632 13308 20634
rect 13169 20576 13174 20632
rect 13230 20576 13308 20632
rect 13169 20574 13308 20576
rect 13169 20571 13235 20574
rect 13302 20572 13308 20574
rect 13372 20572 13378 20636
rect 10501 20498 10567 20501
rect 13077 20498 13143 20501
rect 10501 20496 13143 20498
rect 10501 20440 10506 20496
rect 10562 20440 13082 20496
rect 13138 20440 13143 20496
rect 10501 20438 13143 20440
rect 13494 20498 13554 20707
rect 16849 20634 16915 20637
rect 23933 20634 23999 20637
rect 24902 20634 24962 20710
rect 26785 20707 26851 20710
rect 26969 20770 27035 20773
rect 27102 20770 27108 20772
rect 26969 20768 27108 20770
rect 26969 20712 26974 20768
rect 27030 20712 27108 20768
rect 26969 20710 27108 20712
rect 26969 20707 27035 20710
rect 27102 20708 27108 20710
rect 27172 20708 27178 20772
rect 27470 20708 27476 20772
rect 27540 20770 27546 20772
rect 27705 20770 27771 20773
rect 27540 20768 27771 20770
rect 27540 20712 27710 20768
rect 27766 20712 27771 20768
rect 27540 20710 27771 20712
rect 27540 20708 27546 20710
rect 27705 20707 27771 20710
rect 27889 20770 27955 20773
rect 32213 20770 32279 20773
rect 27889 20768 32279 20770
rect 27889 20712 27894 20768
rect 27950 20712 32218 20768
rect 32274 20712 32279 20768
rect 27889 20710 32279 20712
rect 27889 20707 27955 20710
rect 32213 20707 32279 20710
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 16849 20632 24962 20634
rect 16849 20576 16854 20632
rect 16910 20576 23938 20632
rect 23994 20576 24962 20632
rect 16849 20574 24962 20576
rect 26049 20634 26115 20637
rect 26182 20634 26188 20636
rect 26049 20632 26188 20634
rect 26049 20576 26054 20632
rect 26110 20576 26188 20632
rect 26049 20574 26188 20576
rect 16849 20571 16915 20574
rect 23933 20571 23999 20574
rect 26049 20571 26115 20574
rect 26182 20572 26188 20574
rect 26252 20634 26258 20636
rect 27245 20634 27311 20637
rect 27981 20636 28047 20637
rect 27981 20634 28028 20636
rect 26252 20632 27311 20634
rect 26252 20576 27250 20632
rect 27306 20576 27311 20632
rect 26252 20574 27311 20576
rect 27936 20632 28028 20634
rect 27936 20576 27986 20632
rect 27936 20574 28028 20576
rect 26252 20572 26258 20574
rect 27245 20571 27311 20574
rect 27981 20572 28028 20574
rect 28092 20572 28098 20636
rect 29310 20572 29316 20636
rect 29380 20634 29386 20636
rect 30005 20634 30071 20637
rect 29380 20632 30071 20634
rect 29380 20576 30010 20632
rect 30066 20576 30071 20632
rect 29380 20574 30071 20576
rect 29380 20572 29386 20574
rect 27981 20571 28047 20572
rect 30005 20571 30071 20574
rect 30925 20634 30991 20637
rect 31385 20634 31451 20637
rect 30925 20632 31451 20634
rect 30925 20576 30930 20632
rect 30986 20576 31390 20632
rect 31446 20576 31451 20632
rect 30925 20574 31451 20576
rect 30925 20571 30991 20574
rect 31385 20571 31451 20574
rect 31569 20634 31635 20637
rect 32254 20634 32260 20636
rect 31569 20632 32260 20634
rect 31569 20576 31574 20632
rect 31630 20576 32260 20632
rect 31569 20574 32260 20576
rect 31569 20571 31635 20574
rect 32254 20572 32260 20574
rect 32324 20572 32330 20636
rect 24209 20498 24275 20501
rect 32622 20498 32628 20500
rect 13494 20438 22110 20498
rect 10501 20435 10567 20438
rect 13077 20435 13143 20438
rect 9397 20362 9463 20365
rect 10041 20362 10107 20365
rect 9397 20360 10107 20362
rect 9397 20304 9402 20360
rect 9458 20304 10046 20360
rect 10102 20304 10107 20360
rect 9397 20302 10107 20304
rect 9397 20299 9463 20302
rect 10041 20299 10107 20302
rect 10501 20362 10567 20365
rect 10726 20362 10732 20364
rect 10501 20360 10732 20362
rect 10501 20304 10506 20360
rect 10562 20304 10732 20360
rect 10501 20302 10732 20304
rect 10501 20299 10567 20302
rect 10726 20300 10732 20302
rect 10796 20300 10802 20364
rect 15326 20362 15332 20364
rect 11102 20302 15332 20362
rect 5993 20226 6059 20229
rect 11102 20226 11162 20302
rect 15326 20300 15332 20302
rect 15396 20362 15402 20364
rect 16481 20362 16547 20365
rect 15396 20360 16547 20362
rect 15396 20304 16486 20360
rect 16542 20304 16547 20360
rect 15396 20302 16547 20304
rect 15396 20300 15402 20302
rect 16481 20299 16547 20302
rect 18229 20362 18295 20365
rect 18505 20362 18571 20365
rect 18229 20360 18571 20362
rect 18229 20304 18234 20360
rect 18290 20304 18510 20360
rect 18566 20304 18571 20360
rect 18229 20302 18571 20304
rect 22050 20362 22110 20438
rect 24209 20496 32628 20498
rect 24209 20440 24214 20496
rect 24270 20440 32628 20496
rect 24209 20438 32628 20440
rect 24209 20435 24275 20438
rect 32622 20436 32628 20438
rect 32692 20498 32698 20500
rect 40217 20498 40283 20501
rect 32692 20496 40283 20498
rect 32692 20440 40222 20496
rect 40278 20440 40283 20496
rect 32692 20438 40283 20440
rect 32692 20436 32698 20438
rect 40217 20435 40283 20438
rect 44081 20498 44147 20501
rect 45200 20498 46000 20528
rect 44081 20496 46000 20498
rect 44081 20440 44086 20496
rect 44142 20440 46000 20496
rect 44081 20438 46000 20440
rect 44081 20435 44147 20438
rect 45200 20408 46000 20438
rect 29085 20362 29151 20365
rect 22050 20360 29151 20362
rect 22050 20304 29090 20360
rect 29146 20304 29151 20360
rect 22050 20302 29151 20304
rect 18229 20299 18295 20302
rect 18505 20299 18571 20302
rect 29085 20299 29151 20302
rect 29310 20300 29316 20364
rect 29380 20362 29386 20364
rect 31569 20362 31635 20365
rect 34605 20362 34671 20365
rect 29380 20360 31635 20362
rect 29380 20304 31574 20360
rect 31630 20304 31635 20360
rect 29380 20302 31635 20304
rect 29380 20300 29386 20302
rect 31569 20299 31635 20302
rect 31710 20360 34671 20362
rect 31710 20304 34610 20360
rect 34666 20304 34671 20360
rect 31710 20302 34671 20304
rect 5993 20224 11162 20226
rect 5993 20168 5998 20224
rect 6054 20168 11162 20224
rect 5993 20166 11162 20168
rect 11513 20226 11579 20229
rect 22645 20226 22711 20229
rect 23381 20226 23447 20229
rect 11513 20224 23447 20226
rect 11513 20168 11518 20224
rect 11574 20168 22650 20224
rect 22706 20168 23386 20224
rect 23442 20168 23447 20224
rect 11513 20166 23447 20168
rect 5993 20163 6059 20166
rect 11513 20163 11579 20166
rect 22645 20163 22711 20166
rect 23381 20163 23447 20166
rect 24894 20164 24900 20228
rect 24964 20226 24970 20228
rect 31710 20226 31770 20302
rect 34605 20299 34671 20302
rect 24964 20166 31770 20226
rect 24964 20164 24970 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 9397 20090 9463 20093
rect 18781 20090 18847 20093
rect 9397 20088 18847 20090
rect 9397 20032 9402 20088
rect 9458 20032 18786 20088
rect 18842 20032 18847 20088
rect 9397 20030 18847 20032
rect 9397 20027 9463 20030
rect 18781 20027 18847 20030
rect 18965 20090 19031 20093
rect 28993 20092 29059 20093
rect 25262 20090 25268 20092
rect 18965 20088 25268 20090
rect 18965 20032 18970 20088
rect 19026 20032 25268 20088
rect 18965 20030 25268 20032
rect 18965 20027 19031 20030
rect 25262 20028 25268 20030
rect 25332 20028 25338 20092
rect 28942 20028 28948 20092
rect 29012 20090 29059 20092
rect 29269 20090 29335 20093
rect 33961 20090 34027 20093
rect 29012 20088 29104 20090
rect 29054 20032 29104 20088
rect 29012 20030 29104 20032
rect 29269 20088 34027 20090
rect 29269 20032 29274 20088
rect 29330 20032 33966 20088
rect 34022 20032 34027 20088
rect 29269 20030 34027 20032
rect 29012 20028 29059 20030
rect 28993 20027 29059 20028
rect 29269 20027 29335 20030
rect 33961 20027 34027 20030
rect 9438 19892 9444 19956
rect 9508 19954 9514 19956
rect 9581 19954 9647 19957
rect 9508 19952 9647 19954
rect 9508 19896 9586 19952
rect 9642 19896 9647 19952
rect 9508 19894 9647 19896
rect 9508 19892 9514 19894
rect 9581 19891 9647 19894
rect 9765 19956 9831 19957
rect 10501 19956 10567 19957
rect 9765 19952 9812 19956
rect 9876 19954 9882 19956
rect 10501 19954 10548 19956
rect 9765 19896 9770 19952
rect 9765 19892 9812 19896
rect 9876 19894 9922 19954
rect 10460 19952 10548 19954
rect 10612 19954 10618 19956
rect 20989 19954 21055 19957
rect 10612 19952 21055 19954
rect 10460 19896 10506 19952
rect 10612 19896 20994 19952
rect 21050 19896 21055 19952
rect 10460 19894 10548 19896
rect 9876 19892 9882 19894
rect 10501 19892 10548 19894
rect 10612 19894 21055 19896
rect 10612 19892 10618 19894
rect 9765 19891 9831 19892
rect 10501 19891 10567 19892
rect 20989 19891 21055 19894
rect 21265 19954 21331 19957
rect 25681 19954 25747 19957
rect 37089 19954 37155 19957
rect 21265 19952 37155 19954
rect 21265 19896 21270 19952
rect 21326 19896 25686 19952
rect 25742 19896 37094 19952
rect 37150 19896 37155 19952
rect 21265 19894 37155 19896
rect 21265 19891 21331 19894
rect 25681 19891 25747 19894
rect 37089 19891 37155 19894
rect 8293 19818 8359 19821
rect 33961 19818 34027 19821
rect 34094 19818 34100 19820
rect 8293 19816 31770 19818
rect 8293 19760 8298 19816
rect 8354 19760 31770 19816
rect 8293 19758 31770 19760
rect 8293 19755 8359 19758
rect 22142 19685 22202 19758
rect 5717 19682 5783 19685
rect 18229 19682 18295 19685
rect 5717 19680 18295 19682
rect 5717 19624 5722 19680
rect 5778 19624 18234 19680
rect 18290 19624 18295 19680
rect 5717 19622 18295 19624
rect 5717 19619 5783 19622
rect 18229 19619 18295 19622
rect 22093 19680 22202 19685
rect 22093 19624 22098 19680
rect 22154 19624 22202 19680
rect 22093 19622 22202 19624
rect 23105 19682 23171 19685
rect 26509 19682 26575 19685
rect 23105 19680 26575 19682
rect 23105 19624 23110 19680
rect 23166 19624 26514 19680
rect 26570 19624 26575 19680
rect 23105 19622 26575 19624
rect 22093 19619 22159 19622
rect 23105 19619 23171 19622
rect 26509 19619 26575 19622
rect 27429 19682 27495 19685
rect 29269 19682 29335 19685
rect 30557 19684 30623 19685
rect 30557 19682 30604 19684
rect 27429 19680 29335 19682
rect 27429 19624 27434 19680
rect 27490 19624 29274 19680
rect 29330 19624 29335 19680
rect 27429 19622 29335 19624
rect 30512 19680 30604 19682
rect 30668 19682 30674 19684
rect 31150 19682 31156 19684
rect 30512 19624 30562 19680
rect 30512 19622 30604 19624
rect 27429 19619 27495 19622
rect 29269 19619 29335 19622
rect 30557 19620 30604 19622
rect 30668 19622 31156 19682
rect 30668 19620 30674 19622
rect 31150 19620 31156 19622
rect 31220 19620 31226 19684
rect 30557 19619 30623 19620
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 11830 19484 11836 19548
rect 11900 19546 11906 19548
rect 12893 19546 12959 19549
rect 11900 19544 12959 19546
rect 11900 19488 12898 19544
rect 12954 19488 12959 19544
rect 11900 19486 12959 19488
rect 11900 19484 11906 19486
rect 12893 19483 12959 19486
rect 13261 19546 13327 19549
rect 14089 19546 14155 19549
rect 13261 19544 14155 19546
rect 13261 19488 13266 19544
rect 13322 19488 14094 19544
rect 14150 19488 14155 19544
rect 13261 19486 14155 19488
rect 13261 19483 13327 19486
rect 14089 19483 14155 19486
rect 14365 19546 14431 19549
rect 18505 19546 18571 19549
rect 14365 19544 18571 19546
rect 14365 19488 14370 19544
rect 14426 19488 18510 19544
rect 18566 19488 18571 19544
rect 14365 19486 18571 19488
rect 14365 19483 14431 19486
rect 18505 19483 18571 19486
rect 20161 19546 20227 19549
rect 21950 19546 21956 19548
rect 20161 19544 21956 19546
rect 20161 19488 20166 19544
rect 20222 19488 21956 19544
rect 20161 19486 21956 19488
rect 20161 19483 20227 19486
rect 21950 19484 21956 19486
rect 22020 19484 22026 19548
rect 22645 19546 22711 19549
rect 29310 19546 29316 19548
rect 22645 19544 29316 19546
rect 22645 19488 22650 19544
rect 22706 19488 29316 19544
rect 22645 19486 29316 19488
rect 22645 19483 22711 19486
rect 29310 19484 29316 19486
rect 29380 19484 29386 19548
rect 29729 19546 29795 19549
rect 31385 19546 31451 19549
rect 29729 19544 31451 19546
rect 29729 19488 29734 19544
rect 29790 19488 31390 19544
rect 31446 19488 31451 19544
rect 29729 19486 31451 19488
rect 31710 19546 31770 19758
rect 33961 19816 34100 19818
rect 33961 19760 33966 19816
rect 34022 19760 34100 19816
rect 33961 19758 34100 19760
rect 33961 19755 34027 19758
rect 34094 19756 34100 19758
rect 34164 19756 34170 19820
rect 34513 19818 34579 19821
rect 34646 19818 34652 19820
rect 34513 19816 34652 19818
rect 34513 19760 34518 19816
rect 34574 19760 34652 19816
rect 34513 19758 34652 19760
rect 34513 19755 34579 19758
rect 34646 19756 34652 19758
rect 34716 19756 34722 19820
rect 44449 19818 44515 19821
rect 45200 19818 46000 19848
rect 44449 19816 46000 19818
rect 44449 19760 44454 19816
rect 44510 19760 46000 19816
rect 44449 19758 46000 19760
rect 44449 19755 44515 19758
rect 45200 19728 46000 19758
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 32305 19546 32371 19549
rect 31710 19544 32371 19546
rect 31710 19488 32310 19544
rect 32366 19488 32371 19544
rect 31710 19486 32371 19488
rect 29729 19483 29795 19486
rect 31385 19483 31451 19486
rect 32305 19483 32371 19486
rect 2497 19410 2563 19413
rect 8845 19410 8911 19413
rect 15101 19412 15167 19413
rect 15101 19410 15148 19412
rect 2497 19408 8911 19410
rect 2497 19352 2502 19408
rect 2558 19352 8850 19408
rect 8906 19352 8911 19408
rect 2497 19350 8911 19352
rect 15056 19408 15148 19410
rect 15056 19352 15106 19408
rect 15056 19350 15148 19352
rect 2497 19347 2563 19350
rect 8845 19347 8911 19350
rect 15101 19348 15148 19350
rect 15212 19348 15218 19412
rect 18873 19410 18939 19413
rect 27337 19412 27403 19413
rect 18873 19408 19074 19410
rect 18873 19352 18878 19408
rect 18934 19352 19074 19408
rect 18873 19350 19074 19352
rect 15101 19347 15167 19348
rect 18873 19347 18939 19350
rect 8293 19274 8359 19277
rect 8702 19274 8708 19276
rect 8293 19272 8708 19274
rect 8293 19216 8298 19272
rect 8354 19216 8708 19272
rect 8293 19214 8708 19216
rect 8293 19211 8359 19214
rect 8702 19212 8708 19214
rect 8772 19212 8778 19276
rect 11973 19274 12039 19277
rect 12709 19274 12775 19277
rect 11973 19272 12775 19274
rect 11973 19216 11978 19272
rect 12034 19216 12714 19272
rect 12770 19216 12775 19272
rect 11973 19214 12775 19216
rect 19014 19274 19074 19350
rect 27286 19348 27292 19412
rect 27356 19410 27403 19412
rect 30925 19410 30991 19413
rect 33869 19410 33935 19413
rect 27356 19408 27448 19410
rect 27398 19352 27448 19408
rect 27356 19350 27448 19352
rect 30925 19408 33935 19410
rect 30925 19352 30930 19408
rect 30986 19352 33874 19408
rect 33930 19352 33935 19408
rect 30925 19350 33935 19352
rect 27356 19348 27403 19350
rect 27337 19347 27403 19348
rect 30925 19347 30991 19350
rect 33869 19347 33935 19350
rect 19374 19274 19380 19276
rect 19014 19214 19380 19274
rect 11973 19211 12039 19214
rect 12709 19211 12775 19214
rect 19374 19212 19380 19214
rect 19444 19212 19450 19276
rect 19517 19274 19583 19277
rect 20161 19274 20227 19277
rect 19517 19272 20227 19274
rect 19517 19216 19522 19272
rect 19578 19216 20166 19272
rect 20222 19216 20227 19272
rect 19517 19214 20227 19216
rect 19517 19211 19583 19214
rect 20161 19211 20227 19214
rect 21173 19274 21239 19277
rect 24853 19274 24919 19277
rect 21173 19272 24919 19274
rect 21173 19216 21178 19272
rect 21234 19216 24858 19272
rect 24914 19216 24919 19272
rect 21173 19214 24919 19216
rect 21173 19211 21239 19214
rect 24853 19211 24919 19214
rect 27797 19274 27863 19277
rect 30782 19274 30788 19276
rect 27797 19272 30788 19274
rect 27797 19216 27802 19272
rect 27858 19216 30788 19272
rect 27797 19214 30788 19216
rect 27797 19211 27863 19214
rect 30782 19212 30788 19214
rect 30852 19274 30858 19276
rect 32213 19274 32279 19277
rect 30852 19272 32279 19274
rect 30852 19216 32218 19272
rect 32274 19216 32279 19272
rect 30852 19214 32279 19216
rect 30852 19212 30858 19214
rect 32213 19211 32279 19214
rect 5441 19138 5507 19141
rect 14406 19138 14412 19140
rect 5441 19136 14412 19138
rect 5441 19080 5446 19136
rect 5502 19080 14412 19136
rect 5441 19078 14412 19080
rect 5441 19075 5507 19078
rect 14406 19076 14412 19078
rect 14476 19138 14482 19140
rect 26969 19138 27035 19141
rect 29085 19138 29151 19141
rect 14476 19136 29151 19138
rect 14476 19080 26974 19136
rect 27030 19080 29090 19136
rect 29146 19080 29151 19136
rect 14476 19078 29151 19080
rect 14476 19076 14482 19078
rect 26969 19075 27035 19078
rect 29085 19075 29151 19078
rect 31477 19138 31543 19141
rect 32121 19138 32187 19141
rect 31477 19136 32187 19138
rect 31477 19080 31482 19136
rect 31538 19080 32126 19136
rect 32182 19080 32187 19136
rect 31477 19078 32187 19080
rect 31477 19075 31543 19078
rect 32121 19075 32187 19078
rect 44081 19138 44147 19141
rect 45200 19138 46000 19168
rect 44081 19136 46000 19138
rect 44081 19080 44086 19136
rect 44142 19080 46000 19136
rect 44081 19078 46000 19080
rect 44081 19075 44147 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 45200 19048 46000 19078
rect 34930 19007 35246 19008
rect 9857 19002 9923 19005
rect 12893 19002 12959 19005
rect 9857 19000 12959 19002
rect 9857 18944 9862 19000
rect 9918 18944 12898 19000
rect 12954 18944 12959 19000
rect 9857 18942 12959 18944
rect 9857 18939 9923 18942
rect 12893 18939 12959 18942
rect 19558 18940 19564 19004
rect 19628 19002 19634 19004
rect 20161 19002 20227 19005
rect 22277 19002 22343 19005
rect 19628 19000 22343 19002
rect 19628 18944 20166 19000
rect 20222 18944 22282 19000
rect 22338 18944 22343 19000
rect 19628 18942 22343 18944
rect 19628 18940 19634 18942
rect 20161 18939 20227 18942
rect 22277 18939 22343 18942
rect 22461 19002 22527 19005
rect 28809 19002 28875 19005
rect 22461 19000 28875 19002
rect 22461 18944 22466 19000
rect 22522 18944 28814 19000
rect 28870 18944 28875 19000
rect 22461 18942 28875 18944
rect 22461 18939 22527 18942
rect 28809 18939 28875 18942
rect 8661 18866 8727 18869
rect 9029 18866 9095 18869
rect 11697 18866 11763 18869
rect 17125 18866 17191 18869
rect 8661 18864 11763 18866
rect 8661 18808 8666 18864
rect 8722 18808 9034 18864
rect 9090 18808 11702 18864
rect 11758 18808 11763 18864
rect 8661 18806 11763 18808
rect 8661 18803 8727 18806
rect 9029 18803 9095 18806
rect 11697 18803 11763 18806
rect 12390 18864 17191 18866
rect 12390 18808 17130 18864
rect 17186 18808 17191 18864
rect 12390 18806 17191 18808
rect 7097 18730 7163 18733
rect 7649 18730 7715 18733
rect 12390 18730 12450 18806
rect 17125 18803 17191 18806
rect 17493 18866 17559 18869
rect 31201 18866 31267 18869
rect 17493 18864 31267 18866
rect 17493 18808 17498 18864
rect 17554 18808 31206 18864
rect 31262 18808 31267 18864
rect 17493 18806 31267 18808
rect 17493 18803 17559 18806
rect 31201 18803 31267 18806
rect 7097 18728 12450 18730
rect 7097 18672 7102 18728
rect 7158 18672 7654 18728
rect 7710 18672 12450 18728
rect 7097 18670 12450 18672
rect 7097 18667 7163 18670
rect 7649 18667 7715 18670
rect 15694 18668 15700 18732
rect 15764 18730 15770 18732
rect 22185 18730 22251 18733
rect 15764 18728 22251 18730
rect 15764 18672 22190 18728
rect 22246 18672 22251 18728
rect 15764 18670 22251 18672
rect 15764 18668 15770 18670
rect 22185 18667 22251 18670
rect 25405 18730 25471 18733
rect 36905 18730 36971 18733
rect 25405 18728 36971 18730
rect 25405 18672 25410 18728
rect 25466 18672 36910 18728
rect 36966 18672 36971 18728
rect 25405 18670 36971 18672
rect 25405 18667 25471 18670
rect 36905 18667 36971 18670
rect 7005 18594 7071 18597
rect 17033 18594 17099 18597
rect 28758 18594 28764 18596
rect 7005 18592 28764 18594
rect 7005 18536 7010 18592
rect 7066 18536 17038 18592
rect 17094 18536 28764 18592
rect 7005 18534 28764 18536
rect 7005 18531 7071 18534
rect 17033 18531 17099 18534
rect 28758 18532 28764 18534
rect 28828 18594 28834 18596
rect 29269 18594 29335 18597
rect 28828 18592 29335 18594
rect 28828 18536 29274 18592
rect 29330 18536 29335 18592
rect 28828 18534 29335 18536
rect 28828 18532 28834 18534
rect 29269 18531 29335 18534
rect 31661 18594 31727 18597
rect 31937 18594 32003 18597
rect 31661 18592 32003 18594
rect 31661 18536 31666 18592
rect 31722 18536 31942 18592
rect 31998 18536 32003 18592
rect 31661 18534 32003 18536
rect 31661 18531 31727 18534
rect 31937 18531 32003 18534
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 4613 18458 4679 18461
rect 7925 18458 7991 18461
rect 8937 18458 9003 18461
rect 4613 18456 4722 18458
rect 4613 18400 4618 18456
rect 4674 18400 4722 18456
rect 4613 18395 4722 18400
rect 7925 18456 9003 18458
rect 7925 18400 7930 18456
rect 7986 18400 8942 18456
rect 8998 18400 9003 18456
rect 7925 18398 9003 18400
rect 7925 18395 7991 18398
rect 8937 18395 9003 18398
rect 9213 18458 9279 18461
rect 19374 18458 19380 18460
rect 9213 18456 19380 18458
rect 9213 18400 9218 18456
rect 9274 18400 19380 18456
rect 9213 18398 19380 18400
rect 9213 18395 9279 18398
rect 19374 18396 19380 18398
rect 19444 18458 19450 18460
rect 19793 18458 19859 18461
rect 19444 18456 19859 18458
rect 19444 18400 19798 18456
rect 19854 18400 19859 18456
rect 19444 18398 19859 18400
rect 19444 18396 19450 18398
rect 19793 18395 19859 18398
rect 20713 18458 20779 18461
rect 22461 18458 22527 18461
rect 20713 18456 22527 18458
rect 20713 18400 20718 18456
rect 20774 18400 22466 18456
rect 22522 18400 22527 18456
rect 20713 18398 22527 18400
rect 20713 18395 20779 18398
rect 22461 18395 22527 18398
rect 22829 18458 22895 18461
rect 25405 18458 25471 18461
rect 22829 18456 25471 18458
rect 22829 18400 22834 18456
rect 22890 18400 25410 18456
rect 25466 18400 25471 18456
rect 22829 18398 25471 18400
rect 22829 18395 22895 18398
rect 25405 18395 25471 18398
rect 26918 18396 26924 18460
rect 26988 18458 26994 18460
rect 27061 18458 27127 18461
rect 26988 18456 27127 18458
rect 26988 18400 27066 18456
rect 27122 18400 27127 18456
rect 26988 18398 27127 18400
rect 26988 18396 26994 18398
rect 27061 18395 27127 18398
rect 31017 18458 31083 18461
rect 34237 18458 34303 18461
rect 31017 18456 34303 18458
rect 31017 18400 31022 18456
rect 31078 18400 34242 18456
rect 34298 18400 34303 18456
rect 31017 18398 34303 18400
rect 31017 18395 31083 18398
rect 34237 18395 34303 18398
rect 44449 18458 44515 18461
rect 45200 18458 46000 18488
rect 44449 18456 46000 18458
rect 44449 18400 44454 18456
rect 44510 18400 46000 18456
rect 44449 18398 46000 18400
rect 44449 18395 44515 18398
rect 4662 18322 4722 18395
rect 45200 18368 46000 18398
rect 4889 18322 4955 18325
rect 4662 18320 4955 18322
rect 4662 18264 4894 18320
rect 4950 18264 4955 18320
rect 4662 18262 4955 18264
rect 4889 18259 4955 18262
rect 9949 18324 10015 18325
rect 10685 18324 10751 18325
rect 9949 18320 9996 18324
rect 10060 18322 10066 18324
rect 10685 18322 10732 18324
rect 9949 18264 9954 18320
rect 9949 18260 9996 18264
rect 10060 18262 10106 18322
rect 10640 18320 10732 18322
rect 10640 18264 10690 18320
rect 10640 18262 10732 18264
rect 10060 18260 10066 18262
rect 10685 18260 10732 18262
rect 10796 18260 10802 18324
rect 11697 18322 11763 18325
rect 14917 18322 14983 18325
rect 17493 18322 17559 18325
rect 11697 18320 17559 18322
rect 11697 18264 11702 18320
rect 11758 18264 14922 18320
rect 14978 18264 17498 18320
rect 17554 18264 17559 18320
rect 11697 18262 17559 18264
rect 9949 18259 10015 18260
rect 10685 18259 10751 18260
rect 11697 18259 11763 18262
rect 14917 18259 14983 18262
rect 17493 18259 17559 18262
rect 19609 18322 19675 18325
rect 19742 18322 19748 18324
rect 19609 18320 19748 18322
rect 19609 18264 19614 18320
rect 19670 18264 19748 18320
rect 19609 18262 19748 18264
rect 19609 18259 19675 18262
rect 19742 18260 19748 18262
rect 19812 18260 19818 18324
rect 21081 18322 21147 18325
rect 34697 18322 34763 18325
rect 35341 18322 35407 18325
rect 21081 18320 35407 18322
rect 21081 18264 21086 18320
rect 21142 18264 34702 18320
rect 34758 18264 35346 18320
rect 35402 18264 35407 18320
rect 21081 18262 35407 18264
rect 21081 18259 21147 18262
rect 34697 18259 34763 18262
rect 35341 18259 35407 18262
rect 8477 18186 8543 18189
rect 18597 18186 18663 18189
rect 22502 18186 22508 18188
rect 8477 18184 22508 18186
rect 8477 18128 8482 18184
rect 8538 18128 18602 18184
rect 18658 18128 22508 18184
rect 8477 18126 22508 18128
rect 8477 18123 8543 18126
rect 18597 18123 18663 18126
rect 22502 18124 22508 18126
rect 22572 18124 22578 18188
rect 22645 18186 22711 18189
rect 37457 18186 37523 18189
rect 22645 18184 37523 18186
rect 22645 18128 22650 18184
rect 22706 18128 37462 18184
rect 37518 18128 37523 18184
rect 22645 18126 37523 18128
rect 8845 18050 8911 18053
rect 15101 18050 15167 18053
rect 18045 18050 18111 18053
rect 8845 18048 18111 18050
rect 8845 17992 8850 18048
rect 8906 17992 15106 18048
rect 15162 17992 18050 18048
rect 18106 17992 18111 18048
rect 8845 17990 18111 17992
rect 8845 17987 8911 17990
rect 15101 17987 15167 17990
rect 18045 17987 18111 17990
rect 19793 18050 19859 18053
rect 19926 18050 19932 18052
rect 19793 18048 19932 18050
rect 19793 17992 19798 18048
rect 19854 17992 19932 18048
rect 19793 17990 19932 17992
rect 19793 17987 19859 17990
rect 19926 17988 19932 17990
rect 19996 18050 20002 18052
rect 22510 18050 22570 18124
rect 22645 18123 22711 18126
rect 37457 18123 37523 18126
rect 23381 18050 23447 18053
rect 19996 17990 22386 18050
rect 22510 18048 23447 18050
rect 22510 17992 23386 18048
rect 23442 17992 23447 18048
rect 22510 17990 23447 17992
rect 19996 17988 20002 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 9949 17914 10015 17917
rect 14038 17914 14044 17916
rect 9949 17912 14044 17914
rect 9949 17856 9954 17912
rect 10010 17856 14044 17912
rect 9949 17854 14044 17856
rect 9949 17851 10015 17854
rect 14038 17852 14044 17854
rect 14108 17914 14114 17916
rect 22185 17914 22251 17917
rect 14108 17912 22251 17914
rect 14108 17856 22190 17912
rect 22246 17856 22251 17912
rect 14108 17854 22251 17856
rect 22326 17914 22386 17990
rect 23381 17987 23447 17990
rect 25405 18050 25471 18053
rect 27797 18050 27863 18053
rect 25405 18048 27863 18050
rect 25405 17992 25410 18048
rect 25466 17992 27802 18048
rect 27858 17992 27863 18048
rect 25405 17990 27863 17992
rect 25405 17987 25471 17990
rect 27797 17987 27863 17990
rect 28533 18052 28599 18053
rect 28533 18048 28580 18052
rect 28644 18050 28650 18052
rect 29729 18050 29795 18053
rect 32213 18050 32279 18053
rect 34513 18050 34579 18053
rect 28533 17992 28538 18048
rect 28533 17988 28580 17992
rect 28644 17990 28690 18050
rect 29729 18048 32279 18050
rect 29729 17992 29734 18048
rect 29790 17992 32218 18048
rect 32274 17992 32279 18048
rect 29729 17990 32279 17992
rect 28644 17988 28650 17990
rect 28533 17987 28599 17988
rect 29729 17987 29795 17990
rect 32213 17987 32279 17990
rect 32630 18048 34579 18050
rect 32630 17992 34518 18048
rect 34574 17992 34579 18048
rect 32630 17990 34579 17992
rect 32630 17917 32690 17990
rect 34513 17987 34579 17990
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 24025 17914 24091 17917
rect 22326 17912 24091 17914
rect 22326 17856 24030 17912
rect 24086 17856 24091 17912
rect 22326 17854 24091 17856
rect 14108 17852 14114 17854
rect 22185 17851 22251 17854
rect 24025 17851 24091 17854
rect 26141 17914 26207 17917
rect 27981 17914 28047 17917
rect 26141 17912 28047 17914
rect 26141 17856 26146 17912
rect 26202 17856 27986 17912
rect 28042 17856 28047 17912
rect 26141 17854 28047 17856
rect 26141 17851 26207 17854
rect 27981 17851 28047 17854
rect 29361 17914 29427 17917
rect 31937 17914 32003 17917
rect 29361 17912 32003 17914
rect 29361 17856 29366 17912
rect 29422 17856 31942 17912
rect 31998 17856 32003 17912
rect 29361 17854 32003 17856
rect 29361 17851 29427 17854
rect 31937 17851 32003 17854
rect 32581 17912 32690 17917
rect 32581 17856 32586 17912
rect 32642 17856 32690 17912
rect 32581 17854 32690 17856
rect 32581 17851 32647 17854
rect 6913 17778 6979 17781
rect 7046 17778 7052 17780
rect 6913 17776 7052 17778
rect 6913 17720 6918 17776
rect 6974 17720 7052 17776
rect 6913 17718 7052 17720
rect 6913 17715 6979 17718
rect 7046 17716 7052 17718
rect 7116 17716 7122 17780
rect 7925 17778 7991 17781
rect 8937 17778 9003 17781
rect 10409 17778 10475 17781
rect 7925 17776 10475 17778
rect 7925 17720 7930 17776
rect 7986 17720 8942 17776
rect 8998 17720 10414 17776
rect 10470 17720 10475 17776
rect 7925 17718 10475 17720
rect 7925 17715 7991 17718
rect 8937 17715 9003 17718
rect 10409 17715 10475 17718
rect 10961 17778 11027 17781
rect 12985 17778 13051 17781
rect 10961 17776 13051 17778
rect 10961 17720 10966 17776
rect 11022 17720 12990 17776
rect 13046 17720 13051 17776
rect 10961 17718 13051 17720
rect 10961 17715 11027 17718
rect 12985 17715 13051 17718
rect 13302 17716 13308 17780
rect 13372 17778 13378 17780
rect 13721 17778 13787 17781
rect 26785 17778 26851 17781
rect 28942 17778 28948 17780
rect 13372 17776 28948 17778
rect 13372 17720 13726 17776
rect 13782 17720 26790 17776
rect 26846 17720 28948 17776
rect 13372 17718 28948 17720
rect 13372 17716 13378 17718
rect 13721 17715 13787 17718
rect 26785 17715 26851 17718
rect 28942 17716 28948 17718
rect 29012 17778 29018 17780
rect 29012 17718 31770 17778
rect 29012 17716 29018 17718
rect 10501 17642 10567 17645
rect 12801 17642 12867 17645
rect 10501 17640 12867 17642
rect 10501 17584 10506 17640
rect 10562 17584 12806 17640
rect 12862 17584 12867 17640
rect 10501 17582 12867 17584
rect 10501 17579 10567 17582
rect 12801 17579 12867 17582
rect 15193 17642 15259 17645
rect 23013 17642 23079 17645
rect 29545 17642 29611 17645
rect 15193 17640 22938 17642
rect 15193 17584 15198 17640
rect 15254 17584 22938 17640
rect 15193 17582 22938 17584
rect 15193 17579 15259 17582
rect 6637 17506 6703 17509
rect 15101 17506 15167 17509
rect 22369 17506 22435 17509
rect 22686 17506 22692 17508
rect 6637 17504 22692 17506
rect 6637 17448 6642 17504
rect 6698 17448 15106 17504
rect 15162 17448 22374 17504
rect 22430 17448 22692 17504
rect 6637 17446 22692 17448
rect 6637 17443 6703 17446
rect 15101 17443 15167 17446
rect 22369 17443 22435 17446
rect 22686 17444 22692 17446
rect 22756 17444 22762 17508
rect 22878 17506 22938 17582
rect 23013 17640 29611 17642
rect 23013 17584 23018 17640
rect 23074 17584 29550 17640
rect 29606 17584 29611 17640
rect 23013 17582 29611 17584
rect 31710 17642 31770 17718
rect 32990 17716 32996 17780
rect 33060 17778 33066 17780
rect 33777 17778 33843 17781
rect 33060 17776 33843 17778
rect 33060 17720 33782 17776
rect 33838 17720 33843 17776
rect 33060 17718 33843 17720
rect 33060 17716 33066 17718
rect 33777 17715 33843 17718
rect 35341 17778 35407 17781
rect 38009 17778 38075 17781
rect 35341 17776 38075 17778
rect 35341 17720 35346 17776
rect 35402 17720 38014 17776
rect 38070 17720 38075 17776
rect 35341 17718 38075 17720
rect 35341 17715 35407 17718
rect 38009 17715 38075 17718
rect 44081 17778 44147 17781
rect 45200 17778 46000 17808
rect 44081 17776 46000 17778
rect 44081 17720 44086 17776
rect 44142 17720 46000 17776
rect 44081 17718 46000 17720
rect 44081 17715 44147 17718
rect 45200 17688 46000 17718
rect 38745 17642 38811 17645
rect 31710 17640 38811 17642
rect 31710 17584 38750 17640
rect 38806 17584 38811 17640
rect 31710 17582 38811 17584
rect 23013 17579 23079 17582
rect 29545 17579 29611 17582
rect 38745 17579 38811 17582
rect 30046 17506 30052 17508
rect 22878 17446 30052 17506
rect 30046 17444 30052 17446
rect 30116 17506 30122 17508
rect 32581 17506 32647 17509
rect 30116 17504 32647 17506
rect 30116 17448 32586 17504
rect 32642 17448 32647 17504
rect 30116 17446 32647 17448
rect 30116 17444 30122 17446
rect 32581 17443 32647 17446
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 8109 17370 8175 17373
rect 13261 17370 13327 17373
rect 8109 17368 13327 17370
rect 8109 17312 8114 17368
rect 8170 17312 13266 17368
rect 13322 17312 13327 17368
rect 8109 17310 13327 17312
rect 8109 17307 8175 17310
rect 13261 17307 13327 17310
rect 13537 17370 13603 17373
rect 13670 17370 13676 17372
rect 13537 17368 13676 17370
rect 13537 17312 13542 17368
rect 13598 17312 13676 17368
rect 13537 17310 13676 17312
rect 13537 17307 13603 17310
rect 13670 17308 13676 17310
rect 13740 17370 13746 17372
rect 26969 17370 27035 17373
rect 13740 17368 27035 17370
rect 13740 17312 26974 17368
rect 27030 17312 27035 17368
rect 13740 17310 27035 17312
rect 13740 17308 13746 17310
rect 26969 17307 27035 17310
rect 30189 17370 30255 17373
rect 35065 17370 35131 17373
rect 30189 17368 35131 17370
rect 30189 17312 30194 17368
rect 30250 17312 35070 17368
rect 35126 17312 35131 17368
rect 30189 17310 35131 17312
rect 30189 17307 30255 17310
rect 35065 17307 35131 17310
rect 4981 17234 5047 17237
rect 11053 17234 11119 17237
rect 4981 17232 11119 17234
rect 4981 17176 4986 17232
rect 5042 17176 11058 17232
rect 11114 17176 11119 17232
rect 4981 17174 11119 17176
rect 4981 17171 5047 17174
rect 11053 17171 11119 17174
rect 11329 17234 11395 17237
rect 12525 17234 12591 17237
rect 12985 17234 13051 17237
rect 11329 17232 13051 17234
rect 11329 17176 11334 17232
rect 11390 17176 12530 17232
rect 12586 17176 12990 17232
rect 13046 17176 13051 17232
rect 11329 17174 13051 17176
rect 11329 17171 11395 17174
rect 12525 17171 12591 17174
rect 12985 17171 13051 17174
rect 18873 17234 18939 17237
rect 19149 17234 19215 17237
rect 18873 17232 19215 17234
rect 18873 17176 18878 17232
rect 18934 17176 19154 17232
rect 19210 17176 19215 17232
rect 18873 17174 19215 17176
rect 18873 17171 18939 17174
rect 19149 17171 19215 17174
rect 25262 17172 25268 17236
rect 25332 17234 25338 17236
rect 27521 17234 27587 17237
rect 25332 17232 27587 17234
rect 25332 17176 27526 17232
rect 27582 17176 27587 17232
rect 25332 17174 27587 17176
rect 25332 17172 25338 17174
rect 27521 17171 27587 17174
rect 28073 17234 28139 17237
rect 28349 17234 28415 17237
rect 35341 17234 35407 17237
rect 36629 17234 36695 17237
rect 28073 17232 36695 17234
rect 28073 17176 28078 17232
rect 28134 17176 28354 17232
rect 28410 17176 35346 17232
rect 35402 17176 36634 17232
rect 36690 17176 36695 17232
rect 28073 17174 36695 17176
rect 28073 17171 28139 17174
rect 28349 17171 28415 17174
rect 35341 17171 35407 17174
rect 36629 17171 36695 17174
rect 10409 17098 10475 17101
rect 19333 17098 19399 17101
rect 31886 17098 31892 17100
rect 10409 17096 31892 17098
rect 10409 17040 10414 17096
rect 10470 17040 19338 17096
rect 19394 17040 31892 17096
rect 10409 17038 31892 17040
rect 10409 17035 10475 17038
rect 19333 17035 19399 17038
rect 31886 17036 31892 17038
rect 31956 17098 31962 17100
rect 33317 17098 33383 17101
rect 31956 17096 33383 17098
rect 31956 17040 33322 17096
rect 33378 17040 33383 17096
rect 31956 17038 33383 17040
rect 31956 17036 31962 17038
rect 33317 17035 33383 17038
rect 34145 17098 34211 17101
rect 36537 17098 36603 17101
rect 34145 17096 36603 17098
rect 34145 17040 34150 17096
rect 34206 17040 36542 17096
rect 36598 17040 36603 17096
rect 34145 17038 36603 17040
rect 34145 17035 34211 17038
rect 36537 17035 36603 17038
rect 44449 17098 44515 17101
rect 45200 17098 46000 17128
rect 44449 17096 46000 17098
rect 44449 17040 44454 17096
rect 44510 17040 46000 17096
rect 44449 17038 46000 17040
rect 44449 17035 44515 17038
rect 45200 17008 46000 17038
rect 10961 16962 11027 16965
rect 18873 16962 18939 16965
rect 24761 16964 24827 16965
rect 10961 16960 18939 16962
rect 10961 16904 10966 16960
rect 11022 16904 18878 16960
rect 18934 16904 18939 16960
rect 10961 16902 18939 16904
rect 10961 16899 11027 16902
rect 18873 16899 18939 16902
rect 24710 16900 24716 16964
rect 24780 16962 24827 16964
rect 24780 16960 31770 16962
rect 24822 16904 31770 16960
rect 24780 16902 31770 16904
rect 24780 16900 24827 16902
rect 24761 16899 24827 16900
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 11053 16826 11119 16829
rect 13813 16826 13879 16829
rect 14641 16826 14707 16829
rect 11053 16824 14707 16826
rect 11053 16768 11058 16824
rect 11114 16768 13818 16824
rect 13874 16768 14646 16824
rect 14702 16768 14707 16824
rect 11053 16766 14707 16768
rect 11053 16763 11119 16766
rect 13813 16763 13879 16766
rect 14641 16763 14707 16766
rect 17401 16826 17467 16829
rect 17534 16826 17540 16828
rect 17401 16824 17540 16826
rect 17401 16768 17406 16824
rect 17462 16768 17540 16824
rect 17401 16766 17540 16768
rect 17401 16763 17467 16766
rect 17534 16764 17540 16766
rect 17604 16764 17610 16828
rect 24025 16826 24091 16829
rect 27889 16826 27955 16829
rect 24025 16824 27955 16826
rect 24025 16768 24030 16824
rect 24086 16768 27894 16824
rect 27950 16768 27955 16824
rect 24025 16766 27955 16768
rect 24025 16763 24091 16766
rect 27889 16763 27955 16766
rect 3693 16690 3759 16693
rect 4889 16690 4955 16693
rect 7281 16690 7347 16693
rect 3693 16688 7347 16690
rect 3693 16632 3698 16688
rect 3754 16632 4894 16688
rect 4950 16632 7286 16688
rect 7342 16632 7347 16688
rect 3693 16630 7347 16632
rect 3693 16627 3759 16630
rect 4889 16627 4955 16630
rect 7281 16627 7347 16630
rect 8569 16690 8635 16693
rect 15009 16690 15075 16693
rect 8569 16688 15075 16690
rect 8569 16632 8574 16688
rect 8630 16632 15014 16688
rect 15070 16632 15075 16688
rect 8569 16630 15075 16632
rect 31710 16690 31770 16902
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 32397 16826 32463 16829
rect 33542 16826 33548 16828
rect 32397 16824 33548 16826
rect 32397 16768 32402 16824
rect 32458 16768 33548 16824
rect 32397 16766 33548 16768
rect 32397 16763 32463 16766
rect 33542 16764 33548 16766
rect 33612 16764 33618 16828
rect 39021 16690 39087 16693
rect 31710 16688 39087 16690
rect 31710 16632 39026 16688
rect 39082 16632 39087 16688
rect 31710 16630 39087 16632
rect 8569 16627 8635 16630
rect 15009 16627 15075 16630
rect 39021 16627 39087 16630
rect 841 16554 907 16557
rect 798 16552 907 16554
rect 798 16496 846 16552
rect 902 16496 907 16552
rect 798 16491 907 16496
rect 7557 16554 7623 16557
rect 16389 16554 16455 16557
rect 18321 16554 18387 16557
rect 7557 16552 18387 16554
rect 7557 16496 7562 16552
rect 7618 16496 16394 16552
rect 16450 16496 18326 16552
rect 18382 16496 18387 16552
rect 7557 16494 18387 16496
rect 7557 16491 7623 16494
rect 16389 16491 16455 16494
rect 18321 16491 18387 16494
rect 25814 16492 25820 16556
rect 25884 16554 25890 16556
rect 27337 16554 27403 16557
rect 25884 16552 27403 16554
rect 25884 16496 27342 16552
rect 27398 16496 27403 16552
rect 25884 16494 27403 16496
rect 25884 16492 25890 16494
rect 27337 16491 27403 16494
rect 28901 16554 28967 16557
rect 37089 16554 37155 16557
rect 28901 16552 37155 16554
rect 28901 16496 28906 16552
rect 28962 16496 37094 16552
rect 37150 16496 37155 16552
rect 28901 16494 37155 16496
rect 28901 16491 28967 16494
rect 37089 16491 37155 16494
rect 798 16448 858 16491
rect 0 16358 858 16448
rect 9397 16418 9463 16421
rect 9673 16418 9739 16421
rect 9397 16416 9739 16418
rect 9397 16360 9402 16416
rect 9458 16360 9678 16416
rect 9734 16360 9739 16416
rect 9397 16358 9739 16360
rect 0 16328 800 16358
rect 9397 16355 9463 16358
rect 9673 16355 9739 16358
rect 10593 16418 10659 16421
rect 10726 16418 10732 16420
rect 10593 16416 10732 16418
rect 10593 16360 10598 16416
rect 10654 16360 10732 16416
rect 10593 16358 10732 16360
rect 10593 16355 10659 16358
rect 10726 16356 10732 16358
rect 10796 16356 10802 16420
rect 11513 16418 11579 16421
rect 11973 16418 12039 16421
rect 13905 16418 13971 16421
rect 11513 16416 13971 16418
rect 11513 16360 11518 16416
rect 11574 16360 11978 16416
rect 12034 16360 13910 16416
rect 13966 16360 13971 16416
rect 11513 16358 13971 16360
rect 11513 16355 11579 16358
rect 11973 16355 12039 16358
rect 13905 16355 13971 16358
rect 16021 16418 16087 16421
rect 18689 16418 18755 16421
rect 16021 16416 18755 16418
rect 16021 16360 16026 16416
rect 16082 16360 18694 16416
rect 18750 16360 18755 16416
rect 16021 16358 18755 16360
rect 16021 16355 16087 16358
rect 18689 16355 18755 16358
rect 22870 16356 22876 16420
rect 22940 16418 22946 16420
rect 23013 16418 23079 16421
rect 22940 16416 23079 16418
rect 22940 16360 23018 16416
rect 23074 16360 23079 16416
rect 22940 16358 23079 16360
rect 22940 16356 22946 16358
rect 23013 16355 23079 16358
rect 27102 16356 27108 16420
rect 27172 16418 27178 16420
rect 29637 16418 29703 16421
rect 27172 16416 29703 16418
rect 27172 16360 29642 16416
rect 29698 16360 29703 16416
rect 27172 16358 29703 16360
rect 27172 16356 27178 16358
rect 29637 16355 29703 16358
rect 31385 16418 31451 16421
rect 33409 16418 33475 16421
rect 31385 16416 33475 16418
rect 31385 16360 31390 16416
rect 31446 16360 33414 16416
rect 33470 16360 33475 16416
rect 31385 16358 33475 16360
rect 31385 16355 31451 16358
rect 33409 16355 33475 16358
rect 44449 16418 44515 16421
rect 45200 16418 46000 16448
rect 44449 16416 46000 16418
rect 44449 16360 44454 16416
rect 44510 16360 46000 16416
rect 44449 16358 46000 16360
rect 44449 16355 44515 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 45200 16328 46000 16358
rect 35590 16287 35906 16288
rect 10685 16282 10751 16285
rect 15193 16282 15259 16285
rect 26877 16282 26943 16285
rect 10685 16280 15259 16282
rect 10685 16224 10690 16280
rect 10746 16224 15198 16280
rect 15254 16224 15259 16280
rect 10685 16222 15259 16224
rect 10685 16219 10751 16222
rect 15193 16219 15259 16222
rect 20486 16280 26943 16282
rect 20486 16224 26882 16280
rect 26938 16224 26943 16280
rect 20486 16222 26943 16224
rect 8753 16146 8819 16149
rect 8886 16146 8892 16148
rect 8753 16144 8892 16146
rect 8753 16088 8758 16144
rect 8814 16088 8892 16144
rect 8753 16086 8892 16088
rect 8753 16083 8819 16086
rect 8886 16084 8892 16086
rect 8956 16084 8962 16148
rect 17309 16146 17375 16149
rect 20345 16146 20411 16149
rect 20486 16146 20546 16222
rect 26877 16219 26943 16222
rect 27337 16282 27403 16285
rect 32397 16282 32463 16285
rect 27337 16280 32463 16282
rect 27337 16224 27342 16280
rect 27398 16224 32402 16280
rect 32458 16224 32463 16280
rect 27337 16222 32463 16224
rect 27337 16219 27403 16222
rect 32397 16219 32463 16222
rect 32806 16220 32812 16284
rect 32876 16282 32882 16284
rect 33225 16282 33291 16285
rect 32876 16280 33291 16282
rect 32876 16224 33230 16280
rect 33286 16224 33291 16280
rect 32876 16222 33291 16224
rect 32876 16220 32882 16222
rect 33225 16219 33291 16222
rect 32581 16146 32647 16149
rect 9078 16144 20546 16146
rect 9078 16088 17314 16144
rect 17370 16088 20350 16144
rect 20406 16088 20546 16144
rect 9078 16086 20546 16088
rect 20624 16144 32647 16146
rect 20624 16088 32586 16144
rect 32642 16088 32647 16144
rect 20624 16086 32647 16088
rect 6637 16010 6703 16013
rect 8150 16010 8156 16012
rect 6637 16008 8156 16010
rect 6637 15952 6642 16008
rect 6698 15952 8156 16008
rect 6637 15950 8156 15952
rect 6637 15947 6703 15950
rect 8150 15948 8156 15950
rect 8220 16010 8226 16012
rect 9078 16010 9138 16086
rect 17309 16083 17375 16086
rect 20345 16083 20411 16086
rect 8220 15950 9138 16010
rect 8220 15948 8226 15950
rect 9806 15948 9812 16012
rect 9876 16010 9882 16012
rect 9949 16010 10015 16013
rect 9876 16008 10015 16010
rect 9876 15952 9954 16008
rect 10010 15952 10015 16008
rect 9876 15950 10015 15952
rect 9876 15948 9882 15950
rect 9949 15947 10015 15950
rect 10225 16010 10291 16013
rect 14733 16010 14799 16013
rect 16205 16012 16271 16013
rect 16205 16010 16252 16012
rect 10225 16008 14799 16010
rect 10225 15952 10230 16008
rect 10286 15952 14738 16008
rect 14794 15952 14799 16008
rect 10225 15950 14799 15952
rect 16160 16008 16252 16010
rect 16160 15952 16210 16008
rect 16160 15950 16252 15952
rect 10225 15947 10291 15950
rect 14733 15947 14799 15950
rect 16205 15948 16252 15950
rect 16316 15948 16322 16012
rect 19006 15948 19012 16012
rect 19076 16010 19082 16012
rect 20624 16010 20684 16086
rect 32581 16083 32647 16086
rect 32949 16146 33015 16149
rect 36629 16146 36695 16149
rect 32949 16144 36695 16146
rect 32949 16088 32954 16144
rect 33010 16088 36634 16144
rect 36690 16088 36695 16144
rect 32949 16086 36695 16088
rect 32949 16083 33015 16086
rect 36629 16083 36695 16086
rect 22093 16010 22159 16013
rect 19076 15950 20684 16010
rect 20854 16008 22159 16010
rect 20854 15952 22098 16008
rect 22154 15952 22159 16008
rect 20854 15950 22159 15952
rect 19076 15948 19082 15950
rect 16205 15947 16271 15948
rect 841 15874 907 15877
rect 798 15872 907 15874
rect 798 15816 846 15872
rect 902 15816 907 15872
rect 798 15811 907 15816
rect 10041 15874 10107 15877
rect 12893 15874 12959 15877
rect 10041 15872 12959 15874
rect 10041 15816 10046 15872
rect 10102 15816 12898 15872
rect 12954 15816 12959 15872
rect 10041 15814 12959 15816
rect 10041 15811 10107 15814
rect 12893 15811 12959 15814
rect 13261 15874 13327 15877
rect 13486 15874 13492 15876
rect 13261 15872 13492 15874
rect 13261 15816 13266 15872
rect 13322 15816 13492 15872
rect 13261 15814 13492 15816
rect 13261 15811 13327 15814
rect 13486 15812 13492 15814
rect 13556 15812 13562 15876
rect 18413 15874 18479 15877
rect 20854 15874 20914 15950
rect 22093 15947 22159 15950
rect 22277 16012 22343 16013
rect 22277 16008 22324 16012
rect 22388 16010 22394 16012
rect 26417 16010 26483 16013
rect 29545 16010 29611 16013
rect 29729 16012 29795 16013
rect 22277 15952 22282 16008
rect 22277 15948 22324 15952
rect 22388 15950 22434 16010
rect 26417 16008 29611 16010
rect 26417 15952 26422 16008
rect 26478 15952 29550 16008
rect 29606 15952 29611 16008
rect 26417 15950 29611 15952
rect 22388 15948 22394 15950
rect 22277 15947 22343 15948
rect 26417 15947 26483 15950
rect 29545 15947 29611 15950
rect 29678 15948 29684 16012
rect 29748 16010 29795 16012
rect 29748 16008 29840 16010
rect 29790 15952 29840 16008
rect 29748 15950 29840 15952
rect 29748 15948 29795 15950
rect 29729 15947 29795 15948
rect 18413 15872 20914 15874
rect 18413 15816 18418 15872
rect 18474 15816 20914 15872
rect 18413 15814 20914 15816
rect 20989 15874 21055 15877
rect 21357 15874 21423 15877
rect 22461 15874 22527 15877
rect 20989 15872 22527 15874
rect 20989 15816 20994 15872
rect 21050 15816 21362 15872
rect 21418 15816 22466 15872
rect 22522 15816 22527 15872
rect 20989 15814 22527 15816
rect 18413 15811 18479 15814
rect 20989 15811 21055 15814
rect 21357 15811 21423 15814
rect 22461 15811 22527 15814
rect 22645 15874 22711 15877
rect 26693 15874 26759 15877
rect 22645 15872 26759 15874
rect 22645 15816 22650 15872
rect 22706 15816 26698 15872
rect 26754 15816 26759 15872
rect 22645 15814 26759 15816
rect 22645 15811 22711 15814
rect 26693 15811 26759 15814
rect 26877 15874 26943 15877
rect 32990 15874 32996 15876
rect 26877 15872 32996 15874
rect 26877 15816 26882 15872
rect 26938 15816 32996 15872
rect 26877 15814 32996 15816
rect 26877 15811 26943 15814
rect 32990 15812 32996 15814
rect 33060 15812 33066 15876
rect 798 15768 858 15811
rect 0 15678 858 15768
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 9029 15738 9095 15741
rect 10777 15738 10843 15741
rect 9029 15736 10843 15738
rect 9029 15680 9034 15736
rect 9090 15680 10782 15736
rect 10838 15680 10843 15736
rect 9029 15678 10843 15680
rect 0 15648 800 15678
rect 9029 15675 9095 15678
rect 10777 15675 10843 15678
rect 10961 15738 11027 15741
rect 15510 15738 15516 15740
rect 10961 15736 15516 15738
rect 10961 15680 10966 15736
rect 11022 15680 15516 15736
rect 10961 15678 15516 15680
rect 10961 15675 11027 15678
rect 15510 15676 15516 15678
rect 15580 15676 15586 15740
rect 18137 15738 18203 15741
rect 19241 15738 19307 15741
rect 32857 15738 32923 15741
rect 18137 15736 32923 15738
rect 18137 15680 18142 15736
rect 18198 15680 19246 15736
rect 19302 15680 32862 15736
rect 32918 15680 32923 15736
rect 18137 15678 32923 15680
rect 18137 15675 18203 15678
rect 19241 15675 19307 15678
rect 32857 15675 32923 15678
rect 44449 15738 44515 15741
rect 45200 15738 46000 15768
rect 44449 15736 46000 15738
rect 44449 15680 44454 15736
rect 44510 15680 46000 15736
rect 44449 15678 46000 15680
rect 44449 15675 44515 15678
rect 45200 15648 46000 15678
rect 5533 15602 5599 15605
rect 18505 15602 18571 15605
rect 18873 15602 18939 15605
rect 5533 15600 18939 15602
rect 5533 15544 5538 15600
rect 5594 15544 18510 15600
rect 18566 15544 18878 15600
rect 18934 15544 18939 15600
rect 5533 15542 18939 15544
rect 5533 15539 5599 15542
rect 18505 15539 18571 15542
rect 18873 15539 18939 15542
rect 22093 15602 22159 15605
rect 26417 15602 26483 15605
rect 22093 15600 26483 15602
rect 22093 15544 22098 15600
rect 22154 15544 26422 15600
rect 26478 15544 26483 15600
rect 22093 15542 26483 15544
rect 22093 15539 22159 15542
rect 26417 15539 26483 15542
rect 29310 15540 29316 15604
rect 29380 15602 29386 15604
rect 29545 15602 29611 15605
rect 29380 15600 29611 15602
rect 29380 15544 29550 15600
rect 29606 15544 29611 15600
rect 29380 15542 29611 15544
rect 29380 15540 29386 15542
rect 29545 15539 29611 15542
rect 6729 15466 6795 15469
rect 7373 15466 7439 15469
rect 6729 15464 7439 15466
rect 6729 15408 6734 15464
rect 6790 15408 7378 15464
rect 7434 15408 7439 15464
rect 6729 15406 7439 15408
rect 6729 15403 6795 15406
rect 7373 15403 7439 15406
rect 10133 15466 10199 15469
rect 12709 15466 12775 15469
rect 10133 15464 12775 15466
rect 10133 15408 10138 15464
rect 10194 15408 12714 15464
rect 12770 15408 12775 15464
rect 10133 15406 12775 15408
rect 10133 15403 10199 15406
rect 12709 15403 12775 15406
rect 12985 15466 13051 15469
rect 18781 15466 18847 15469
rect 20989 15466 21055 15469
rect 12985 15464 21055 15466
rect 12985 15408 12990 15464
rect 13046 15408 18786 15464
rect 18842 15408 20994 15464
rect 21050 15408 21055 15464
rect 12985 15406 21055 15408
rect 12985 15403 13051 15406
rect 18781 15403 18847 15406
rect 20989 15403 21055 15406
rect 22277 15466 22343 15469
rect 25589 15466 25655 15469
rect 22277 15464 25655 15466
rect 22277 15408 22282 15464
rect 22338 15408 25594 15464
rect 25650 15408 25655 15464
rect 22277 15406 25655 15408
rect 22277 15403 22343 15406
rect 25589 15403 25655 15406
rect 32857 15466 32923 15469
rect 33593 15466 33659 15469
rect 32857 15464 33659 15466
rect 32857 15408 32862 15464
rect 32918 15408 33598 15464
rect 33654 15408 33659 15464
rect 32857 15406 33659 15408
rect 32857 15403 32923 15406
rect 33593 15403 33659 15406
rect 10777 15330 10843 15333
rect 19977 15330 20043 15333
rect 10777 15328 20043 15330
rect 10777 15272 10782 15328
rect 10838 15272 19982 15328
rect 20038 15272 20043 15328
rect 10777 15270 20043 15272
rect 10777 15267 10843 15270
rect 19977 15267 20043 15270
rect 22093 15330 22159 15333
rect 23381 15330 23447 15333
rect 26693 15330 26759 15333
rect 22093 15328 26759 15330
rect 22093 15272 22098 15328
rect 22154 15272 23386 15328
rect 23442 15272 26698 15328
rect 26754 15272 26759 15328
rect 22093 15270 26759 15272
rect 22093 15267 22159 15270
rect 23381 15267 23447 15270
rect 26693 15267 26759 15270
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 11053 15196 11119 15197
rect 11053 15194 11100 15196
rect 11008 15192 11100 15194
rect 11164 15194 11170 15196
rect 12801 15194 12867 15197
rect 16757 15194 16823 15197
rect 11008 15136 11058 15192
rect 11008 15134 11100 15136
rect 11053 15132 11100 15134
rect 11164 15134 12450 15194
rect 11164 15132 11170 15134
rect 11053 15131 11119 15132
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 11145 15058 11211 15061
rect 12157 15058 12223 15061
rect 11145 15056 12223 15058
rect 11145 15000 11150 15056
rect 11206 15000 12162 15056
rect 12218 15000 12223 15056
rect 11145 14998 12223 15000
rect 11145 14995 11211 14998
rect 12157 14995 12223 14998
rect 12390 14922 12450 15134
rect 12801 15192 16823 15194
rect 12801 15136 12806 15192
rect 12862 15136 16762 15192
rect 16818 15136 16823 15192
rect 12801 15134 16823 15136
rect 12801 15131 12867 15134
rect 16757 15131 16823 15134
rect 18045 15194 18111 15197
rect 18873 15194 18939 15197
rect 18045 15192 18939 15194
rect 18045 15136 18050 15192
rect 18106 15136 18878 15192
rect 18934 15136 18939 15192
rect 18045 15134 18939 15136
rect 18045 15131 18111 15134
rect 18873 15131 18939 15134
rect 27337 15194 27403 15197
rect 27470 15194 27476 15196
rect 27337 15192 27476 15194
rect 27337 15136 27342 15192
rect 27398 15136 27476 15192
rect 27337 15134 27476 15136
rect 27337 15131 27403 15134
rect 27470 15132 27476 15134
rect 27540 15132 27546 15196
rect 30833 15194 30899 15197
rect 30966 15194 30972 15196
rect 30833 15192 30972 15194
rect 30833 15136 30838 15192
rect 30894 15136 30972 15192
rect 30833 15134 30972 15136
rect 30833 15131 30899 15134
rect 30966 15132 30972 15134
rect 31036 15132 31042 15196
rect 17350 14996 17356 15060
rect 17420 15058 17426 15060
rect 30598 15058 30604 15060
rect 17420 14998 30604 15058
rect 17420 14996 17426 14998
rect 30598 14996 30604 14998
rect 30668 15058 30674 15060
rect 31017 15058 31083 15061
rect 31569 15058 31635 15061
rect 30668 15056 31635 15058
rect 30668 15000 31022 15056
rect 31078 15000 31574 15056
rect 31630 15000 31635 15056
rect 30668 14998 31635 15000
rect 30668 14996 30674 14998
rect 31017 14995 31083 14998
rect 31569 14995 31635 14998
rect 33685 15058 33751 15061
rect 36118 15058 36124 15060
rect 33685 15056 36124 15058
rect 33685 15000 33690 15056
rect 33746 15000 36124 15056
rect 33685 14998 36124 15000
rect 33685 14995 33751 14998
rect 36118 14996 36124 14998
rect 36188 14996 36194 15060
rect 44081 15058 44147 15061
rect 45200 15058 46000 15088
rect 44081 15056 46000 15058
rect 44081 15000 44086 15056
rect 44142 15000 46000 15056
rect 44081 14998 46000 15000
rect 44081 14995 44147 14998
rect 45200 14968 46000 14998
rect 26325 14922 26391 14925
rect 12390 14920 26391 14922
rect 12390 14864 26330 14920
rect 26386 14864 26391 14920
rect 12390 14862 26391 14864
rect 26325 14859 26391 14862
rect 30649 14922 30715 14925
rect 33501 14922 33567 14925
rect 30649 14920 33567 14922
rect 30649 14864 30654 14920
rect 30710 14864 33506 14920
rect 33562 14864 33567 14920
rect 30649 14862 33567 14864
rect 30649 14859 30715 14862
rect 33501 14859 33567 14862
rect 9121 14786 9187 14789
rect 16205 14786 16271 14789
rect 9121 14784 16271 14786
rect 9121 14728 9126 14784
rect 9182 14728 16210 14784
rect 16266 14728 16271 14784
rect 9121 14726 16271 14728
rect 9121 14723 9187 14726
rect 16205 14723 16271 14726
rect 25405 14786 25471 14789
rect 27797 14786 27863 14789
rect 31569 14788 31635 14789
rect 25405 14784 27863 14786
rect 25405 14728 25410 14784
rect 25466 14728 27802 14784
rect 27858 14728 27863 14784
rect 25405 14726 27863 14728
rect 25405 14723 25471 14726
rect 27797 14723 27863 14726
rect 31518 14724 31524 14788
rect 31588 14786 31635 14788
rect 31588 14784 31680 14786
rect 31630 14728 31680 14784
rect 31588 14726 31680 14728
rect 31588 14724 31635 14726
rect 31569 14723 31635 14724
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 6177 14650 6243 14653
rect 15193 14650 15259 14653
rect 6177 14648 15259 14650
rect 6177 14592 6182 14648
rect 6238 14592 15198 14648
rect 15254 14592 15259 14648
rect 6177 14590 15259 14592
rect 6177 14587 6243 14590
rect 15193 14587 15259 14590
rect 16665 14650 16731 14653
rect 17350 14650 17356 14652
rect 16665 14648 17356 14650
rect 16665 14592 16670 14648
rect 16726 14592 17356 14648
rect 16665 14590 17356 14592
rect 16665 14587 16731 14590
rect 17350 14588 17356 14590
rect 17420 14588 17426 14652
rect 20345 14650 20411 14653
rect 27705 14650 27771 14653
rect 20345 14648 27771 14650
rect 20345 14592 20350 14648
rect 20406 14592 27710 14648
rect 27766 14592 27771 14648
rect 20345 14590 27771 14592
rect 20345 14587 20411 14590
rect 27705 14587 27771 14590
rect 30925 14650 30991 14653
rect 32673 14650 32739 14653
rect 30925 14648 32739 14650
rect 30925 14592 30930 14648
rect 30986 14592 32678 14648
rect 32734 14592 32739 14648
rect 30925 14590 32739 14592
rect 30925 14587 30991 14590
rect 32673 14587 32739 14590
rect 841 14514 907 14517
rect 798 14512 907 14514
rect 798 14456 846 14512
rect 902 14456 907 14512
rect 798 14451 907 14456
rect 13261 14514 13327 14517
rect 22461 14514 22527 14517
rect 13261 14512 22527 14514
rect 13261 14456 13266 14512
rect 13322 14456 22466 14512
rect 22522 14456 22527 14512
rect 13261 14454 22527 14456
rect 13261 14451 13327 14454
rect 22461 14451 22527 14454
rect 24209 14514 24275 14517
rect 37457 14514 37523 14517
rect 24209 14512 37523 14514
rect 24209 14456 24214 14512
rect 24270 14456 37462 14512
rect 37518 14456 37523 14512
rect 24209 14454 37523 14456
rect 24209 14451 24275 14454
rect 37457 14451 37523 14454
rect 798 14408 858 14451
rect 0 14318 858 14408
rect 20529 14378 20595 14381
rect 17910 14376 20595 14378
rect 17910 14320 20534 14376
rect 20590 14320 20595 14376
rect 17910 14318 20595 14320
rect 0 14288 800 14318
rect 9121 14242 9187 14245
rect 17910 14242 17970 14318
rect 20529 14315 20595 14318
rect 22001 14378 22067 14381
rect 34789 14378 34855 14381
rect 22001 14376 34855 14378
rect 22001 14320 22006 14376
rect 22062 14320 34794 14376
rect 34850 14320 34855 14376
rect 22001 14318 34855 14320
rect 22001 14315 22067 14318
rect 34789 14315 34855 14318
rect 44449 14378 44515 14381
rect 45200 14378 46000 14408
rect 44449 14376 46000 14378
rect 44449 14320 44454 14376
rect 44510 14320 46000 14376
rect 44449 14318 46000 14320
rect 44449 14315 44515 14318
rect 45200 14288 46000 14318
rect 9121 14240 17970 14242
rect 9121 14184 9126 14240
rect 9182 14184 17970 14240
rect 9121 14182 17970 14184
rect 9121 14179 9187 14182
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 7925 14106 7991 14109
rect 9673 14106 9739 14109
rect 7925 14104 9739 14106
rect 7925 14048 7930 14104
rect 7986 14048 9678 14104
rect 9734 14048 9739 14104
rect 7925 14046 9739 14048
rect 7925 14043 7991 14046
rect 9673 14043 9739 14046
rect 12433 14106 12499 14109
rect 17401 14106 17467 14109
rect 12433 14104 17467 14106
rect 12433 14048 12438 14104
rect 12494 14048 17406 14104
rect 17462 14048 17467 14104
rect 12433 14046 17467 14048
rect 12433 14043 12499 14046
rect 17401 14043 17467 14046
rect 23105 14106 23171 14109
rect 23974 14106 23980 14108
rect 23105 14104 23980 14106
rect 23105 14048 23110 14104
rect 23166 14048 23980 14104
rect 23105 14046 23980 14048
rect 23105 14043 23171 14046
rect 23974 14044 23980 14046
rect 24044 14044 24050 14108
rect 28073 14106 28139 14109
rect 28206 14106 28212 14108
rect 28073 14104 28212 14106
rect 28073 14048 28078 14104
rect 28134 14048 28212 14104
rect 28073 14046 28212 14048
rect 28073 14043 28139 14046
rect 28206 14044 28212 14046
rect 28276 14044 28282 14108
rect 8845 13970 8911 13973
rect 11973 13970 12039 13973
rect 8845 13968 12039 13970
rect 8845 13912 8850 13968
rect 8906 13912 11978 13968
rect 12034 13912 12039 13968
rect 8845 13910 12039 13912
rect 8845 13907 8911 13910
rect 11973 13907 12039 13910
rect 13077 13970 13143 13973
rect 26509 13970 26575 13973
rect 13077 13968 26575 13970
rect 13077 13912 13082 13968
rect 13138 13912 26514 13968
rect 26570 13912 26575 13968
rect 13077 13910 26575 13912
rect 13077 13907 13143 13910
rect 26509 13907 26575 13910
rect 12065 13834 12131 13837
rect 12198 13834 12204 13836
rect 12065 13832 12204 13834
rect 12065 13776 12070 13832
rect 12126 13776 12204 13832
rect 12065 13774 12204 13776
rect 12065 13771 12131 13774
rect 12198 13772 12204 13774
rect 12268 13834 12274 13836
rect 20161 13834 20227 13837
rect 12268 13832 20227 13834
rect 12268 13776 20166 13832
rect 20222 13776 20227 13832
rect 12268 13774 20227 13776
rect 12268 13772 12274 13774
rect 20161 13771 20227 13774
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 7925 13700 7991 13701
rect 7925 13698 7972 13700
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 7880 13696 7972 13698
rect 7880 13640 7930 13696
rect 7880 13638 7972 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 7925 13636 7972 13638
rect 8036 13636 8042 13700
rect 11789 13698 11855 13701
rect 20345 13698 20411 13701
rect 11789 13696 20411 13698
rect 11789 13640 11794 13696
rect 11850 13640 20350 13696
rect 20406 13640 20411 13696
rect 11789 13638 20411 13640
rect 7925 13635 7991 13636
rect 11789 13635 11855 13638
rect 20345 13635 20411 13638
rect 23841 13698 23907 13701
rect 25446 13698 25452 13700
rect 23841 13696 25452 13698
rect 23841 13640 23846 13696
rect 23902 13640 25452 13696
rect 23841 13638 25452 13640
rect 23841 13635 23907 13638
rect 25446 13636 25452 13638
rect 25516 13698 25522 13700
rect 30925 13698 30991 13701
rect 25516 13696 30991 13698
rect 25516 13640 30930 13696
rect 30986 13640 30991 13696
rect 25516 13638 30991 13640
rect 25516 13636 25522 13638
rect 30925 13635 30991 13638
rect 44081 13698 44147 13701
rect 45200 13698 46000 13728
rect 44081 13696 46000 13698
rect 44081 13640 44086 13696
rect 44142 13640 46000 13696
rect 44081 13638 46000 13640
rect 44081 13635 44147 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 45200 13608 46000 13638
rect 34930 13567 35246 13568
rect 7782 13500 7788 13564
rect 7852 13562 7858 13564
rect 8661 13562 8727 13565
rect 7852 13560 8727 13562
rect 7852 13504 8666 13560
rect 8722 13504 8727 13560
rect 7852 13502 8727 13504
rect 7852 13500 7858 13502
rect 8661 13499 8727 13502
rect 9121 13562 9187 13565
rect 9254 13562 9260 13564
rect 9121 13560 9260 13562
rect 9121 13504 9126 13560
rect 9182 13504 9260 13560
rect 9121 13502 9260 13504
rect 9121 13499 9187 13502
rect 9254 13500 9260 13502
rect 9324 13562 9330 13564
rect 22277 13562 22343 13565
rect 9324 13560 22343 13562
rect 9324 13504 22282 13560
rect 22338 13504 22343 13560
rect 9324 13502 22343 13504
rect 9324 13500 9330 13502
rect 22277 13499 22343 13502
rect 24393 13562 24459 13565
rect 29821 13562 29887 13565
rect 31017 13562 31083 13565
rect 24393 13560 31083 13562
rect 24393 13504 24398 13560
rect 24454 13504 29826 13560
rect 29882 13504 31022 13560
rect 31078 13504 31083 13560
rect 24393 13502 31083 13504
rect 24393 13499 24459 13502
rect 29821 13499 29887 13502
rect 31017 13499 31083 13502
rect 5073 13426 5139 13429
rect 7465 13426 7531 13429
rect 5073 13424 7531 13426
rect 5073 13368 5078 13424
rect 5134 13368 7470 13424
rect 7526 13368 7531 13424
rect 5073 13366 7531 13368
rect 5073 13363 5139 13366
rect 7465 13363 7531 13366
rect 12249 13426 12315 13429
rect 17677 13426 17743 13429
rect 18505 13426 18571 13429
rect 12249 13424 18571 13426
rect 12249 13368 12254 13424
rect 12310 13368 17682 13424
rect 17738 13368 18510 13424
rect 18566 13368 18571 13424
rect 12249 13366 18571 13368
rect 12249 13363 12315 13366
rect 17677 13363 17743 13366
rect 18505 13363 18571 13366
rect 21766 13364 21772 13428
rect 21836 13426 21842 13428
rect 34421 13426 34487 13429
rect 21836 13424 34487 13426
rect 21836 13368 34426 13424
rect 34482 13368 34487 13424
rect 21836 13366 34487 13368
rect 21836 13364 21842 13366
rect 34421 13363 34487 13366
rect 3141 13290 3207 13293
rect 13261 13290 13327 13293
rect 3141 13288 13327 13290
rect 3141 13232 3146 13288
rect 3202 13232 13266 13288
rect 13322 13232 13327 13288
rect 3141 13230 13327 13232
rect 3141 13227 3207 13230
rect 13261 13227 13327 13230
rect 17217 13290 17283 13293
rect 23197 13290 23263 13293
rect 17217 13288 23263 13290
rect 17217 13232 17222 13288
rect 17278 13232 23202 13288
rect 23258 13232 23263 13288
rect 17217 13230 23263 13232
rect 17217 13227 17283 13230
rect 23197 13227 23263 13230
rect 10685 13154 10751 13157
rect 13629 13154 13695 13157
rect 15193 13154 15259 13157
rect 16389 13154 16455 13157
rect 10685 13152 16455 13154
rect 10685 13096 10690 13152
rect 10746 13096 13634 13152
rect 13690 13096 15198 13152
rect 15254 13096 16394 13152
rect 16450 13096 16455 13152
rect 10685 13094 16455 13096
rect 10685 13091 10751 13094
rect 13629 13091 13695 13094
rect 15193 13091 15259 13094
rect 16389 13091 16455 13094
rect 17902 13092 17908 13156
rect 17972 13154 17978 13156
rect 28349 13154 28415 13157
rect 17972 13152 28415 13154
rect 17972 13096 28354 13152
rect 28410 13096 28415 13152
rect 17972 13094 28415 13096
rect 17972 13092 17978 13094
rect 28349 13091 28415 13094
rect 4870 13088 5186 13089
rect 0 13018 800 13048
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 1393 13018 1459 13021
rect 11605 13020 11671 13021
rect 11605 13018 11652 13020
rect 0 13016 1459 13018
rect 0 12960 1398 13016
rect 1454 12960 1459 13016
rect 0 12958 1459 12960
rect 11560 13016 11652 13018
rect 11560 12960 11610 13016
rect 11560 12958 11652 12960
rect 0 12928 800 12958
rect 1393 12955 1459 12958
rect 11605 12956 11652 12958
rect 11716 12956 11722 13020
rect 18229 13018 18295 13021
rect 23933 13018 23999 13021
rect 25630 13018 25636 13020
rect 18229 13016 25636 13018
rect 18229 12960 18234 13016
rect 18290 12960 23938 13016
rect 23994 12960 25636 13016
rect 18229 12958 25636 12960
rect 11605 12955 11671 12956
rect 18229 12955 18295 12958
rect 23933 12955 23999 12958
rect 25630 12956 25636 12958
rect 25700 13018 25706 13020
rect 26049 13018 26115 13021
rect 25700 13016 26115 13018
rect 25700 12960 26054 13016
rect 26110 12960 26115 13016
rect 25700 12958 26115 12960
rect 25700 12956 25706 12958
rect 26049 12955 26115 12958
rect 8661 12882 8727 12885
rect 24393 12882 24459 12885
rect 8661 12880 24459 12882
rect 8661 12824 8666 12880
rect 8722 12824 24398 12880
rect 24454 12824 24459 12880
rect 8661 12822 24459 12824
rect 8661 12819 8727 12822
rect 24393 12819 24459 12822
rect 11145 12746 11211 12749
rect 12525 12746 12591 12749
rect 12985 12746 13051 12749
rect 11145 12744 13051 12746
rect 11145 12688 11150 12744
rect 11206 12688 12530 12744
rect 12586 12688 12990 12744
rect 13046 12688 13051 12744
rect 11145 12686 13051 12688
rect 11145 12683 11211 12686
rect 12525 12683 12591 12686
rect 12985 12683 13051 12686
rect 13445 12746 13511 12749
rect 14733 12746 14799 12749
rect 13445 12744 14799 12746
rect 13445 12688 13450 12744
rect 13506 12688 14738 12744
rect 14794 12688 14799 12744
rect 13445 12686 14799 12688
rect 13445 12683 13511 12686
rect 14733 12683 14799 12686
rect 17677 12746 17743 12749
rect 17902 12746 17908 12748
rect 17677 12744 17908 12746
rect 17677 12688 17682 12744
rect 17738 12688 17908 12744
rect 17677 12686 17908 12688
rect 17677 12683 17743 12686
rect 17902 12684 17908 12686
rect 17972 12684 17978 12748
rect 10777 12610 10843 12613
rect 16481 12610 16547 12613
rect 23197 12610 23263 12613
rect 10777 12608 23263 12610
rect 10777 12552 10782 12608
rect 10838 12552 16486 12608
rect 16542 12552 23202 12608
rect 23258 12552 23263 12608
rect 10777 12550 23263 12552
rect 10777 12547 10843 12550
rect 16481 12547 16547 12550
rect 23197 12547 23263 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 11605 12474 11671 12477
rect 25681 12474 25747 12477
rect 11605 12472 25747 12474
rect 11605 12416 11610 12472
rect 11666 12416 25686 12472
rect 25742 12416 25747 12472
rect 11605 12414 25747 12416
rect 11605 12411 11671 12414
rect 25681 12411 25747 12414
rect 0 12338 800 12368
rect 0 12248 858 12338
rect 7046 12276 7052 12340
rect 7116 12338 7122 12340
rect 27153 12338 27219 12341
rect 7116 12336 27219 12338
rect 7116 12280 27158 12336
rect 27214 12280 27219 12336
rect 7116 12278 27219 12280
rect 7116 12276 7122 12278
rect 27153 12275 27219 12278
rect 798 12205 858 12248
rect 798 12200 907 12205
rect 798 12144 846 12200
rect 902 12144 907 12200
rect 798 12142 907 12144
rect 841 12139 907 12142
rect 15510 12140 15516 12204
rect 15580 12202 15586 12204
rect 29085 12202 29151 12205
rect 15580 12200 29151 12202
rect 15580 12144 29090 12200
rect 29146 12144 29151 12200
rect 15580 12142 29151 12144
rect 15580 12140 15586 12142
rect 29085 12139 29151 12142
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 841 11794 907 11797
rect 798 11792 907 11794
rect 798 11736 846 11792
rect 902 11736 907 11792
rect 798 11731 907 11736
rect 798 11688 858 11731
rect 0 11598 858 11688
rect 0 11568 800 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 8702 10916 8708 10980
rect 8772 10978 8778 10980
rect 27613 10978 27679 10981
rect 8772 10976 27679 10978
rect 8772 10920 27618 10976
rect 27674 10920 27679 10976
rect 8772 10918 27679 10920
rect 8772 10916 8778 10918
rect 27613 10915 27679 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 25084 33220 25148 33284
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 23244 32056 23308 32060
rect 23244 32000 23294 32056
rect 23294 32000 23308 32056
rect 23244 31996 23308 32000
rect 28028 32132 28092 32196
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 28212 31996 28276 32060
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 19196 31180 19260 31244
rect 19932 31044 19996 31108
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 33364 30696 33428 30700
rect 33364 30640 33414 30696
rect 33414 30640 33428 30696
rect 19748 30500 19812 30564
rect 33364 30636 33428 30640
rect 29684 30500 29748 30564
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 15332 29956 15396 30020
rect 17540 30152 17604 30156
rect 17540 30096 17590 30152
rect 17590 30096 17604 30152
rect 17540 30092 17604 30096
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 21588 29548 21652 29612
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 15700 29140 15764 29204
rect 13308 29064 13372 29068
rect 13308 29008 13322 29064
rect 13322 29008 13372 29064
rect 13308 29004 13372 29008
rect 13492 29064 13556 29068
rect 13492 29008 13542 29064
rect 13542 29008 13556 29064
rect 13492 29004 13556 29008
rect 17356 29064 17420 29068
rect 17356 29008 17370 29064
rect 17370 29008 17420 29064
rect 17356 29004 17420 29008
rect 23980 29004 24044 29068
rect 36124 29140 36188 29204
rect 28580 29004 28644 29068
rect 31524 29064 31588 29068
rect 31524 29008 31538 29064
rect 31538 29008 31588 29064
rect 31524 29004 31588 29008
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19564 28732 19628 28796
rect 32260 28324 32324 28388
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 10732 28188 10796 28252
rect 28948 28188 29012 28252
rect 15516 28112 15580 28116
rect 15516 28056 15530 28112
rect 15530 28056 15580 28112
rect 15516 28052 15580 28056
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 32812 27704 32876 27708
rect 32812 27648 32826 27704
rect 32826 27648 32876 27704
rect 32812 27644 32876 27648
rect 34468 27644 34532 27708
rect 35388 27644 35452 27708
rect 37228 27508 37292 27572
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 9260 27100 9324 27164
rect 34652 27100 34716 27164
rect 27108 26828 27172 26892
rect 20668 26752 20732 26756
rect 20668 26696 20682 26752
rect 20682 26696 20732 26752
rect 20668 26692 20732 26696
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 22692 26556 22756 26620
rect 34284 26692 34348 26756
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 32444 26556 32508 26620
rect 18276 26284 18340 26348
rect 25636 26284 25700 26348
rect 25820 26344 25884 26348
rect 25820 26288 25834 26344
rect 25834 26288 25884 26344
rect 25820 26284 25884 26288
rect 30788 26284 30852 26348
rect 21956 26148 22020 26212
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 11836 26012 11900 26076
rect 33548 26012 33612 26076
rect 36308 26012 36372 26076
rect 8156 25664 8220 25668
rect 8156 25608 8206 25664
rect 8206 25608 8220 25664
rect 8156 25604 8220 25608
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 25452 25604 25516 25668
rect 33548 25604 33612 25668
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 16252 25256 16316 25260
rect 16252 25200 16302 25256
rect 16302 25200 16316 25256
rect 16252 25196 16316 25200
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 7972 24984 8036 24988
rect 7972 24928 7986 24984
rect 7986 24928 8036 24984
rect 7972 24924 8036 24928
rect 10548 24984 10612 24988
rect 10548 24928 10598 24984
rect 10598 24928 10612 24984
rect 10548 24924 10612 24928
rect 19380 24924 19444 24988
rect 24716 24924 24780 24988
rect 26556 24924 26620 24988
rect 27292 24924 27356 24988
rect 28764 24924 28828 24988
rect 30052 24924 30116 24988
rect 34100 24924 34164 24988
rect 26372 24848 26436 24852
rect 26372 24792 26422 24848
rect 26422 24792 26436 24848
rect 26372 24788 26436 24792
rect 26924 24788 26988 24852
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 8708 24712 8772 24716
rect 8708 24656 8758 24712
rect 8758 24656 8772 24712
rect 8708 24652 8772 24656
rect 14412 24712 14476 24716
rect 14412 24656 14426 24712
rect 14426 24656 14476 24712
rect 14412 24652 14476 24656
rect 9996 24576 10060 24580
rect 9996 24520 10010 24576
rect 10010 24520 10060 24576
rect 9996 24516 10060 24520
rect 11100 24516 11164 24580
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 21772 24380 21836 24444
rect 22876 24576 22940 24580
rect 22876 24520 22926 24576
rect 22926 24520 22940 24576
rect 22876 24516 22940 24520
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 13676 24304 13740 24308
rect 13676 24248 13690 24304
rect 13690 24248 13740 24304
rect 13676 24244 13740 24248
rect 22508 24244 22572 24308
rect 26004 24244 26068 24308
rect 26188 24244 26252 24308
rect 14044 24108 14108 24172
rect 15148 24168 15212 24172
rect 15148 24112 15162 24168
rect 15162 24112 15212 24168
rect 15148 24108 15212 24112
rect 22692 24108 22756 24172
rect 24900 24108 24964 24172
rect 26556 24108 26620 24172
rect 34468 24032 34532 24036
rect 34468 23976 34482 24032
rect 34482 23976 34532 24032
rect 34468 23972 34532 23976
rect 34652 23972 34716 24036
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 30972 23700 31036 23764
rect 37228 23700 37292 23764
rect 7052 23564 7116 23628
rect 19012 23564 19076 23628
rect 7788 23488 7852 23492
rect 7788 23432 7838 23488
rect 7838 23432 7852 23488
rect 7788 23428 7852 23432
rect 12204 23428 12268 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 11652 23292 11716 23356
rect 29316 23428 29380 23492
rect 31892 23428 31956 23492
rect 32996 23488 33060 23492
rect 32996 23432 33010 23488
rect 33010 23432 33060 23488
rect 32996 23428 33060 23432
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 9996 23156 10060 23220
rect 22692 23156 22756 23220
rect 29684 23156 29748 23220
rect 34284 23156 34348 23220
rect 35388 23020 35452 23084
rect 10732 22944 10796 22948
rect 10732 22888 10782 22944
rect 10782 22888 10796 22944
rect 10732 22884 10796 22888
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 13308 22808 13372 22812
rect 13308 22752 13358 22808
rect 13358 22752 13372 22808
rect 13308 22748 13372 22752
rect 19380 22748 19444 22812
rect 25636 22884 25700 22948
rect 31156 22884 31220 22948
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 8892 22476 8956 22540
rect 17908 22476 17972 22540
rect 10732 22340 10796 22404
rect 18276 22340 18340 22404
rect 26556 22340 26620 22404
rect 28948 22400 29012 22404
rect 28948 22344 28998 22400
rect 28998 22344 29012 22400
rect 28948 22340 29012 22344
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 32628 22264 32692 22268
rect 32628 22208 32678 22264
rect 32678 22208 32692 22264
rect 32628 22204 32692 22208
rect 24716 22068 24780 22132
rect 12940 21932 13004 21996
rect 25268 21932 25332 21996
rect 32444 21932 32508 21996
rect 17908 21796 17972 21860
rect 34652 21932 34716 21996
rect 36308 21932 36372 21996
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 21588 21660 21652 21724
rect 33180 21720 33244 21724
rect 33180 21664 33230 21720
rect 33230 21664 33244 21720
rect 33180 21660 33244 21664
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 22324 21524 22388 21588
rect 26004 21584 26068 21588
rect 26004 21528 26018 21584
rect 26018 21528 26068 21584
rect 26004 21524 26068 21528
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 25084 21176 25148 21180
rect 25084 21120 25134 21176
rect 25134 21120 25148 21176
rect 25084 21116 25148 21120
rect 26372 21176 26436 21180
rect 26372 21120 26422 21176
rect 26422 21120 26436 21176
rect 26372 21116 26436 21120
rect 27292 21116 27356 21180
rect 20668 20844 20732 20908
rect 12940 20708 13004 20772
rect 17908 20708 17972 20772
rect 21588 20708 21652 20772
rect 23244 20768 23308 20772
rect 23244 20712 23294 20768
rect 23294 20712 23308 20768
rect 23244 20708 23308 20712
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 9444 20572 9508 20636
rect 13308 20572 13372 20636
rect 27108 20708 27172 20772
rect 27476 20708 27540 20772
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 26188 20572 26252 20636
rect 28028 20632 28092 20636
rect 28028 20576 28042 20632
rect 28042 20576 28092 20632
rect 28028 20572 28092 20576
rect 29316 20572 29380 20636
rect 32260 20572 32324 20636
rect 10732 20300 10796 20364
rect 15332 20300 15396 20364
rect 32628 20436 32692 20500
rect 29316 20300 29380 20364
rect 24900 20164 24964 20228
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 25268 20028 25332 20092
rect 28948 20088 29012 20092
rect 28948 20032 28998 20088
rect 28998 20032 29012 20088
rect 28948 20028 29012 20032
rect 9444 19892 9508 19956
rect 9812 19952 9876 19956
rect 9812 19896 9826 19952
rect 9826 19896 9876 19952
rect 9812 19892 9876 19896
rect 10548 19952 10612 19956
rect 10548 19896 10562 19952
rect 10562 19896 10612 19952
rect 10548 19892 10612 19896
rect 30604 19680 30668 19684
rect 30604 19624 30618 19680
rect 30618 19624 30668 19680
rect 30604 19620 30668 19624
rect 31156 19620 31220 19684
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 11836 19484 11900 19548
rect 21956 19484 22020 19548
rect 29316 19484 29380 19548
rect 34100 19756 34164 19820
rect 34652 19756 34716 19820
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 15148 19408 15212 19412
rect 15148 19352 15162 19408
rect 15162 19352 15212 19408
rect 15148 19348 15212 19352
rect 8708 19212 8772 19276
rect 27292 19408 27356 19412
rect 27292 19352 27342 19408
rect 27342 19352 27356 19408
rect 27292 19348 27356 19352
rect 19380 19212 19444 19276
rect 30788 19212 30852 19276
rect 14412 19076 14476 19140
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19564 18940 19628 19004
rect 15700 18668 15764 18732
rect 28764 18532 28828 18596
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 19380 18396 19444 18460
rect 26924 18396 26988 18460
rect 9996 18320 10060 18324
rect 9996 18264 10010 18320
rect 10010 18264 10060 18320
rect 9996 18260 10060 18264
rect 10732 18320 10796 18324
rect 10732 18264 10746 18320
rect 10746 18264 10796 18320
rect 10732 18260 10796 18264
rect 19748 18260 19812 18324
rect 22508 18124 22572 18188
rect 19932 17988 19996 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 14044 17852 14108 17916
rect 28580 18048 28644 18052
rect 28580 17992 28594 18048
rect 28594 17992 28644 18048
rect 28580 17988 28644 17992
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 7052 17716 7116 17780
rect 13308 17716 13372 17780
rect 28948 17716 29012 17780
rect 22692 17444 22756 17508
rect 32996 17716 33060 17780
rect 30052 17444 30116 17508
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 13676 17308 13740 17372
rect 25268 17172 25332 17236
rect 31892 17036 31956 17100
rect 24716 16960 24780 16964
rect 24716 16904 24766 16960
rect 24766 16904 24780 16960
rect 24716 16900 24780 16904
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 17540 16764 17604 16828
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 33548 16764 33612 16828
rect 25820 16492 25884 16556
rect 10732 16356 10796 16420
rect 22876 16356 22940 16420
rect 27108 16356 27172 16420
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 8892 16084 8956 16148
rect 32812 16220 32876 16284
rect 8156 15948 8220 16012
rect 9812 15948 9876 16012
rect 16252 16008 16316 16012
rect 16252 15952 16266 16008
rect 16266 15952 16316 16008
rect 16252 15948 16316 15952
rect 19012 15948 19076 16012
rect 13492 15812 13556 15876
rect 22324 16008 22388 16012
rect 22324 15952 22338 16008
rect 22338 15952 22388 16008
rect 22324 15948 22388 15952
rect 29684 16008 29748 16012
rect 29684 15952 29734 16008
rect 29734 15952 29748 16008
rect 29684 15948 29748 15952
rect 32996 15812 33060 15876
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 15516 15676 15580 15740
rect 29316 15540 29380 15604
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 11100 15192 11164 15196
rect 11100 15136 11114 15192
rect 11114 15136 11164 15192
rect 11100 15132 11164 15136
rect 27476 15132 27540 15196
rect 30972 15132 31036 15196
rect 17356 14996 17420 15060
rect 30604 14996 30668 15060
rect 36124 14996 36188 15060
rect 31524 14784 31588 14788
rect 31524 14728 31574 14784
rect 31574 14728 31588 14784
rect 31524 14724 31588 14728
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 17356 14588 17420 14652
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 23980 14044 24044 14108
rect 28212 14044 28276 14108
rect 12204 13772 12268 13836
rect 7972 13696 8036 13700
rect 7972 13640 7986 13696
rect 7986 13640 8036 13696
rect 7972 13636 8036 13640
rect 25452 13636 25516 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 7788 13500 7852 13564
rect 9260 13500 9324 13564
rect 21772 13364 21836 13428
rect 17908 13092 17972 13156
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 11652 13016 11716 13020
rect 11652 12960 11666 13016
rect 11666 12960 11716 13016
rect 11652 12956 11716 12960
rect 25636 12956 25700 13020
rect 17908 12684 17972 12748
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 7052 12276 7116 12340
rect 15516 12140 15580 12204
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 8708 10916 8772 10980
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 37024 5188 37584
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 35936 5188 36960
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 25083 33284 25149 33285
rect 25083 33220 25084 33284
rect 25148 33220 25149 33284
rect 25083 33219 25149 33220
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 23243 32060 23309 32061
rect 23243 31996 23244 32060
rect 23308 31996 23309 32060
rect 23243 31995 23309 31996
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 19195 31244 19261 31245
rect 19195 31180 19196 31244
rect 19260 31180 19261 31244
rect 19195 31179 19261 31180
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 17539 30156 17605 30157
rect 17539 30092 17540 30156
rect 17604 30092 17605 30156
rect 17539 30091 17605 30092
rect 15331 30020 15397 30021
rect 15331 29956 15332 30020
rect 15396 29956 15397 30020
rect 15331 29955 15397 29956
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 13307 29068 13373 29069
rect 13307 29004 13308 29068
rect 13372 29004 13373 29068
rect 13307 29003 13373 29004
rect 13491 29068 13557 29069
rect 13491 29004 13492 29068
rect 13556 29004 13557 29068
rect 13491 29003 13557 29004
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 10731 28252 10797 28253
rect 10731 28188 10732 28252
rect 10796 28188 10797 28252
rect 10731 28187 10797 28188
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 9259 27164 9325 27165
rect 9259 27100 9260 27164
rect 9324 27100 9325 27164
rect 9259 27099 9325 27100
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 8155 25668 8221 25669
rect 8155 25604 8156 25668
rect 8220 25604 8221 25668
rect 8155 25603 8221 25604
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 7971 24988 8037 24989
rect 7971 24924 7972 24988
rect 8036 24924 8037 24988
rect 7971 24923 8037 24924
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 7051 23628 7117 23629
rect 7051 23564 7052 23628
rect 7116 23564 7117 23628
rect 7051 23563 7117 23564
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 7054 17781 7114 23563
rect 7787 23492 7853 23493
rect 7787 23428 7788 23492
rect 7852 23428 7853 23492
rect 7787 23427 7853 23428
rect 7051 17780 7117 17781
rect 7051 17716 7052 17780
rect 7116 17716 7117 17780
rect 7051 17715 7117 17716
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 7054 12341 7114 17715
rect 7790 13565 7850 23427
rect 7974 13701 8034 24923
rect 8158 16013 8218 25603
rect 8707 24716 8773 24717
rect 8707 24652 8708 24716
rect 8772 24652 8773 24716
rect 8707 24651 8773 24652
rect 8710 19277 8770 24651
rect 8891 22540 8957 22541
rect 8891 22476 8892 22540
rect 8956 22476 8957 22540
rect 8891 22475 8957 22476
rect 8707 19276 8773 19277
rect 8707 19212 8708 19276
rect 8772 19212 8773 19276
rect 8707 19211 8773 19212
rect 8155 16012 8221 16013
rect 8155 15948 8156 16012
rect 8220 15948 8221 16012
rect 8155 15947 8221 15948
rect 7971 13700 8037 13701
rect 7971 13636 7972 13700
rect 8036 13636 8037 13700
rect 7971 13635 8037 13636
rect 7787 13564 7853 13565
rect 7787 13500 7788 13564
rect 7852 13500 7853 13564
rect 7787 13499 7853 13500
rect 7051 12340 7117 12341
rect 7051 12276 7052 12340
rect 7116 12276 7117 12340
rect 7051 12275 7117 12276
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 8710 10981 8770 19211
rect 8894 16149 8954 22475
rect 8891 16148 8957 16149
rect 8891 16084 8892 16148
rect 8956 16084 8957 16148
rect 8891 16083 8957 16084
rect 9262 13565 9322 27099
rect 10547 24988 10613 24989
rect 10547 24924 10548 24988
rect 10612 24924 10613 24988
rect 10547 24923 10613 24924
rect 9995 24580 10061 24581
rect 9995 24516 9996 24580
rect 10060 24516 10061 24580
rect 9995 24515 10061 24516
rect 9998 23221 10058 24515
rect 9995 23220 10061 23221
rect 9995 23156 9996 23220
rect 10060 23156 10061 23220
rect 9995 23155 10061 23156
rect 9443 20636 9509 20637
rect 9443 20572 9444 20636
rect 9508 20572 9509 20636
rect 9443 20571 9509 20572
rect 9446 19957 9506 20571
rect 9443 19956 9509 19957
rect 9443 19892 9444 19956
rect 9508 19892 9509 19956
rect 9443 19891 9509 19892
rect 9811 19956 9877 19957
rect 9811 19892 9812 19956
rect 9876 19892 9877 19956
rect 9811 19891 9877 19892
rect 9814 16013 9874 19891
rect 9998 18325 10058 23155
rect 10550 19957 10610 24923
rect 10734 22949 10794 28187
rect 11835 26076 11901 26077
rect 11835 26012 11836 26076
rect 11900 26012 11901 26076
rect 11835 26011 11901 26012
rect 11099 24580 11165 24581
rect 11099 24516 11100 24580
rect 11164 24516 11165 24580
rect 11099 24515 11165 24516
rect 10731 22948 10797 22949
rect 10731 22884 10732 22948
rect 10796 22884 10797 22948
rect 10731 22883 10797 22884
rect 10731 22404 10797 22405
rect 10731 22340 10732 22404
rect 10796 22340 10797 22404
rect 10731 22339 10797 22340
rect 10734 20365 10794 22339
rect 10731 20364 10797 20365
rect 10731 20300 10732 20364
rect 10796 20300 10797 20364
rect 10731 20299 10797 20300
rect 10547 19956 10613 19957
rect 10547 19892 10548 19956
rect 10612 19892 10613 19956
rect 10547 19891 10613 19892
rect 9995 18324 10061 18325
rect 9995 18260 9996 18324
rect 10060 18260 10061 18324
rect 9995 18259 10061 18260
rect 10731 18324 10797 18325
rect 10731 18260 10732 18324
rect 10796 18260 10797 18324
rect 10731 18259 10797 18260
rect 10734 16421 10794 18259
rect 10731 16420 10797 16421
rect 10731 16356 10732 16420
rect 10796 16356 10797 16420
rect 10731 16355 10797 16356
rect 9811 16012 9877 16013
rect 9811 15948 9812 16012
rect 9876 15948 9877 16012
rect 9811 15947 9877 15948
rect 11102 15197 11162 24515
rect 11651 23356 11717 23357
rect 11651 23292 11652 23356
rect 11716 23292 11717 23356
rect 11651 23291 11717 23292
rect 11099 15196 11165 15197
rect 11099 15132 11100 15196
rect 11164 15132 11165 15196
rect 11099 15131 11165 15132
rect 9259 13564 9325 13565
rect 9259 13500 9260 13564
rect 9324 13500 9325 13564
rect 9259 13499 9325 13500
rect 11654 13021 11714 23291
rect 11838 19549 11898 26011
rect 12203 23492 12269 23493
rect 12203 23428 12204 23492
rect 12268 23428 12269 23492
rect 12203 23427 12269 23428
rect 11835 19548 11901 19549
rect 11835 19484 11836 19548
rect 11900 19484 11901 19548
rect 11835 19483 11901 19484
rect 12206 13837 12266 23427
rect 13310 22813 13370 29003
rect 13307 22812 13373 22813
rect 13307 22748 13308 22812
rect 13372 22748 13373 22812
rect 13307 22747 13373 22748
rect 12939 21996 13005 21997
rect 12939 21932 12940 21996
rect 13004 21932 13005 21996
rect 12939 21931 13005 21932
rect 12942 20773 13002 21931
rect 12939 20772 13005 20773
rect 12939 20708 12940 20772
rect 13004 20708 13005 20772
rect 12939 20707 13005 20708
rect 13307 20636 13373 20637
rect 13307 20572 13308 20636
rect 13372 20572 13373 20636
rect 13307 20571 13373 20572
rect 13310 17781 13370 20571
rect 13307 17780 13373 17781
rect 13307 17716 13308 17780
rect 13372 17716 13373 17780
rect 13307 17715 13373 17716
rect 13494 15877 13554 29003
rect 14411 24716 14477 24717
rect 14411 24652 14412 24716
rect 14476 24652 14477 24716
rect 14411 24651 14477 24652
rect 13675 24308 13741 24309
rect 13675 24244 13676 24308
rect 13740 24244 13741 24308
rect 13675 24243 13741 24244
rect 13678 17373 13738 24243
rect 14043 24172 14109 24173
rect 14043 24108 14044 24172
rect 14108 24108 14109 24172
rect 14043 24107 14109 24108
rect 14046 17917 14106 24107
rect 14414 19141 14474 24651
rect 15147 24172 15213 24173
rect 15147 24108 15148 24172
rect 15212 24108 15213 24172
rect 15147 24107 15213 24108
rect 15150 19413 15210 24107
rect 15334 20365 15394 29955
rect 15699 29204 15765 29205
rect 15699 29140 15700 29204
rect 15764 29140 15765 29204
rect 15699 29139 15765 29140
rect 15515 28116 15581 28117
rect 15515 28052 15516 28116
rect 15580 28052 15581 28116
rect 15515 28051 15581 28052
rect 15331 20364 15397 20365
rect 15331 20300 15332 20364
rect 15396 20300 15397 20364
rect 15331 20299 15397 20300
rect 15147 19412 15213 19413
rect 15147 19348 15148 19412
rect 15212 19348 15213 19412
rect 15147 19347 15213 19348
rect 14411 19140 14477 19141
rect 14411 19076 14412 19140
rect 14476 19076 14477 19140
rect 14411 19075 14477 19076
rect 14043 17916 14109 17917
rect 14043 17852 14044 17916
rect 14108 17852 14109 17916
rect 14043 17851 14109 17852
rect 13675 17372 13741 17373
rect 13675 17308 13676 17372
rect 13740 17308 13741 17372
rect 13675 17307 13741 17308
rect 13491 15876 13557 15877
rect 13491 15812 13492 15876
rect 13556 15812 13557 15876
rect 13491 15811 13557 15812
rect 15518 15741 15578 28051
rect 15702 18733 15762 29139
rect 17355 29068 17421 29069
rect 17355 29004 17356 29068
rect 17420 29004 17421 29068
rect 17355 29003 17421 29004
rect 16251 25260 16317 25261
rect 16251 25196 16252 25260
rect 16316 25196 16317 25260
rect 16251 25195 16317 25196
rect 15699 18732 15765 18733
rect 15699 18668 15700 18732
rect 15764 18668 15765 18732
rect 15699 18667 15765 18668
rect 16254 16013 16314 25195
rect 16251 16012 16317 16013
rect 16251 15948 16252 16012
rect 16316 15948 16317 16012
rect 16251 15947 16317 15948
rect 15515 15740 15581 15741
rect 15515 15676 15516 15740
rect 15580 15676 15581 15740
rect 15515 15675 15581 15676
rect 12203 13836 12269 13837
rect 12203 13772 12204 13836
rect 12268 13772 12269 13836
rect 12203 13771 12269 13772
rect 11651 13020 11717 13021
rect 11651 12956 11652 13020
rect 11716 12956 11717 13020
rect 11651 12955 11717 12956
rect 15518 12205 15578 15675
rect 17358 15061 17418 29003
rect 17542 16829 17602 30091
rect 18275 26348 18341 26349
rect 18275 26284 18276 26348
rect 18340 26284 18341 26348
rect 18275 26283 18341 26284
rect 17907 22540 17973 22541
rect 17907 22476 17908 22540
rect 17972 22476 17973 22540
rect 17907 22475 17973 22476
rect 17910 21861 17970 22475
rect 18278 22405 18338 26283
rect 19198 24850 19258 31179
rect 19931 31108 19997 31109
rect 19931 31044 19932 31108
rect 19996 31044 19997 31108
rect 19931 31043 19997 31044
rect 19747 30564 19813 30565
rect 19747 30500 19748 30564
rect 19812 30500 19813 30564
rect 19747 30499 19813 30500
rect 19563 28796 19629 28797
rect 19563 28732 19564 28796
rect 19628 28732 19629 28796
rect 19563 28731 19629 28732
rect 19379 24988 19445 24989
rect 19379 24924 19380 24988
rect 19444 24924 19445 24988
rect 19379 24923 19445 24924
rect 19382 24850 19442 24923
rect 19198 24790 19442 24850
rect 19011 23628 19077 23629
rect 19011 23564 19012 23628
rect 19076 23564 19077 23628
rect 19011 23563 19077 23564
rect 18275 22404 18341 22405
rect 18275 22340 18276 22404
rect 18340 22340 18341 22404
rect 18275 22339 18341 22340
rect 17907 21860 17973 21861
rect 17907 21796 17908 21860
rect 17972 21796 17973 21860
rect 17907 21795 17973 21796
rect 17907 20772 17973 20773
rect 17907 20708 17908 20772
rect 17972 20708 17973 20772
rect 17907 20707 17973 20708
rect 17539 16828 17605 16829
rect 17539 16764 17540 16828
rect 17604 16764 17605 16828
rect 17539 16763 17605 16764
rect 17355 15060 17421 15061
rect 17355 14996 17356 15060
rect 17420 14996 17421 15060
rect 17355 14995 17421 14996
rect 17358 14653 17418 14995
rect 17355 14652 17421 14653
rect 17355 14588 17356 14652
rect 17420 14588 17421 14652
rect 17355 14587 17421 14588
rect 17910 13157 17970 20707
rect 19014 16013 19074 23563
rect 19382 22813 19442 24790
rect 19379 22812 19445 22813
rect 19379 22748 19380 22812
rect 19444 22748 19445 22812
rect 19379 22747 19445 22748
rect 19379 19276 19445 19277
rect 19379 19212 19380 19276
rect 19444 19212 19445 19276
rect 19379 19211 19445 19212
rect 19382 18461 19442 19211
rect 19566 19005 19626 28731
rect 19563 19004 19629 19005
rect 19563 18940 19564 19004
rect 19628 18940 19629 19004
rect 19563 18939 19629 18940
rect 19379 18460 19445 18461
rect 19379 18396 19380 18460
rect 19444 18396 19445 18460
rect 19379 18395 19445 18396
rect 19750 18325 19810 30499
rect 19747 18324 19813 18325
rect 19747 18260 19748 18324
rect 19812 18260 19813 18324
rect 19747 18259 19813 18260
rect 19934 18053 19994 31043
rect 21587 29612 21653 29613
rect 21587 29548 21588 29612
rect 21652 29548 21653 29612
rect 21587 29547 21653 29548
rect 20667 26756 20733 26757
rect 20667 26692 20668 26756
rect 20732 26692 20733 26756
rect 20667 26691 20733 26692
rect 20670 20909 20730 26691
rect 21590 21725 21650 29547
rect 22691 26620 22757 26621
rect 22691 26556 22692 26620
rect 22756 26556 22757 26620
rect 22691 26555 22757 26556
rect 21955 26212 22021 26213
rect 21955 26148 21956 26212
rect 22020 26148 22021 26212
rect 21955 26147 22021 26148
rect 21771 24444 21837 24445
rect 21771 24380 21772 24444
rect 21836 24380 21837 24444
rect 21771 24379 21837 24380
rect 21587 21724 21653 21725
rect 21587 21660 21588 21724
rect 21652 21660 21653 21724
rect 21587 21659 21653 21660
rect 20667 20908 20733 20909
rect 20667 20844 20668 20908
rect 20732 20844 20733 20908
rect 20667 20843 20733 20844
rect 21590 20773 21650 21659
rect 21587 20772 21653 20773
rect 21587 20708 21588 20772
rect 21652 20708 21653 20772
rect 21587 20707 21653 20708
rect 19931 18052 19997 18053
rect 19931 17988 19932 18052
rect 19996 17988 19997 18052
rect 19931 17987 19997 17988
rect 19011 16012 19077 16013
rect 19011 15948 19012 16012
rect 19076 15948 19077 16012
rect 19011 15947 19077 15948
rect 21774 13429 21834 24379
rect 21958 19549 22018 26147
rect 22507 24308 22573 24309
rect 22507 24244 22508 24308
rect 22572 24244 22573 24308
rect 22507 24243 22573 24244
rect 22323 21588 22389 21589
rect 22323 21524 22324 21588
rect 22388 21524 22389 21588
rect 22323 21523 22389 21524
rect 21955 19548 22021 19549
rect 21955 19484 21956 19548
rect 22020 19484 22021 19548
rect 21955 19483 22021 19484
rect 22326 16013 22386 21523
rect 22510 18189 22570 24243
rect 22694 24173 22754 26555
rect 22875 24580 22941 24581
rect 22875 24516 22876 24580
rect 22940 24516 22941 24580
rect 22875 24515 22941 24516
rect 22691 24172 22757 24173
rect 22691 24108 22692 24172
rect 22756 24108 22757 24172
rect 22691 24107 22757 24108
rect 22694 23221 22754 24107
rect 22691 23220 22757 23221
rect 22691 23156 22692 23220
rect 22756 23156 22757 23220
rect 22691 23155 22757 23156
rect 22507 18188 22573 18189
rect 22507 18124 22508 18188
rect 22572 18124 22573 18188
rect 22507 18123 22573 18124
rect 22694 17509 22754 23155
rect 22691 17508 22757 17509
rect 22691 17444 22692 17508
rect 22756 17444 22757 17508
rect 22691 17443 22757 17444
rect 22878 16421 22938 24515
rect 23246 20773 23306 31995
rect 23979 29068 24045 29069
rect 23979 29004 23980 29068
rect 24044 29004 24045 29068
rect 23979 29003 24045 29004
rect 23243 20772 23309 20773
rect 23243 20708 23244 20772
rect 23308 20708 23309 20772
rect 23243 20707 23309 20708
rect 22875 16420 22941 16421
rect 22875 16356 22876 16420
rect 22940 16356 22941 16420
rect 22875 16355 22941 16356
rect 22323 16012 22389 16013
rect 22323 15948 22324 16012
rect 22388 15948 22389 16012
rect 22323 15947 22389 15948
rect 23982 14109 24042 29003
rect 24715 24988 24781 24989
rect 24715 24924 24716 24988
rect 24780 24924 24781 24988
rect 24715 24923 24781 24924
rect 24718 22133 24778 24923
rect 24899 24172 24965 24173
rect 24899 24108 24900 24172
rect 24964 24108 24965 24172
rect 24899 24107 24965 24108
rect 24715 22132 24781 22133
rect 24715 22068 24716 22132
rect 24780 22068 24781 22132
rect 24715 22067 24781 22068
rect 24718 16965 24778 22067
rect 24902 20229 24962 24107
rect 25086 21181 25146 33219
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 28027 32196 28093 32197
rect 28027 32132 28028 32196
rect 28092 32132 28093 32196
rect 28027 32131 28093 32132
rect 27107 26892 27173 26893
rect 27107 26828 27108 26892
rect 27172 26828 27173 26892
rect 27107 26827 27173 26828
rect 25635 26348 25701 26349
rect 25635 26284 25636 26348
rect 25700 26284 25701 26348
rect 25635 26283 25701 26284
rect 25819 26348 25885 26349
rect 25819 26284 25820 26348
rect 25884 26284 25885 26348
rect 25819 26283 25885 26284
rect 25451 25668 25517 25669
rect 25451 25604 25452 25668
rect 25516 25604 25517 25668
rect 25451 25603 25517 25604
rect 25267 21996 25333 21997
rect 25267 21932 25268 21996
rect 25332 21932 25333 21996
rect 25267 21931 25333 21932
rect 25083 21180 25149 21181
rect 25083 21116 25084 21180
rect 25148 21116 25149 21180
rect 25083 21115 25149 21116
rect 24899 20228 24965 20229
rect 24899 20164 24900 20228
rect 24964 20164 24965 20228
rect 24899 20163 24965 20164
rect 25270 20093 25330 21931
rect 25267 20092 25333 20093
rect 25267 20028 25268 20092
rect 25332 20028 25333 20092
rect 25267 20027 25333 20028
rect 25270 17237 25330 20027
rect 25267 17236 25333 17237
rect 25267 17172 25268 17236
rect 25332 17172 25333 17236
rect 25267 17171 25333 17172
rect 24715 16964 24781 16965
rect 24715 16900 24716 16964
rect 24780 16900 24781 16964
rect 24715 16899 24781 16900
rect 23979 14108 24045 14109
rect 23979 14044 23980 14108
rect 24044 14044 24045 14108
rect 23979 14043 24045 14044
rect 25454 13701 25514 25603
rect 25638 22949 25698 26283
rect 25635 22948 25701 22949
rect 25635 22884 25636 22948
rect 25700 22884 25701 22948
rect 25635 22883 25701 22884
rect 25451 13700 25517 13701
rect 25451 13636 25452 13700
rect 25516 13636 25517 13700
rect 25451 13635 25517 13636
rect 21771 13428 21837 13429
rect 21771 13364 21772 13428
rect 21836 13364 21837 13428
rect 21771 13363 21837 13364
rect 17907 13156 17973 13157
rect 17907 13092 17908 13156
rect 17972 13092 17973 13156
rect 17907 13091 17973 13092
rect 17910 12749 17970 13091
rect 25638 13021 25698 22883
rect 25822 16557 25882 26283
rect 26555 24988 26621 24989
rect 26555 24924 26556 24988
rect 26620 24924 26621 24988
rect 26555 24923 26621 24924
rect 26371 24852 26437 24853
rect 26371 24788 26372 24852
rect 26436 24788 26437 24852
rect 26371 24787 26437 24788
rect 26003 24308 26069 24309
rect 26003 24244 26004 24308
rect 26068 24244 26069 24308
rect 26003 24243 26069 24244
rect 26187 24308 26253 24309
rect 26187 24244 26188 24308
rect 26252 24244 26253 24308
rect 26187 24243 26253 24244
rect 26006 21589 26066 24243
rect 26003 21588 26069 21589
rect 26003 21524 26004 21588
rect 26068 21524 26069 21588
rect 26003 21523 26069 21524
rect 26190 20637 26250 24243
rect 26374 21181 26434 24787
rect 26558 24173 26618 24923
rect 26923 24852 26989 24853
rect 26923 24788 26924 24852
rect 26988 24788 26989 24852
rect 26923 24787 26989 24788
rect 26555 24172 26621 24173
rect 26555 24108 26556 24172
rect 26620 24108 26621 24172
rect 26555 24107 26621 24108
rect 26558 22405 26618 24107
rect 26555 22404 26621 22405
rect 26555 22340 26556 22404
rect 26620 22340 26621 22404
rect 26555 22339 26621 22340
rect 26371 21180 26437 21181
rect 26371 21116 26372 21180
rect 26436 21116 26437 21180
rect 26371 21115 26437 21116
rect 26187 20636 26253 20637
rect 26187 20572 26188 20636
rect 26252 20572 26253 20636
rect 26187 20571 26253 20572
rect 26926 18461 26986 24787
rect 27110 20773 27170 26827
rect 27291 24988 27357 24989
rect 27291 24924 27292 24988
rect 27356 24924 27357 24988
rect 27291 24923 27357 24924
rect 27294 21181 27354 24923
rect 27291 21180 27357 21181
rect 27291 21116 27292 21180
rect 27356 21116 27357 21180
rect 27291 21115 27357 21116
rect 27107 20772 27173 20773
rect 27107 20708 27108 20772
rect 27172 20708 27173 20772
rect 27107 20707 27173 20708
rect 26923 18460 26989 18461
rect 26923 18396 26924 18460
rect 26988 18396 26989 18460
rect 26923 18395 26989 18396
rect 25819 16556 25885 16557
rect 25819 16492 25820 16556
rect 25884 16492 25885 16556
rect 25819 16491 25885 16492
rect 27110 16421 27170 20707
rect 27294 19413 27354 21115
rect 27475 20772 27541 20773
rect 27475 20708 27476 20772
rect 27540 20708 27541 20772
rect 27475 20707 27541 20708
rect 27291 19412 27357 19413
rect 27291 19348 27292 19412
rect 27356 19348 27357 19412
rect 27291 19347 27357 19348
rect 27107 16420 27173 16421
rect 27107 16356 27108 16420
rect 27172 16356 27173 16420
rect 27107 16355 27173 16356
rect 27478 15197 27538 20707
rect 28030 20637 28090 32131
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 28211 32060 28277 32061
rect 28211 31996 28212 32060
rect 28276 31996 28277 32060
rect 28211 31995 28277 31996
rect 28027 20636 28093 20637
rect 28027 20572 28028 20636
rect 28092 20572 28093 20636
rect 28027 20571 28093 20572
rect 27475 15196 27541 15197
rect 27475 15132 27476 15196
rect 27540 15132 27541 15196
rect 27475 15131 27541 15132
rect 28214 14109 28274 31995
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 33363 30700 33429 30701
rect 33363 30636 33364 30700
rect 33428 30636 33429 30700
rect 33363 30635 33429 30636
rect 29683 30564 29749 30565
rect 29683 30500 29684 30564
rect 29748 30500 29749 30564
rect 29683 30499 29749 30500
rect 28579 29068 28645 29069
rect 28579 29004 28580 29068
rect 28644 29004 28645 29068
rect 28579 29003 28645 29004
rect 28582 18053 28642 29003
rect 28947 28252 29013 28253
rect 28947 28188 28948 28252
rect 29012 28188 29013 28252
rect 28947 28187 29013 28188
rect 28763 24988 28829 24989
rect 28763 24924 28764 24988
rect 28828 24924 28829 24988
rect 28763 24923 28829 24924
rect 28766 18597 28826 24923
rect 28950 22405 29010 28187
rect 29315 23492 29381 23493
rect 29315 23428 29316 23492
rect 29380 23428 29381 23492
rect 29315 23427 29381 23428
rect 28947 22404 29013 22405
rect 28947 22340 28948 22404
rect 29012 22340 29013 22404
rect 28947 22339 29013 22340
rect 29318 20637 29378 23427
rect 29686 23221 29746 30499
rect 31523 29068 31589 29069
rect 31523 29004 31524 29068
rect 31588 29004 31589 29068
rect 31523 29003 31589 29004
rect 30787 26348 30853 26349
rect 30787 26284 30788 26348
rect 30852 26284 30853 26348
rect 30787 26283 30853 26284
rect 30051 24988 30117 24989
rect 30051 24924 30052 24988
rect 30116 24924 30117 24988
rect 30051 24923 30117 24924
rect 29683 23220 29749 23221
rect 29683 23156 29684 23220
rect 29748 23156 29749 23220
rect 29683 23155 29749 23156
rect 29315 20636 29381 20637
rect 29315 20572 29316 20636
rect 29380 20572 29381 20636
rect 29315 20571 29381 20572
rect 29315 20364 29381 20365
rect 29315 20300 29316 20364
rect 29380 20300 29381 20364
rect 29315 20299 29381 20300
rect 28947 20092 29013 20093
rect 28947 20028 28948 20092
rect 29012 20028 29013 20092
rect 28947 20027 29013 20028
rect 28763 18596 28829 18597
rect 28763 18532 28764 18596
rect 28828 18532 28829 18596
rect 28763 18531 28829 18532
rect 28579 18052 28645 18053
rect 28579 17988 28580 18052
rect 28644 17988 28645 18052
rect 28579 17987 28645 17988
rect 28950 17781 29010 20027
rect 29318 19549 29378 20299
rect 29315 19548 29381 19549
rect 29315 19484 29316 19548
rect 29380 19484 29381 19548
rect 29315 19483 29381 19484
rect 28947 17780 29013 17781
rect 28947 17716 28948 17780
rect 29012 17716 29013 17780
rect 28947 17715 29013 17716
rect 29318 15605 29378 19483
rect 29686 16013 29746 23155
rect 30054 17509 30114 24923
rect 30603 19684 30669 19685
rect 30603 19620 30604 19684
rect 30668 19620 30669 19684
rect 30603 19619 30669 19620
rect 30051 17508 30117 17509
rect 30051 17444 30052 17508
rect 30116 17444 30117 17508
rect 30051 17443 30117 17444
rect 29683 16012 29749 16013
rect 29683 15948 29684 16012
rect 29748 15948 29749 16012
rect 29683 15947 29749 15948
rect 29315 15604 29381 15605
rect 29315 15540 29316 15604
rect 29380 15540 29381 15604
rect 29315 15539 29381 15540
rect 30606 15061 30666 19619
rect 30790 19277 30850 26283
rect 30971 23764 31037 23765
rect 30971 23700 30972 23764
rect 31036 23700 31037 23764
rect 30971 23699 31037 23700
rect 30787 19276 30853 19277
rect 30787 19212 30788 19276
rect 30852 19212 30853 19276
rect 30787 19211 30853 19212
rect 30974 15197 31034 23699
rect 31155 22948 31221 22949
rect 31155 22884 31156 22948
rect 31220 22884 31221 22948
rect 31155 22883 31221 22884
rect 31158 19685 31218 22883
rect 31155 19684 31221 19685
rect 31155 19620 31156 19684
rect 31220 19620 31221 19684
rect 31155 19619 31221 19620
rect 30971 15196 31037 15197
rect 30971 15132 30972 15196
rect 31036 15132 31037 15196
rect 30971 15131 31037 15132
rect 30603 15060 30669 15061
rect 30603 14996 30604 15060
rect 30668 14996 30669 15060
rect 30603 14995 30669 14996
rect 31526 14789 31586 29003
rect 32259 28388 32325 28389
rect 32259 28324 32260 28388
rect 32324 28324 32325 28388
rect 32259 28323 32325 28324
rect 31891 23492 31957 23493
rect 31891 23428 31892 23492
rect 31956 23428 31957 23492
rect 31891 23427 31957 23428
rect 31894 17101 31954 23427
rect 32262 20637 32322 28323
rect 32811 27708 32877 27709
rect 32811 27644 32812 27708
rect 32876 27644 32877 27708
rect 32811 27643 32877 27644
rect 32443 26620 32509 26621
rect 32443 26556 32444 26620
rect 32508 26556 32509 26620
rect 32443 26555 32509 26556
rect 32446 21997 32506 26555
rect 32627 22268 32693 22269
rect 32627 22204 32628 22268
rect 32692 22204 32693 22268
rect 32627 22203 32693 22204
rect 32443 21996 32509 21997
rect 32443 21932 32444 21996
rect 32508 21932 32509 21996
rect 32443 21931 32509 21932
rect 32259 20636 32325 20637
rect 32259 20572 32260 20636
rect 32324 20572 32325 20636
rect 32259 20571 32325 20572
rect 32630 20501 32690 22203
rect 32627 20500 32693 20501
rect 32627 20436 32628 20500
rect 32692 20436 32693 20500
rect 32627 20435 32693 20436
rect 31891 17100 31957 17101
rect 31891 17036 31892 17100
rect 31956 17036 31957 17100
rect 31891 17035 31957 17036
rect 32814 16285 32874 27643
rect 32995 23492 33061 23493
rect 32995 23428 32996 23492
rect 33060 23428 33061 23492
rect 32995 23427 33061 23428
rect 32998 17781 33058 23427
rect 33366 22110 33426 30635
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34467 27708 34533 27709
rect 34467 27644 34468 27708
rect 34532 27644 34533 27708
rect 34467 27643 34533 27644
rect 34283 26756 34349 26757
rect 34283 26692 34284 26756
rect 34348 26692 34349 26756
rect 34283 26691 34349 26692
rect 33547 26076 33613 26077
rect 33547 26012 33548 26076
rect 33612 26012 33613 26076
rect 33547 26011 33613 26012
rect 33550 25669 33610 26011
rect 33547 25668 33613 25669
rect 33547 25604 33548 25668
rect 33612 25604 33613 25668
rect 33547 25603 33613 25604
rect 33182 22050 33426 22110
rect 33182 21725 33242 22050
rect 33179 21724 33245 21725
rect 33179 21660 33180 21724
rect 33244 21660 33245 21724
rect 33179 21659 33245 21660
rect 32995 17780 33061 17781
rect 32995 17716 32996 17780
rect 33060 17716 33061 17780
rect 32995 17715 33061 17716
rect 32811 16284 32877 16285
rect 32811 16220 32812 16284
rect 32876 16220 32877 16284
rect 32811 16219 32877 16220
rect 32998 15877 33058 17715
rect 33550 16829 33610 25603
rect 34099 24988 34165 24989
rect 34099 24924 34100 24988
rect 34164 24924 34165 24988
rect 34099 24923 34165 24924
rect 34102 19821 34162 24923
rect 34286 23221 34346 26691
rect 34470 24037 34530 27643
rect 34651 27164 34717 27165
rect 34651 27100 34652 27164
rect 34716 27100 34717 27164
rect 34651 27099 34717 27100
rect 34654 24037 34714 27099
rect 34928 26688 35248 27712
rect 35588 37024 35908 37584
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 35936 35908 36960
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 36123 29204 36189 29205
rect 36123 29140 36124 29204
rect 36188 29140 36189 29204
rect 36123 29139 36189 29140
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35387 27708 35453 27709
rect 35387 27644 35388 27708
rect 35452 27644 35453 27708
rect 35387 27643 35453 27644
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34467 24036 34533 24037
rect 34467 23972 34468 24036
rect 34532 23972 34533 24036
rect 34467 23971 34533 23972
rect 34651 24036 34717 24037
rect 34651 23972 34652 24036
rect 34716 23972 34717 24036
rect 34651 23971 34717 23972
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34283 23220 34349 23221
rect 34283 23156 34284 23220
rect 34348 23156 34349 23220
rect 34283 23155 34349 23156
rect 34928 22336 35248 23360
rect 35390 23085 35450 27643
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35387 23084 35453 23085
rect 35387 23020 35388 23084
rect 35452 23020 35453 23084
rect 35387 23019 35453 23020
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34651 21996 34717 21997
rect 34651 21932 34652 21996
rect 34716 21932 34717 21996
rect 34651 21931 34717 21932
rect 34654 19821 34714 21931
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34099 19820 34165 19821
rect 34099 19756 34100 19820
rect 34164 19756 34165 19820
rect 34099 19755 34165 19756
rect 34651 19820 34717 19821
rect 34651 19756 34652 19820
rect 34716 19756 34717 19820
rect 34651 19755 34717 19756
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 33547 16828 33613 16829
rect 33547 16764 33548 16828
rect 33612 16764 33613 16828
rect 33547 16763 33613 16764
rect 32995 15876 33061 15877
rect 32995 15812 32996 15876
rect 33060 15812 33061 15876
rect 32995 15811 33061 15812
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 31523 14788 31589 14789
rect 31523 14724 31524 14788
rect 31588 14724 31589 14788
rect 31523 14723 31589 14724
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 28211 14108 28277 14109
rect 28211 14044 28212 14108
rect 28276 14044 28277 14108
rect 28211 14043 28277 14044
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 25635 13020 25701 13021
rect 25635 12956 25636 13020
rect 25700 12956 25701 13020
rect 25635 12955 25701 12956
rect 17907 12748 17973 12749
rect 17907 12684 17908 12748
rect 17972 12684 17973 12748
rect 17907 12683 17973 12684
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 15515 12204 15581 12205
rect 15515 12140 15516 12204
rect 15580 12140 15581 12204
rect 15515 12139 15581 12140
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 8707 10980 8773 10981
rect 8707 10916 8708 10980
rect 8772 10916 8773 10980
rect 8707 10915 8773 10916
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 36126 15061 36186 29139
rect 37227 27572 37293 27573
rect 37227 27508 37228 27572
rect 37292 27508 37293 27572
rect 37227 27507 37293 27508
rect 36307 26076 36373 26077
rect 36307 26012 36308 26076
rect 36372 26012 36373 26076
rect 36307 26011 36373 26012
rect 36310 21997 36370 26011
rect 37230 23765 37290 27507
rect 37227 23764 37293 23765
rect 37227 23700 37228 23764
rect 37292 23700 37293 23764
rect 37227 23699 37293 23700
rect 36307 21996 36373 21997
rect 36307 21932 36308 21996
rect 36372 21932 36373 21996
rect 36307 21931 36373 21932
rect 36123 15060 36189 15061
rect 36123 14996 36124 15060
rect 36188 14996 36189 15060
rect 36123 14995 36189 14996
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 5472 35908 6496
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1
transform -1 0 38732 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _0715_
timestamp 1
transform 1 0 4600 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _0716_
timestamp 1
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0717_
timestamp 1
transform 1 0 5244 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_1  _0718_
timestamp 1
transform -1 0 8280 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0719_
timestamp 1
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0720_
timestamp 1
transform 1 0 3772 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _0721_
timestamp 1
transform 1 0 2576 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0722_
timestamp 1
transform -1 0 15732 0 -1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__and4_1  _0723_
timestamp 1
transform 1 0 3036 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0724_
timestamp 1
transform -1 0 6992 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0725_
timestamp 1
transform -1 0 4416 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0726_
timestamp 1
transform -1 0 6256 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0727_
timestamp 1
transform 1 0 12972 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0728_
timestamp 1
transform 1 0 5244 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _0729_
timestamp 1
transform 1 0 8188 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_2  _0730_
timestamp 1
transform -1 0 15180 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0731_
timestamp 1
transform 1 0 28980 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0732_
timestamp 1
transform 1 0 9108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0733_
timestamp 1
transform 1 0 18492 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0734_
timestamp 1
transform 1 0 6808 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0735_
timestamp 1
transform 1 0 4416 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0736_
timestamp 1
transform 1 0 9476 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0737_
timestamp 1
transform 1 0 19412 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0738_
timestamp 1
transform 1 0 7544 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _0739_
timestamp 1
transform 1 0 7452 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0740_
timestamp 1
transform 1 0 14812 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0741_
timestamp 1
transform 1 0 8188 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0742_
timestamp 1
transform 1 0 1564 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0743_
timestamp 1
transform 1 0 1932 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0744_
timestamp 1
transform 1 0 12328 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0745_
timestamp 1
transform 1 0 20976 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0746_
timestamp 1
transform 1 0 7912 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0747_
timestamp 1
transform 1 0 7912 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _0748_
timestamp 1
transform 1 0 9936 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_1  _0749_
timestamp 1
transform 1 0 1656 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0750_
timestamp 1
transform 1 0 2300 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _0751_
timestamp 1
transform 1 0 10304 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0752_
timestamp 1
transform 1 0 10028 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0753_
timestamp 1
transform 1 0 23552 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _0754_
timestamp 1
transform 1 0 4232 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__nor4b_1  _0755_
timestamp 1
transform -1 0 2484 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0756_
timestamp 1
transform 1 0 1656 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_2  _0757_
timestamp 1
transform -1 0 5428 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0758_
timestamp 1
transform 1 0 5612 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0759_
timestamp 1
transform 1 0 7544 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0760_
timestamp 1
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0761_
timestamp 1
transform 1 0 2116 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0762_
timestamp 1
transform 1 0 6624 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0763_
timestamp 1
transform 1 0 7084 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0764_
timestamp 1
transform 1 0 7084 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0765_
timestamp 1
transform 1 0 4784 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0766_
timestamp 1
transform -1 0 3588 0 -1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0767_
timestamp 1
transform 1 0 2944 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0768_
timestamp 1
transform 1 0 5704 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0769_
timestamp 1
transform 1 0 2760 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nor4b_1  _0770_
timestamp 1
transform -1 0 3128 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0771_
timestamp 1
transform 1 0 11592 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0772_
timestamp 1
transform 1 0 5428 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0773_
timestamp 1
transform -1 0 16560 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0774_
timestamp 1
transform 1 0 5060 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _0775_
timestamp 1
transform -1 0 6808 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0776_
timestamp 1
transform 1 0 6348 0 -1 16320
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0777_
timestamp 1
transform -1 0 4600 0 -1 16320
box -38 -48 1326 592
use sky130_fd_sc_hd__and4bb_1  _0778_
timestamp 1
transform 1 0 6164 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nor4b_1  _0779_
timestamp 1
transform -1 0 6164 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0780_
timestamp 1
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_2  _0781_
timestamp 1
transform 1 0 8004 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _0782_
timestamp 1
transform 1 0 17112 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0783_
timestamp 1
transform 1 0 28336 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0784_
timestamp 1
transform 1 0 6072 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0785_
timestamp 1
transform 1 0 33488 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0786_
timestamp 1
transform 1 0 16100 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0787_
timestamp 1
transform 1 0 28244 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0788_
timestamp 1
transform 1 0 8832 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0789_
timestamp 1
transform 1 0 9108 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0790_
timestamp 1
transform -1 0 10304 0 -1 16320
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_2  _0791_
timestamp 1
transform 1 0 15732 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0792_
timestamp 1
transform -1 0 30912 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0793_
timestamp 1
transform 1 0 15732 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0794_
timestamp 1
transform -1 0 12512 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0795_
timestamp 1
transform 1 0 23000 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0796_
timestamp 1
transform 1 0 6348 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0797_
timestamp 1
transform 1 0 5152 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0798_
timestamp 1
transform 1 0 5428 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0799_
timestamp 1
transform 1 0 16560 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0800_
timestamp 1
transform 1 0 16100 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_2  _0801_
timestamp 1
transform -1 0 14812 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0802_
timestamp 1
transform -1 0 11408 0 -1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_2  _0803_
timestamp 1
transform 1 0 13708 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0804_
timestamp 1
transform 1 0 29440 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_4  _0805_
timestamp 1
transform 1 0 7728 0 -1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0806_
timestamp 1
transform -1 0 8740 0 1 11968
box -38 -48 1326 592
use sky130_fd_sc_hd__o21ba_2  _0807_
timestamp 1
transform 1 0 14628 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0808_
timestamp 1
transform -1 0 31740 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0809_
timestamp 1
transform -1 0 24012 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0810_
timestamp 1
transform 1 0 14536 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0811_
timestamp 1
transform 1 0 10028 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0812_
timestamp 1
transform 1 0 18768 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0813_
timestamp 1
transform 1 0 18032 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0814_
timestamp 1
transform -1 0 23552 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0815_
timestamp 1
transform 1 0 11224 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0816_
timestamp 1
transform 1 0 20516 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0817_
timestamp 1
transform 1 0 13800 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0818_
timestamp 1
transform 1 0 15732 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _0819_
timestamp 1
transform 1 0 7912 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0820_
timestamp 1
transform 1 0 8464 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0821_
timestamp 1
transform 1 0 17020 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0822_
timestamp 1
transform 1 0 11868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0823_
timestamp 1
transform 1 0 3864 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0824_
timestamp 1
transform 1 0 30912 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0825_
timestamp 1
transform 1 0 8096 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0826_
timestamp 1
transform 1 0 12512 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0827_
timestamp 1
transform 1 0 18676 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0828_
timestamp 1
transform 1 0 17388 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0829_
timestamp 1
transform 1 0 12328 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0830_
timestamp 1
transform -1 0 5612 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0831_
timestamp 1
transform 1 0 9200 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_2  _0832_
timestamp 1
transform -1 0 10212 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0833_
timestamp 1
transform 1 0 9292 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0834_
timestamp 1
transform 1 0 15364 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0835_
timestamp 1
transform 1 0 10120 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0836_
timestamp 1
transform -1 0 10672 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0837_
timestamp 1
transform 1 0 12972 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0838_
timestamp 1
transform 1 0 11776 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0839_
timestamp 1
transform 1 0 13064 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0840_
timestamp 1
transform -1 0 23828 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0841_
timestamp 1
transform 1 0 12236 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0842_
timestamp 1
transform 1 0 14444 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0843_
timestamp 1
transform 1 0 15456 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0844_
timestamp 1
transform 1 0 9936 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0845_
timestamp 1
transform 1 0 9200 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0846_
timestamp 1
transform 1 0 18124 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0847_
timestamp 1
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0848_
timestamp 1
transform -1 0 14812 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0849_
timestamp 1
transform 1 0 12880 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0850_
timestamp 1
transform 1 0 10856 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0851_
timestamp 1
transform 1 0 14444 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0852_
timestamp 1
transform 1 0 19228 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0853_
timestamp 1
transform 1 0 23552 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0854_
timestamp 1
transform -1 0 24380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0855_
timestamp 1
transform 1 0 22264 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0856_
timestamp 1
transform 1 0 22724 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0857_
timestamp 1
transform 1 0 28336 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0858_
timestamp 1
transform -1 0 26864 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0859_
timestamp 1
transform 1 0 25300 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0860_
timestamp 1
transform 1 0 26220 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0861_
timestamp 1
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0862_
timestamp 1
transform 1 0 27692 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0863_
timestamp 1
transform 1 0 23828 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_4  _0864_
timestamp 1
transform 1 0 11500 0 -1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_2  _0865_
timestamp 1
transform 1 0 6808 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0866_
timestamp 1
transform 1 0 25024 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0867_
timestamp 1
transform 1 0 25392 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0868_
timestamp 1
transform 1 0 2668 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0869_
timestamp 1
transform 1 0 14720 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0870_
timestamp 1
transform 1 0 15640 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0871_
timestamp 1
transform 1 0 28060 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_4  _0872_
timestamp 1
transform -1 0 7176 0 1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_1  _0873_
timestamp 1
transform 1 0 13984 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_4  _0874_
timestamp 1
transform -1 0 7268 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_2  _0875_
timestamp 1
transform 1 0 6164 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0876_
timestamp 1
transform 1 0 32292 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0877_
timestamp 1
transform -1 0 29440 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0878_
timestamp 1
transform 1 0 2208 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0879_
timestamp 1
transform 1 0 18308 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0880_
timestamp 1
transform 1 0 18032 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0881_
timestamp 1
transform 1 0 27968 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0882_
timestamp 1
transform 1 0 17112 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0883_
timestamp 1
transform -1 0 31372 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0884_
timestamp 1
transform -1 0 31188 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0885_
timestamp 1
transform 1 0 31004 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0886_
timestamp 1
transform 1 0 16836 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0887_
timestamp 1
transform 1 0 13248 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0888_
timestamp 1
transform 1 0 25944 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0889_
timestamp 1
transform 1 0 15916 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0890_
timestamp 1
transform 1 0 26680 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0891_
timestamp 1
transform 1 0 31556 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0892_
timestamp 1
transform 1 0 36340 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0893_
timestamp 1
transform -1 0 5152 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0894_
timestamp 1
transform 1 0 4140 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0895_
timestamp 1
transform 1 0 5152 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0896_
timestamp 1
transform 1 0 7820 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0897_
timestamp 1
transform 1 0 5796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0898_
timestamp 1
transform 1 0 5060 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0899_
timestamp 1
transform 1 0 8372 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0900_
timestamp 1
transform 1 0 12236 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0901_
timestamp 1
transform 1 0 31004 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0902_
timestamp 1
transform -1 0 13892 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0903_
timestamp 1
transform 1 0 35420 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0904_
timestamp 1
transform 1 0 7268 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0905_
timestamp 1
transform 1 0 6440 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0906_
timestamp 1
transform 1 0 28336 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0907_
timestamp 1
transform -1 0 29164 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0908_
timestamp 1
transform 1 0 8004 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0909_
timestamp 1
transform 1 0 28520 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0910_
timestamp 1
transform 1 0 11684 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0911_
timestamp 1
transform -1 0 7544 0 1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_1  _0912_
timestamp 1
transform -1 0 29900 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0913_
timestamp 1
transform 1 0 13248 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0914_
timestamp 1
transform 1 0 29900 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0915_
timestamp 1
transform 1 0 37076 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0916_
timestamp 1
transform 1 0 18400 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0917_
timestamp 1
transform -1 0 35880 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0918_
timestamp 1
transform 1 0 14628 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0919_
timestamp 1
transform -1 0 25760 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0920_
timestamp 1
transform 1 0 10304 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0921_
timestamp 1
transform 1 0 17480 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0922_
timestamp 1
transform 1 0 11592 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0923_
timestamp 1
transform 1 0 21436 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0924_
timestamp 1
transform -1 0 22908 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_2  _0925_
timestamp 1
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0926_
timestamp 1
transform -1 0 11960 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0927_
timestamp 1
transform 1 0 9844 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0928_
timestamp 1
transform 1 0 18216 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_4  _0929_
timestamp 1
transform -1 0 10488 0 1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0930_
timestamp 1
transform -1 0 11132 0 1 16320
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_1  _0931_
timestamp 1
transform -1 0 15548 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0932_
timestamp 1
transform 1 0 10488 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0933_
timestamp 1
transform 1 0 9200 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0934_
timestamp 1
transform 1 0 22908 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0935_
timestamp 1
transform 1 0 22816 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0936_
timestamp 1
transform -1 0 10120 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0937_
timestamp 1
transform 1 0 9200 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0938_
timestamp 1
transform 1 0 17020 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0939_
timestamp 1
transform 1 0 10120 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0940_
timestamp 1
transform 1 0 14720 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0941_
timestamp 1
transform 1 0 21160 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0942_
timestamp 1
transform 1 0 21436 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0943_
timestamp 1
transform 1 0 20884 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0944_
timestamp 1
transform 1 0 9936 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_2  _0945_
timestamp 1
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0946_
timestamp 1
transform 1 0 34316 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0947_
timestamp 1
transform 1 0 10672 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0948_
timestamp 1
transform 1 0 10212 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0949_
timestamp 1
transform 1 0 20884 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0950_
timestamp 1
transform -1 0 32568 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0951_
timestamp 1
transform -1 0 22356 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_4  _0952_
timestamp 1
transform 1 0 10488 0 1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_2  _0953_
timestamp 1
transform 1 0 17664 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0954_
timestamp 1
transform -1 0 29348 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0955_
timestamp 1
transform 1 0 19320 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0956_
timestamp 1
transform 1 0 8096 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0957_
timestamp 1
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0958_
timestamp 1
transform 1 0 14720 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0959_
timestamp 1
transform 1 0 20424 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0960_
timestamp 1
transform -1 0 17204 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0961_
timestamp 1
transform 1 0 8924 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0962_
timestamp 1
transform 1 0 18584 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0963_
timestamp 1
transform 1 0 21528 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0964_
timestamp 1
transform 1 0 11500 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0965_
timestamp 1
transform 1 0 22172 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0966_
timestamp 1
transform 1 0 12512 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0967_
timestamp 1
transform -1 0 12512 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0968_
timestamp 1
transform 1 0 26312 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0969_
timestamp 1
transform 1 0 26036 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0970_
timestamp 1
transform 1 0 12696 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0971_
timestamp 1
transform 1 0 13708 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0972_
timestamp 1
transform 1 0 14076 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0973_
timestamp 1
transform 1 0 14904 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0974_
timestamp 1
transform 1 0 12236 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0975_
timestamp 1
transform 1 0 22816 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0976_
timestamp 1
transform 1 0 23368 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0977_
timestamp 1
transform 1 0 34500 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0978_
timestamp 1
transform 1 0 9384 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0979_
timestamp 1
transform 1 0 14352 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0980_
timestamp 1
transform -1 0 29992 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0981_
timestamp 1
transform 1 0 29532 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0982_
timestamp 1
transform -1 0 9752 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0983_
timestamp 1
transform 1 0 26956 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0984_
timestamp 1
transform 1 0 19504 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0985_
timestamp 1
transform 1 0 12512 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0986_
timestamp 1
transform 1 0 26404 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0987_
timestamp 1
transform 1 0 34040 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0988_
timestamp 1
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0989_
timestamp 1
transform -1 0 27508 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0990_
timestamp 1
transform 1 0 10672 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0991_
timestamp 1
transform 1 0 20700 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0992_
timestamp 1
transform -1 0 20424 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0993_
timestamp 1
transform 1 0 18676 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0994_
timestamp 1
transform 1 0 21804 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0995_
timestamp 1
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0996_
timestamp 1
transform 1 0 20884 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0997_
timestamp 1
transform 1 0 21344 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0998_
timestamp 1
transform 1 0 15916 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0999_
timestamp 1
transform -1 0 27784 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_2  _1000_
timestamp 1
transform 1 0 14536 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1001_
timestamp 1
transform 1 0 26312 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1002_
timestamp 1
transform 1 0 31464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _1003_
timestamp 1
transform 1 0 14076 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1004_
timestamp 1
transform 1 0 37260 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _1005_
timestamp 1
transform 1 0 2576 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1006_
timestamp 1
transform 1 0 4692 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1007_
timestamp 1
transform 1 0 33672 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1008_
timestamp 1
transform 1 0 34960 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1009_
timestamp 1
transform 1 0 32292 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1010_
timestamp 1
transform 1 0 33580 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1011_
timestamp 1
transform 1 0 34684 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _1012_
timestamp 1
transform 1 0 37352 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1013_
timestamp 1
transform 1 0 37352 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1014_
timestamp 1
transform 1 0 38640 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1015_
timestamp 1
transform -1 0 33028 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1016_
timestamp 1
transform -1 0 32016 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1017_
timestamp 1
transform 1 0 22356 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1018_
timestamp 1
transform 1 0 19780 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1019_
timestamp 1
transform 1 0 22080 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1020_
timestamp 1
transform 1 0 22632 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1021_
timestamp 1
transform 1 0 18584 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1022_
timestamp 1
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1
transform 1 0 31188 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1024_
timestamp 1
transform 1 0 31096 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1025_
timestamp 1
transform 1 0 30820 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1026_
timestamp 1
transform 1 0 14904 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1027_
timestamp 1
transform 1 0 13984 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1028_
timestamp 1
transform 1 0 14812 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1029_
timestamp 1
transform 1 0 9936 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1030_
timestamp 1
transform 1 0 10488 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1031_
timestamp 1
transform -1 0 16100 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1032_
timestamp 1
transform 1 0 15180 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1033_
timestamp 1
transform 1 0 31464 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1034_
timestamp 1
transform 1 0 41584 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1035_
timestamp 1
transform 1 0 23276 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1036_
timestamp 1
transform -1 0 25760 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1037_
timestamp 1
transform 1 0 23368 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1038_
timestamp 1
transform -1 0 13616 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1039_
timestamp 1
transform 1 0 25668 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1040_
timestamp 1
transform 1 0 26128 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1041_
timestamp 1
transform 1 0 26956 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1042_
timestamp 1
transform 1 0 12972 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1043_
timestamp 1
transform 1 0 20608 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1044_
timestamp 1
transform 1 0 21804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1045_
timestamp 1
transform 1 0 5060 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1046_
timestamp 1
transform 1 0 28520 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1047_
timestamp 1
transform -1 0 28980 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1048_
timestamp 1
transform -1 0 24840 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1049_
timestamp 1
transform 1 0 9844 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1050_
timestamp 1
transform 1 0 13156 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1051_
timestamp 1
transform 1 0 26956 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1052_
timestamp 1
transform 1 0 24472 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1053_
timestamp 1
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1054_
timestamp 1
transform 1 0 24380 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1055_
timestamp 1
transform 1 0 24380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1056_
timestamp 1
transform 1 0 26956 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1057_
timestamp 1
transform 1 0 27692 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1058_
timestamp 1
transform -1 0 11408 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1059_
timestamp 1
transform -1 0 18216 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1060_
timestamp 1
transform 1 0 32108 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1061_
timestamp 1
transform 1 0 27968 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1062_
timestamp 1
transform 1 0 29348 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1063_
timestamp 1
transform 1 0 13156 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1064_
timestamp 1
transform 1 0 18676 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1065_
timestamp 1
transform 1 0 19320 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1066_
timestamp 1
transform 1 0 14720 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1067_
timestamp 1
transform 1 0 11960 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1068_
timestamp 1
transform 1 0 13524 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1069_
timestamp 1
transform 1 0 37260 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1070_
timestamp 1
transform -1 0 24012 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1071_
timestamp 1
transform -1 0 22540 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1072_
timestamp 1
transform 1 0 14628 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1073_
timestamp 1
transform 1 0 13064 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1074_
timestamp 1
transform -1 0 22724 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1075_
timestamp 1
transform 1 0 21896 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1076_
timestamp 1
transform -1 0 23368 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1077_
timestamp 1
transform 1 0 22816 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1078_
timestamp 1
transform 1 0 31740 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1079_
timestamp 1
transform 1 0 21896 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1080_
timestamp 1
transform -1 0 23552 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1081_
timestamp 1
transform 1 0 16100 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1082_
timestamp 1
transform 1 0 19228 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1083_
timestamp 1
transform -1 0 32016 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1084_
timestamp 1
transform 1 0 20240 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1085_
timestamp 1
transform 1 0 24288 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1086_
timestamp 1
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1087_
timestamp 1
transform 1 0 24472 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1088_
timestamp 1
transform 1 0 16928 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1089_
timestamp 1
transform -1 0 18952 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1090_
timestamp 1
transform 1 0 16008 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1091_
timestamp 1
transform 1 0 17020 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1092_
timestamp 1
transform 1 0 16744 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1093_
timestamp 1
transform 1 0 17296 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1094_
timestamp 1
transform -1 0 30084 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1095_
timestamp 1
transform 1 0 23920 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1096_
timestamp 1
transform 1 0 24472 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1097_
timestamp 1
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1098_
timestamp 1
transform -1 0 25760 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1099_
timestamp 1
transform 1 0 31372 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1100_
timestamp 1
transform 1 0 37260 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1101_
timestamp 1
transform 1 0 26680 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1102_
timestamp 1
transform -1 0 10856 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1103_
timestamp 1
transform 1 0 17848 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1104_
timestamp 1
transform 1 0 35788 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1105_
timestamp 1
transform 1 0 31280 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1106_
timestamp 1
transform 1 0 37904 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1107_
timestamp 1
transform 1 0 36524 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1108_
timestamp 1
transform 1 0 38364 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1109_
timestamp 1
transform -1 0 13432 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1110_
timestamp 1
transform -1 0 16192 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1111_
timestamp 1
transform -1 0 11500 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1112_
timestamp 1
transform 1 0 10948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1113_
timestamp 1
transform 1 0 13156 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1114_
timestamp 1
transform 1 0 37904 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1115_
timestamp 1
transform 1 0 38180 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1116_
timestamp 1
transform 1 0 39008 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1117_
timestamp 1
transform 1 0 43332 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1118_
timestamp 1
transform -1 0 26864 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1119_
timestamp 1
transform 1 0 25852 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1120_
timestamp 1
transform 1 0 34408 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1121_
timestamp 1
transform 1 0 32660 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1122_
timestamp 1
transform 1 0 34684 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1123_
timestamp 1
transform 1 0 27784 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1124_
timestamp 1
transform 1 0 34408 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1
transform 1 0 20424 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1126_
timestamp 1
transform 1 0 17756 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1127_
timestamp 1
transform 1 0 19136 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1128_
timestamp 1
transform -1 0 6256 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1129_
timestamp 1
transform 1 0 20056 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1
transform 1 0 20240 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1131_
timestamp 1
transform 1 0 19780 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1132_
timestamp 1
transform 1 0 8464 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1133_
timestamp 1
transform 1 0 7728 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1134_
timestamp 1
transform 1 0 8924 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1135_
timestamp 1
transform 1 0 20332 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1136_
timestamp 1
transform -1 0 20976 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1137_
timestamp 1
transform 1 0 20424 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1138_
timestamp 1
transform -1 0 41768 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1139_
timestamp 1
transform 1 0 34960 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1140_
timestamp 1
transform 1 0 35144 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1141_
timestamp 1
transform 1 0 32844 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1142_
timestamp 1
transform 1 0 28336 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1143_
timestamp 1
transform 1 0 31096 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1144_
timestamp 1
transform -1 0 18676 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1145_
timestamp 1
transform 1 0 18400 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1146_
timestamp 1
transform -1 0 34040 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1147_
timestamp 1
transform 1 0 17204 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1148_
timestamp 1
transform 1 0 35052 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1149_
timestamp 1
transform 1 0 33672 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1150_
timestamp 1
transform 1 0 35604 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1151_
timestamp 1
transform 1 0 33764 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1152_
timestamp 1
transform 1 0 23276 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1153_
timestamp 1
transform 1 0 22540 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1154_
timestamp 1
transform 1 0 12144 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1155_
timestamp 1
transform 1 0 12880 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1156_
timestamp 1
transform 1 0 23828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1157_
timestamp 1
transform 1 0 34776 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1158_
timestamp 1
transform 1 0 41584 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1159_
timestamp 1
transform 1 0 19228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1160_
timestamp 1
transform 1 0 23276 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1161_
timestamp 1
transform 1 0 23736 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _1162_
timestamp 1
transform 1 0 6348 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1163_
timestamp 1
transform 1 0 27600 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1164_
timestamp 1
transform 1 0 28336 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 1
transform 1 0 28796 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1166_
timestamp 1
transform 1 0 29900 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1167_
timestamp 1
transform 1 0 17204 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1168_
timestamp 1
transform 1 0 29992 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1169_
timestamp 1
transform 1 0 30452 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1170_
timestamp 1
transform 1 0 30728 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1171_
timestamp 1
transform 1 0 30912 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1172_
timestamp 1
transform -1 0 31556 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1173_
timestamp 1
transform 1 0 29532 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1174_
timestamp 1
transform 1 0 15732 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1175_
timestamp 1
transform 1 0 19596 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1176_
timestamp 1
transform -1 0 12236 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1177_
timestamp 1
transform 1 0 28060 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1178_
timestamp 1
transform -1 0 26496 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1179_
timestamp 1
transform -1 0 8004 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1180_
timestamp 1
transform 1 0 7636 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1181_
timestamp 1
transform 1 0 15824 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1182_
timestamp 1
transform -1 0 35052 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1183_
timestamp 1
transform -1 0 5796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1184_
timestamp 1
transform 1 0 6348 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1185_
timestamp 1
transform -1 0 23460 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1186_
timestamp 1
transform 1 0 21436 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1187_
timestamp 1
transform 1 0 21804 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1188_
timestamp 1
transform -1 0 22908 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1189_
timestamp 1
transform 1 0 32844 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1190_
timestamp 1
transform 1 0 26312 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1191_
timestamp 1
transform 1 0 8004 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1192_
timestamp 1
transform 1 0 20056 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1193_
timestamp 1
transform -1 0 27048 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1194_
timestamp 1
transform 1 0 26956 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1195_
timestamp 1
transform 1 0 25760 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1196_
timestamp 1
transform 1 0 37260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1197_
timestamp 1
transform 1 0 36432 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1198_
timestamp 1
transform -1 0 37628 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1199_
timestamp 1
transform -1 0 27968 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1200_
timestamp 1
transform -1 0 26496 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1201_
timestamp 1
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1202_
timestamp 1
transform 1 0 19780 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1203_
timestamp 1
transform -1 0 29348 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1204_
timestamp 1
transform 1 0 26036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1205_
timestamp 1
transform 1 0 26128 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1206_
timestamp 1
transform 1 0 19596 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1207_
timestamp 1
transform 1 0 13064 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1208_
timestamp 1
transform 1 0 16100 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1209_
timestamp 1
transform -1 0 32568 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1210_
timestamp 1
transform -1 0 31556 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1211_
timestamp 1
transform -1 0 22632 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1212_
timestamp 1
transform 1 0 10580 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1213_
timestamp 1
transform -1 0 22264 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1214_
timestamp 1
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1215_
timestamp 1
transform 1 0 21712 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1216_
timestamp 1
transform 1 0 31556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1217_
timestamp 1
transform 1 0 29532 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1218_
timestamp 1
transform 1 0 31004 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1219_
timestamp 1
transform 1 0 32108 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1220_
timestamp 1
transform 1 0 39560 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1221_
timestamp 1
transform -1 0 33764 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1222_
timestamp 1
transform 1 0 25852 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1223_
timestamp 1
transform 1 0 30636 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1224_
timestamp 1
transform 1 0 31556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1225_
timestamp 1
transform 1 0 17664 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1226_
timestamp 1
transform 1 0 19688 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1227_
timestamp 1
transform -1 0 35788 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1228_
timestamp 1
transform -1 0 33488 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1229_
timestamp 1
transform 1 0 32844 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1230_
timestamp 1
transform 1 0 33028 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1231_
timestamp 1
transform 1 0 40296 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1232_
timestamp 1
transform -1 0 30084 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1233_
timestamp 1
transform 1 0 29716 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1234_
timestamp 1
transform 1 0 14444 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1235_
timestamp 1
transform 1 0 20516 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1236_
timestamp 1
transform -1 0 23828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1237_
timestamp 1
transform 1 0 24380 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1238_
timestamp 1
transform 1 0 38364 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1239_
timestamp 1
transform 1 0 37168 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1240_
timestamp 1
transform 1 0 39100 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1241_
timestamp 1
transform 1 0 18584 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1242_
timestamp 1
transform 1 0 14536 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1243_
timestamp 1
transform 1 0 14628 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1244_
timestamp 1
transform 1 0 15180 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1245_
timestamp 1
transform 1 0 19320 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1246_
timestamp 1
transform 1 0 40388 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1247_
timestamp 1
transform 1 0 28980 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1248_
timestamp 1
transform 1 0 33212 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1249_
timestamp 1
transform 1 0 28888 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1250_
timestamp 1
transform 1 0 33028 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1251_
timestamp 1
transform 1 0 28612 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1252_
timestamp 1
transform 1 0 29072 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1253_
timestamp 1
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1254_
timestamp 1
transform 1 0 33304 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1255_
timestamp 1
transform 1 0 34040 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1256_
timestamp 1
transform 1 0 34684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1257_
timestamp 1
transform 1 0 38456 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1258_
timestamp 1
transform 1 0 26496 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1259_
timestamp 1
transform 1 0 6900 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1260_
timestamp 1
transform -1 0 9384 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1261_
timestamp 1
transform 1 0 7176 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1262_
timestamp 1
transform 1 0 26680 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1263_
timestamp 1
transform 1 0 25760 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1264_
timestamp 1
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1265_
timestamp 1
transform 1 0 24012 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1266_
timestamp 1
transform 1 0 17204 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1267_
timestamp 1
transform -1 0 27048 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1268_
timestamp 1
transform -1 0 26588 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1269_
timestamp 1
transform 1 0 26036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1270_
timestamp 1
transform 1 0 27324 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1271_
timestamp 1
transform 1 0 27692 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1272_
timestamp 1
transform 1 0 22540 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1273_
timestamp 1
transform -1 0 37260 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1274_
timestamp 1
transform 1 0 11500 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1275_
timestamp 1
transform 1 0 33672 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1276_
timestamp 1
transform 1 0 34040 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1277_
timestamp 1
transform -1 0 19688 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1278_
timestamp 1
transform 1 0 17848 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1279_
timestamp 1
transform 1 0 17388 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1280_
timestamp 1
transform 1 0 18032 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1281_
timestamp 1
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1282_
timestamp 1
transform 1 0 34500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1283_
timestamp 1
transform -1 0 42320 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1284_
timestamp 1
transform 1 0 29532 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1285_
timestamp 1
transform 1 0 29532 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1286_
timestamp 1
transform 1 0 24380 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1287_
timestamp 1
transform -1 0 29532 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1288_
timestamp 1
transform 1 0 26956 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1289_
timestamp 1
transform 1 0 27692 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1290_
timestamp 1
transform 1 0 19044 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1291_
timestamp 1
transform -1 0 26312 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1292_
timestamp 1
transform 1 0 24564 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1293_
timestamp 1
transform 1 0 18584 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1294_
timestamp 1
transform 1 0 27508 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1295_
timestamp 1
transform 1 0 27784 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1296_
timestamp 1
transform 1 0 28428 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1297_
timestamp 1
transform -1 0 41492 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _1298_
timestamp 1
transform 1 0 17756 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1299_
timestamp 1
transform 1 0 25576 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1300_
timestamp 1
transform 1 0 15364 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1301_
timestamp 1
transform 1 0 20056 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1302_
timestamp 1
transform 1 0 20884 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1303_
timestamp 1
transform 1 0 24748 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1304_
timestamp 1
transform 1 0 17664 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1305_
timestamp 1
transform 1 0 24840 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1306_
timestamp 1
transform 1 0 31188 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1307_
timestamp 1
transform 1 0 37260 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1308_
timestamp 1
transform 1 0 38456 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1309_
timestamp 1
transform 1 0 40112 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1310_
timestamp 1
transform 1 0 22448 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1311_
timestamp 1
transform -1 0 17112 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1312_
timestamp 1
transform 1 0 16652 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1313_
timestamp 1
transform 1 0 22816 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1314_
timestamp 1
transform 1 0 22816 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1315_
timestamp 1
transform -1 0 36248 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1316_
timestamp 1
transform -1 0 24012 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1317_
timestamp 1
transform -1 0 24288 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1318_
timestamp 1
transform 1 0 23092 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1319_
timestamp 1
transform 1 0 23644 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1320_
timestamp 1
transform 1 0 32752 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1321_
timestamp 1
transform 1 0 34684 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1322_
timestamp 1
transform 1 0 34868 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1323_
timestamp 1
transform 1 0 35236 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1324_
timestamp 1
transform 1 0 35512 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1325_
timestamp 1
transform 1 0 33488 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1326_
timestamp 1
transform -1 0 37076 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1327_
timestamp 1
transform 1 0 34960 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1328_
timestamp 1
transform 1 0 35972 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1329_
timestamp 1
transform 1 0 36248 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1330_
timestamp 1
transform 1 0 43148 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1331_
timestamp 1
transform -1 0 34500 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1332_
timestamp 1
transform 1 0 24840 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1333_
timestamp 1
transform 1 0 26312 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1334_
timestamp 1
transform 1 0 26956 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1335_
timestamp 1
transform 1 0 10028 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1336_
timestamp 1
transform 1 0 31648 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1337_
timestamp 1
transform 1 0 32108 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1338_
timestamp 1
transform 1 0 25024 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1339_
timestamp 1
transform 1 0 24748 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1340_
timestamp 1
transform 1 0 25300 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1341_
timestamp 1
transform -1 0 33028 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1342_
timestamp 1
transform -1 0 14628 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1343_
timestamp 1
transform 1 0 12696 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1344_
timestamp 1
transform 1 0 13340 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1345_
timestamp 1
transform 1 0 32568 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1346_
timestamp 1
transform -1 0 37076 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1347_
timestamp 1
transform 1 0 34684 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1348_
timestamp 1
transform 1 0 20792 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1349_
timestamp 1
transform 1 0 26956 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1350_
timestamp 1
transform 1 0 29532 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1351_
timestamp 1
transform 1 0 34960 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1352_
timestamp 1
transform 1 0 18032 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1353_
timestamp 1
transform 1 0 15180 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1354_
timestamp 1
transform 1 0 22264 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1355_
timestamp 1
transform 1 0 27508 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1356_
timestamp 1
transform 1 0 42044 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1357_
timestamp 1
transform 1 0 29256 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1358_
timestamp 1
transform -1 0 30820 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1359_
timestamp 1
transform 1 0 35052 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1360_
timestamp 1
transform 1 0 29532 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1361_
timestamp 1
transform 1 0 28428 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1362_
timestamp 1
transform 1 0 29532 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1363_
timestamp 1
transform 1 0 24840 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1364_
timestamp 1
transform 1 0 25392 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1365_
timestamp 1
transform 1 0 26588 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1366_
timestamp 1
transform 1 0 29808 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1367_
timestamp 1
transform 1 0 35604 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1368_
timestamp 1
transform 1 0 31648 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1369_
timestamp 1
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1370_
timestamp 1
transform 1 0 20608 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1371_
timestamp 1
transform 1 0 21896 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1372_
timestamp 1
transform 1 0 26036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1373_
timestamp 1
transform 1 0 27784 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1374_
timestamp 1
transform 1 0 32108 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1375_
timestamp 1
transform 1 0 32660 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1376_
timestamp 1
transform 1 0 10396 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1377_
timestamp 1
transform 1 0 10856 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1378_
timestamp 1
transform 1 0 35604 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1379_
timestamp 1
transform 1 0 41032 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1380_
timestamp 1
transform 1 0 35328 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1381_
timestamp 1
transform 1 0 34684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1382_
timestamp 1
transform 1 0 39836 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1383_
timestamp 1
transform 1 0 38548 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1384_
timestamp 1
transform 1 0 37352 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1385_
timestamp 1
transform 1 0 38180 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1386_
timestamp 1
transform 1 0 12144 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1387_
timestamp 1
transform 1 0 39100 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1388_
timestamp 1
transform 1 0 40296 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1389_
timestamp 1
transform 1 0 31648 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1390_
timestamp 1
transform -1 0 32660 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1391_
timestamp 1
transform 1 0 26772 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1392_
timestamp 1
transform -1 0 26772 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1393_
timestamp 1
transform 1 0 25484 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1394_
timestamp 1
transform 1 0 26312 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1395_
timestamp 1
transform 1 0 25760 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1396_
timestamp 1
transform 1 0 19504 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1397_
timestamp 1
transform 1 0 26956 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1398_
timestamp 1
transform 1 0 27508 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1399_
timestamp 1
transform 1 0 31004 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1400_
timestamp 1
transform 1 0 32292 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1401_
timestamp 1
transform 1 0 22908 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1402_
timestamp 1
transform 1 0 23552 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1403_
timestamp 1
transform 1 0 24932 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1404_
timestamp 1
transform 1 0 31372 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1405_
timestamp 1
transform 1 0 17020 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1406_
timestamp 1
transform 1 0 31188 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1407_
timestamp 1
transform 1 0 32108 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1408_
timestamp 1
transform -1 0 42688 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1409_
timestamp 1
transform -1 0 34500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1410_
timestamp 1
transform 1 0 33948 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1411_
timestamp 1
transform 1 0 32108 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1412_
timestamp 1
transform 1 0 28980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1413_
timestamp 1
transform 1 0 31096 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1414_
timestamp 1
transform 1 0 32200 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1415_
timestamp 1
transform 1 0 32936 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1416_
timestamp 1
transform -1 0 39284 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1417_
timestamp 1
transform 1 0 35328 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1418_
timestamp 1
transform 1 0 36432 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1419_
timestamp 1
transform 1 0 35604 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1420_
timestamp 1
transform 1 0 36156 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1421_
timestamp 1
transform 1 0 37260 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1422_
timestamp 1
transform 1 0 39836 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1423_
timestamp 1
transform 1 0 36616 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1424_
timestamp 1
transform 1 0 37444 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1425_
timestamp 1
transform -1 0 42044 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1426_
timestamp 1
transform -1 0 40480 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1427_
timestamp 1
transform -1 0 38548 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1428_
timestamp 1
transform 1 0 37628 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1429_
timestamp 1
transform 1 0 41032 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1430_
timestamp 1
transform 1 0 27508 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1431_
timestamp 1
transform -1 0 23276 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1432_
timestamp 1
transform 1 0 24012 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1433_
timestamp 1
transform 1 0 41492 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1434_
timestamp 1
transform 1 0 42136 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1435_
timestamp 1
transform 1 0 41124 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1436_
timestamp 1
transform -1 0 30268 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1437_
timestamp 1
transform 1 0 22172 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1438_
timestamp 1
transform 1 0 25668 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1439_
timestamp 1
transform 1 0 39836 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1440_
timestamp 1
transform 1 0 40664 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1441_
timestamp 1
transform 1 0 40480 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1442_
timestamp 1
transform 1 0 38456 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1443_
timestamp 1
transform 1 0 26956 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1444_
timestamp 1
transform 1 0 42412 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1445_
timestamp 1
transform 1 0 41492 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1446_
timestamp 1
transform 1 0 40296 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1447_
timestamp 1
transform 1 0 22264 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1448_
timestamp 1
transform 1 0 41584 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1449_
timestamp 1
transform 1 0 37076 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1450_
timestamp 1
transform 1 0 41216 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1451_
timestamp 1
transform 1 0 35604 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1452_
timestamp 1
transform 1 0 40572 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1453_
timestamp 1
transform 1 0 40296 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1454_
timestamp 1
transform 1 0 30636 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1455_
timestamp 1
transform 1 0 42412 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1456_
timestamp 1
transform 1 0 39284 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1457_
timestamp 1
transform 1 0 39836 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1458_
timestamp 1
transform 1 0 42412 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1459_
timestamp 1
transform 1 0 38548 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform 1 0 22724 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1
transform 1 0 9384 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1
transform 1 0 33488 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1
transform 1 0 32660 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1
transform -1 0 37904 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1
transform 1 0 24840 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1
transform 1 0 25760 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1
transform 1 0 28704 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1
transform 1 0 26772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1
transform 1 0 29072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1
transform 1 0 28336 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1
transform 1 0 37076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1
transform -1 0 14444 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1
transform -1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1
transform 1 0 27508 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1
transform 1 0 27784 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1
transform 1 0 36248 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1
transform 1 0 26128 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1
transform -1 0 37904 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1
transform 1 0 23828 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1
transform 1 0 38916 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1
transform 1 0 24656 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1
transform -1 0 32568 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1
transform -1 0 33212 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1
transform -1 0 39100 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1
transform 1 0 33120 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1
transform 1 0 20424 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1
transform 1 0 33396 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1
transform 1 0 19136 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1
transform 1 0 32384 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk0
timestamp 1
transform -1 0 34224 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk0
timestamp 1
transform 1 0 36064 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk0
timestamp 1
transform -1 0 29440 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk0
timestamp 1
transform -1 0 39744 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk0
timestamp 1
transform 1 0 40480 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__bufinv_16  clkload0
timestamp 1
transform 1 0 36064 0 1 29376
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_2  clkload1
timestamp 1
transform -1 0 28428 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  clkload2
timestamp 1
transform -1 0 40480 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp 1
transform 1 0 37812 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout43
timestamp 1
transform -1 0 38548 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout44
timestamp 1
transform 1 0 38088 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout45
timestamp 1
transform 1 0 38088 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 1
transform -1 0 7268 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout50
timestamp 1
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout52
timestamp 1
transform -1 0 7820 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout53
timestamp 1
transform 1 0 12788 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout54
timestamp 1
transform -1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout55
timestamp 1
transform 1 0 11960 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout56
timestamp 1
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout57
timestamp 1
transform 1 0 11592 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout58
timestamp 1
transform -1 0 12328 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout59
timestamp 1
transform 1 0 3588 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout60
timestamp 1
transform 1 0 4324 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout61
timestamp 1
transform 1 0 12788 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout62
timestamp 1
transform -1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout63
timestamp 1
transform 1 0 5612 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout64
timestamp 1
transform 1 0 3588 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout65
timestamp 1
transform 1 0 3404 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout67
timestamp 1
transform -1 0 3496 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout68
timestamp 1
transform 1 0 13156 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout69
timestamp 1
transform 1 0 2300 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout70
timestamp 1
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout78
timestamp 1
transform 1 0 8740 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout79
timestamp 1
transform 1 0 9660 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout80
timestamp 1
transform 1 0 9108 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout81
timestamp 1
transform 1 0 9936 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout82
timestamp 1
transform 1 0 7728 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout83
timestamp 1
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout84
timestamp 1
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout85
timestamp 1
transform 1 0 2944 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout86
timestamp 1
transform -1 0 8096 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout87
timestamp 1
transform 1 0 12420 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout88
timestamp 1
transform 1 0 8556 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout89
timestamp 1
transform 1 0 13248 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout90
timestamp 1
transform -1 0 11224 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout91
timestamp 1
transform 1 0 5704 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout92
timestamp 1
transform -1 0 11776 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout93
timestamp 1
transform -1 0 6164 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout94
timestamp 1
transform -1 0 12880 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout95
timestamp 1
transform 1 0 14812 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout96
timestamp 1
transform -1 0 10948 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout97
timestamp 1
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout98
timestamp 1
transform -1 0 5612 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout99
timestamp 1
transform 1 0 16928 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout100
timestamp 1
transform 1 0 4140 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout101
timestamp 1
transform 1 0 12420 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout103
timestamp 1
transform 1 0 5612 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout104
timestamp 1
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout110
timestamp 1
transform -1 0 5152 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout111
timestamp 1
transform 1 0 12236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout112
timestamp 1
transform 1 0 14168 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout113
timestamp 1
transform 1 0 4600 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout114
timestamp 1
transform 1 0 15272 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout115
timestamp 1
transform -1 0 4324 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout116
timestamp 1
transform -1 0 9752 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout117
timestamp 1
transform 1 0 15088 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout119
timestamp 1
transform -1 0 11316 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout120
timestamp 1
transform 1 0 10304 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout121
timestamp 1
transform -1 0 9476 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout122
timestamp 1
transform 1 0 15456 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout123
timestamp 1
transform -1 0 10672 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout124
timestamp 1
transform 1 0 9936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout125
timestamp 1
transform -1 0 37812 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout126
timestamp 1
transform -1 0 42872 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout127
timestamp 1
transform -1 0 44160 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout128
timestamp 1
transform 1 0 43148 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout129
timestamp 1
transform -1 0 42320 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout130
timestamp 1
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout131
timestamp 1
transform 1 0 2392 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout132
timestamp 1
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout133
timestamp 1
transform 1 0 2668 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout134
timestamp 1
transform 1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout135
timestamp 1
transform 1 0 2116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout136
timestamp 1
transform 1 0 7176 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout137
timestamp 1
transform 1 0 2576 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout138
timestamp 1
transform -1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout139
timestamp 1
transform 1 0 3956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout140
timestamp 1
transform 1 0 2852 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout141
timestamp 1
transform 1 0 4140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout142
timestamp 1
transform -1 0 2484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout143
timestamp 1
transform 1 0 5060 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout144
timestamp 1
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout145
timestamp 1
transform 1 0 4692 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1636968456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1636968456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1636968456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1636968456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1636968456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1636968456
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1636968456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1636968456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1636968456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1636968456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1636968456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1636968456
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1636968456
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1636968456
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1636968456
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1636968456
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1636968456
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1636968456
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 1636968456
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_405
timestamp 1636968456
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_417
timestamp 1
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 1636968456
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_433
timestamp 1636968456
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 1
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_449
timestamp 1636968456
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_461
timestamp 1636968456
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1636968456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1636968456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1636968456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1636968456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1636968456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1636968456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1636968456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1636968456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1636968456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1636968456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1636968456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1636968456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1636968456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1636968456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1636968456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1636968456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1636968456
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1636968456
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1636968456
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1636968456
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1636968456
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_405
timestamp 1636968456
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_417
timestamp 1636968456
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_429
timestamp 1636968456
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_441
timestamp 1
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1636968456
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_461
timestamp 1636968456
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1636968456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1636968456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1636968456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1636968456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1636968456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1636968456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1636968456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1636968456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1636968456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1636968456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1636968456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1636968456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1636968456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1636968456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1636968456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1636968456
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1636968456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1636968456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1636968456
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1636968456
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1636968456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1636968456
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1636968456
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1636968456
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 1
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1636968456
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1636968456
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1636968456
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_457
timestamp 1636968456
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_469
timestamp 1
transform 1 0 44252 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1636968456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1636968456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1636968456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1636968456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1636968456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1636968456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1636968456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1636968456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1636968456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1636968456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1636968456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1636968456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1636968456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1636968456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1636968456
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1636968456
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1636968456
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1636968456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1636968456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1636968456
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1636968456
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1636968456
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1636968456
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1636968456
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1636968456
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1636968456
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1636968456
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1636968456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1636968456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1636968456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1636968456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1636968456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1636968456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1636968456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1636968456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1636968456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1636968456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1636968456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1636968456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1636968456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1636968456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1636968456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1636968456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1636968456
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1636968456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1636968456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1636968456
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1636968456
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1636968456
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1636968456
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1636968456
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1636968456
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1636968456
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1636968456
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1636968456
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 1636968456
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_469
timestamp 1
transform 1 0 44252 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636968456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1636968456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1636968456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1636968456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636968456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1636968456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1636968456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1636968456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1636968456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1636968456
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1636968456
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1636968456
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1636968456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1636968456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1636968456
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1636968456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1636968456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1636968456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1636968456
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1636968456
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1636968456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1636968456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1636968456
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1636968456
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1636968456
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1636968456
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1636968456
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1636968456
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1636968456
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1636968456
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1636968456
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1636968456
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1636968456
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 1636968456
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1636968456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1636968456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1636968456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1636968456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1636968456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1636968456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1636968456
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1636968456
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1636968456
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1636968456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1636968456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1636968456
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1636968456
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1636968456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1636968456
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1636968456
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1636968456
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1636968456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1636968456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1636968456
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1636968456
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1636968456
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1636968456
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1636968456
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1636968456
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1636968456
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1636968456
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1636968456
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1636968456
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1636968456
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1636968456
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1636968456
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_457
timestamp 1636968456
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_469
timestamp 1
transform 1 0 44252 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1636968456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1636968456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1636968456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1636968456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1636968456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1636968456
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1636968456
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1636968456
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1636968456
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1636968456
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1636968456
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1636968456
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1636968456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1636968456
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1636968456
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1636968456
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1636968456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1636968456
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1636968456
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1636968456
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1636968456
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1636968456
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1636968456
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1636968456
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1636968456
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1636968456
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1636968456
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1636968456
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1636968456
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1636968456
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1636968456
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1636968456
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1636968456
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_461
timestamp 1636968456
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1636968456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1636968456
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1636968456
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1636968456
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1636968456
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1636968456
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1636968456
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1636968456
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1636968456
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1636968456
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1636968456
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1636968456
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1636968456
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1636968456
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1636968456
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1636968456
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1636968456
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1636968456
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1636968456
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1636968456
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1636968456
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1636968456
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1636968456
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1636968456
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1636968456
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1636968456
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1636968456
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1636968456
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1636968456
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1636968456
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1636968456
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_457
timestamp 1636968456
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_469
timestamp 1
transform 1 0 44252 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1636968456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1636968456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1636968456
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1636968456
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1636968456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1636968456
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1636968456
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1636968456
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1636968456
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1636968456
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1636968456
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1636968456
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1636968456
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1636968456
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1636968456
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1636968456
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1636968456
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1636968456
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1636968456
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1636968456
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1636968456
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1636968456
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1636968456
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1636968456
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1636968456
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1636968456
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1636968456
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1636968456
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1636968456
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1636968456
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1636968456
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1636968456
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1636968456
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_461
timestamp 1636968456
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1636968456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1636968456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1636968456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1636968456
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1636968456
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1636968456
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1636968456
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1636968456
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1636968456
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1636968456
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1636968456
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1636968456
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1636968456
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1636968456
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1636968456
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1636968456
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1636968456
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1636968456
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1636968456
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1636968456
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1636968456
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1636968456
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1636968456
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1636968456
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1636968456
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1636968456
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1636968456
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1636968456
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1636968456
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1636968456
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1636968456
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1636968456
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1636968456
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_457
timestamp 1636968456
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_469
timestamp 1
transform 1 0 44252 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1636968456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1636968456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1636968456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1636968456
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1636968456
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1636968456
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1636968456
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1636968456
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1636968456
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1636968456
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1636968456
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1636968456
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1636968456
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1636968456
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1636968456
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1636968456
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1636968456
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1636968456
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1636968456
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1636968456
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1636968456
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1636968456
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1636968456
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1636968456
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1636968456
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1636968456
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1636968456
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1636968456
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1636968456
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1636968456
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1636968456
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1636968456
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 1636968456
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_461
timestamp 1636968456
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1636968456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1636968456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1636968456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1636968456
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1636968456
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1636968456
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1636968456
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1636968456
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1636968456
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1636968456
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1636968456
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1636968456
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1636968456
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1636968456
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1636968456
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1636968456
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1636968456
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1636968456
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1636968456
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1636968456
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1636968456
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1636968456
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1636968456
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1636968456
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1636968456
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1636968456
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1636968456
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1636968456
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1636968456
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 1636968456
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 1
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1636968456
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1636968456
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1636968456
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_457
timestamp 1636968456
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_469
timestamp 1
transform 1 0 44252 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1636968456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1636968456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1636968456
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1636968456
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1636968456
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1636968456
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1636968456
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1636968456
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1636968456
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1636968456
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1636968456
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1636968456
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1636968456
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1636968456
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1636968456
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1636968456
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1636968456
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1636968456
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1636968456
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1636968456
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1636968456
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1636968456
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1636968456
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 1
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 1636968456
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 1636968456
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_361
timestamp 1636968456
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_373
timestamp 1636968456
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_385
timestamp 1
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 1636968456
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_405
timestamp 1636968456
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_417
timestamp 1636968456
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_429
timestamp 1636968456
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_441
timestamp 1
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 1
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_449
timestamp 1636968456
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_461
timestamp 1636968456
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1636968456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1636968456
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1636968456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1636968456
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1636968456
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1636968456
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1636968456
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1636968456
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1636968456
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1636968456
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1636968456
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1636968456
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1636968456
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1636968456
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1636968456
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1636968456
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1636968456
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1636968456
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1636968456
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1636968456
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1636968456
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1636968456
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1636968456
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 1636968456
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_333
timestamp 1636968456
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_345
timestamp 1636968456
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_357
timestamp 1
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 1636968456
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 1636968456
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 1636968456
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_401
timestamp 1636968456
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_413
timestamp 1
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_419
timestamp 1
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_421
timestamp 1636968456
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_433
timestamp 1636968456
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_445
timestamp 1636968456
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_457
timestamp 1636968456
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_469
timestamp 1
transform 1 0 44252 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1636968456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1636968456
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1636968456
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1636968456
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1636968456
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1636968456
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1636968456
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1636968456
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1636968456
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1636968456
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1636968456
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1636968456
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1636968456
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1636968456
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1636968456
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1636968456
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1636968456
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1636968456
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1636968456
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 1636968456
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 1
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1636968456
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1636968456
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1636968456
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1636968456
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 1
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 1636968456
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 1636968456
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_361
timestamp 1636968456
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_373
timestamp 1636968456
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_385
timestamp 1
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_391
timestamp 1
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_393
timestamp 1636968456
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_405
timestamp 1636968456
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_417
timestamp 1636968456
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_429
timestamp 1636968456
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_441
timestamp 1
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_447
timestamp 1
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_449
timestamp 1636968456
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_461
timestamp 1636968456
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1636968456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1636968456
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1636968456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1636968456
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1636968456
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1636968456
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1636968456
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1636968456
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1636968456
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1636968456
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1636968456
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1636968456
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1636968456
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1636968456
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1636968456
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1636968456
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1636968456
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1636968456
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1636968456
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1636968456
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1636968456
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1636968456
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1636968456
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1636968456
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_333
timestamp 1636968456
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_345
timestamp 1636968456
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_357
timestamp 1
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 1636968456
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_377
timestamp 1636968456
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_389
timestamp 1636968456
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_401
timestamp 1636968456
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_413
timestamp 1
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_419
timestamp 1
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_421
timestamp 1636968456
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_433
timestamp 1636968456
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_445
timestamp 1636968456
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_457
timestamp 1636968456
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_469
timestamp 1
transform 1 0 44252 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_6
timestamp 1636968456
transform 1 0 1656 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_18
timestamp 1636968456
transform 1 0 2760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_30
timestamp 1636968456
transform 1 0 3864 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_42
timestamp 1636968456
transform 1 0 4968 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1636968456
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1636968456
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1636968456
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1636968456
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1636968456
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1636968456
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1636968456
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1636968456
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1636968456
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1636968456
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1636968456
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1636968456
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1636968456
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1636968456
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1636968456
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1636968456
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1636968456
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1636968456
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1636968456
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1636968456
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1636968456
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 1636968456
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_361
timestamp 1636968456
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_373
timestamp 1636968456
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_385
timestamp 1
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 1
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_393
timestamp 1636968456
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_405
timestamp 1636968456
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_417
timestamp 1636968456
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_429
timestamp 1636968456
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_441
timestamp 1
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_447
timestamp 1
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_449
timestamp 1636968456
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_461
timestamp 1636968456
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_9
timestamp 1636968456
transform 1 0 1932 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_21
timestamp 1
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_29
timestamp 1
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_37
timestamp 1
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_56
timestamp 1636968456
transform 1 0 6256 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_68
timestamp 1
transform 1 0 7360 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1636968456
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_97
timestamp 1
transform 1 0 10028 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_104
timestamp 1636968456
transform 1 0 10672 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_116
timestamp 1
transform 1 0 11776 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_120
timestamp 1
transform 1 0 12144 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_129
timestamp 1
transform 1 0 12972 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_137
timestamp 1
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_141
timestamp 1
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_146
timestamp 1
transform 1 0 14536 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_155
timestamp 1636968456
transform 1 0 15364 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_167
timestamp 1
transform 1 0 16468 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_173
timestamp 1
transform 1 0 17020 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_182
timestamp 1636968456
transform 1 0 17848 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_205
timestamp 1636968456
transform 1 0 19964 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_217
timestamp 1636968456
transform 1 0 21068 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_229
timestamp 1636968456
transform 1 0 22172 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_241
timestamp 1
transform 1 0 23276 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_249
timestamp 1
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1636968456
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1636968456
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1636968456
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1636968456
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1636968456
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1636968456
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 1636968456
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 1636968456
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_357
timestamp 1
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 1
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 1636968456
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 1636968456
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 1636968456
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_401
timestamp 1636968456
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_413
timestamp 1
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_419
timestamp 1
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_421
timestamp 1636968456
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_433
timestamp 1636968456
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_445
timestamp 1636968456
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_457
timestamp 1636968456
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_469
timestamp 1
transform 1 0 44252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_3
timestamp 1
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_26
timestamp 1
transform 1 0 3496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_30
timestamp 1
transform 1 0 3864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_64
timestamp 1
transform 1 0 6992 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_86
timestamp 1
transform 1 0 9016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_94
timestamp 1
transform 1 0 9752 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_135
timestamp 1
transform 1 0 13524 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_158
timestamp 1
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_169
timestamp 1
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_173
timestamp 1
transform 1 0 17020 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_182
timestamp 1
transform 1 0 17848 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_207
timestamp 1636968456
transform 1 0 20148 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_219
timestamp 1
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1636968456
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_237
timestamp 1
transform 1 0 22908 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1636968456
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_261
timestamp 1
transform 1 0 25116 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_272
timestamp 1
transform 1 0 26128 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1636968456
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1636968456
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1636968456
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_317
timestamp 1
transform 1 0 30268 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_331
timestamp 1
transform 1 0 31556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 1
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 1636968456
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1636968456
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_361
timestamp 1636968456
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_373
timestamp 1636968456
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_385
timestamp 1
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 1
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 1636968456
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_405
timestamp 1636968456
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_417
timestamp 1636968456
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_429
timestamp 1636968456
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_441
timestamp 1
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_447
timestamp 1
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_449
timestamp 1636968456
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_461
timestamp 1636968456
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_3
timestamp 1
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_85
timestamp 1
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_94
timestamp 1
transform 1 0 9752 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_141
timestamp 1
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_145
timestamp 1
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_154
timestamp 1636968456
transform 1 0 15272 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_166
timestamp 1
transform 1 0 16376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_170
timestamp 1
transform 1 0 16744 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_179
timestamp 1636968456
transform 1 0 17572 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_191
timestamp 1
transform 1 0 18676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1636968456
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1636968456
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_221
timestamp 1
transform 1 0 21436 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_227
timestamp 1
transform 1 0 21988 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 1636968456
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 1
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_253
timestamp 1
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_261
timestamp 1
transform 1 0 25116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_268
timestamp 1
transform 1 0 25760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_276
timestamp 1
transform 1 0 26496 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_284
timestamp 1636968456
transform 1 0 27232 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1636968456
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_321
timestamp 1
transform 1 0 30636 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_327
timestamp 1
transform 1 0 31188 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 1636968456
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 1636968456
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_357
timestamp 1
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 1636968456
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_377
timestamp 1636968456
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 1636968456
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_401
timestamp 1636968456
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_413
timestamp 1
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_419
timestamp 1
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_421
timestamp 1636968456
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_433
timestamp 1636968456
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_445
timestamp 1636968456
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_457
timestamp 1636968456
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_469
timestamp 1
transform 1 0 44252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_24
timestamp 1
transform 1 0 3312 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_32
timestamp 1
transform 1 0 4048 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 1
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1636968456
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_69
timestamp 1
transform 1 0 7452 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_91
timestamp 1
transform 1 0 9476 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_99
timestamp 1
transform 1 0 10212 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_104
timestamp 1
transform 1 0 10672 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_121
timestamp 1636968456
transform 1 0 12236 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_133
timestamp 1636968456
transform 1 0 13340 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 1
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_169
timestamp 1
transform 1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_176
timestamp 1
transform 1 0 17296 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_184
timestamp 1
transform 1 0 18032 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_190
timestamp 1
transform 1 0 18584 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_199
timestamp 1636968456
transform 1 0 19412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_211
timestamp 1
transform 1 0 20516 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_220
timestamp 1
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_230
timestamp 1
transform 1 0 22264 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_239
timestamp 1636968456
transform 1 0 23092 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_251
timestamp 1636968456
transform 1 0 24196 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_263
timestamp 1
transform 1 0 25300 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_297
timestamp 1
transform 1 0 28428 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_304
timestamp 1636968456
transform 1 0 29072 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_316
timestamp 1636968456
transform 1 0 30176 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_328
timestamp 1
transform 1 0 31280 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_342
timestamp 1636968456
transform 1 0 32568 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_354
timestamp 1636968456
transform 1 0 33672 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_366
timestamp 1636968456
transform 1 0 34776 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_378
timestamp 1636968456
transform 1 0 35880 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_390
timestamp 1
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 1636968456
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_405
timestamp 1636968456
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_417
timestamp 1636968456
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_429
timestamp 1636968456
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_441
timestamp 1
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_447
timestamp 1
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_449
timestamp 1636968456
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_461
timestamp 1
transform 1 0 43516 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_6
timestamp 1
transform 1 0 1656 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_10
timestamp 1
transform 1 0 2024 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1636968456
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1636968456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_41
timestamp 1
transform 1 0 4876 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_46
timestamp 1
transform 1 0 5336 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_65
timestamp 1
transform 1 0 7084 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_96
timestamp 1636968456
transform 1 0 9936 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_108
timestamp 1636968456
transform 1 0 11040 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_120
timestamp 1636968456
transform 1 0 12144 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_132
timestamp 1
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_149
timestamp 1
transform 1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_160
timestamp 1
transform 1 0 15824 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_169
timestamp 1636968456
transform 1 0 16652 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_181
timestamp 1636968456
transform 1 0 17756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_193
timestamp 1
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_197
timestamp 1
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_210
timestamp 1
transform 1 0 20424 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_218
timestamp 1
transform 1 0 21160 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_228
timestamp 1
transform 1 0 22080 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_238
timestamp 1
transform 1 0 23000 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 1
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1636968456
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1636968456
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1636968456
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1636968456
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1636968456
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_321
timestamp 1
transform 1 0 30636 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_327
timestamp 1636968456
transform 1 0 31188 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_339
timestamp 1636968456
transform 1 0 32292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_351
timestamp 1636968456
transform 1 0 33396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 1
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 1636968456
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 1636968456
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 1636968456
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_401
timestamp 1636968456
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_413
timestamp 1
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_419
timestamp 1
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_421
timestamp 1636968456
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_433
timestamp 1636968456
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_445
timestamp 1636968456
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_457
timestamp 1636968456
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1636968456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_25
timestamp 1636968456
transform 1 0 3404 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_37
timestamp 1636968456
transform 1 0 4508 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_49
timestamp 1
transform 1 0 5612 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_70
timestamp 1
transform 1 0 7544 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_76
timestamp 1
transform 1 0 8096 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_95
timestamp 1
transform 1 0 9844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_113
timestamp 1
transform 1 0 11500 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1636968456
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_137
timestamp 1
transform 1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_145
timestamp 1
transform 1 0 14444 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_155
timestamp 1636968456
transform 1 0 15364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1636968456
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_181
timestamp 1
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_189
timestamp 1
transform 1 0 18492 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_199
timestamp 1636968456
transform 1 0 19412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_211
timestamp 1636968456
transform 1 0 20516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1636968456
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_237
timestamp 1
transform 1 0 22908 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_245
timestamp 1
transform 1 0 23644 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_253
timestamp 1636968456
transform 1 0 24380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_265
timestamp 1
transform 1 0 25484 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_271
timestamp 1
transform 1 0 26036 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_278
timestamp 1
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_286
timestamp 1
transform 1 0 27416 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_292
timestamp 1636968456
transform 1 0 27968 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_304
timestamp 1636968456
transform 1 0 29072 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_316
timestamp 1
transform 1 0 30176 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1636968456
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_349
timestamp 1
transform 1 0 33212 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_358
timestamp 1636968456
transform 1 0 34040 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_370
timestamp 1636968456
transform 1 0 35144 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_382
timestamp 1
transform 1 0 36248 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_390
timestamp 1
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_393
timestamp 1
transform 1 0 37260 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_413
timestamp 1636968456
transform 1 0 39100 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_425
timestamp 1636968456
transform 1 0 40204 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_437
timestamp 1
transform 1 0 41308 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_445
timestamp 1
transform 1 0 42044 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_457
timestamp 1636968456
transform 1 0 43148 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_469
timestamp 1
transform 1 0 44252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_6
timestamp 1
transform 1 0 1656 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1636968456
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_41
timestamp 1
transform 1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_73
timestamp 1
transform 1 0 7820 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_122
timestamp 1
transform 1 0 12328 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_132
timestamp 1
transform 1 0 13248 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_148
timestamp 1
transform 1 0 14720 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_159
timestamp 1
transform 1 0 15732 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_169
timestamp 1
transform 1 0 16652 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_177
timestamp 1
transform 1 0 17388 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1636968456
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1636968456
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_221
timestamp 1
transform 1 0 21436 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_229
timestamp 1
transform 1 0 22172 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_236
timestamp 1
transform 1 0 22816 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_244
timestamp 1
transform 1 0 23552 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_253
timestamp 1
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_261
timestamp 1
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_268
timestamp 1
transform 1 0 25760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_276
timestamp 1
transform 1 0 26496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_283
timestamp 1
transform 1 0 27140 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_289
timestamp 1
transform 1 0 27692 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_296
timestamp 1636968456
transform 1 0 28336 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_314
timestamp 1636968456
transform 1 0 29992 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_326
timestamp 1636968456
transform 1 0 31096 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_338
timestamp 1
transform 1 0 32200 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_371
timestamp 1
transform 1 0 35236 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_407
timestamp 1636968456
transform 1 0 38548 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_419
timestamp 1
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_421
timestamp 1
transform 1 0 39836 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_429
timestamp 1
transform 1 0 40572 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_455
timestamp 1636968456
transform 1 0 42964 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_467
timestamp 1
transform 1 0 44068 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_6
timestamp 1
transform 1 0 1656 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_15
timestamp 1
transform 1 0 2484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_21
timestamp 1
transform 1 0 3036 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_42
timestamp 1
transform 1 0 4968 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_71
timestamp 1
transform 1 0 7636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_82
timestamp 1
transform 1 0 8648 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_107
timestamp 1
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_113
timestamp 1
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_128
timestamp 1
transform 1 0 12880 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_135
timestamp 1636968456
transform 1 0 13524 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_147
timestamp 1
transform 1 0 14628 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_151
timestamp 1
transform 1 0 14996 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_156
timestamp 1
transform 1 0 15456 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_166
timestamp 1
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_169
timestamp 1
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_179
timestamp 1
transform 1 0 17572 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_187
timestamp 1
transform 1 0 18308 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_196
timestamp 1
transform 1 0 19136 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_204
timestamp 1
transform 1 0 19872 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_212
timestamp 1636968456
transform 1 0 20608 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_225
timestamp 1
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_241
timestamp 1636968456
transform 1 0 23276 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_253
timestamp 1
transform 1 0 24380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_259
timestamp 1
transform 1 0 24932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_265
timestamp 1
transform 1 0 25484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 1
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1636968456
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_293
timestamp 1
transform 1 0 28060 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_301
timestamp 1
transform 1 0 28796 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_314
timestamp 1636968456
transform 1 0 29992 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_326
timestamp 1
transform 1 0 31096 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_334
timestamp 1
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_337
timestamp 1
transform 1 0 32108 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1636968456
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_361
timestamp 1
transform 1 0 34316 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 1
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_417
timestamp 1636968456
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_429
timestamp 1636968456
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_441
timestamp 1
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_447
timestamp 1
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_449
timestamp 1636968456
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_461
timestamp 1
transform 1 0 43516 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_20
timestamp 1
transform 1 0 2944 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_36
timestamp 1
transform 1 0 4416 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_73
timestamp 1
transform 1 0 7820 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_85
timestamp 1
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_109
timestamp 1
transform 1 0 11132 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_118
timestamp 1636968456
transform 1 0 11960 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_130
timestamp 1
transform 1 0 13064 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1636968456
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_153
timestamp 1
transform 1 0 15180 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_166
timestamp 1
transform 1 0 16376 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_172
timestamp 1
transform 1 0 16928 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_183
timestamp 1636968456
transform 1 0 17940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1636968456
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_209
timestamp 1
transform 1 0 20332 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_226
timestamp 1
transform 1 0 21896 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_237
timestamp 1636968456
transform 1 0 22908 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_249
timestamp 1
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_253
timestamp 1
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_275
timestamp 1636968456
transform 1 0 26404 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_287
timestamp 1
transform 1 0 27508 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_295
timestamp 1
transform 1 0 28244 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_303
timestamp 1
transform 1 0 28980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1636968456
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_321
timestamp 1
transform 1 0 30636 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_329
timestamp 1
transform 1 0 31372 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_342
timestamp 1636968456
transform 1 0 32568 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_354
timestamp 1
transform 1 0 33672 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_362
timestamp 1
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 1636968456
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_377
timestamp 1636968456
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_389
timestamp 1
transform 1 0 36892 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_393
timestamp 1
transform 1 0 37260 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_409
timestamp 1
transform 1 0 38732 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_417
timestamp 1
transform 1 0 39468 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_421
timestamp 1636968456
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_433
timestamp 1636968456
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_445
timestamp 1636968456
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_457
timestamp 1636968456
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_3
timestamp 1
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1636968456
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_41
timestamp 1
transform 1 0 4876 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_49
timestamp 1
transform 1 0 5612 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_57
timestamp 1
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_61
timestamp 1
transform 1 0 6716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_80
timestamp 1
transform 1 0 8464 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_99
timestamp 1
transform 1 0 10212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_107
timestamp 1
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_125
timestamp 1
transform 1 0 12604 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_153
timestamp 1636968456
transform 1 0 15180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_165
timestamp 1
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1636968456
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_181
timestamp 1
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_203
timestamp 1636968456
transform 1 0 19780 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_215
timestamp 1
transform 1 0 20884 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1636968456
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_237
timestamp 1
transform 1 0 22908 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_243
timestamp 1636968456
transform 1 0 23460 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_255
timestamp 1
transform 1 0 24564 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_263
timestamp 1636968456
transform 1 0 25300 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_275
timestamp 1
transform 1 0 26404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_286
timestamp 1
transform 1 0 27416 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_295
timestamp 1636968456
transform 1 0 28244 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_307
timestamp 1
transform 1 0 29348 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_313
timestamp 1636968456
transform 1 0 29900 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_325
timestamp 1
transform 1 0 31004 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_342
timestamp 1636968456
transform 1 0 32568 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_354
timestamp 1636968456
transform 1 0 33672 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_366
timestamp 1
transform 1 0 34776 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_374
timestamp 1
transform 1 0 35512 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_381
timestamp 1
transform 1 0 36156 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_389
timestamp 1
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_431
timestamp 1636968456
transform 1 0 40756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_443
timestamp 1
transform 1 0 41860 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_447
timestamp 1
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_465
timestamp 1
transform 1 0 43884 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_3
timestamp 1
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_11
timestamp 1
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_17
timestamp 1
transform 1 0 2668 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_29
timestamp 1
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_33
timestamp 1
transform 1 0 4140 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_37
timestamp 1
transform 1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_53
timestamp 1
transform 1 0 5980 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_63
timestamp 1
transform 1 0 6900 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_85
timestamp 1
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_89
timestamp 1
transform 1 0 9292 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_98
timestamp 1636968456
transform 1 0 10120 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_110
timestamp 1
transform 1 0 11224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_114
timestamp 1
transform 1 0 11592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_141
timestamp 1
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_149
timestamp 1
transform 1 0 14812 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_155
timestamp 1636968456
transform 1 0 15364 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_167
timestamp 1
transform 1 0 16468 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_175
timestamp 1636968456
transform 1 0 17204 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_187
timestamp 1
transform 1 0 18308 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_197
timestamp 1
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_204
timestamp 1636968456
transform 1 0 19872 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_216
timestamp 1636968456
transform 1 0 20976 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_228
timestamp 1
transform 1 0 22080 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_236
timestamp 1
transform 1 0 22816 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_243
timestamp 1
transform 1 0 23460 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1636968456
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_265
timestamp 1
transform 1 0 25484 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_271
timestamp 1
transform 1 0 26036 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_287
timestamp 1
transform 1 0 27508 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_295
timestamp 1636968456
transform 1 0 28244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_316
timestamp 1
transform 1 0 30176 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_324
timestamp 1
transform 1 0 30912 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_344
timestamp 1
transform 1 0 32752 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_362
timestamp 1
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_365
timestamp 1
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_377
timestamp 1
transform 1 0 35788 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_387
timestamp 1
transform 1 0 36708 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_399
timestamp 1
transform 1 0 37812 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_413
timestamp 1
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_419
timestamp 1
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_437
timestamp 1
transform 1 0 41308 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_452
timestamp 1
transform 1 0 42688 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_464
timestamp 1
transform 1 0 43792 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_472
timestamp 1
transform 1 0 44528 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_3
timestamp 1
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_11
timestamp 1
transform 1 0 2116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_39
timestamp 1
transform 1 0 4692 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_57
timestamp 1
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_66
timestamp 1
transform 1 0 7176 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_74
timestamp 1
transform 1 0 7912 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_92
timestamp 1636968456
transform 1 0 9568 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_104
timestamp 1
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_113
timestamp 1
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_125
timestamp 1
transform 1 0 12604 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_144
timestamp 1
transform 1 0 14352 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_155
timestamp 1636968456
transform 1 0 15364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_169
timestamp 1
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_179
timestamp 1
transform 1 0 17572 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_186
timestamp 1
transform 1 0 18216 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_194
timestamp 1
transform 1 0 18952 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1636968456
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_225
timestamp 1
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_242
timestamp 1
transform 1 0 23368 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_250
timestamp 1636968456
transform 1 0 24104 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_262
timestamp 1
transform 1 0 25208 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_268
timestamp 1636968456
transform 1 0 25760 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_287
timestamp 1636968456
transform 1 0 27508 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_299
timestamp 1
transform 1 0 28612 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_303
timestamp 1
transform 1 0 28980 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_312
timestamp 1636968456
transform 1 0 29808 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_324
timestamp 1
transform 1 0 30912 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_333
timestamp 1
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_343
timestamp 1636968456
transform 1 0 32660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_355
timestamp 1
transform 1 0 33764 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_368
timestamp 1636968456
transform 1 0 34960 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_380
timestamp 1
transform 1 0 36064 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_393
timestamp 1
transform 1 0 37260 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_399
timestamp 1636968456
transform 1 0 37812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_411
timestamp 1
transform 1 0 38916 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_427
timestamp 1
transform 1 0 40388 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_431
timestamp 1
transform 1 0 40756 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_447
timestamp 1
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_449
timestamp 1636968456
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_461
timestamp 1
transform 1 0 43516 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_3
timestamp 1
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_11
timestamp 1
transform 1 0 2116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_19
timestamp 1
transform 1 0 2852 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_24
timestamp 1
transform 1 0 3312 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_29
timestamp 1
transform 1 0 3772 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_66
timestamp 1
transform 1 0 7176 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_85
timestamp 1
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_111
timestamp 1
transform 1 0 11316 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_119
timestamp 1
transform 1 0 12052 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_136
timestamp 1
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_141
timestamp 1
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_152
timestamp 1636968456
transform 1 0 15088 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_164
timestamp 1
transform 1 0 16192 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_174
timestamp 1636968456
transform 1 0 17112 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_186
timestamp 1
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_202
timestamp 1636968456
transform 1 0 19688 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_214
timestamp 1
transform 1 0 20792 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_228
timestamp 1636968456
transform 1 0 22080 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_240
timestamp 1636968456
transform 1 0 23184 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_253
timestamp 1
transform 1 0 24380 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_264
timestamp 1636968456
transform 1 0 25392 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_276
timestamp 1636968456
transform 1 0 26496 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_288
timestamp 1
transform 1 0 27600 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_299
timestamp 1
transform 1 0 28612 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1636968456
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_321
timestamp 1
transform 1 0 30636 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_335
timestamp 1636968456
transform 1 0 31924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_347
timestamp 1636968456
transform 1 0 33028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_359
timestamp 1
transform 1 0 34132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_365
timestamp 1636968456
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_377
timestamp 1636968456
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_389
timestamp 1
transform 1 0 36892 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_407
timestamp 1636968456
transform 1 0 38548 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_419
timestamp 1
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_429
timestamp 1
transform 1 0 40572 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_433
timestamp 1
transform 1 0 40940 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_466
timestamp 1
transform 1 0 43976 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_3
timestamp 1
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_11
timestamp 1
transform 1 0 2116 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_26
timestamp 1636968456
transform 1 0 3496 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_38
timestamp 1636968456
transform 1 0 4600 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_50
timestamp 1
transform 1 0 5704 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_64
timestamp 1636968456
transform 1 0 6992 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_76
timestamp 1
transform 1 0 8096 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_80
timestamp 1
transform 1 0 8464 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_85
timestamp 1636968456
transform 1 0 8924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_97
timestamp 1
transform 1 0 10028 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_107
timestamp 1
transform 1 0 10948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_113
timestamp 1
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_121
timestamp 1
transform 1 0 12236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_127
timestamp 1
transform 1 0 12788 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_138
timestamp 1
transform 1 0 13800 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_146
timestamp 1
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1636968456
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_181
timestamp 1
transform 1 0 17756 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_189
timestamp 1
transform 1 0 18492 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_208
timestamp 1
transform 1 0 20240 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_214
timestamp 1
transform 1 0 20792 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_220
timestamp 1
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_231
timestamp 1636968456
transform 1 0 22356 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_243
timestamp 1636968456
transform 1 0 23460 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_255
timestamp 1636968456
transform 1 0 24564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_267
timestamp 1636968456
transform 1 0 25668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1636968456
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1636968456
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1636968456
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1636968456
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_334
timestamp 1
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_342
timestamp 1636968456
transform 1 0 32568 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_354
timestamp 1
transform 1 0 33672 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_364
timestamp 1636968456
transform 1 0 34592 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_376
timestamp 1636968456
transform 1 0 35696 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_388
timestamp 1
transform 1 0 36800 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 1636968456
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_405
timestamp 1
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_428
timestamp 1636968456
transform 1 0 40480 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_440
timestamp 1
transform 1 0 41584 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_465
timestamp 1
transform 1 0 43884 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1636968456
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_15
timestamp 1
transform 1 0 2484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_19
timestamp 1
transform 1 0 2852 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_29
timestamp 1
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_37
timestamp 1
transform 1 0 4508 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_48
timestamp 1
transform 1 0 5520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_70
timestamp 1
transform 1 0 7544 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_93
timestamp 1636968456
transform 1 0 9660 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_105
timestamp 1636968456
transform 1 0 10764 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_117
timestamp 1
transform 1 0 11868 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_125
timestamp 1
transform 1 0 12604 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_136
timestamp 1
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_147
timestamp 1
transform 1 0 14628 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_155
timestamp 1
transform 1 0 15364 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_163
timestamp 1636968456
transform 1 0 16100 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_175
timestamp 1
transform 1 0 17204 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_183
timestamp 1
transform 1 0 17940 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_190
timestamp 1
transform 1 0 18584 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1636968456
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1636968456
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1636968456
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_233
timestamp 1
transform 1 0 22540 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_247
timestamp 1
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_258
timestamp 1
transform 1 0 24840 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_264
timestamp 1
transform 1 0 25392 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_271
timestamp 1
transform 1 0 26036 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_280
timestamp 1636968456
transform 1 0 26864 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_292
timestamp 1
transform 1 0 27968 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_300
timestamp 1
transform 1 0 28704 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_315
timestamp 1636968456
transform 1 0 30084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_327
timestamp 1
transform 1 0 31188 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_333
timestamp 1
transform 1 0 31740 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_345
timestamp 1
transform 1 0 32844 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_349
timestamp 1
transform 1 0 33212 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_356
timestamp 1
transform 1 0 33856 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 1
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_365
timestamp 1
transform 1 0 34684 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_378
timestamp 1636968456
transform 1 0 35880 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_390
timestamp 1
transform 1 0 36984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_396
timestamp 1
transform 1 0 37536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_421
timestamp 1
transform 1 0 39836 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_433
timestamp 1636968456
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_445
timestamp 1636968456
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_457
timestamp 1636968456
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1636968456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_15
timestamp 1
transform 1 0 2484 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_23
timestamp 1
transform 1 0 3220 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_35
timestamp 1636968456
transform 1 0 4324 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_47
timestamp 1
transform 1 0 5428 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1636968456
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1636968456
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_81
timestamp 1
transform 1 0 8556 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_104
timestamp 1
transform 1 0 10672 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_113
timestamp 1
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_121
timestamp 1
transform 1 0 12236 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_130
timestamp 1
transform 1 0 13064 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_142
timestamp 1
transform 1 0 14168 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_151
timestamp 1
transform 1 0 14996 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_161
timestamp 1
transform 1 0 15916 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1636968456
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_181
timestamp 1
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_191
timestamp 1
transform 1 0 18676 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_199
timestamp 1
transform 1 0 19412 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_206
timestamp 1
transform 1 0 20056 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_214
timestamp 1
transform 1 0 20792 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_225
timestamp 1
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_233
timestamp 1
transform 1 0 22540 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_242
timestamp 1
transform 1 0 23368 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_253
timestamp 1636968456
transform 1 0 24380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_265
timestamp 1
transform 1 0 25484 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_298
timestamp 1
transform 1 0 28520 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_302
timestamp 1
transform 1 0 28888 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_318
timestamp 1636968456
transform 1 0 30360 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_330
timestamp 1
transform 1 0 31464 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1636968456
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1636968456
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_361
timestamp 1
transform 1 0 34316 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_370
timestamp 1636968456
transform 1 0 35144 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_382
timestamp 1
transform 1 0 36248 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 1
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_393
timestamp 1636968456
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_411
timestamp 1636968456
transform 1 0 38916 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_423
timestamp 1636968456
transform 1 0 40020 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_435
timestamp 1
transform 1 0 41124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_439
timestamp 1
transform 1 0 41492 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_447
timestamp 1
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_449
timestamp 1636968456
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_461
timestamp 1636968456
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_3
timestamp 1
transform 1 0 1380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_18
timestamp 1
transform 1 0 2760 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_26
timestamp 1
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_37
timestamp 1636968456
transform 1 0 4508 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_49
timestamp 1636968456
transform 1 0 5612 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_61
timestamp 1
transform 1 0 6716 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_72
timestamp 1
transform 1 0 7728 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_76
timestamp 1
transform 1 0 8096 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_85
timestamp 1
transform 1 0 8924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_114
timestamp 1
transform 1 0 11592 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_137
timestamp 1
transform 1 0 13708 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_156
timestamp 1636968456
transform 1 0 15456 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_168
timestamp 1
transform 1 0 16560 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_176
timestamp 1
transform 1 0 17296 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_183
timestamp 1
transform 1 0 17940 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_190
timestamp 1
transform 1 0 18584 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_203
timestamp 1636968456
transform 1 0 19780 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_226
timestamp 1636968456
transform 1 0 21896 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_238
timestamp 1
transform 1 0 23000 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_244
timestamp 1
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_253
timestamp 1
transform 1 0 24380 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_260
timestamp 1636968456
transform 1 0 25024 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_272
timestamp 1
transform 1 0 26128 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_284
timestamp 1636968456
transform 1 0 27232 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_296
timestamp 1636968456
transform 1 0 28336 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1636968456
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 1636968456
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 1636968456
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_345
timestamp 1636968456
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_357
timestamp 1
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 1
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_365
timestamp 1
transform 1 0 34684 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_374
timestamp 1
transform 1 0 35512 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_378
timestamp 1
transform 1 0 35880 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_385
timestamp 1636968456
transform 1 0 36524 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_397
timestamp 1
transform 1 0 37628 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_408
timestamp 1636968456
transform 1 0 38640 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_421
timestamp 1636968456
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_433
timestamp 1
transform 1 0 40940 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_466
timestamp 1
transform 1 0 43976 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1636968456
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_15
timestamp 1
transform 1 0 2484 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_24
timestamp 1636968456
transform 1 0 3312 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_36
timestamp 1636968456
transform 1 0 4416 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_48
timestamp 1
transform 1 0 5520 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1636968456
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1636968456
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1636968456
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_103
timestamp 1
transform 1 0 10580 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_113
timestamp 1
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_121
timestamp 1
transform 1 0 12236 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_129
timestamp 1636968456
transform 1 0 12972 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_141
timestamp 1636968456
transform 1 0 14076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_153
timestamp 1636968456
transform 1 0 15180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_165
timestamp 1
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1636968456
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1636968456
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 1636968456
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_205
timestamp 1
transform 1 0 19964 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_209
timestamp 1
transform 1 0 20332 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_215
timestamp 1
transform 1 0 20884 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1636968456
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_237
timestamp 1
transform 1 0 22908 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_245
timestamp 1
transform 1 0 23644 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_260
timestamp 1636968456
transform 1 0 25024 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_272
timestamp 1
transform 1 0 26128 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1636968456
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 1636968456
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_305
timestamp 1
transform 1 0 29164 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_311
timestamp 1
transform 1 0 29716 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_323
timestamp 1
transform 1 0 30820 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_333
timestamp 1
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_342
timestamp 1
transform 1 0 32568 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_355
timestamp 1
transform 1 0 33764 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_366
timestamp 1636968456
transform 1 0 34776 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_378
timestamp 1636968456
transform 1 0 35880 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_390
timestamp 1
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_399
timestamp 1
transform 1 0 37812 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_417
timestamp 1
transform 1 0 39468 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_425
timestamp 1
transform 1 0 40204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_442
timestamp 1
transform 1 0 41768 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_449
timestamp 1
transform 1 0 42412 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_454
timestamp 1
transform 1 0 42872 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_463
timestamp 1
transform 1 0 43700 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1636968456
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1636968456
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1636968456
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_41
timestamp 1
transform 1 0 4876 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_50
timestamp 1
transform 1 0 5704 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_58
timestamp 1
transform 1 0 6440 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_75
timestamp 1
transform 1 0 8004 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1636968456
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1636968456
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_109
timestamp 1
transform 1 0 11132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_113
timestamp 1
transform 1 0 11500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_128
timestamp 1636968456
transform 1 0 12880 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_141
timestamp 1
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_147
timestamp 1
transform 1 0 14628 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_154
timestamp 1
transform 1 0 15272 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_165
timestamp 1
transform 1 0 16284 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_173
timestamp 1
transform 1 0 17020 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_192
timestamp 1
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_203
timestamp 1636968456
transform 1 0 19780 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_215
timestamp 1636968456
transform 1 0 20884 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_227
timestamp 1636968456
transform 1 0 21988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_239
timestamp 1636968456
transform 1 0 23092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_270
timestamp 1
transform 1 0 25944 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_282
timestamp 1
transform 1 0 27048 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_301
timestamp 1
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1636968456
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 1636968456
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_333
timestamp 1
transform 1 0 31740 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_341
timestamp 1
transform 1 0 32476 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_354
timestamp 1
transform 1 0 33672 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_362
timestamp 1
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_371
timestamp 1
transform 1 0 35236 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_380
timestamp 1636968456
transform 1 0 36064 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_392
timestamp 1636968456
transform 1 0 37168 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_404
timestamp 1636968456
transform 1 0 38272 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_416
timestamp 1
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_421
timestamp 1
transform 1 0 39836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_432
timestamp 1
transform 1 0 40848 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_438
timestamp 1
transform 1 0 41400 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_463
timestamp 1
transform 1 0 43700 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1636968456
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1636968456
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1636968456
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_54
timestamp 1
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1636968456
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_69
timestamp 1
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_77
timestamp 1
transform 1 0 8188 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_86
timestamp 1
transform 1 0 9016 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_96
timestamp 1
transform 1 0 9936 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 1
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_113
timestamp 1
transform 1 0 11500 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_124
timestamp 1
transform 1 0 12512 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_135
timestamp 1
transform 1 0 13524 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_139
timestamp 1
transform 1 0 13892 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_146
timestamp 1636968456
transform 1 0 14536 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_158
timestamp 1
transform 1 0 15640 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_162
timestamp 1
transform 1 0 16008 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1636968456
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 1636968456
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 1636968456
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_205
timestamp 1
transform 1 0 19964 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_211
timestamp 1
transform 1 0 20516 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_225
timestamp 1
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_232
timestamp 1636968456
transform 1 0 22448 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_244
timestamp 1
transform 1 0 23552 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_257
timestamp 1636968456
transform 1 0 24748 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_269
timestamp 1
transform 1 0 25852 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1636968456
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_293
timestamp 1
transform 1 0 28060 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_301
timestamp 1
transform 1 0 28796 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_309
timestamp 1636968456
transform 1 0 29532 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_321
timestamp 1
transform 1 0 30636 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 1636968456
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 1636968456
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_361
timestamp 1636968456
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_373
timestamp 1636968456
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_385
timestamp 1
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 1
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_393
timestamp 1636968456
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_405
timestamp 1636968456
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_417
timestamp 1
transform 1 0 39468 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_425
timestamp 1
transform 1 0 40204 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_442
timestamp 1
transform 1 0 41768 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_449
timestamp 1636968456
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_461
timestamp 1
transform 1 0 43516 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1636968456
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_15
timestamp 1
transform 1 0 2484 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_24
timestamp 1
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_29
timestamp 1
transform 1 0 3772 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_35
timestamp 1
transform 1 0 4324 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_51
timestamp 1636968456
transform 1 0 5796 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_63
timestamp 1
transform 1 0 6900 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_75
timestamp 1
transform 1 0 8004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_85
timestamp 1
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_99
timestamp 1
transform 1 0 10212 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_108
timestamp 1636968456
transform 1 0 11040 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_120
timestamp 1
transform 1 0 12144 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_128
timestamp 1636968456
transform 1 0 12880 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_154
timestamp 1636968456
transform 1 0 15272 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_166
timestamp 1636968456
transform 1 0 16376 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_178
timestamp 1
transform 1 0 17480 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_186
timestamp 1
transform 1 0 18216 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 1
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_197
timestamp 1
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_205
timestamp 1
transform 1 0 19964 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_216
timestamp 1636968456
transform 1 0 20976 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_228
timestamp 1636968456
transform 1 0 22080 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_240
timestamp 1
transform 1 0 23184 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_249
timestamp 1
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1636968456
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_265
timestamp 1
transform 1 0 25484 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_276
timestamp 1
transform 1 0 26496 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_284
timestamp 1
transform 1 0 27232 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_290
timestamp 1636968456
transform 1 0 27784 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_302
timestamp 1
transform 1 0 28888 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_315
timestamp 1636968456
transform 1 0 30084 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_327
timestamp 1636968456
transform 1 0 31188 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_339
timestamp 1
transform 1 0 32292 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_347
timestamp 1
transform 1 0 33028 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_353
timestamp 1
transform 1 0 33580 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_360
timestamp 1
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_371
timestamp 1636968456
transform 1 0 35236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_383
timestamp 1
transform 1 0 36340 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_387
timestamp 1
transform 1 0 36708 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_393
timestamp 1
transform 1 0 37260 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_399
timestamp 1
transform 1 0 37812 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_409
timestamp 1
transform 1 0 38732 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_417
timestamp 1
transform 1 0 39468 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_450
timestamp 1636968456
transform 1 0 42504 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_462
timestamp 1
transform 1 0 43608 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_470
timestamp 1
transform 1 0 44344 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1636968456
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1636968456
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_27
timestamp 1
transform 1 0 3588 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_41
timestamp 1636968456
transform 1 0 4876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_53
timestamp 1
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_57
timestamp 1
transform 1 0 6348 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_75
timestamp 1636968456
transform 1 0 8004 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_87
timestamp 1
transform 1 0 9108 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_102
timestamp 1
transform 1 0 10488 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_110
timestamp 1
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1636968456
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_125
timestamp 1
transform 1 0 12604 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_133
timestamp 1
transform 1 0 13340 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_139
timestamp 1636968456
transform 1 0 13892 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_151
timestamp 1
transform 1 0 14996 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_159
timestamp 1
transform 1 0 15732 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1636968456
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1636968456
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 1636968456
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_205
timestamp 1
transform 1 0 19964 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_213
timestamp 1
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_221
timestamp 1
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_225
timestamp 1
transform 1 0 21804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_233
timestamp 1
transform 1 0 22540 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_247
timestamp 1
transform 1 0 23828 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_255
timestamp 1
transform 1 0 24564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_263
timestamp 1
transform 1 0 25300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_267
timestamp 1
transform 1 0 25668 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_281
timestamp 1
transform 1 0 26956 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_289
timestamp 1
transform 1 0 27692 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_297
timestamp 1636968456
transform 1 0 28428 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_309
timestamp 1
transform 1 0 29532 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_317
timestamp 1
transform 1 0 30268 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_328
timestamp 1
transform 1 0 31280 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_337
timestamp 1
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_346
timestamp 1636968456
transform 1 0 32936 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_369
timestamp 1636968456
transform 1 0 35052 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_381
timestamp 1
transform 1 0 36156 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_390
timestamp 1
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_393
timestamp 1636968456
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_405
timestamp 1
transform 1 0 38364 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_419
timestamp 1
transform 1 0 39652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_464
timestamp 1
transform 1 0 43792 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_468
timestamp 1
transform 1 0 44160 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1636968456
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1636968456
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1636968456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1636968456
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1636968456
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_65
timestamp 1
transform 1 0 7084 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_76
timestamp 1
transform 1 0 8096 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_85
timestamp 1
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_93
timestamp 1
transform 1 0 9660 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_108
timestamp 1636968456
transform 1 0 11040 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_120
timestamp 1
transform 1 0 12144 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_131
timestamp 1
transform 1 0 13156 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_141
timestamp 1
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_149
timestamp 1
transform 1 0 14812 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_156
timestamp 1
transform 1 0 15456 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_168
timestamp 1
transform 1 0 16560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_176
timestamp 1
transform 1 0 17296 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_191
timestamp 1
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1636968456
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1636968456
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 1636968456
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_239
timestamp 1
transform 1 0 23092 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_247
timestamp 1
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1636968456
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1636968456
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 1636968456
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_289
timestamp 1
transform 1 0 27692 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 1
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_314
timestamp 1
transform 1 0 29992 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_322
timestamp 1
transform 1 0 30728 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_336
timestamp 1636968456
transform 1 0 32016 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_348
timestamp 1
transform 1 0 33120 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_356
timestamp 1
transform 1 0 33856 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_387
timestamp 1636968456
transform 1 0 36708 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_399
timestamp 1636968456
transform 1 0 37812 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_411
timestamp 1
transform 1 0 38916 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_419
timestamp 1
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_421
timestamp 1
transform 1 0 39836 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_445
timestamp 1
transform 1 0 42044 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_453
timestamp 1
transform 1 0 42780 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_463
timestamp 1
transform 1 0 43700 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1636968456
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1636968456
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1636968456
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1636968456
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1636968456
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_69
timestamp 1
transform 1 0 7452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_77
timestamp 1
transform 1 0 8188 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_88
timestamp 1
transform 1 0 9200 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_96
timestamp 1
transform 1 0 9936 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_103
timestamp 1
transform 1 0 10580 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_113
timestamp 1
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_121
timestamp 1636968456
transform 1 0 12236 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_133
timestamp 1
transform 1 0 13340 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_139
timestamp 1
transform 1 0 13892 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_145
timestamp 1636968456
transform 1 0 14444 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_157
timestamp 1
transform 1 0 15548 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_165
timestamp 1
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_169
timestamp 1
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_175
timestamp 1
transform 1 0 17204 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_188
timestamp 1636968456
transform 1 0 18400 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_200
timestamp 1
transform 1 0 19504 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_206
timestamp 1
transform 1 0 20056 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_218
timestamp 1
transform 1 0 21160 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_225
timestamp 1
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_239
timestamp 1636968456
transform 1 0 23092 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_251
timestamp 1636968456
transform 1 0 24196 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_263
timestamp 1
transform 1 0 25300 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_276
timestamp 1
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1636968456
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1636968456
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 1636968456
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_317
timestamp 1636968456
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 1
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_342
timestamp 1
transform 1 0 32568 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_350
timestamp 1636968456
transform 1 0 33304 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_362
timestamp 1636968456
transform 1 0 34408 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_374
timestamp 1636968456
transform 1 0 35512 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_386
timestamp 1
transform 1 0 36616 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 1636968456
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_405
timestamp 1
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_413
timestamp 1636968456
transform 1 0 39100 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_425
timestamp 1636968456
transform 1 0 40204 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_437
timestamp 1
transform 1 0 41308 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_465
timestamp 1
transform 1 0 43884 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1636968456
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1636968456
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1636968456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_41
timestamp 1
transform 1 0 4876 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_51
timestamp 1636968456
transform 1 0 5796 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_63
timestamp 1636968456
transform 1 0 6900 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_75
timestamp 1
transform 1 0 8004 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1636968456
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_97
timestamp 1
transform 1 0 10028 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_104
timestamp 1636968456
transform 1 0 10672 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_116
timestamp 1636968456
transform 1 0 11776 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_128
timestamp 1636968456
transform 1 0 12880 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1636968456
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_153
timestamp 1
transform 1 0 15180 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_161
timestamp 1
transform 1 0 15916 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_168
timestamp 1636968456
transform 1 0 16560 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_180
timestamp 1636968456
transform 1 0 17664 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_192
timestamp 1
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_203
timestamp 1
transform 1 0 19780 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_215
timestamp 1636968456
transform 1 0 20884 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_227
timestamp 1636968456
transform 1 0 21988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_239
timestamp 1
transform 1 0 23092 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_247
timestamp 1
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_253
timestamp 1
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_257
timestamp 1
transform 1 0 24748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_266
timestamp 1
transform 1 0 25576 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_274
timestamp 1636968456
transform 1 0 26312 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_286
timestamp 1
transform 1 0 27416 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_294
timestamp 1
transform 1 0 28152 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_305
timestamp 1
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_315
timestamp 1
transform 1 0 30084 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_326
timestamp 1
transform 1 0 31096 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_330
timestamp 1
transform 1 0 31464 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_337
timestamp 1
transform 1 0 32108 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_360
timestamp 1
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_365
timestamp 1
transform 1 0 34684 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_371
timestamp 1636968456
transform 1 0 35236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_383
timestamp 1
transform 1 0 36340 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_390
timestamp 1636968456
transform 1 0 36984 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_402
timestamp 1636968456
transform 1 0 38088 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_414
timestamp 1
transform 1 0 39192 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_421
timestamp 1
transform 1 0 39836 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_435
timestamp 1
transform 1 0 41124 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_439
timestamp 1
transform 1 0 41492 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_468
timestamp 1
transform 1 0 44160 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1636968456
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1636968456
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1636968456
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_39
timestamp 1
transform 1 0 4692 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_48
timestamp 1
transform 1 0 5520 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1636968456
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_69
timestamp 1
transform 1 0 7452 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_78
timestamp 1
transform 1 0 8280 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_84
timestamp 1
transform 1 0 8832 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_91
timestamp 1
transform 1 0 9476 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_97
timestamp 1
transform 1 0 10028 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_109
timestamp 1
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_113
timestamp 1
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_117
timestamp 1
transform 1 0 11868 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_124
timestamp 1
transform 1 0 12512 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_133
timestamp 1636968456
transform 1 0 13340 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_145
timestamp 1
transform 1 0 14444 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_153
timestamp 1
transform 1 0 15180 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_161
timestamp 1
transform 1 0 15916 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1636968456
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1636968456
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 1636968456
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 1636968456
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 1
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_230
timestamp 1
transform 1 0 22264 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_253
timestamp 1
transform 1 0 24380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_260
timestamp 1636968456
transform 1 0 25024 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_272
timestamp 1
transform 1 0 26128 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1636968456
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_293
timestamp 1
transform 1 0 28060 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_303
timestamp 1636968456
transform 1 0 28980 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_315
timestamp 1636968456
transform 1 0 30084 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_327
timestamp 1
transform 1 0 31188 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 1
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_337
timestamp 1
transform 1 0 32108 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_350
timestamp 1
transform 1 0 33304 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_354
timestamp 1
transform 1 0 33672 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_360
timestamp 1
transform 1 0 34224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_367
timestamp 1
transform 1 0 34868 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_371
timestamp 1
transform 1 0 35236 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_377
timestamp 1636968456
transform 1 0 35788 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_389
timestamp 1
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_400
timestamp 1
transform 1 0 37904 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_404
timestamp 1
transform 1 0 38272 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_419
timestamp 1
transform 1 0 39652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_427
timestamp 1
transform 1 0 40388 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_444
timestamp 1
transform 1 0 41952 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_457
timestamp 1636968456
transform 1 0 43148 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_469
timestamp 1
transform 1 0 44252 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1636968456
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1636968456
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1636968456
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1636968456
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1636968456
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_65
timestamp 1
transform 1 0 7084 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_78
timestamp 1
transform 1 0 8280 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1636968456
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_97
timestamp 1
transform 1 0 10028 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_118
timestamp 1
transform 1 0 11960 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_127
timestamp 1636968456
transform 1 0 12788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_141
timestamp 1
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_159
timestamp 1636968456
transform 1 0 15732 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_171
timestamp 1
transform 1 0 16836 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_177
timestamp 1
transform 1 0 17388 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_181
timestamp 1
transform 1 0 17756 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_194
timestamp 1
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1636968456
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_209
timestamp 1
transform 1 0 20332 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_217
timestamp 1
transform 1 0 21068 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_223
timestamp 1
transform 1 0 21620 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_230
timestamp 1636968456
transform 1 0 22264 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_242
timestamp 1
transform 1 0 23368 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_250
timestamp 1
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_253
timestamp 1
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_261
timestamp 1
transform 1 0 25116 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_268
timestamp 1
transform 1 0 25760 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_279
timestamp 1636968456
transform 1 0 26772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_291
timestamp 1636968456
transform 1 0 27876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_303
timestamp 1
transform 1 0 28980 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_315
timestamp 1
transform 1 0 30084 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_323
timestamp 1
transform 1 0 30820 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_337
timestamp 1
transform 1 0 32108 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_345
timestamp 1
transform 1 0 32844 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_352
timestamp 1636968456
transform 1 0 33488 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 1636968456
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 1636968456
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_389
timestamp 1
transform 1 0 36892 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_398
timestamp 1636968456
transform 1 0 37720 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_410
timestamp 1
transform 1 0 38824 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_418
timestamp 1
transform 1 0 39560 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_421
timestamp 1
transform 1 0 39836 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_429
timestamp 1
transform 1 0 40572 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_462
timestamp 1
transform 1 0 43608 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_468
timestamp 1
transform 1 0 44160 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1636968456
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1636968456
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1636968456
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1636968456
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1636968456
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_69
timestamp 1
transform 1 0 7452 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_80
timestamp 1636968456
transform 1 0 8464 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_92
timestamp 1636968456
transform 1 0 9568 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_104
timestamp 1
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1636968456
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_125
timestamp 1
transform 1 0 12604 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_129
timestamp 1
transform 1 0 12972 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_136
timestamp 1636968456
transform 1 0 13616 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_148
timestamp 1
transform 1 0 14720 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_154
timestamp 1
transform 1 0 15272 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_160
timestamp 1
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1636968456
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 1636968456
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_193
timestamp 1
transform 1 0 18860 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_197
timestamp 1
transform 1 0 19228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_204
timestamp 1
transform 1 0 19872 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_216
timestamp 1
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_225
timestamp 1
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_233
timestamp 1636968456
transform 1 0 22540 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_245
timestamp 1636968456
transform 1 0 23644 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_269
timestamp 1
transform 1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_287
timestamp 1
transform 1 0 27508 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_295
timestamp 1
transform 1 0 28244 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1636968456
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 1636968456
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 1
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_343
timestamp 1636968456
transform 1 0 32660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_355
timestamp 1
transform 1 0 33764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_361
timestamp 1
transform 1 0 34316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_373
timestamp 1636968456
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_385
timestamp 1
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 1
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_399
timestamp 1636968456
transform 1 0 37812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_411
timestamp 1
transform 1 0 38916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_417
timestamp 1
transform 1 0 39468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_442
timestamp 1
transform 1 0 41768 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_465
timestamp 1
transform 1 0 43884 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1636968456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1636968456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1636968456
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_41
timestamp 1
transform 1 0 4876 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_49
timestamp 1
transform 1 0 5612 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_63
timestamp 1636968456
transform 1 0 6900 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_75
timestamp 1
transform 1 0 8004 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_85
timestamp 1
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_93
timestamp 1
transform 1 0 9660 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_101
timestamp 1636968456
transform 1 0 10396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_113
timestamp 1636968456
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_125
timestamp 1
transform 1 0 12604 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_129
timestamp 1
transform 1 0 12972 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_136
timestamp 1
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1636968456
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_153
timestamp 1
transform 1 0 15180 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_164
timestamp 1
transform 1 0 16192 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_172
timestamp 1
transform 1 0 16928 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_178
timestamp 1636968456
transform 1 0 17480 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_190
timestamp 1
transform 1 0 18584 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_197
timestamp 1
transform 1 0 19228 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1636968456
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_221
timestamp 1
transform 1 0 21436 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_225
timestamp 1
transform 1 0 21804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_232
timestamp 1636968456
transform 1 0 22448 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_244
timestamp 1
transform 1 0 23552 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_258
timestamp 1636968456
transform 1 0 24840 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_270
timestamp 1
transform 1 0 25944 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_286
timestamp 1636968456
transform 1 0 27416 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_298
timestamp 1
transform 1 0 28520 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_306
timestamp 1
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_315
timestamp 1
transform 1 0 30084 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_323
timestamp 1
transform 1 0 30820 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_329
timestamp 1
transform 1 0 31372 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_338
timestamp 1
transform 1 0 32200 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_352
timestamp 1636968456
transform 1 0 33488 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 1636968456
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_389
timestamp 1
transform 1 0 36892 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_397
timestamp 1636968456
transform 1 0 37628 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_409
timestamp 1
transform 1 0 38732 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_417
timestamp 1
transform 1 0 39468 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_452
timestamp 1636968456
transform 1 0 42688 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_464
timestamp 1
transform 1 0 43792 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_468
timestamp 1
transform 1 0 44160 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1636968456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1636968456
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1636968456
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1636968456
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_63
timestamp 1636968456
transform 1 0 6900 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_80
timestamp 1636968456
transform 1 0 8464 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_92
timestamp 1
transform 1 0 9568 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_100
timestamp 1
transform 1 0 10304 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_107
timestamp 1
transform 1 0 10948 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1636968456
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_125
timestamp 1
transform 1 0 12604 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_137
timestamp 1
transform 1 0 13708 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_145
timestamp 1
transform 1 0 14444 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_159
timestamp 1
transform 1 0 15732 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_166
timestamp 1
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1636968456
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_181
timestamp 1
transform 1 0 17756 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_189
timestamp 1
transform 1 0 18492 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_201
timestamp 1
transform 1 0 19596 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_209
timestamp 1
transform 1 0 20332 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_215
timestamp 1
transform 1 0 20884 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1636968456
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_237
timestamp 1
transform 1 0 22908 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_246
timestamp 1
transform 1 0 23736 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_252
timestamp 1
transform 1 0 24288 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_259
timestamp 1636968456
transform 1 0 24932 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_271
timestamp 1
transform 1 0 26036 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_292
timestamp 1
transform 1 0 27968 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_300
timestamp 1
transform 1 0 28704 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_306
timestamp 1
transform 1 0 29256 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_314
timestamp 1636968456
transform 1 0 29992 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_326
timestamp 1
transform 1 0 31096 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_334
timestamp 1
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_337
timestamp 1
transform 1 0 32108 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_348
timestamp 1636968456
transform 1 0 33120 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_360
timestamp 1636968456
transform 1 0 34224 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_372
timestamp 1636968456
transform 1 0 35328 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_384
timestamp 1
transform 1 0 36432 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_390
timestamp 1
transform 1 0 36984 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_398
timestamp 1636968456
transform 1 0 37720 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_410
timestamp 1636968456
transform 1 0 38824 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_422
timestamp 1636968456
transform 1 0 39928 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_434
timestamp 1
transform 1 0 41032 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_463
timestamp 1
transform 1 0 43700 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1636968456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1636968456
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1636968456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1636968456
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1636968456
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1636968456
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_90
timestamp 1
transform 1 0 9384 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_98
timestamp 1
transform 1 0 10120 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_113
timestamp 1636968456
transform 1 0 11500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_125
timestamp 1636968456
transform 1 0 12604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_137
timestamp 1
transform 1 0 13708 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1636968456
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1636968456
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1636968456
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_177
timestamp 1
transform 1 0 17388 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_191
timestamp 1
transform 1 0 18676 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1636968456
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 1636968456
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 1636968456
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_233
timestamp 1
transform 1 0 22540 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_243
timestamp 1
transform 1 0 23460 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1636968456
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1636968456
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_277
timestamp 1
transform 1 0 26588 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_293
timestamp 1
transform 1 0 28060 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1636968456
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_321
timestamp 1
transform 1 0 30636 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_332
timestamp 1
transform 1 0 31648 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_340
timestamp 1
transform 1 0 32384 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_350
timestamp 1636968456
transform 1 0 33304 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_362
timestamp 1
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_365
timestamp 1
transform 1 0 34684 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_373
timestamp 1
transform 1 0 35420 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_414
timestamp 1
transform 1 0 39192 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_421
timestamp 1636968456
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_433
timestamp 1
transform 1 0 40940 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_452
timestamp 1636968456
transform 1 0 42688 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_464
timestamp 1
transform 1 0 43792 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_472
timestamp 1
transform 1 0 44528 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1636968456
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1636968456
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1636968456
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1636968456
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_57
timestamp 1
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_65
timestamp 1
transform 1 0 7084 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_72
timestamp 1636968456
transform 1 0 7728 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_84
timestamp 1636968456
transform 1 0 8832 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_96
timestamp 1
transform 1 0 9936 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_108
timestamp 1
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_119
timestamp 1
transform 1 0 12052 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_127
timestamp 1
transform 1 0 12788 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_134
timestamp 1636968456
transform 1 0 13432 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_146
timestamp 1636968456
transform 1 0 14536 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_158
timestamp 1
transform 1 0 15640 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_166
timestamp 1
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_169
timestamp 1
transform 1 0 16652 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_180
timestamp 1636968456
transform 1 0 17664 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_192
timestamp 1
transform 1 0 18768 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_201
timestamp 1636968456
transform 1 0 19596 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_213
timestamp 1
transform 1 0 20700 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_221
timestamp 1
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_236
timestamp 1636968456
transform 1 0 22816 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_248
timestamp 1
transform 1 0 23920 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_254
timestamp 1
transform 1 0 24472 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 1636968456
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_273
timestamp 1
transform 1 0 26220 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1636968456
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_298
timestamp 1
transform 1 0 28520 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_308
timestamp 1636968456
transform 1 0 29440 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_320
timestamp 1
transform 1 0 30544 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_332
timestamp 1
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 1636968456
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_349
timestamp 1
transform 1 0 33212 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_353
timestamp 1
transform 1 0 33580 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_359
timestamp 1
transform 1 0 34132 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_381
timestamp 1
transform 1 0 36156 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_389
timestamp 1
transform 1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_400
timestamp 1
transform 1 0 37904 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_430
timestamp 1636968456
transform 1 0 40664 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_442
timestamp 1
transform 1 0 41768 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_449
timestamp 1636968456
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_461
timestamp 1
transform 1 0 43516 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1636968456
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1636968456
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1636968456
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1636968456
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1636968456
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1636968456
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_91
timestamp 1636968456
transform 1 0 9476 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_103
timestamp 1
transform 1 0 10580 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_111
timestamp 1
transform 1 0 11316 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_118
timestamp 1636968456
transform 1 0 11960 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_130
timestamp 1
transform 1 0 13064 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_134
timestamp 1
transform 1 0 13432 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_147
timestamp 1636968456
transform 1 0 14628 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_159
timestamp 1
transform 1 0 15732 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_175
timestamp 1
transform 1 0 17204 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_186
timestamp 1
transform 1 0 18216 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_190
timestamp 1
transform 1 0 18584 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_208
timestamp 1
transform 1 0 20240 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_220
timestamp 1636968456
transform 1 0 21344 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_232
timestamp 1636968456
transform 1 0 22448 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_244
timestamp 1
transform 1 0 23552 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1636968456
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_265
timestamp 1
transform 1 0 25484 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_274
timestamp 1
transform 1 0 26312 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_283
timestamp 1636968456
transform 1 0 27140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_295
timestamp 1
transform 1 0 28244 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_305
timestamp 1
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_309
timestamp 1
transform 1 0 29532 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_313
timestamp 1
transform 1 0 29900 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_319
timestamp 1636968456
transform 1 0 30452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_331
timestamp 1
transform 1 0 31556 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_338
timestamp 1
transform 1 0 32200 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_344
timestamp 1636968456
transform 1 0 32752 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_356
timestamp 1
transform 1 0 33856 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_365
timestamp 1
transform 1 0 34684 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_369
timestamp 1
transform 1 0 35052 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_375
timestamp 1
transform 1 0 35604 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_379
timestamp 1
transform 1 0 35972 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_404
timestamp 1636968456
transform 1 0 38272 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_416
timestamp 1
transform 1 0 39376 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_421
timestamp 1636968456
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_433
timestamp 1636968456
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_445
timestamp 1636968456
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_457
timestamp 1636968456
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_469
timestamp 1
transform 1 0 44252 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1636968456
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1636968456
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1636968456
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1636968456
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1636968456
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1636968456
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_81
timestamp 1
transform 1 0 8556 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_89
timestamp 1
transform 1 0 9292 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_98
timestamp 1636968456
transform 1 0 10120 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_110
timestamp 1
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1636968456
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_125
timestamp 1
transform 1 0 12604 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_129
timestamp 1
transform 1 0 12972 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_135
timestamp 1636968456
transform 1 0 13524 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_147
timestamp 1636968456
transform 1 0 14628 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_164
timestamp 1
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_169
timestamp 1
transform 1 0 16652 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_181
timestamp 1
transform 1 0 17756 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_195
timestamp 1636968456
transform 1 0 19044 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_207
timestamp 1636968456
transform 1 0 20148 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_219
timestamp 1
transform 1 0 21252 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_225
timestamp 1
transform 1 0 21804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_231
timestamp 1
transform 1 0 22356 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_237
timestamp 1
transform 1 0 22908 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_241
timestamp 1
transform 1 0 23276 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_255
timestamp 1636968456
transform 1 0 24564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_267
timestamp 1636968456
transform 1 0 25668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1636968456
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_293
timestamp 1
transform 1 0 28060 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_301
timestamp 1
transform 1 0 28796 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_310
timestamp 1
transform 1 0 29624 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_331
timestamp 1
transform 1 0 31556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_343
timestamp 1636968456
transform 1 0 32660 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_355
timestamp 1636968456
transform 1 0 33764 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_367
timestamp 1
transform 1 0 34868 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_373
timestamp 1636968456
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_385
timestamp 1
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 1
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_393
timestamp 1636968456
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_405
timestamp 1636968456
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_417
timestamp 1636968456
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_429
timestamp 1636968456
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_441
timestamp 1
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_447
timestamp 1
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_449
timestamp 1636968456
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_461
timestamp 1636968456
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1636968456
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1636968456
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1636968456
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1636968456
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1636968456
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1636968456
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1636968456
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1636968456
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_109
timestamp 1
transform 1 0 11132 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_117
timestamp 1
transform 1 0 11868 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_126
timestamp 1636968456
transform 1 0 12696 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_138
timestamp 1
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_141
timestamp 1
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_150
timestamp 1636968456
transform 1 0 14904 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_162
timestamp 1636968456
transform 1 0 16008 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_174
timestamp 1636968456
transform 1 0 17112 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_186
timestamp 1
transform 1 0 18216 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_194
timestamp 1
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1636968456
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_209
timestamp 1
transform 1 0 20332 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_217
timestamp 1636968456
transform 1 0 21068 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_229
timestamp 1
transform 1 0 22172 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_236
timestamp 1
transform 1 0 22816 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_242
timestamp 1
transform 1 0 23368 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_249
timestamp 1
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1636968456
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_265
timestamp 1
transform 1 0 25484 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_282
timestamp 1
transform 1 0 27048 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_290
timestamp 1
transform 1 0 27784 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_303
timestamp 1
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1636968456
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1636968456
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 1636968456
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_345
timestamp 1
transform 1 0 32844 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_351
timestamp 1
transform 1 0 33396 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_360
timestamp 1
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_365
timestamp 1
transform 1 0 34684 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_373
timestamp 1
transform 1 0 35420 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_382
timestamp 1636968456
transform 1 0 36248 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_394
timestamp 1636968456
transform 1 0 37352 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_406
timestamp 1636968456
transform 1 0 38456 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_418
timestamp 1
transform 1 0 39560 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_421
timestamp 1636968456
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_433
timestamp 1636968456
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_445
timestamp 1636968456
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_457
timestamp 1636968456
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_469
timestamp 1
transform 1 0 44252 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1636968456
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1636968456
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1636968456
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1636968456
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1636968456
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1636968456
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1636968456
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1636968456
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_105
timestamp 1
transform 1 0 10764 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1636968456
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1636968456
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_137
timestamp 1
transform 1 0 13708 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_145
timestamp 1
transform 1 0 14444 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_157
timestamp 1
transform 1 0 15548 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_165
timestamp 1
transform 1 0 16284 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1636968456
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 1636968456
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_193
timestamp 1
transform 1 0 18860 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_216
timestamp 1
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_225
timestamp 1
transform 1 0 21804 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_234
timestamp 1636968456
transform 1 0 22632 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_246
timestamp 1
transform 1 0 23736 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_252
timestamp 1
transform 1 0 24288 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_258
timestamp 1636968456
transform 1 0 24840 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_270
timestamp 1
transform 1 0 25944 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_277
timestamp 1
transform 1 0 26588 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1636968456
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_297
timestamp 1
transform 1 0 28428 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_303
timestamp 1636968456
transform 1 0 28980 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_315
timestamp 1
transform 1 0 30084 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_323
timestamp 1
transform 1 0 30820 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_337
timestamp 1
transform 1 0 32108 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_358
timestamp 1636968456
transform 1 0 34040 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_370
timestamp 1
transform 1 0 35144 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_378
timestamp 1636968456
transform 1 0 35880 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_390
timestamp 1
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_393
timestamp 1636968456
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_405
timestamp 1636968456
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_417
timestamp 1636968456
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_429
timestamp 1636968456
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_441
timestamp 1
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_447
timestamp 1
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_449
timestamp 1636968456
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_461
timestamp 1636968456
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1636968456
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1636968456
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1636968456
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1636968456
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1636968456
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1636968456
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1636968456
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_97
timestamp 1
transform 1 0 10028 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_105
timestamp 1
transform 1 0 10764 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_113
timestamp 1636968456
transform 1 0 11500 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_125
timestamp 1
transform 1 0 12604 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_136
timestamp 1
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1636968456
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1636968456
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_165
timestamp 1
transform 1 0 16284 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_173
timestamp 1
transform 1 0 17020 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_181
timestamp 1636968456
transform 1 0 17756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_193
timestamp 1
transform 1 0 18860 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_208
timestamp 1636968456
transform 1 0 20240 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_220
timestamp 1
transform 1 0 21344 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_231
timestamp 1
transform 1 0 22356 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_235
timestamp 1
transform 1 0 22724 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_241
timestamp 1
transform 1 0 23276 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_245
timestamp 1
transform 1 0 23644 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1636968456
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_265
timestamp 1
transform 1 0 25484 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_282
timestamp 1
transform 1 0 27048 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1636968456
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_321
timestamp 1
transform 1 0 30636 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_325
timestamp 1
transform 1 0 31004 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_331
timestamp 1636968456
transform 1 0 31556 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_343
timestamp 1636968456
transform 1 0 32660 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_355
timestamp 1
transform 1 0 33764 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 1
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 1636968456
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_377
timestamp 1636968456
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_389
timestamp 1636968456
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_401
timestamp 1636968456
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_413
timestamp 1
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_419
timestamp 1
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_421
timestamp 1636968456
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_433
timestamp 1636968456
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_445
timestamp 1636968456
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_457
timestamp 1636968456
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_469
timestamp 1
transform 1 0 44252 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1636968456
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1636968456
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1636968456
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1636968456
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1636968456
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1636968456
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1636968456
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1636968456
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1636968456
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_125
timestamp 1
transform 1 0 12604 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_138
timestamp 1636968456
transform 1 0 13800 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_150
timestamp 1
transform 1 0 14904 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_164
timestamp 1
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1636968456
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 1636968456
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_193
timestamp 1
transform 1 0 18860 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_197
timestamp 1
transform 1 0 19228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_203
timestamp 1636968456
transform 1 0 19780 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_215
timestamp 1
transform 1 0 20884 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_230
timestamp 1
transform 1 0 22264 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_238
timestamp 1
transform 1 0 23000 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1636968456
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_261
timestamp 1
transform 1 0 25116 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_267
timestamp 1
transform 1 0 25668 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_278
timestamp 1
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1636968456
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_293
timestamp 1
transform 1 0 28060 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_312
timestamp 1636968456
transform 1 0 29808 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_324
timestamp 1
transform 1 0 30912 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_333
timestamp 1
transform 1 0 31740 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1636968456
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1636968456
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_361
timestamp 1636968456
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_373
timestamp 1636968456
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_385
timestamp 1
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 1
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 1636968456
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_405
timestamp 1636968456
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_417
timestamp 1636968456
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_429
timestamp 1636968456
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_441
timestamp 1
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_447
timestamp 1
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_449
timestamp 1636968456
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_461
timestamp 1636968456
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1636968456
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1636968456
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1636968456
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1636968456
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1636968456
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1636968456
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1636968456
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1636968456
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1636968456
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1636968456
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1636968456
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1636968456
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1636968456
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1636968456
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1636968456
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1636968456
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1636968456
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1636968456
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1636968456
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1636968456
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1636968456
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_296
timestamp 1636968456
transform 1 0 28336 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_317
timestamp 1
transform 1 0 30268 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 1636968456
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 1
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 1636968456
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_377
timestamp 1636968456
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_389
timestamp 1636968456
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_401
timestamp 1636968456
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_413
timestamp 1
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_419
timestamp 1
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_421
timestamp 1636968456
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_433
timestamp 1636968456
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_445
timestamp 1636968456
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_457
timestamp 1636968456
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_469
timestamp 1
transform 1 0 44252 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1636968456
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1636968456
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1636968456
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1636968456
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1636968456
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1636968456
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1636968456
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 1636968456
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 1
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1636968456
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1636968456
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1636968456
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1636968456
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1636968456
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1636968456
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1636968456
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1636968456
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_225
timestamp 1
transform 1 0 21804 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_233
timestamp 1
transform 1 0 22540 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_250
timestamp 1636968456
transform 1 0 24104 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_262
timestamp 1
transform 1 0 25208 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_270
timestamp 1
transform 1 0 25944 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_296
timestamp 1
transform 1 0 28336 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_300
timestamp 1
transform 1 0 28704 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_325
timestamp 1
transform 1 0 31004 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_333
timestamp 1
transform 1 0 31740 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1636968456
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1636968456
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_361
timestamp 1636968456
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_373
timestamp 1636968456
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_385
timestamp 1
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_391
timestamp 1
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 1636968456
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_405
timestamp 1636968456
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_417
timestamp 1636968456
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_429
timestamp 1636968456
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_441
timestamp 1
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_447
timestamp 1
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_449
timestamp 1636968456
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_461
timestamp 1636968456
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1636968456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1636968456
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1636968456
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1636968456
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1636968456
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1636968456
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1636968456
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1636968456
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1636968456
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1636968456
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1636968456
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1636968456
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1636968456
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1636968456
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1636968456
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1636968456
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_261
timestamp 1
transform 1 0 25116 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_283
timestamp 1
transform 1 0 27140 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_303
timestamp 1
transform 1 0 28980 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_317
timestamp 1636968456
transform 1 0 30268 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_329
timestamp 1636968456
transform 1 0 31372 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_341
timestamp 1636968456
transform 1 0 32476 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_353
timestamp 1
transform 1 0 33580 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_361
timestamp 1
transform 1 0 34316 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1636968456
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 1636968456
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 1636968456
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_401
timestamp 1636968456
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_413
timestamp 1
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_419
timestamp 1
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_421
timestamp 1636968456
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_433
timestamp 1636968456
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_445
timestamp 1636968456
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_457
timestamp 1636968456
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_469
timestamp 1
transform 1 0 44252 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1636968456
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1636968456
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1636968456
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1636968456
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1636968456
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1636968456
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1636968456
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1636968456
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1636968456
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1636968456
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1636968456
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1636968456
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1636968456
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1636968456
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1636968456
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 1636968456
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 1
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_225
timestamp 1
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_229
timestamp 1
transform 1 0 22172 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_246
timestamp 1
transform 1 0 23736 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1636968456
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1636968456
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1636968456
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1636968456
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 1636968456
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 1636968456
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 1
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 1
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 1636968456
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_405
timestamp 1636968456
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_417
timestamp 1636968456
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_429
timestamp 1636968456
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_441
timestamp 1
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_447
timestamp 1
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_449
timestamp 1636968456
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_461
timestamp 1636968456
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1636968456
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1636968456
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1636968456
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1636968456
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1636968456
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1636968456
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1636968456
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1636968456
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1636968456
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1636968456
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1636968456
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1636968456
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1636968456
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 1636968456
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 1
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1636968456
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1636968456
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_221
timestamp 1
transform 1 0 21436 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_241
timestamp 1
transform 1 0 23276 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_249
timestamp 1
transform 1 0 24012 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_261
timestamp 1636968456
transform 1 0 25116 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_273
timestamp 1636968456
transform 1 0 26220 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_285
timestamp 1636968456
transform 1 0 27324 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_297
timestamp 1
transform 1 0 28428 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_305
timestamp 1
transform 1 0 29164 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1636968456
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1636968456
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1636968456
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1636968456
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 1
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1636968456
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1636968456
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1636968456
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_401
timestamp 1636968456
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_413
timestamp 1
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_419
timestamp 1
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_421
timestamp 1636968456
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_433
timestamp 1636968456
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_445
timestamp 1636968456
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_457
timestamp 1636968456
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_469
timestamp 1
transform 1 0 44252 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1636968456
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1636968456
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1636968456
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1636968456
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1636968456
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1636968456
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1636968456
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1636968456
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1636968456
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1636968456
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1636968456
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1636968456
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1636968456
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1636968456
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1636968456
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1636968456
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_225
timestamp 1
transform 1 0 21804 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_229
timestamp 1
transform 1 0 22172 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_238
timestamp 1636968456
transform 1 0 23000 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_250
timestamp 1636968456
transform 1 0 24104 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_262
timestamp 1636968456
transform 1 0 25208 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_274
timestamp 1
transform 1 0 26312 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1636968456
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1636968456
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1636968456
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1636968456
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 1
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1636968456
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1636968456
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 1636968456
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 1636968456
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 1
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 1
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1636968456
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_405
timestamp 1636968456
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_417
timestamp 1636968456
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_429
timestamp 1636968456
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_441
timestamp 1
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_447
timestamp 1
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_449
timestamp 1636968456
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_461
timestamp 1636968456
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1636968456
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1636968456
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1636968456
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1636968456
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1636968456
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1636968456
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1636968456
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1636968456
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 1636968456
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 1636968456
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 1
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 1
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1636968456
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1636968456
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 1636968456
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 1636968456
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 1
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 1
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1636968456
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1636968456
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 1636968456
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_233
timestamp 1636968456
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 1
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 1
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1636968456
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1636968456
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 1636968456
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 1636968456
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 1
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 1
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1636968456
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1636968456
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 1636968456
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 1636968456
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 1
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 1
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1636968456
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1636968456
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1636968456
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_401
timestamp 1636968456
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_413
timestamp 1
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_419
timestamp 1
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_421
timestamp 1636968456
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_433
timestamp 1636968456
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_445
timestamp 1636968456
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_457
timestamp 1636968456
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_469
timestamp 1
transform 1 0 44252 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1636968456
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1636968456
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1636968456
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1636968456
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1636968456
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1636968456
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1636968456
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 1636968456
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 1
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1636968456
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1636968456
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1636968456
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1636968456
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 1
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1636968456
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1636968456
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1636968456
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 1636968456
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 1
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 1
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 1636968456
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_237
timestamp 1636968456
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_249
timestamp 1636968456
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_261
timestamp 1636968456
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_273
timestamp 1
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 1
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 1636968456
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 1636968456
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 1636968456
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 1636968456
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 1
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1636968456
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 1636968456
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 1636968456
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 1636968456
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 1
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 1
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 1636968456
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_405
timestamp 1636968456
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_417
timestamp 1636968456
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_429
timestamp 1636968456
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_441
timestamp 1
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_447
timestamp 1
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_449
timestamp 1636968456
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_461
timestamp 1636968456
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1636968456
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1636968456
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1636968456
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1636968456
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_53
timestamp 1
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_57
timestamp 1636968456
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_69
timestamp 1636968456
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_81
timestamp 1
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1636968456
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1636968456
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_109
timestamp 1
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_113
timestamp 1636968456
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_125
timestamp 1636968456
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_137
timestamp 1
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1636968456
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1636968456
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_165
timestamp 1
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_169
timestamp 1636968456
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_181
timestamp 1636968456
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_193
timestamp 1
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1636968456
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 1636968456
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_221
timestamp 1
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_225
timestamp 1
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_233
timestamp 1
transform 1 0 22540 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_240
timestamp 1
transform 1 0 23184 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_247
timestamp 1
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 1
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_253
timestamp 1
transform 1 0 24380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_261
timestamp 1
transform 1 0 25116 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_268
timestamp 1
transform 1 0 25760 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_275
timestamp 1
transform 1 0 26404 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_279
timestamp 1
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_281
timestamp 1
transform 1 0 26956 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_289
timestamp 1
transform 1 0 27692 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_296
timestamp 1636968456
transform 1 0 28336 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1636968456
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_333
timestamp 1
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_343
timestamp 1636968456
transform 1 0 32660 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_355
timestamp 1
transform 1 0 33764 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 1
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1636968456
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1636968456
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_389
timestamp 1
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_393
timestamp 1636968456
transform 1 0 37260 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_405
timestamp 1636968456
transform 1 0 38364 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_417
timestamp 1
transform 1 0 39468 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_421
timestamp 1636968456
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_433
timestamp 1636968456
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_445
timestamp 1
transform 1 0 42044 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_449
timestamp 1636968456
transform 1 0 42412 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_461
timestamp 1636968456
transform 1 0 43516 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 43792 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform -1 0 43332 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 43240 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 42504 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform 1 0 42964 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform -1 0 26220 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform -1 0 43148 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 43792 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform -1 0 43148 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform -1 0 43148 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform 1 0 42964 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform -1 0 42044 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform -1 0 27692 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform -1 0 43148 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform -1 0 43884 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 25116 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 41584 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform -1 0 24104 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform -1 0 43700 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform -1 0 32844 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform -1 0 40664 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform -1 0 30268 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform -1 0 39468 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform 1 0 22264 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform -1 0 40388 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 29164 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform -1 0 43976 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform -1 0 31004 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform -1 0 43148 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform -1 0 38732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform -1 0 37996 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1
transform -1 0 40940 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform -1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform -1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform -1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1
transform -1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1
transform 1 0 44344 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap46
timestamp 1
transform 1 0 8740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap47
timestamp 1
transform -1 0 29072 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap48
timestamp 1
transform -1 0 28428 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap51
timestamp 1
transform -1 0 7544 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap66
timestamp 1
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap77
timestamp 1
transform -1 0 2576 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap102
timestamp 1
transform -1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap109
timestamp 1
transform -1 0 5704 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap118
timestamp 1
transform -1 0 9936 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1
transform 1 0 44252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 1
transform -1 0 26404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1
transform 1 0 44252 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1
transform 1 0 44252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1
transform 1 0 44252 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1
transform 1 0 44252 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1
transform -1 0 28336 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1
transform 1 0 44252 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1
transform 1 0 44252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1
transform 1 0 44252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1
transform -1 0 23828 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1
transform 1 0 44252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1
transform 1 0 44252 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1
transform 1 0 44252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1
transform 1 0 44252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1
transform 1 0 44252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1
transform 1 0 44252 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1
transform 1 0 44252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1
transform 1 0 32108 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1
transform 1 0 44252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1
transform 1 0 44252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1
transform 1 0 44252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1
transform 1 0 29532 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1
transform 1 0 44252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1
transform 1 0 44252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1
transform -1 0 22540 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1
transform -1 0 25760 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1
transform 1 0 44252 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1
transform 1 0 44252 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1
transform 1 0 44252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1
transform -1 0 30636 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1
transform -1 0 23184 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_65
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 44896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_66
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 44896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_67
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 44896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_68
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 44896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_69
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 44896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_70
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 44896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_71
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 44896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_72
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 44896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_73
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 44896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_74
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 44896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_75
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 44896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_76
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 44896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_77
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 44896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_78
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 44896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_79
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 44896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_80
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 44896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_81
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 44896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_82
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 44896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_83
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 44896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_84
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 44896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_85
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 44896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_86
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 44896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_87
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 44896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_88
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 44896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_89
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 44896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_90
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 44896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_91
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 44896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_92
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 44896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_93
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 44896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_94
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 44896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_95
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 44896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_96
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 44896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_97
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 44896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_98
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 44896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_99
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 44896 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_100
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 44896 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_101
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 44896 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_102
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 44896 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_103
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 44896 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_104
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1
transform -1 0 44896 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_105
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1
transform -1 0 44896 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_106
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1
transform -1 0 44896 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_107
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1
transform -1 0 44896 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_108
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1
transform -1 0 44896 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_109
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1
transform -1 0 44896 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_110
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1
transform -1 0 44896 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_111
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1
transform -1 0 44896 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_112
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1
transform -1 0 44896 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_113
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1
transform -1 0 44896 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_114
timestamp 1
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1
transform -1 0 44896 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_115
timestamp 1
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1
transform -1 0 44896 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_116
timestamp 1
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1
transform -1 0 44896 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_117
timestamp 1
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1
transform -1 0 44896 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_118
timestamp 1
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1
transform -1 0 44896 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_119
timestamp 1
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1
transform -1 0 44896 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_120
timestamp 1
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1
transform -1 0 44896 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_121
timestamp 1
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 1
transform -1 0 44896 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_122
timestamp 1
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 1
transform -1 0 44896 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_123
timestamp 1
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 1
transform -1 0 44896 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_124
timestamp 1
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 1
transform -1 0 44896 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_125
timestamp 1
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 1
transform -1 0 44896 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_126
timestamp 1
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 1
transform -1 0 44896 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_127
timestamp 1
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 1
transform -1 0 44896 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_128
timestamp 1
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 1
transform -1 0 44896 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_129
timestamp 1
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 1
transform -1 0 44896 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_130
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_131
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_132
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_133
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_134
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_135
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_136
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_137
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_138
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_139
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_140
timestamp 1
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_141
timestamp 1
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_142
timestamp 1
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_143
timestamp 1
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_144
timestamp 1
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_145
timestamp 1
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_146
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_147
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_148
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_149
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_150
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_151
timestamp 1
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_152
timestamp 1
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_153
timestamp 1
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_154
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_155
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_156
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_157
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_158
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_159
timestamp 1
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_160
timestamp 1
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_161
timestamp 1
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_162
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_163
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_164
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_165
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_166
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_167
timestamp 1
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_168
timestamp 1
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_169
timestamp 1
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_170
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_171
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_172
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_173
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_174
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_175
timestamp 1
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_176
timestamp 1
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_177
timestamp 1
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_178
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_179
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_180
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_181
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_182
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_183
timestamp 1
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_184
timestamp 1
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_185
timestamp 1
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_186
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_187
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_188
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_189
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_190
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_191
timestamp 1
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_192
timestamp 1
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_193
timestamp 1
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_194
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_195
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_196
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_197
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_198
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_199
timestamp 1
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_200
timestamp 1
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_201
timestamp 1
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_202
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_203
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_204
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_205
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_206
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_207
timestamp 1
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_208
timestamp 1
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_209
timestamp 1
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_210
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_211
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_212
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_213
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_214
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_215
timestamp 1
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_216
timestamp 1
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_217
timestamp 1
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_218
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_219
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_220
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_221
timestamp 1
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_222
timestamp 1
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_223
timestamp 1
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_224
timestamp 1
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_225
timestamp 1
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_226
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_227
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_228
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_229
timestamp 1
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_230
timestamp 1
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_231
timestamp 1
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_232
timestamp 1
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_233
timestamp 1
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_234
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_235
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_236
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_237
timestamp 1
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_238
timestamp 1
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_239
timestamp 1
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_240
timestamp 1
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_241
timestamp 1
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_242
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_243
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_244
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_245
timestamp 1
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_246
timestamp 1
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_247
timestamp 1
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_248
timestamp 1
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_249
timestamp 1
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_250
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_251
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_252
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_253
timestamp 1
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_254
timestamp 1
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_255
timestamp 1
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_256
timestamp 1
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_257
timestamp 1
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_258
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_259
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_260
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_261
timestamp 1
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_262
timestamp 1
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_263
timestamp 1
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_264
timestamp 1
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_265
timestamp 1
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_266
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_267
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_268
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_269
timestamp 1
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_270
timestamp 1
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_271
timestamp 1
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_272
timestamp 1
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_273
timestamp 1
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_274
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_275
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_276
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_277
timestamp 1
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_278
timestamp 1
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_279
timestamp 1
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_280
timestamp 1
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_281
timestamp 1
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_282
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_283
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_284
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_285
timestamp 1
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_286
timestamp 1
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_287
timestamp 1
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_288
timestamp 1
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_289
timestamp 1
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_290
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_291
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_292
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_293
timestamp 1
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_294
timestamp 1
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_295
timestamp 1
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_296
timestamp 1
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_297
timestamp 1
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_298
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_299
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_300
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_301
timestamp 1
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_302
timestamp 1
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_303
timestamp 1
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_304
timestamp 1
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_305
timestamp 1
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_306
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_307
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_308
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_309
timestamp 1
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_310
timestamp 1
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_311
timestamp 1
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_312
timestamp 1
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_313
timestamp 1
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_314
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_315
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_316
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_317
timestamp 1
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_318
timestamp 1
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_319
timestamp 1
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_320
timestamp 1
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_321
timestamp 1
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_322
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_323
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_324
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_325
timestamp 1
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_326
timestamp 1
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_327
timestamp 1
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_328
timestamp 1
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_329
timestamp 1
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_330
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_331
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_332
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_333
timestamp 1
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_334
timestamp 1
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_335
timestamp 1
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_336
timestamp 1
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_337
timestamp 1
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_338
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_339
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_340
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_341
timestamp 1
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_342
timestamp 1
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_343
timestamp 1
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_344
timestamp 1
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_345
timestamp 1
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_346
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_347
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_348
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_349
timestamp 1
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_350
timestamp 1
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_351
timestamp 1
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_352
timestamp 1
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_353
timestamp 1
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_354
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_355
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_356
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_357
timestamp 1
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_358
timestamp 1
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_359
timestamp 1
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_360
timestamp 1
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_361
timestamp 1
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_362
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_363
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_364
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_365
timestamp 1
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_366
timestamp 1
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_367
timestamp 1
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_368
timestamp 1
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_369
timestamp 1
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_370
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_371
timestamp 1
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_372
timestamp 1
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_373
timestamp 1
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_374
timestamp 1
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_375
timestamp 1
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_376
timestamp 1
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_377
timestamp 1
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_378
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_379
timestamp 1
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_380
timestamp 1
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_381
timestamp 1
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_382
timestamp 1
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_383
timestamp 1
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_384
timestamp 1
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_385
timestamp 1
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_386
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_387
timestamp 1
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_388
timestamp 1
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_389
timestamp 1
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_390
timestamp 1
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_391
timestamp 1
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_392
timestamp 1
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_393
timestamp 1
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_394
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_395
timestamp 1
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_396
timestamp 1
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_397
timestamp 1
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_398
timestamp 1
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_399
timestamp 1
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_400
timestamp 1
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_401
timestamp 1
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_402
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_403
timestamp 1
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_404
timestamp 1
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_405
timestamp 1
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_406
timestamp 1
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_407
timestamp 1
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_408
timestamp 1
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_409
timestamp 1
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_410
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_411
timestamp 1
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_412
timestamp 1
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_413
timestamp 1
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_414
timestamp 1
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_415
timestamp 1
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_416
timestamp 1
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_417
timestamp 1
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_418
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_419
timestamp 1
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_420
timestamp 1
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_421
timestamp 1
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_422
timestamp 1
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_423
timestamp 1
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_424
timestamp 1
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_425
timestamp 1
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_426
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_427
timestamp 1
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_428
timestamp 1
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_429
timestamp 1
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_430
timestamp 1
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_431
timestamp 1
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_432
timestamp 1
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_433
timestamp 1
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_434
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_435
timestamp 1
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_436
timestamp 1
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_437
timestamp 1
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_438
timestamp 1
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_439
timestamp 1
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_440
timestamp 1
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_441
timestamp 1
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_442
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_443
timestamp 1
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_444
timestamp 1
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_445
timestamp 1
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_446
timestamp 1
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_447
timestamp 1
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_448
timestamp 1
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_449
timestamp 1
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_450
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_451
timestamp 1
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_452
timestamp 1
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_453
timestamp 1
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_454
timestamp 1
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_455
timestamp 1
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_456
timestamp 1
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_457
timestamp 1
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_458
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_459
timestamp 1
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_460
timestamp 1
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_461
timestamp 1
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_462
timestamp 1
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_463
timestamp 1
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_464
timestamp 1
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_465
timestamp 1
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_466
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_467
timestamp 1
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_468
timestamp 1
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_469
timestamp 1
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_470
timestamp 1
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_471
timestamp 1
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_472
timestamp 1
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_473
timestamp 1
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_474
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_475
timestamp 1
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_476
timestamp 1
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_477
timestamp 1
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_478
timestamp 1
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_479
timestamp 1
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_480
timestamp 1
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_481
timestamp 1
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_482
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_483
timestamp 1
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_484
timestamp 1
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_485
timestamp 1
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_486
timestamp 1
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_487
timestamp 1
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_488
timestamp 1
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_489
timestamp 1
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_490
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_491
timestamp 1
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_492
timestamp 1
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_493
timestamp 1
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_494
timestamp 1
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_495
timestamp 1
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_496
timestamp 1
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_497
timestamp 1
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_498
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_499
timestamp 1
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_500
timestamp 1
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_501
timestamp 1
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_502
timestamp 1
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_503
timestamp 1
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_504
timestamp 1
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_505
timestamp 1
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_506
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_507
timestamp 1
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_508
timestamp 1
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_509
timestamp 1
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_510
timestamp 1
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_511
timestamp 1
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_512
timestamp 1
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_513
timestamp 1
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_514
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_515
timestamp 1
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_516
timestamp 1
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_517
timestamp 1
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_518
timestamp 1
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_519
timestamp 1
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_520
timestamp 1
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_521
timestamp 1
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_522
timestamp 1
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_523
timestamp 1
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_524
timestamp 1
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_525
timestamp 1
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_526
timestamp 1
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_527
timestamp 1
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_528
timestamp 1
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_529
timestamp 1
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_530
timestamp 1
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_531
timestamp 1
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_532
timestamp 1
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_533
timestamp 1
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_534
timestamp 1
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_535
timestamp 1
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_536
timestamp 1
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_537
timestamp 1
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_538
timestamp 1
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_539
timestamp 1
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_540
timestamp 1
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_541
timestamp 1
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_542
timestamp 1
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_543
timestamp 1
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_544
timestamp 1
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_545
timestamp 1
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_546
timestamp 1
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_547
timestamp 1
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_548
timestamp 1
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_549
timestamp 1
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_550
timestamp 1
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_551
timestamp 1
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_552
timestamp 1
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_553
timestamp 1
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_554
timestamp 1
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_555
timestamp 1
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_556
timestamp 1
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_557
timestamp 1
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_558
timestamp 1
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_559
timestamp 1
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_560
timestamp 1
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_561
timestamp 1
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_562
timestamp 1
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_563
timestamp 1
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_564
timestamp 1
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_565
timestamp 1
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_566
timestamp 1
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_567
timestamp 1
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_568
timestamp 1
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_569
timestamp 1
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_570
timestamp 1
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_571
timestamp 1
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_572
timestamp 1
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_573
timestamp 1
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_574
timestamp 1
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_575
timestamp 1
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_576
timestamp 1
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_577
timestamp 1
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_578
timestamp 1
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_579
timestamp 1
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_580
timestamp 1
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_581
timestamp 1
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_582
timestamp 1
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_583
timestamp 1
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_584
timestamp 1
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_585
timestamp 1
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_586
timestamp 1
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_587
timestamp 1
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_588
timestamp 1
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_589
timestamp 1
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_590
timestamp 1
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_591
timestamp 1
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_592
timestamp 1
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_593
timestamp 1
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_594
timestamp 1
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_595
timestamp 1
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_596
timestamp 1
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_597
timestamp 1
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_598
timestamp 1
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_599
timestamp 1
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_600
timestamp 1
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_601
timestamp 1
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_602
timestamp 1
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_603
timestamp 1
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_604
timestamp 1
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_605
timestamp 1
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_606
timestamp 1
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_607
timestamp 1
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_608
timestamp 1
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_609
timestamp 1
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_610
timestamp 1
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_611
timestamp 1
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_612
timestamp 1
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_613
timestamp 1
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_614
timestamp 1
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_615
timestamp 1
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_616
timestamp 1
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_617
timestamp 1
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_618
timestamp 1
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_619
timestamp 1
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_620
timestamp 1
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_621
timestamp 1
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_622
timestamp 1
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_623
timestamp 1
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_624
timestamp 1
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_625
timestamp 1
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_626
timestamp 1
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_627
timestamp 1
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_628
timestamp 1
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_629
timestamp 1
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_630
timestamp 1
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_631
timestamp 1
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_632
timestamp 1
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_633
timestamp 1
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_634
timestamp 1
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_635
timestamp 1
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_636
timestamp 1
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_637
timestamp 1
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_638
timestamp 1
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_639
timestamp 1
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_640
timestamp 1
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_641
timestamp 1
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_642
timestamp 1
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_643
timestamp 1
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_644
timestamp 1
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_645
timestamp 1
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_646
timestamp 1
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_647
timestamp 1
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_648
timestamp 1
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_649
timestamp 1
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_650
timestamp 1
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_651
timestamp 1
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_652
timestamp 1
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_653
timestamp 1
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_654
timestamp 1
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_655
timestamp 1
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_656
timestamp 1
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_657
timestamp 1
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_658
timestamp 1
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_659
timestamp 1
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_660
timestamp 1
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_661
timestamp 1
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_662
timestamp 1
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_663
timestamp 1
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_664
timestamp 1
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_665
timestamp 1
transform 1 0 42320 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire71
timestamp 1
transform 1 0 2392 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire72
timestamp 1
transform 1 0 3128 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire73
timestamp 1
transform -1 0 10672 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire74
timestamp 1
transform -1 0 7728 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire75
timestamp 1
transform -1 0 5244 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire76
timestamp 1
transform -1 0 3496 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire105
timestamp 1
transform -1 0 5428 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire106
timestamp 1
transform -1 0 12604 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire107
timestamp 1
transform -1 0 9200 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire108
timestamp 1
transform -1 0 7820 0 1 15232
box -38 -48 314 592
<< labels >>
flabel metal4 s 4868 2128 5188 37584 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 37584 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 addr0[0]
port 2 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 addr0[1]
port 3 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 addr0[2]
port 4 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 addr0[3]
port 5 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 addr0[4]
port 6 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 addr0[5]
port 7 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 addr0[6]
port 8 nsew signal input
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 addr0[7]
port 9 nsew signal input
flabel metal3 s 45200 29928 46000 30048 0 FreeSans 480 0 0 0 clk0
port 10 nsew signal input
flabel metal3 s 45200 29248 46000 29368 0 FreeSans 480 0 0 0 cs0
port 11 nsew signal input
flabel metal3 s 45200 15648 46000 15768 0 FreeSans 480 0 0 0 dout0[0]
port 12 nsew signal output
flabel metal2 s 25778 39200 25834 40000 0 FreeSans 224 90 0 0 dout0[10]
port 13 nsew signal output
flabel metal3 s 45200 27208 46000 27328 0 FreeSans 480 0 0 0 dout0[11]
port 14 nsew signal output
flabel metal3 s 45200 26528 46000 26648 0 FreeSans 480 0 0 0 dout0[12]
port 15 nsew signal output
flabel metal3 s 45200 20408 46000 20528 0 FreeSans 480 0 0 0 dout0[13]
port 16 nsew signal output
flabel metal3 s 45200 28568 46000 28688 0 FreeSans 480 0 0 0 dout0[14]
port 17 nsew signal output
flabel metal2 s 27710 39200 27766 40000 0 FreeSans 224 90 0 0 dout0[15]
port 18 nsew signal output
flabel metal3 s 45200 25848 46000 25968 0 FreeSans 480 0 0 0 dout0[16]
port 19 nsew signal output
flabel metal3 s 45200 13608 46000 13728 0 FreeSans 480 0 0 0 dout0[17]
port 20 nsew signal output
flabel metal3 s 45200 23128 46000 23248 0 FreeSans 480 0 0 0 dout0[18]
port 21 nsew signal output
flabel metal2 s 23202 39200 23258 40000 0 FreeSans 224 90 0 0 dout0[19]
port 22 nsew signal output
flabel metal3 s 45200 17688 46000 17808 0 FreeSans 480 0 0 0 dout0[1]
port 23 nsew signal output
flabel metal3 s 45200 24488 46000 24608 0 FreeSans 480 0 0 0 dout0[20]
port 24 nsew signal output
flabel metal3 s 45200 14968 46000 15088 0 FreeSans 480 0 0 0 dout0[21]
port 25 nsew signal output
flabel metal3 s 45200 27888 46000 28008 0 FreeSans 480 0 0 0 dout0[22]
port 26 nsew signal output
flabel metal3 s 45200 14288 46000 14408 0 FreeSans 480 0 0 0 dout0[23]
port 27 nsew signal output
flabel metal3 s 45200 23808 46000 23928 0 FreeSans 480 0 0 0 dout0[24]
port 28 nsew signal output
flabel metal3 s 45200 22448 46000 22568 0 FreeSans 480 0 0 0 dout0[25]
port 29 nsew signal output
flabel metal2 s 31574 39200 31630 40000 0 FreeSans 224 90 0 0 dout0[26]
port 30 nsew signal output
flabel metal3 s 45200 17008 46000 17128 0 FreeSans 480 0 0 0 dout0[27]
port 31 nsew signal output
flabel metal3 s 45200 16328 46000 16448 0 FreeSans 480 0 0 0 dout0[28]
port 32 nsew signal output
flabel metal3 s 45200 18368 46000 18488 0 FreeSans 480 0 0 0 dout0[29]
port 33 nsew signal output
flabel metal2 s 28998 39200 29054 40000 0 FreeSans 224 90 0 0 dout0[2]
port 34 nsew signal output
flabel metal3 s 45200 19048 46000 19168 0 FreeSans 480 0 0 0 dout0[30]
port 35 nsew signal output
flabel metal3 s 45200 21088 46000 21208 0 FreeSans 480 0 0 0 dout0[31]
port 36 nsew signal output
flabel metal2 s 21914 39200 21970 40000 0 FreeSans 224 90 0 0 dout0[3]
port 37 nsew signal output
flabel metal2 s 25134 39200 25190 40000 0 FreeSans 224 90 0 0 dout0[4]
port 38 nsew signal output
flabel metal3 s 45200 21768 46000 21888 0 FreeSans 480 0 0 0 dout0[5]
port 39 nsew signal output
flabel metal3 s 45200 25168 46000 25288 0 FreeSans 480 0 0 0 dout0[6]
port 40 nsew signal output
flabel metal3 s 45200 19728 46000 19848 0 FreeSans 480 0 0 0 dout0[7]
port 41 nsew signal output
flabel metal2 s 29642 39200 29698 40000 0 FreeSans 224 90 0 0 dout0[8]
port 42 nsew signal output
flabel metal2 s 22558 39200 22614 40000 0 FreeSans 224 90 0 0 dout0[9]
port 43 nsew signal output
rlabel metal1 23000 36992 23000 36992 0 VGND
rlabel metal1 23000 37536 23000 37536 0 VPWR
rlabel metal1 37658 15062 37658 15062 0 _0000_
rlabel metal2 41630 18530 41630 18530 0 _0001_
rlabel metal1 27784 33082 27784 33082 0 _0002_
rlabel metal2 23322 34306 23322 34306 0 _0003_
rlabel metal1 24380 34170 24380 34170 0 _0004_
rlabel metal2 43378 21488 43378 21488 0 _0005_
rlabel metal1 42356 26350 42356 26350 0 _0006_
rlabel metal2 41630 20706 41630 20706 0 _0007_
rlabel metal2 29578 33286 29578 33286 0 _0008_
rlabel metal1 21781 33830 21781 33830 0 _0009_
rlabel metal2 26174 33762 26174 33762 0 _0010_
rlabel metal2 39606 27234 39606 27234 0 _0011_
rlabel metal1 40654 26350 40654 26350 0 _0012_
rlabel metal1 40526 25466 40526 25466 0 _0013_
rlabel metal1 38640 28730 38640 28730 0 _0014_
rlabel metal2 27738 34102 27738 34102 0 _0015_
rlabel metal1 42494 24786 42494 24786 0 _0016_
rlabel metal1 41614 15402 41614 15402 0 _0017_
rlabel metal1 40372 21590 40372 21590 0 _0018_
rlabel metal2 23690 34374 23690 34374 0 _0019_
rlabel metal2 43194 24514 43194 24514 0 _0020_
rlabel metal1 37290 15402 37290 15402 0 _0021_
rlabel metal2 42090 28050 42090 28050 0 _0022_
rlabel viali 35921 15470 35921 15470 0 _0023_
rlabel metal2 41078 23664 41078 23664 0 _0024_
rlabel metal1 40516 22610 40516 22610 0 _0025_
rlabel metal2 31050 32674 31050 32674 0 _0026_
rlabel via1 42729 17170 42729 17170 0 _0027_
rlabel metal1 39504 17170 39504 17170 0 _0028_
rlabel via1 40153 17646 40153 17646 0 _0029_
rlabel metal1 42366 17782 42366 17782 0 _0030_
rlabel metal1 38594 18938 38594 18938 0 _0031_
rlabel metal1 15226 21046 15226 21046 0 _0032_
rlabel metal1 8832 21114 8832 21114 0 _0033_
rlabel metal2 2898 15572 2898 15572 0 _0034_
rlabel metal1 3082 12954 3082 12954 0 _0035_
rlabel metal1 20976 20978 20976 20978 0 _0036_
rlabel metal1 21735 20230 21735 20230 0 _0037_
rlabel metal1 8878 16218 8878 16218 0 _0038_
rlabel metal2 8786 19346 8786 19346 0 _0039_
rlabel metal1 10534 29138 10534 29138 0 _0040_
rlabel metal1 2024 13906 2024 13906 0 _0041_
rlabel metal2 13294 13073 13294 13073 0 _0042_
rlabel metal1 18308 24718 18308 24718 0 _0043_
rlabel metal1 10810 29818 10810 29818 0 _0044_
rlabel metal1 24288 14382 24288 14382 0 _0045_
rlabel metal2 14766 12347 14766 12347 0 _0046_
rlabel metal1 3588 18258 3588 18258 0 _0047_
rlabel metal2 3266 17748 3266 17748 0 _0048_
rlabel metal2 18906 15827 18906 15827 0 _0049_
rlabel metal1 6900 21930 6900 21930 0 _0050_
rlabel metal1 16330 24140 16330 24140 0 _0051_
rlabel metal1 7222 23528 7222 23528 0 _0052_
rlabel metal1 7130 20808 7130 20808 0 _0053_
rlabel metal2 7038 21539 7038 21539 0 _0054_
rlabel metal1 13202 27438 13202 27438 0 _0055_
rlabel metal1 16514 19210 16514 19210 0 _0056_
rlabel metal1 13340 30158 13340 30158 0 _0057_
rlabel metal1 18676 20026 18676 20026 0 _0058_
rlabel metal2 18262 19737 18262 19737 0 _0059_
rlabel metal1 20378 20774 20378 20774 0 _0060_
rlabel metal1 4968 17170 4968 17170 0 _0061_
rlabel metal1 3358 15062 3358 15062 0 _0062_
rlabel metal1 17848 22678 17848 22678 0 _0063_
rlabel metal2 6026 23630 6026 23630 0 _0064_
rlabel metal2 16330 23392 16330 23392 0 _0065_
rlabel metal1 8418 14042 8418 14042 0 _0066_
rlabel metal2 6118 13498 6118 13498 0 _0067_
rlabel metal2 15134 17527 15134 17527 0 _0068_
rlabel metal2 18354 21233 18354 21233 0 _0069_
rlabel metal2 7038 13430 7038 13430 0 _0070_
rlabel metal2 7130 14790 7130 14790 0 _0071_
rlabel via2 16238 15963 16238 15963 0 _0072_
rlabel metal1 16560 12308 16560 12308 0 _0073_
rlabel via2 17710 12699 17710 12699 0 _0074_
rlabel metal1 33672 17578 33672 17578 0 _0075_
rlabel via2 17342 16099 17342 16099 0 _0076_
rlabel metal1 32890 19822 32890 19822 0 _0077_
rlabel metal2 16514 25024 16514 25024 0 _0078_
rlabel metal2 35374 16643 35374 16643 0 _0079_
rlabel metal2 9798 28475 9798 28475 0 _0080_
rlabel metal3 22333 12172 22333 12172 0 _0081_
rlabel metal1 33534 14824 33534 14824 0 _0082_
rlabel metal2 15870 32283 15870 32283 0 _0083_
rlabel metal1 24334 14824 24334 14824 0 _0084_
rlabel metal1 16928 17646 16928 17646 0 _0085_
rlabel metal1 20378 13974 20378 13974 0 _0086_
rlabel metal2 26266 17544 26266 17544 0 _0087_
rlabel metal1 7682 19482 7682 19482 0 _0088_
rlabel metal1 16514 17850 16514 17850 0 _0089_
rlabel metal3 17388 16524 17388 16524 0 _0090_
rlabel metal3 19297 21692 19297 21692 0 _0091_
rlabel metal3 24932 20672 24932 20672 0 _0092_
rlabel metal1 18262 20876 18262 20876 0 _0093_
rlabel via2 11086 15147 11086 15147 0 _0094_
rlabel metal1 14260 17034 14260 17034 0 _0095_
rlabel metal1 27968 16966 27968 16966 0 _0096_
rlabel metal1 11914 11662 11914 11662 0 _0097_
rlabel via2 33718 15011 33718 15011 0 _0098_
rlabel metal1 17664 12342 17664 12342 0 _0099_
rlabel metal2 36110 15011 36110 15011 0 _0100_
rlabel metal1 23966 14926 23966 14926 0 _0101_
rlabel metal2 17250 12971 17250 12971 0 _0102_
rlabel metal2 16100 21318 16100 21318 0 _0103_
rlabel metal1 20056 14586 20056 14586 0 _0104_
rlabel metal1 18768 12614 18768 12614 0 _0105_
rlabel metal1 22908 14382 22908 14382 0 _0106_
rlabel metal1 20286 31280 20286 31280 0 _0107_
rlabel metal2 36938 18479 36938 18479 0 _0108_
rlabel metal1 14306 12614 14306 12614 0 _0109_
rlabel metal1 17204 16490 17204 16490 0 _0110_
rlabel metal1 8464 15470 8464 15470 0 _0111_
rlabel via2 8786 16099 8786 16099 0 _0112_
rlabel metal2 17434 16745 17434 16745 0 _0113_
rlabel metal2 29578 18530 29578 18530 0 _0114_
rlabel metal3 18193 10948 18193 10948 0 _0115_
rlabel metal1 34546 27438 34546 27438 0 _0116_
rlabel via2 18906 19363 18906 19363 0 _0117_
rlabel metal2 18814 15657 18814 15657 0 _0118_
rlabel metal2 23506 26044 23506 26044 0 _0119_
rlabel metal1 18676 16014 18676 16014 0 _0120_
rlabel metal1 22172 29138 22172 29138 0 _0121_
rlabel metal1 14306 24786 14306 24786 0 _0122_
rlabel metal2 10166 24140 10166 24140 0 _0123_
rlabel metal2 17250 26690 17250 26690 0 _0124_
rlabel metal1 11638 20230 11638 20230 0 _0125_
rlabel metal1 18584 26350 18584 26350 0 _0126_
rlabel metal1 17664 18054 17664 18054 0 _0127_
rlabel metal2 9246 25500 9246 25500 0 _0128_
rlabel metal2 13570 17187 13570 17187 0 _0129_
rlabel metal1 12926 30702 12926 30702 0 _0130_
rlabel metal1 31372 19346 31372 19346 0 _0131_
rlabel metal1 23230 24310 23230 24310 0 _0132_
rlabel metal1 15180 29138 15180 29138 0 _0133_
rlabel metal1 18492 20230 18492 20230 0 _0134_
rlabel metal1 17296 19346 17296 19346 0 _0135_
rlabel metal1 12742 21318 12742 21318 0 _0136_
rlabel metal1 18538 21998 18538 21998 0 _0137_
rlabel metal2 20010 19822 20010 19822 0 _0138_
rlabel metal1 14674 20026 14674 20026 0 _0139_
rlabel metal1 17296 21114 17296 21114 0 _0140_
rlabel metal1 17710 31790 17710 31790 0 _0141_
rlabel metal1 11500 21114 11500 21114 0 _0142_
rlabel metal1 19274 18768 19274 18768 0 _0143_
rlabel metal1 22494 18292 22494 18292 0 _0144_
rlabel metal1 24196 14586 24196 14586 0 _0145_
rlabel metal2 23874 15402 23874 15402 0 _0146_
rlabel metal1 22678 15674 22678 15674 0 _0147_
rlabel metal1 23552 15470 23552 15470 0 _0148_
rlabel metal1 26910 20434 26910 20434 0 _0149_
rlabel metal1 26404 17646 26404 17646 0 _0150_
rlabel metal1 25990 17646 25990 17646 0 _0151_
rlabel metal1 27600 17170 27600 17170 0 _0152_
rlabel metal2 27738 17646 27738 17646 0 _0153_
rlabel metal2 29394 16830 29394 16830 0 _0154_
rlabel metal2 37490 15623 37490 15623 0 _0155_
rlabel metal1 14260 32470 14260 32470 0 _0156_
rlabel metal1 17480 18190 17480 18190 0 _0157_
rlabel metal1 25300 16218 25300 16218 0 _0158_
rlabel metal1 35098 15912 35098 15912 0 _0159_
rlabel metal1 15272 21930 15272 21930 0 _0160_
rlabel via2 20562 23035 20562 23035 0 _0161_
rlabel metal1 17112 21862 17112 21862 0 _0162_
rlabel metal1 27830 20400 27830 20400 0 _0163_
rlabel metal1 13340 30226 13340 30226 0 _0164_
rlabel metal1 15134 24344 15134 24344 0 _0165_
rlabel via2 17618 20893 17618 20893 0 _0166_
rlabel metal3 17135 12308 17135 12308 0 _0167_
rlabel metal1 38318 28730 38318 28730 0 _0168_
rlabel metal1 29348 19822 29348 19822 0 _0169_
rlabel via1 2814 19346 2814 19346 0 _0170_
rlabel metal1 18400 22066 18400 22066 0 _0171_
rlabel metal2 19274 19006 19274 19006 0 _0172_
rlabel metal2 36478 17289 36478 17289 0 _0173_
rlabel metal1 24012 12410 24012 12410 0 _0174_
rlabel metal1 22586 30736 22586 30736 0 _0175_
rlabel metal1 31786 29784 31786 29784 0 _0176_
rlabel metal1 31786 17136 31786 17136 0 _0177_
rlabel metal2 17434 13600 17434 13600 0 _0178_
rlabel metal1 13892 13158 13892 13158 0 _0179_
rlabel metal1 26910 16626 26910 16626 0 _0180_
rlabel metal1 36386 16490 36386 16490 0 _0181_
rlabel metal2 27094 15062 27094 15062 0 _0182_
rlabel metal1 36064 17238 36064 17238 0 _0183_
rlabel metal1 37536 18190 37536 18190 0 _0184_
rlabel metal2 8694 23494 8694 23494 0 _0185_
rlabel metal1 9430 31790 9430 31790 0 _0186_
rlabel metal1 7636 24786 7636 24786 0 _0187_
rlabel metal1 16974 18054 16974 18054 0 _0188_
rlabel metal1 6578 27302 6578 27302 0 _0189_
rlabel metal2 38870 25007 38870 25007 0 _0190_
rlabel metal1 34362 19822 34362 19822 0 _0191_
rlabel metal1 13386 22066 13386 22066 0 _0192_
rlabel metal1 33948 20026 33948 20026 0 _0193_
rlabel metal2 14306 29257 14306 29257 0 _0194_
rlabel metal1 37996 19890 37996 19890 0 _0195_
rlabel metal1 7912 28118 7912 28118 0 _0196_
rlabel metal2 17066 18751 17066 18751 0 _0197_
rlabel metal2 38318 23052 38318 23052 0 _0198_
rlabel metal1 24426 25874 24426 25874 0 _0199_
rlabel metal2 23230 27744 23230 27744 0 _0200_
rlabel metal1 36386 26962 36386 26962 0 _0201_
rlabel via2 13754 17765 13754 17765 0 _0202_
rlabel metal1 17342 20910 17342 20910 0 _0203_
rlabel metal2 20010 31841 20010 31841 0 _0204_
rlabel metal1 13570 21114 13570 21114 0 _0205_
rlabel metal1 37122 19890 37122 19890 0 _0206_
rlabel metal2 37490 19312 37490 19312 0 _0207_
rlabel metal1 35236 31314 35236 31314 0 _0208_
rlabel metal1 24288 30702 24288 30702 0 _0209_
rlabel metal1 17158 16082 17158 16082 0 _0210_
rlabel metal2 25254 15130 25254 15130 0 _0211_
rlabel metal1 17572 16490 17572 16490 0 _0212_
rlabel metal2 17894 17102 17894 17102 0 _0213_
rlabel metal2 13018 16286 13018 16286 0 _0214_
rlabel metal2 22310 17731 22310 17731 0 _0215_
rlabel metal2 22402 17850 22402 17850 0 _0216_
rlabel metal1 19872 17170 19872 17170 0 _0217_
rlabel metal2 11822 29308 11822 29308 0 _0218_
rlabel metal2 10810 26146 10810 26146 0 _0219_
rlabel metal1 20930 26792 20930 26792 0 _0220_
rlabel metal2 19366 17017 19366 17017 0 _0221_
rlabel metal1 19228 17170 19228 17170 0 _0222_
rlabel metal1 14858 31144 14858 31144 0 _0223_
rlabel metal1 11316 29002 11316 29002 0 _0224_
rlabel metal1 22816 20434 22816 20434 0 _0225_
rlabel metal1 31464 18258 31464 18258 0 _0226_
rlabel metal1 24518 25976 24518 25976 0 _0227_
rlabel metal2 7222 28390 7222 28390 0 _0228_
rlabel metal1 17112 29138 17112 29138 0 _0229_
rlabel metal1 17480 27506 17480 27506 0 _0230_
rlabel metal1 11500 29138 11500 29138 0 _0231_
rlabel metal1 16928 18734 16928 18734 0 _0232_
rlabel metal2 21574 21182 21574 21182 0 _0233_
rlabel metal1 24610 21488 24610 21488 0 _0234_
rlabel metal1 21620 20774 21620 20774 0 _0235_
rlabel metal2 10534 19431 10534 19431 0 _0236_
rlabel metal2 32338 20417 32338 20417 0 _0237_
rlabel metal1 35052 21658 35052 21658 0 _0238_
rlabel metal1 21068 19346 21068 19346 0 _0239_
rlabel metal1 14674 21930 14674 21930 0 _0240_
rlabel metal2 37122 20179 37122 20179 0 _0241_
rlabel metal2 27554 27166 27554 27166 0 _0242_
rlabel metal1 26358 18938 26358 18938 0 _0243_
rlabel metal1 19734 18190 19734 18190 0 _0244_
rlabel via1 32890 31331 32890 31331 0 _0245_
rlabel metal1 27876 32334 27876 32334 0 _0246_
rlabel metal2 35006 18360 35006 18360 0 _0247_
rlabel metal2 18630 18649 18630 18649 0 _0248_
rlabel metal2 18814 19703 18814 19703 0 _0249_
rlabel metal1 15686 19278 15686 19278 0 _0250_
rlabel metal2 34454 23885 34454 23885 0 _0251_
rlabel metal2 16790 30107 16790 30107 0 _0252_
rlabel metal2 21666 28016 21666 28016 0 _0253_
rlabel metal1 19918 19380 19918 19380 0 _0254_
rlabel metal2 22402 18428 22402 18428 0 _0255_
rlabel metal4 15732 23936 15732 23936 0 _0256_
rlabel metal1 37536 18054 37536 18054 0 _0257_
rlabel metal1 13054 22406 13054 22406 0 _0258_
rlabel metal1 12788 22610 12788 22610 0 _0259_
rlabel metal1 30958 23596 30958 23596 0 _0260_
rlabel metal1 29670 23630 29670 23630 0 _0261_
rlabel metal2 21114 19788 21114 19788 0 _0262_
rlabel metal1 22586 18088 22586 18088 0 _0263_
rlabel metal1 15456 15674 15456 15674 0 _0264_
rlabel metal2 15226 18547 15226 18547 0 _0265_
rlabel metal1 21620 23698 21620 23698 0 _0266_
rlabel metal2 35558 24514 35558 24514 0 _0267_
rlabel metal1 24058 23494 24058 23494 0 _0268_
rlabel metal1 34822 18054 34822 18054 0 _0269_
rlabel via2 9982 17867 9982 17867 0 _0270_
rlabel metal1 15502 24106 15502 24106 0 _0271_
rlabel metal1 29348 29070 29348 29070 0 _0272_
rlabel metal2 28842 15912 28842 15912 0 _0273_
rlabel via3 32821 27676 32821 27676 0 _0274_
rlabel metal1 17066 18224 17066 18224 0 _0275_
rlabel metal1 22126 13260 22126 13260 0 _0276_
rlabel metal2 13110 13719 13110 13719 0 _0277_
rlabel metal1 33902 15402 33902 15402 0 _0278_
rlabel metal2 34822 15844 34822 15844 0 _0279_
rlabel via1 12102 14042 12102 14042 0 _0280_
rlabel metal1 26772 26350 26772 26350 0 _0281_
rlabel metal2 20378 13991 20378 13991 0 _0282_
rlabel metal1 35374 23630 35374 23630 0 _0283_
rlabel metal2 16606 15487 16606 15487 0 _0284_
rlabel metal1 19512 13906 19512 13906 0 _0285_
rlabel metal2 22218 15198 22218 15198 0 _0286_
rlabel via2 20562 14365 20562 14365 0 _0287_
rlabel metal1 24978 17034 24978 17034 0 _0288_
rlabel metal2 22034 14297 22034 14297 0 _0289_
rlabel metal1 16606 14518 16606 14518 0 _0290_
rlabel metal1 27094 23222 27094 23222 0 _0291_
rlabel metal1 14536 13158 14536 13158 0 _0292_
rlabel metal2 26726 27370 26726 27370 0 _0293_
rlabel metal2 33810 15266 33810 15266 0 _0294_
rlabel metal2 14674 26690 14674 26690 0 _0295_
rlabel metal1 37996 29002 37996 29002 0 _0296_
rlabel metal2 21942 29988 21942 29988 0 _0297_
rlabel metal4 17940 22168 17940 22168 0 _0298_
rlabel metal1 34316 29138 34316 29138 0 _0299_
rlabel metal2 35374 27948 35374 27948 0 _0300_
rlabel metal1 28106 15436 28106 15436 0 _0301_
rlabel metal1 34362 15402 34362 15402 0 _0302_
rlabel metal1 35880 15674 35880 15674 0 _0303_
rlabel metal2 38226 17884 38226 17884 0 _0304_
rlabel metal2 39054 17119 39054 17119 0 _0305_
rlabel metal1 32936 23086 32936 23086 0 _0306_
rlabel metal1 31234 24276 31234 24276 0 _0307_
rlabel metal1 25576 19822 25576 19822 0 _0308_
rlabel via1 20194 28934 20194 28934 0 _0309_
rlabel metal1 22586 13906 22586 13906 0 _0310_
rlabel metal1 23092 14042 23092 14042 0 _0311_
rlabel metal1 19274 31824 19274 31824 0 _0312_
rlabel metal1 30820 23698 30820 23698 0 _0313_
rlabel metal1 31648 28730 31648 28730 0 _0314_
rlabel metal2 31602 26248 31602 26248 0 _0315_
rlabel metal1 31602 23596 31602 23596 0 _0316_
rlabel metal2 15502 24038 15502 24038 0 _0317_
rlabel metal1 14674 22746 14674 22746 0 _0318_
rlabel metal2 15226 23392 15226 23392 0 _0319_
rlabel metal1 10534 24072 10534 24072 0 _0320_
rlabel metal2 10994 23834 10994 23834 0 _0321_
rlabel metal1 15548 20026 15548 20026 0 _0322_
rlabel via2 15686 23851 15686 23851 0 _0323_
rlabel metal2 31970 23069 31970 23069 0 _0324_
rlabel metal1 24794 28050 24794 28050 0 _0325_
rlabel metal1 26220 20230 26220 20230 0 _0326_
rlabel metal1 23920 30090 23920 30090 0 _0327_
rlabel metal2 13294 27744 13294 27744 0 _0328_
rlabel via1 26174 13974 26174 13974 0 _0329_
rlabel metal1 26818 14994 26818 14994 0 _0330_
rlabel via2 27370 15147 27370 15147 0 _0331_
rlabel metal1 13340 15878 13340 15878 0 _0332_
rlabel metal1 21436 30566 21436 30566 0 _0333_
rlabel metal2 23322 28288 23322 28288 0 _0334_
rlabel metal2 21114 22022 21114 22022 0 _0335_
rlabel metal2 28934 30906 28934 30906 0 _0336_
rlabel metal1 26358 30736 26358 30736 0 _0337_
rlabel metal2 24426 27166 24426 27166 0 _0338_
rlabel metal1 10718 27574 10718 27574 0 _0339_
rlabel via2 13662 27829 13662 27829 0 _0340_
rlabel metal2 27462 27506 27462 27506 0 _0341_
rlabel metal1 25024 26010 25024 26010 0 _0342_
rlabel metal1 27002 27608 27002 27608 0 _0343_
rlabel metal1 24702 22066 24702 22066 0 _0344_
rlabel metal1 27002 27472 27002 27472 0 _0345_
rlabel metal1 27830 32810 27830 32810 0 _0346_
rlabel metal1 10672 31110 10672 31110 0 _0347_
rlabel metal1 16376 28390 16376 28390 0 _0348_
rlabel metal2 34592 18156 34592 18156 0 _0349_
rlabel metal2 29210 22950 29210 22950 0 _0350_
rlabel metal2 29762 32062 29762 32062 0 _0351_
rlabel metal1 13478 32368 13478 32368 0 _0352_
rlabel metal1 19228 32402 19228 32402 0 _0353_
rlabel metal2 23046 32232 23046 32232 0 _0354_
rlabel metal1 14858 28084 14858 28084 0 _0355_
rlabel metal1 12788 26010 12788 26010 0 _0356_
rlabel metal2 14490 28900 14490 28900 0 _0357_
rlabel metal1 37490 25738 37490 25738 0 _0358_
rlabel metal2 23598 32946 23598 32946 0 _0359_
rlabel metal2 22218 27268 22218 27268 0 _0360_
rlabel metal2 21942 27778 21942 27778 0 _0361_
rlabel metal2 19734 27710 19734 27710 0 _0362_
rlabel metal2 21988 19244 21988 19244 0 _0363_
rlabel metal1 22678 27574 22678 27574 0 _0364_
rlabel metal1 23736 21318 23736 21318 0 _0365_
rlabel metal2 18814 26843 18814 26843 0 _0366_
rlabel metal2 22586 30634 22586 30634 0 _0367_
rlabel metal1 22448 20978 22448 20978 0 _0368_
rlabel metal2 16514 26180 16514 26180 0 _0369_
rlabel metal1 19504 20910 19504 20910 0 _0370_
rlabel metal1 31556 22406 31556 22406 0 _0371_
rlabel metal2 20976 27030 20976 27030 0 _0372_
rlabel metal1 24334 22406 24334 22406 0 _0373_
rlabel metal1 29670 13498 29670 13498 0 _0374_
rlabel metal1 24840 21114 24840 21114 0 _0375_
rlabel metal1 18998 26282 18998 26282 0 _0376_
rlabel metal2 17618 25636 17618 25636 0 _0377_
rlabel metal2 16514 24480 16514 24480 0 _0378_
rlabel metal1 17158 16218 17158 16218 0 _0379_
rlabel metal2 17250 24582 17250 24582 0 _0380_
rlabel metal2 17802 29138 17802 29138 0 _0381_
rlabel metal1 27600 19958 27600 19958 0 _0382_
rlabel metal1 24472 20910 24472 20910 0 _0383_
rlabel metal3 24955 33252 24955 33252 0 _0384_
rlabel metal2 25346 26996 25346 26996 0 _0385_
rlabel metal1 35144 20298 35144 20298 0 _0386_
rlabel metal2 38042 29750 38042 29750 0 _0387_
rlabel metal1 38226 20366 38226 20366 0 _0388_
rlabel metal2 13754 28441 13754 28441 0 _0389_
rlabel via2 18262 24667 18262 24667 0 _0390_
rlabel metal1 39330 23154 39330 23154 0 _0391_
rlabel metal1 32430 19822 32430 19822 0 _0392_
rlabel metal1 38456 21318 38456 21318 0 _0393_
rlabel metal2 37306 21835 37306 21835 0 _0394_
rlabel metal1 39008 20570 39008 20570 0 _0395_
rlabel metal1 12972 29274 12972 29274 0 _0396_
rlabel metal1 13386 32300 13386 32300 0 _0397_
rlabel metal2 10994 29172 10994 29172 0 _0398_
rlabel metal2 11454 32198 11454 32198 0 _0399_
rlabel metal2 13662 32249 13662 32249 0 _0400_
rlabel metal1 38318 28390 38318 28390 0 _0401_
rlabel metal1 38732 21114 38732 21114 0 _0402_
rlabel metal1 43654 21012 43654 21012 0 _0403_
rlabel metal1 31142 26384 31142 26384 0 _0404_
rlabel via2 33994 19771 33994 19771 0 _0405_
rlabel metal1 34776 26962 34776 26962 0 _0406_
rlabel metal2 33166 27200 33166 27200 0 _0407_
rlabel metal2 35190 27302 35190 27302 0 _0408_
rlabel metal2 28290 24480 28290 24480 0 _0409_
rlabel metal2 35006 26826 35006 26826 0 _0410_
rlabel metal1 20792 25262 20792 25262 0 _0411_
rlabel metal2 19182 28764 19182 28764 0 _0412_
rlabel metal1 19090 28118 19090 28118 0 _0413_
rlabel metal2 5658 25126 5658 25126 0 _0414_
rlabel metal1 20424 23154 20424 23154 0 _0415_
rlabel metal1 21229 25194 21229 25194 0 _0416_
rlabel metal2 20746 26826 20746 26826 0 _0417_
rlabel metal1 9016 22746 9016 22746 0 _0418_
rlabel metal1 8970 25976 8970 25976 0 _0419_
rlabel metal2 12558 26078 12558 26078 0 _0420_
rlabel metal1 20746 25466 20746 25466 0 _0421_
rlabel metal2 20470 26554 20470 26554 0 _0422_
rlabel metal2 20930 26639 20930 26639 0 _0423_
rlabel metal1 35696 30294 35696 30294 0 _0424_
rlabel metal1 35926 29172 35926 29172 0 _0425_
rlabel metal1 33488 31178 33488 31178 0 _0426_
rlabel metal1 39836 23290 39836 23290 0 _0427_
rlabel metal1 31878 26418 31878 26418 0 _0428_
rlabel metal1 18630 29138 18630 29138 0 _0429_
rlabel metal1 19642 31382 19642 31382 0 _0430_
rlabel metal2 33810 31110 33810 31110 0 _0431_
rlabel metal1 20746 29546 20746 29546 0 _0432_
rlabel metal1 35650 29070 35650 29070 0 _0433_
rlabel metal1 35558 29138 35558 29138 0 _0434_
rlabel metal1 35604 25262 35604 25262 0 _0435_
rlabel metal1 34500 25466 34500 25466 0 _0436_
rlabel metal2 23782 25568 23782 25568 0 _0437_
rlabel metal1 23736 24922 23736 24922 0 _0438_
rlabel metal2 12926 28220 12926 28220 0 _0439_
rlabel via2 13294 25653 13294 25653 0 _0440_
rlabel metal2 31970 25279 31970 25279 0 _0441_
rlabel metal1 41952 20434 41952 20434 0 _0442_
rlabel metal1 25981 29512 25981 29512 0 _0443_
rlabel metal1 23782 19754 23782 19754 0 _0444_
rlabel via3 32683 22236 32683 22236 0 _0445_
rlabel metal2 17250 27880 17250 27880 0 _0446_
rlabel via2 28106 14059 28106 14059 0 _0447_
rlabel metal1 29348 32538 29348 32538 0 _0448_
rlabel metal2 33994 26214 33994 26214 0 _0449_
rlabel metal1 31050 30022 31050 30022 0 _0450_
rlabel via2 17710 32011 17710 32011 0 _0451_
rlabel metal2 30406 30022 30406 30022 0 _0452_
rlabel metal1 31142 30158 31142 30158 0 _0453_
rlabel metal2 31142 14790 31142 14790 0 _0454_
rlabel via3 31533 29036 31533 29036 0 _0455_
rlabel metal1 31096 30090 31096 30090 0 _0456_
rlabel metal2 16146 28254 16146 28254 0 _0457_
rlabel metal1 30820 21454 30820 21454 0 _0458_
rlabel metal1 11040 24582 11040 24582 0 _0459_
rlabel metal1 29256 28594 29256 28594 0 _0460_
rlabel metal2 16054 27200 16054 27200 0 _0461_
rlabel metal2 7498 24004 7498 24004 0 _0462_
rlabel metal2 15870 27727 15870 27727 0 _0463_
rlabel metal1 19044 34034 19044 34034 0 _0464_
rlabel metal1 23368 28594 23368 28594 0 _0465_
rlabel metal2 5290 26758 5290 26758 0 _0466_
rlabel via2 6854 27931 6854 27931 0 _0467_
rlabel metal1 21965 34034 21965 34034 0 _0468_
rlabel metal1 25346 31790 25346 31790 0 _0469_
rlabel metal1 22954 30022 22954 30022 0 _0470_
rlabel metal1 27094 28628 27094 28628 0 _0471_
rlabel metal1 26864 28526 26864 28526 0 _0472_
rlabel metal2 27002 20927 27002 20927 0 _0473_
rlabel metal1 26312 31110 26312 31110 0 _0474_
rlabel metal2 26634 32198 26634 32198 0 _0475_
rlabel metal2 27738 28220 27738 28220 0 _0476_
rlabel metal1 27462 27846 27462 27846 0 _0477_
rlabel metal1 37582 27098 37582 27098 0 _0478_
rlabel metal1 37260 25466 37260 25466 0 _0479_
rlabel metal1 36524 27302 36524 27302 0 _0480_
rlabel metal1 26956 33354 26956 33354 0 _0481_
rlabel metal2 26082 32096 26082 32096 0 _0482_
rlabel metal1 20194 21862 20194 21862 0 _0483_
rlabel metal1 23736 31858 23736 31858 0 _0484_
rlabel metal1 27968 31790 27968 31790 0 _0485_
rlabel metal2 26542 32708 26542 32708 0 _0486_
rlabel metal2 29394 30736 29394 30736 0 _0487_
rlabel metal2 14582 29818 14582 29818 0 _0488_
rlabel metal1 19642 29784 19642 29784 0 _0489_
rlabel metal2 31786 25806 31786 25806 0 _0490_
rlabel metal2 21114 26894 21114 26894 0 _0491_
rlabel metal2 22126 28832 22126 28832 0 _0492_
rlabel via2 15134 25755 15134 25755 0 _0493_
rlabel metal2 21850 26214 21850 26214 0 _0494_
rlabel metal2 19734 25874 19734 25874 0 _0495_
rlabel via2 39882 26979 39882 26979 0 _0496_
rlabel metal2 32062 26724 32062 26724 0 _0497_
rlabel metal1 30498 24106 30498 24106 0 _0498_
rlabel metal1 31832 24310 31832 24310 0 _0499_
rlabel metal2 39974 26656 39974 26656 0 _0500_
rlabel metal1 33258 22032 33258 22032 0 _0501_
rlabel metal1 26404 25330 26404 25330 0 _0502_
rlabel metal1 31556 21522 31556 21522 0 _0503_
rlabel metal2 32062 25636 32062 25636 0 _0504_
rlabel metal2 18170 18802 18170 18802 0 _0505_
rlabel via2 20194 19499 20194 19499 0 _0506_
rlabel metal1 33442 27506 33442 27506 0 _0507_
rlabel metal2 32890 26588 32890 26588 0 _0508_
rlabel metal1 33350 25670 33350 25670 0 _0509_
rlabel metal2 40710 26724 40710 26724 0 _0510_
rlabel metal2 29578 23460 29578 23460 0 _0511_
rlabel metal2 39882 23324 39882 23324 0 _0512_
rlabel via2 14582 31331 14582 31331 0 _0513_
rlabel metal1 27922 17782 27922 17782 0 _0514_
rlabel metal2 19550 26350 19550 26350 0 _0515_
rlabel metal1 36846 25942 36846 25942 0 _0516_
rlabel metal1 39238 25772 39238 25772 0 _0517_
rlabel metal2 39146 26214 39146 26214 0 _0518_
rlabel metal2 40710 25534 40710 25534 0 _0519_
rlabel metal1 19228 26758 19228 26758 0 _0520_
rlabel metal2 15318 28764 15318 28764 0 _0521_
rlabel metal1 15180 26350 15180 26350 0 _0522_
rlabel metal2 15686 26758 15686 26758 0 _0523_
rlabel via2 19734 27115 19734 27115 0 _0524_
rlabel metal1 29256 20570 29256 20570 0 _0525_
rlabel metal1 34270 21862 34270 21862 0 _0526_
rlabel metal2 27738 29920 27738 29920 0 _0527_
rlabel metal2 33534 17408 33534 17408 0 _0528_
rlabel metal2 29118 29988 29118 29988 0 _0529_
rlabel metal1 38686 28594 38686 28594 0 _0530_
rlabel metal2 34270 19516 34270 19516 0 _0531_
rlabel metal2 34086 19550 34086 19550 0 _0532_
rlabel metal1 34638 19482 34638 19482 0 _0533_
rlabel metal1 35558 21862 35558 21862 0 _0534_
rlabel metal2 26910 28730 26910 28730 0 _0535_
rlabel metal2 7406 26452 7406 26452 0 _0536_
rlabel metal2 8970 28968 8970 28968 0 _0537_
rlabel metal2 7682 29359 7682 29359 0 _0538_
rlabel metal1 27278 29818 27278 29818 0 _0539_
rlabel metal1 26404 16218 26404 16218 0 _0540_
rlabel metal1 26726 22712 26726 22712 0 _0541_
rlabel metal2 24518 30634 24518 30634 0 _0542_
rlabel metal2 17710 30464 17710 30464 0 _0543_
rlabel metal1 26404 30906 26404 30906 0 _0544_
rlabel metal2 26082 30872 26082 30872 0 _0545_
rlabel metal1 26956 30702 26956 30702 0 _0546_
rlabel metal1 27876 30906 27876 30906 0 _0547_
rlabel via2 28106 24293 28106 24293 0 _0548_
rlabel metal1 35328 23086 35328 23086 0 _0549_
rlabel metal1 14582 26316 14582 26316 0 _0550_
rlabel metal1 34362 23290 34362 23290 0 _0551_
rlabel metal1 34684 23698 34684 23698 0 _0552_
rlabel metal1 19228 19482 19228 19482 0 _0553_
rlabel metal1 18906 20978 18906 20978 0 _0554_
rlabel metal1 18078 20808 18078 20808 0 _0555_
rlabel metal1 19274 20808 19274 20808 0 _0556_
rlabel metal2 19734 22287 19734 22287 0 _0557_
rlabel metal1 41901 24786 41901 24786 0 _0558_
rlabel metal1 33396 22950 33396 22950 0 _0559_
rlabel metal1 31142 15878 31142 15878 0 _0560_
rlabel metal2 26266 29818 26266 29818 0 _0561_
rlabel metal2 29026 16388 29026 16388 0 _0562_
rlabel metal1 27738 17544 27738 17544 0 _0563_
rlabel metal2 28474 17136 28474 17136 0 _0564_
rlabel metal1 20815 29002 20815 29002 0 _0565_
rlabel metal1 25254 29206 25254 29206 0 _0566_
rlabel metal3 26841 29036 26841 29036 0 _0567_
rlabel metal2 19090 15742 19090 15742 0 _0568_
rlabel metal1 27876 15130 27876 15130 0 _0569_
rlabel metal2 28290 16082 28290 16082 0 _0570_
rlabel metal1 41170 15436 41170 15436 0 _0571_
rlabel metal2 18170 21726 18170 21726 0 _0572_
rlabel metal2 27002 19788 27002 19788 0 _0573_
rlabel metal1 20286 16626 20286 16626 0 _0574_
rlabel metal2 20562 16354 20562 16354 0 _0575_
rlabel metal1 24886 16728 24886 16728 0 _0576_
rlabel metal2 25070 16796 25070 16796 0 _0577_
rlabel metal1 18630 24310 18630 24310 0 _0578_
rlabel metal1 29118 16524 29118 16524 0 _0579_
rlabel metal1 39238 21454 39238 21454 0 _0580_
rlabel metal1 38318 21590 38318 21590 0 _0581_
rlabel metal2 38962 21794 38962 21794 0 _0582_
rlabel metal2 22954 16388 22954 16388 0 _0583_
rlabel metal1 16652 17646 16652 17646 0 _0584_
rlabel metal2 22862 18054 22862 18054 0 _0585_
rlabel metal2 23322 19567 23322 19567 0 _0586_
rlabel metal2 23230 32096 23230 32096 0 _0587_
rlabel metal1 35098 30906 35098 30906 0 _0588_
rlabel metal2 23506 31314 23506 31314 0 _0589_
rlabel metal2 23782 32164 23782 32164 0 _0590_
rlabel metal2 23506 33218 23506 33218 0 _0591_
rlabel metal1 33166 30158 33166 30158 0 _0592_
rlabel metal1 36386 24276 36386 24276 0 _0593_
rlabel metal1 35788 17782 35788 17782 0 _0594_
rlabel metal1 36018 24378 36018 24378 0 _0595_
rlabel metal2 36018 21488 36018 21488 0 _0596_
rlabel metal1 35098 15130 35098 15130 0 _0597_
rlabel metal1 36386 20570 36386 20570 0 _0598_
rlabel metal1 36018 20808 36018 20808 0 _0599_
rlabel metal1 36386 21114 36386 21114 0 _0600_
rlabel metal2 41906 23902 41906 23902 0 _0601_
rlabel metal1 32154 17850 32154 17850 0 _0602_
rlabel metal2 25300 23562 25300 23562 0 _0603_
rlabel metal2 31786 18258 31786 18258 0 _0604_
rlabel metal2 31970 17034 31970 17034 0 _0605_
rlabel metal2 13386 24514 13386 24514 0 _0606_
rlabel metal2 32154 17374 32154 17374 0 _0607_
rlabel metal2 36754 16490 36754 16490 0 _0608_
rlabel metal2 25530 26180 25530 26180 0 _0609_
rlabel metal1 25346 27064 25346 27064 0 _0610_
rlabel via2 32430 16235 32430 16235 0 _0611_
rlabel metal2 32614 15776 32614 15776 0 _0612_
rlabel metal1 13846 24242 13846 24242 0 _0613_
rlabel metal1 13386 24072 13386 24072 0 _0614_
rlabel metal3 19849 15980 19849 15980 0 _0615_
rlabel metal2 36662 16065 36662 16065 0 _0616_
rlabel metal2 34868 16762 34868 16762 0 _0617_
rlabel metal2 22034 28696 22034 28696 0 _0618_
rlabel metal2 27462 28458 27462 28458 0 _0619_
rlabel metal1 35006 26996 35006 26996 0 _0620_
rlabel metal1 34960 27098 34960 27098 0 _0621_
rlabel metal2 18538 30566 18538 30566 0 _0622_
rlabel metal2 15686 29274 15686 29274 0 _0623_
rlabel metal1 27324 28458 27324 28458 0 _0624_
rlabel metal2 28014 28237 28014 28237 0 _0625_
rlabel metal1 31096 18734 31096 18734 0 _0626_
rlabel metal1 30176 21454 30176 21454 0 _0627_
rlabel metal1 35742 15946 35742 15946 0 _0628_
rlabel metal2 29762 25738 29762 25738 0 _0629_
rlabel metal2 29578 25466 29578 25466 0 _0630_
rlabel metal2 30038 23222 30038 23222 0 _0631_
rlabel metal1 25392 21930 25392 21930 0 _0632_
rlabel metal1 26174 21862 26174 21862 0 _0633_
rlabel metal2 27002 21692 27002 21692 0 _0634_
rlabel metal2 30222 21148 30222 21148 0 _0635_
rlabel metal1 32706 16558 32706 16558 0 _0636_
rlabel metal1 22034 22508 22034 22508 0 _0637_
rlabel metal1 21942 22712 21942 22712 0 _0638_
rlabel via2 28474 22219 28474 22219 0 _0639_
rlabel metal1 26542 21896 26542 21896 0 _0640_
rlabel metal1 32315 21998 32315 21998 0 _0641_
rlabel metal2 32522 19346 32522 19346 0 _0642_
rlabel metal2 39974 22576 39974 22576 0 _0643_
rlabel metal2 10902 28322 10902 28322 0 _0644_
rlabel via2 35650 28475 35650 28475 0 _0645_
rlabel metal2 41170 25908 41170 25908 0 _0646_
rlabel metal1 33810 14960 33810 14960 0 _0647_
rlabel metal1 37030 24786 37030 24786 0 _0648_
rlabel metal1 37306 23222 37306 23222 0 _0649_
rlabel metal1 40434 23222 40434 23222 0 _0650_
rlabel metal2 39146 24038 39146 24038 0 _0651_
rlabel metal1 38226 22984 38226 22984 0 _0652_
rlabel metal1 38962 23290 38962 23290 0 _0653_
rlabel metal2 12650 27047 12650 27047 0 _0654_
rlabel metal2 40710 23324 40710 23324 0 _0655_
rlabel metal1 32016 29818 32016 29818 0 _0656_
rlabel metal2 5474 11934 5474 11934 0 _0657_
rlabel metal2 32154 31178 32154 31178 0 _0658_
rlabel metal2 27646 20502 27646 20502 0 _0659_
rlabel metal2 26450 20757 26450 20757 0 _0660_
rlabel metal1 26174 20026 26174 20026 0 _0661_
rlabel metal1 27646 20332 27646 20332 0 _0662_
rlabel metal1 26910 20366 26910 20366 0 _0663_
rlabel metal1 23506 20502 23506 20502 0 _0664_
rlabel metal1 27554 20536 27554 20536 0 _0665_
rlabel via2 28014 20587 28014 20587 0 _0666_
rlabel metal1 12604 14518 12604 14518 0 _0667_
rlabel metal1 32614 18258 32614 18258 0 _0668_
rlabel metal1 23506 17850 23506 17850 0 _0669_
rlabel metal2 24058 18564 24058 18564 0 _0670_
rlabel metal2 28566 18462 28566 18462 0 _0671_
rlabel metal2 32338 18428 32338 18428 0 _0672_
rlabel metal1 17388 18054 17388 18054 0 _0673_
rlabel metal1 31694 18360 31694 18360 0 _0674_
rlabel viali 42290 17646 42290 17646 0 _0675_
rlabel metal2 33994 17850 33994 17850 0 _0676_
rlabel metal1 8096 12954 8096 12954 0 _0677_
rlabel metal1 33810 17782 33810 17782 0 _0678_
rlabel metal2 32430 18598 32430 18598 0 _0679_
rlabel metal1 32545 22678 32545 22678 0 _0680_
rlabel metal1 31970 17544 31970 17544 0 _0681_
rlabel metal1 32982 17544 32982 17544 0 _0682_
rlabel via2 36570 17085 36570 17085 0 _0683_
rlabel metal1 35972 17850 35972 17850 0 _0684_
rlabel metal1 36570 17714 36570 17714 0 _0685_
rlabel metal2 36110 17442 36110 17442 0 _0686_
rlabel metal2 9706 14229 9706 14229 0 _0687_
rlabel metal1 36984 17578 36984 17578 0 _0688_
rlabel metal1 38272 17850 38272 17850 0 _0689_
rlabel metal2 37122 18564 37122 18564 0 _0690_
rlabel metal1 41722 17612 41722 17612 0 _0691_
rlabel metal1 38042 18768 38042 18768 0 _0692_
rlabel metal1 19964 14382 19964 14382 0 _0693_
rlabel metal1 4692 13498 4692 13498 0 _0694_
rlabel metal1 3956 14042 3956 14042 0 _0695_
rlabel metal1 15732 14042 15732 14042 0 _0696_
rlabel metal1 5060 18666 5060 18666 0 _0697_
rlabel metal1 5474 15436 5474 15436 0 _0698_
rlabel metal1 4462 17646 4462 17646 0 _0699_
rlabel metal1 5934 12410 5934 12410 0 _0700_
rlabel metal2 13478 20791 13478 20791 0 _0701_
rlabel metal1 14582 19754 14582 19754 0 _0702_
rlabel metal2 15226 16201 15226 16201 0 _0703_
rlabel metal1 14950 17170 14950 17170 0 _0704_
rlabel metal2 29394 20060 29394 20060 0 _0705_
rlabel metal1 12696 16082 12696 16082 0 _0706_
rlabel via2 19642 18275 19642 18275 0 _0707_
rlabel metal1 7176 13498 7176 13498 0 _0708_
rlabel metal1 5198 13906 5198 13906 0 _0709_
rlabel metal2 19366 17816 19366 17816 0 _0710_
rlabel metal1 11224 31790 11224 31790 0 _0711_
rlabel metal1 13294 20332 13294 20332 0 _0712_
rlabel metal2 8050 19074 8050 19074 0 _0713_
rlabel metal3 751 11628 751 11628 0 addr0[0]
rlabel metal3 1050 13668 1050 13668 0 addr0[1]
rlabel metal3 751 12308 751 12308 0 addr0[2]
rlabel metal3 1050 12988 1050 12988 0 addr0[3]
rlabel metal3 751 16388 751 16388 0 addr0[4]
rlabel metal3 751 15708 751 15708 0 addr0[5]
rlabel metal3 1050 15028 1050 15028 0 addr0[6]
rlabel metal3 751 14348 751 14348 0 addr0[7]
rlabel metal3 41546 29988 41546 29988 0 clk0
rlabel metal1 40112 23698 40112 23698 0 clknet_0_clk0
rlabel metal1 32246 32844 32246 32844 0 clknet_2_0__leaf_clk0
rlabel metal1 27002 34612 27002 34612 0 clknet_2_1__leaf_clk0
rlabel metal1 42458 19380 42458 19380 0 clknet_2_2__leaf_clk0
rlabel metal2 40342 21216 40342 21216 0 clknet_2_3__leaf_clk0
rlabel metal2 44574 29461 44574 29461 0 cs0
rlabel metal2 44482 15793 44482 15793 0 dout0[0]
rlabel metal1 25898 37434 25898 37434 0 dout0[10]
rlabel via2 44482 27285 44482 27285 0 dout0[11]
rlabel metal2 44482 26673 44482 26673 0 dout0[12]
rlabel metal1 44298 20774 44298 20774 0 dout0[13]
rlabel metal1 44298 29002 44298 29002 0 dout0[14]
rlabel metal1 27830 37434 27830 37434 0 dout0[15]
rlabel metal1 44298 26486 44298 26486 0 dout0[16]
rlabel metal1 44298 14042 44298 14042 0 dout0[17]
rlabel metal1 44298 23494 44298 23494 0 dout0[18]
rlabel metal1 23322 37434 23322 37434 0 dout0[19]
rlabel metal1 44298 18054 44298 18054 0 dout0[1]
rlabel via2 44482 24565 44482 24565 0 dout0[20]
rlabel metal1 44298 15334 44298 15334 0 dout0[21]
rlabel via2 44482 27931 44482 27931 0 dout0[22]
rlabel metal2 44482 14297 44482 14297 0 dout0[23]
rlabel metal2 44482 23953 44482 23953 0 dout0[24]
rlabel via2 44482 22491 44482 22491 0 dout0[25]
rlabel metal2 31602 38328 31602 38328 0 dout0[26]
rlabel via2 44482 17051 44482 17051 0 dout0[27]
rlabel via2 44482 16405 44482 16405 0 dout0[28]
rlabel metal2 44482 18513 44482 18513 0 dout0[29]
rlabel metal1 29440 37366 29440 37366 0 dout0[2]
rlabel metal1 44298 19482 44298 19482 0 dout0[30]
rlabel metal2 44482 21233 44482 21233 0 dout0[31]
rlabel metal2 21942 38328 21942 38328 0 dout0[3]
rlabel metal1 25254 37434 25254 37434 0 dout0[4]
rlabel via2 44482 21845 44482 21845 0 dout0[5]
rlabel metal2 44482 25177 44482 25177 0 dout0[6]
rlabel metal2 44482 19737 44482 19737 0 dout0[7]
rlabel metal1 29946 37434 29946 37434 0 dout0[8]
rlabel metal1 22678 37434 22678 37434 0 dout0[9]
rlabel metal1 2208 11866 2208 11866 0 net1
rlabel metal2 39054 15606 39054 15606 0 net10
rlabel via1 6856 18258 6856 18258 0 net100
rlabel metal1 12972 19414 12972 19414 0 net101
rlabel metal1 4462 17748 4462 17748 0 net102
rlabel metal1 6762 18224 6762 18224 0 net103
rlabel metal2 14398 17034 14398 17034 0 net104
rlabel metal1 5566 15674 5566 15674 0 net105
rlabel metal1 13156 15130 13156 15130 0 net106
rlabel metal1 12374 15028 12374 15028 0 net107
rlabel metal1 8970 15436 8970 15436 0 net108
rlabel metal1 7590 15504 7590 15504 0 net109
rlabel metal2 27094 35666 27094 35666 0 net11
rlabel metal1 13294 18632 13294 18632 0 net110
rlabel metal1 12604 17238 12604 17238 0 net111
rlabel metal1 14858 14994 14858 14994 0 net112
rlabel metal1 10074 12138 10074 12138 0 net113
rlabel metal1 13202 19210 13202 19210 0 net114
rlabel metal1 7682 12172 7682 12172 0 net115
rlabel metal2 18814 12886 18814 12886 0 net116
rlabel metal1 19734 12784 19734 12784 0 net117
rlabel metal1 13892 14314 13892 14314 0 net118
rlabel metal1 10580 12886 10580 12886 0 net119
rlabel metal1 41262 27336 41262 27336 0 net12
rlabel metal1 19688 12138 19688 12138 0 net120
rlabel metal2 18722 13294 18722 13294 0 net121
rlabel via1 19644 12206 19644 12206 0 net122
rlabel metal1 10028 12410 10028 12410 0 net123
rlabel metal2 17434 11934 17434 11934 0 net124
rlabel metal1 18446 32334 18446 32334 0 net125
rlabel metal1 43286 21386 43286 21386 0 net126
rlabel metal1 43792 23698 43792 23698 0 net127
rlabel metal2 42826 18836 42826 18836 0 net128
rlabel metal2 21942 33660 21942 33660 0 net129
rlabel metal1 42550 26894 42550 26894 0 net13
rlabel metal1 6302 14348 6302 14348 0 net130
rlabel metal1 8326 13872 8326 13872 0 net131
rlabel metal1 6348 14450 6348 14450 0 net132
rlabel metal1 6026 14960 6026 14960 0 net133
rlabel metal1 7406 17238 7406 17238 0 net134
rlabel metal1 6992 14518 6992 14518 0 net135
rlabel metal1 7590 17034 7590 17034 0 net136
rlabel metal1 2070 16116 2070 16116 0 net137
rlabel via1 5737 12138 5737 12138 0 net138
rlabel metal1 6394 13396 6394 13396 0 net139
rlabel metal2 44298 21495 44298 21495 0 net14
rlabel metal1 5658 12206 5658 12206 0 net140
rlabel metal1 6578 13362 6578 13362 0 net141
rlabel metal1 5428 12138 5428 12138 0 net142
rlabel metal2 4830 13617 4830 13617 0 net143
rlabel metal1 6394 12274 6394 12274 0 net144
rlabel metal1 6565 13226 6565 13226 0 net145
rlabel metal1 42642 17714 42642 17714 0 net146
rlabel metal1 42366 20366 42366 20366 0 net147
rlabel metal1 42320 18190 42320 18190 0 net148
rlabel metal1 40986 23018 40986 23018 0 net149
rlabel metal1 40250 29002 40250 29002 0 net15
rlabel metal2 43838 21216 43838 21216 0 net150
rlabel metal1 25300 33966 25300 33966 0 net151
rlabel metal2 41722 23290 41722 23290 0 net152
rlabel metal1 42458 24582 42458 24582 0 net153
rlabel via2 40986 26979 40986 26979 0 net154
rlabel metal1 42504 27642 42504 27642 0 net155
rlabel metal2 43654 23834 43654 23834 0 net156
rlabel metal1 40342 26962 40342 26962 0 net157
rlabel metal1 26910 33490 26910 33490 0 net158
rlabel metal1 41952 15130 41952 15130 0 net159
rlabel metal1 28290 34714 28290 34714 0 net16
rlabel via1 41077 26962 41077 26962 0 net160
rlabel metal2 24150 34544 24150 34544 0 net161
rlabel metal2 40894 18564 40894 18564 0 net162
rlabel metal2 23414 33796 23414 33796 0 net163
rlabel metal1 41906 21998 41906 21998 0 net164
rlabel metal2 32154 32572 32154 32572 0 net165
rlabel metal1 39560 28526 39560 28526 0 net166
rlabel metal1 28612 33082 28612 33082 0 net167
rlabel metal2 38778 16422 38778 16422 0 net168
rlabel metal2 22678 34476 22678 34476 0 net169
rlabel metal2 43746 25840 43746 25840 0 net17
rlabel metal1 38640 17170 38640 17170 0 net170
rlabel metal1 28336 33422 28336 33422 0 net171
rlabel metal1 42412 17850 42412 17850 0 net172
rlabel metal2 30222 33082 30222 33082 0 net173
rlabel metal2 41538 25500 41538 25500 0 net174
rlabel metal1 36570 16082 36570 16082 0 net175
rlabel metal1 36294 16116 36294 16116 0 net176
rlabel metal2 40434 19516 40434 19516 0 net177
rlabel metal2 43102 14416 43102 14416 0 net18
rlabel metal2 43562 21828 43562 21828 0 net19
rlabel metal2 2346 14178 2346 14178 0 net2
rlabel metal2 23690 35938 23690 35938 0 net20
rlabel metal2 43194 18496 43194 18496 0 net21
rlabel metal2 43010 24684 43010 24684 0 net22
rlabel metal1 41906 15368 41906 15368 0 net23
rlabel metal2 43010 28220 43010 28220 0 net24
rlabel metal2 44298 15164 44298 15164 0 net25
rlabel metal2 43010 23834 43010 23834 0 net26
rlabel metal2 42458 22848 42458 22848 0 net27
rlabel metal1 32154 33082 32154 33082 0 net28
rlabel metal2 43838 17476 43838 17476 0 net29
rlabel metal1 2484 12410 2484 12410 0 net3
rlabel metal1 40526 17306 40526 17306 0 net30
rlabel metal1 41630 18258 41630 18258 0 net31
rlabel metal1 29900 34034 29900 34034 0 net32
rlabel metal1 43838 19278 43838 19278 0 net33
rlabel metal2 44206 20706 44206 20706 0 net34
rlabel metal2 22402 36414 22402 36414 0 net35
rlabel metal1 25530 34714 25530 34714 0 net36
rlabel metal1 43608 21862 43608 21862 0 net37
rlabel metal1 43930 26554 43930 26554 0 net38
rlabel metal2 43286 20366 43286 20366 0 net39
rlabel metal1 1702 12818 1702 12818 0 net4
rlabel metal1 30682 33490 30682 33490 0 net40
rlabel metal1 23506 34170 23506 34170 0 net41
rlabel metal2 41814 20638 41814 20638 0 net42
rlabel metal1 40296 21998 40296 21998 0 net43
rlabel metal1 38870 16694 38870 16694 0 net44
rlabel metal1 36685 32538 36685 32538 0 net45
rlabel metal1 21666 16456 21666 16456 0 net46
rlabel metal2 29026 13770 29026 13770 0 net47
rlabel metal1 28612 13906 28612 13906 0 net48
rlabel metal1 8418 12852 8418 12852 0 net49
rlabel metal1 2162 16558 2162 16558 0 net5
rlabel metal2 13018 12138 13018 12138 0 net50
rlabel metal1 11914 12138 11914 12138 0 net51
rlabel metal1 8970 12784 8970 12784 0 net52
rlabel via1 17528 12206 17528 12206 0 net53
rlabel metal2 10442 19584 10442 19584 0 net54
rlabel metal1 13432 19958 13432 19958 0 net55
rlabel metal1 12742 20400 12742 20400 0 net56
rlabel metal1 15686 16014 15686 16014 0 net57
rlabel metal1 11592 21930 11592 21930 0 net58
rlabel metal2 6946 16116 6946 16116 0 net59
rlabel metal1 1932 16218 1932 16218 0 net6
rlabel metal1 8924 17646 8924 17646 0 net60
rlabel metal2 12650 23018 12650 23018 0 net61
rlabel metal1 4922 16524 4922 16524 0 net62
rlabel metal2 5934 17068 5934 17068 0 net63
rlabel via1 2624 19346 2624 19346 0 net64
rlabel metal1 4580 20910 4580 20910 0 net65
rlabel metal2 3450 19652 3450 19652 0 net66
rlabel metal2 2714 21012 2714 21012 0 net67
rlabel metal1 12282 23120 12282 23120 0 net68
rlabel metal1 2392 19278 2392 19278 0 net69
rlabel metal2 2806 15878 2806 15878 0 net7
rlabel via1 12262 20910 12262 20910 0 net70
rlabel metal2 2438 18258 2438 18258 0 net71
rlabel metal2 2622 16388 2622 16388 0 net72
rlabel metal1 11500 12206 11500 12206 0 net73
rlabel metal1 9062 13498 9062 13498 0 net74
rlabel metal2 7498 13345 7498 13345 0 net75
rlabel metal1 4140 12954 4140 12954 0 net76
rlabel metal2 2530 14518 2530 14518 0 net77
rlabel metal1 10212 19346 10212 19346 0 net78
rlabel metal1 10028 20502 10028 20502 0 net79
rlabel metal1 2024 14586 2024 14586 0 net8
rlabel metal1 9522 15980 9522 15980 0 net80
rlabel metal1 10304 20978 10304 20978 0 net81
rlabel metal2 8142 12954 8142 12954 0 net82
rlabel metal1 2346 18258 2346 18258 0 net83
rlabel via1 12928 15470 12928 15470 0 net84
rlabel metal1 2668 23086 2668 23086 0 net85
rlabel metal1 15042 20808 15042 20808 0 net86
rlabel metal1 12558 19822 12558 19822 0 net87
rlabel metal1 12790 18734 12790 18734 0 net88
rlabel metal1 13662 20434 13662 20434 0 net89
rlabel metal1 42504 28118 42504 28118 0 net9
rlabel metal1 12282 13192 12282 13192 0 net90
rlabel metal1 9062 16558 9062 16558 0 net91
rlabel metal1 9430 16524 9430 16524 0 net92
rlabel metal1 6348 15470 6348 15470 0 net93
rlabel metal2 12834 15283 12834 15283 0 net94
rlabel metal2 18722 16320 18722 16320 0 net95
rlabel metal1 9522 16456 9522 16456 0 net96
rlabel metal2 17986 16286 17986 16286 0 net97
rlabel metal1 5290 18360 5290 18360 0 net98
rlabel metal1 14260 17238 14260 17238 0 net99
<< properties >>
string FIXED_BBOX 0 0 46000 40000
<< end >>
