assign table1[0] = 32'h7fffffff;
assign table1[1] = 32'h7fff6215;
assign table1[2] = 32'h7ffd8859;
assign table1[3] = 32'h7ffa72d0;
assign table1[4] = 32'h7ff62181;
assign table1[5] = 32'h7ff09477;
assign table1[6] = 32'h7fe9cbbf;
assign table1[7] = 32'h7fe1c76a;
assign table1[8] = 32'h7fd8878d;
assign table1[9] = 32'h7fce0c3d;
assign table1[10] = 32'h7fc25595;
assign table1[11] = 32'h7fb563b2;
assign table1[12] = 32'h7fa736b3;
assign table1[13] = 32'h7f97cebc;
assign table1[14] = 32'h7f872bf2;
assign table1[15] = 32'h7f754e7f;
assign table1[16] = 32'h7f62368e;
assign table1[17] = 32'h7f4de450;
assign table1[18] = 32'h7f3857f5;
assign table1[19] = 32'h7f2191b3;
assign table1[20] = 32'h7f0991c3;
assign table1[21] = 32'h7ef0585f;
assign table1[22] = 32'h7ed5e5c5;
assign table1[23] = 32'h7eba3a38;
assign table1[24] = 32'h7e9d55fb;
assign table1[25] = 32'h7e7f3956;
assign table1[26] = 32'h7e5fe492;
assign table1[27] = 32'h7e3f57fe;
assign table1[28] = 32'h7e1d93e9;
assign table1[29] = 32'h7dfa98a7;
assign table1[30] = 32'h7dd6668e;
assign table1[31] = 32'h7db0fdf7;
assign table1[32] = 32'h7d8a5f3f;
assign table1[33] = 32'h7d628ac5;
assign table1[34] = 32'h7d3980eb;
assign table1[35] = 32'h7d0f4217;
assign table1[36] = 32'h7ce3ceb1;
assign table1[37] = 32'h7cb72723;
assign table1[38] = 32'h7c894bdd;
assign table1[39] = 32'h7c5a3d4f;
assign table1[40] = 32'h7c29fbed;
assign table1[41] = 32'h7bf8882f;
assign table1[42] = 32'h7bc5e28f;
assign table1[43] = 32'h7b920b88;
assign table1[44] = 32'h7b5d039d;
assign table1[45] = 32'h7b26cb4e;
assign table1[46] = 32'h7aef6323;
assign table1[47] = 32'h7ab6cba3;
assign table1[48] = 32'h7a7d055a;
assign table1[49] = 32'h7a4210d8;
assign table1[50] = 32'h7a05eeac;
assign table1[51] = 32'h79c89f6d;
assign table1[52] = 32'h798a23b0;
assign table1[53] = 32'h794a7c11;
assign table1[54] = 32'h7909a92c;
assign table1[55] = 32'h78c7aba1;
assign table1[56] = 32'h78848413;
assign table1[57] = 32'h78403328;
assign table1[58] = 32'h77fab988;
assign table1[59] = 32'h77b417df;
assign table1[60] = 32'h776c4eda;
assign table1[61] = 32'h77235f2c;
assign table1[62] = 32'h76d94988;
assign table1[63] = 32'h768e0ea5;
assign table1[64] = 32'h7641af3c;
assign table1[65] = 32'h75f42c0a;
assign table1[66] = 32'h75a585ce;
assign table1[67] = 32'h7555bd4b;
assign table1[68] = 32'h7504d344;
assign table1[69] = 32'h74b2c883;
assign table1[70] = 32'h745f9dd0;
assign table1[71] = 32'h740b53fa;
assign table1[72] = 32'h73b5ebd0;
assign table1[73] = 32'h735f6625;
assign table1[74] = 32'h7307c3cf;
assign table1[75] = 32'h72af05a6;
assign table1[76] = 32'h72552c84;
assign table1[77] = 32'h71fa3948;
assign table1[78] = 32'h719e2cd1;
assign table1[79] = 32'h71410804;
assign table1[80] = 32'h70e2cbc5;
assign table1[81] = 32'h708378fe;
assign table1[82] = 32'h70231099;
assign table1[83] = 32'h6fc19384;
assign table1[84] = 32'h6f5f02b1;
assign table1[85] = 32'h6efb5f11;
assign table1[86] = 32'h6e96a99c;
assign table1[87] = 32'h6e30e349;
assign table1[88] = 32'h6dca0d14;
assign table1[89] = 32'h6d6227f9;
assign table1[90] = 32'h6cf934fb;
assign table1[91] = 32'h6c8f351b;
assign table1[92] = 32'h6c24295f;
assign table1[93] = 32'h6bb812d0;
assign table1[94] = 32'h6b4af278;
assign table1[95] = 32'h6adcc964;
assign table1[96] = 32'h6a6d98a3;
assign table1[97] = 32'h69fd614a;
assign table1[98] = 32'h698c246b;
assign table1[99] = 32'h6919e31f;
assign table1[100] = 32'h68a69e80;
assign table1[101] = 32'h683257aa;
assign table1[102] = 32'h67bd0fbc;
assign table1[103] = 32'h6746c7d7;
assign table1[104] = 32'h66cf811f;
assign table1[105] = 32'h66573cbb;
assign table1[106] = 32'h65ddfbd2;
assign table1[107] = 32'h6563bf91;
assign table1[108] = 32'h64e88925;
assign table1[109] = 32'h646c59bf;
assign table1[110] = 32'h63ef328f;
assign table1[111] = 32'h637114cc;
assign table1[112] = 32'h62f201ac;
assign table1[113] = 32'h6271fa68;
assign table1[114] = 32'h61f1003e;
assign table1[115] = 32'h616f146b;
assign table1[116] = 32'h60ec382f;
assign table1[117] = 32'h60686cce;
assign table1[118] = 32'h5fe3b38d;
assign table1[119] = 32'h5f5e0db2;
assign table1[120] = 32'h5ed77c89;
assign table1[121] = 32'h5e50015d;
assign table1[122] = 32'h5dc79d7b;
assign table1[123] = 32'h5d3e5236;
assign table1[124] = 32'h5cb420df;
assign table1[125] = 32'h5c290acc;
assign table1[126] = 32'h5b9d1153;
assign table1[127] = 32'h5b1035ce;
assign table1[128] = 32'h5a827999;
assign table1[129] = 32'h59f3de12;
assign table1[130] = 32'h59646497;
assign table1[131] = 32'h58d40e8c;
assign table1[132] = 32'h5842dd54;
assign table1[133] = 32'h57b0d255;
assign table1[134] = 32'h571deef9;
assign table1[135] = 32'h568a34a9;
assign table1[136] = 32'h55f5a4d2;
assign table1[137] = 32'h556040e2;
assign table1[138] = 32'h54ca0a4a;
assign table1[139] = 32'h5433027d;
assign table1[140] = 32'h539b2aef;
assign table1[141] = 32'h53028517;
assign table1[142] = 32'h5269126e;
assign table1[143] = 32'h51ced46e;
assign table1[144] = 32'h5133cc94;
assign table1[145] = 32'h5097fc5e;
assign table1[146] = 32'h4ffb654c;
assign table1[147] = 32'h4f5e08e2;
assign table1[148] = 32'h4ebfe8a4;
assign table1[149] = 32'h4e210617;
assign table1[150] = 32'h4d8162c3;
assign table1[151] = 32'h4ce10034;
assign table1[152] = 32'h4c3fdff3;
assign table1[153] = 32'h4b9e038f;
assign table1[154] = 32'h4afb6c97;
assign table1[155] = 32'h4a581c9d;
assign table1[156] = 32'h49b41533;
assign table1[157] = 32'h490f57ee;
assign table1[158] = 32'h4869e664;
assign table1[159] = 32'h47c3c22e;
assign table1[160] = 32'h471cece6;
assign table1[161] = 32'h46756827;
assign table1[162] = 32'h45cd358f;
assign table1[163] = 32'h452456bc;
assign table1[164] = 32'h447acd50;
assign table1[165] = 32'h43d09aec;
assign table1[166] = 32'h4325c135;
assign table1[167] = 32'h427a41d0;
assign table1[168] = 32'h41ce1e64;
assign table1[169] = 32'h4121589a;
assign table1[170] = 32'h4073f21d;
assign table1[171] = 32'h3fc5ec97;
assign table1[172] = 32'h3f1749b7;
assign table1[173] = 32'h3e680b2c;
assign table1[174] = 32'h3db832a5;
assign table1[175] = 32'h3d07c1d5;
assign table1[176] = 32'h3c56ba70;
assign table1[177] = 32'h3ba51e29;
assign table1[178] = 32'h3af2eeb7;
assign table1[179] = 32'h3a402dd1;
assign table1[180] = 32'h398cdd32;
assign table1[181] = 32'h38d8fe93;
assign table1[182] = 32'h382493b0;
assign table1[183] = 32'h376f9e46;
assign table1[184] = 32'h36ba2013;
assign table1[185] = 32'h36041ad9;
assign table1[186] = 32'h354d9056;
assign table1[187] = 32'h3496824f;
assign table1[188] = 32'h33def287;
assign table1[189] = 32'h3326e2c2;
assign table1[190] = 32'h326e54c7;
assign table1[191] = 32'h31b54a5d;
assign table1[192] = 32'h30fbc54d;
assign table1[193] = 32'h3041c760;
assign table1[194] = 32'h2f875262;
assign table1[195] = 32'h2ecc681e;
assign table1[196] = 32'h2e110a62;
assign table1[197] = 32'h2d553afb;
assign table1[198] = 32'h2c98fbba;
assign table1[199] = 32'h2bdc4e6f;
assign table1[200] = 32'h2b1f34eb;
assign table1[201] = 32'h2a61b101;
assign table1[202] = 32'h29a3c485;
assign table1[203] = 32'h28e5714a;
assign table1[204] = 32'h2826b928;
assign table1[205] = 32'h27679df4;
assign table1[206] = 32'h26a82185;
assign table1[207] = 32'h25e845b6;
assign table1[208] = 32'h25280c5d;
assign table1[209] = 32'h24677757;
assign table1[210] = 32'h23a6887e;
assign table1[211] = 32'h22e541af;
assign table1[212] = 32'h2223a4c5;
assign table1[213] = 32'h2161b39f;
assign table1[214] = 32'h209f701c;
assign table1[215] = 32'h1fdcdc1b;
assign table1[216] = 32'h1f19f97b;
assign table1[217] = 32'h1e56ca1e;
assign table1[218] = 32'h1d934fe5;
assign table1[219] = 32'h1ccf8cb3;
assign table1[220] = 32'h1c0b826a;
assign table1[221] = 32'h1b4732ef;
assign table1[222] = 32'h1a82a025;
assign table1[223] = 32'h19bdcbf3;
assign table1[224] = 32'h18f8b83c;
assign table1[225] = 32'h183366e8;
assign table1[226] = 32'h176dd9de;
assign table1[227] = 32'h16a81305;
assign table1[228] = 32'h15e21444;
assign table1[229] = 32'h151bdf85;
assign table1[230] = 32'h145576b1;
assign table1[231] = 32'h138edbb1;
assign table1[232] = 32'h12c8106e;
assign table1[233] = 32'h120116d5;
assign table1[234] = 32'h1139f0cf;
assign table1[235] = 32'h1072a048;
assign table1[236] = 32'h0fab272b;
assign table1[237] = 32'h0ee38766;
assign table1[238] = 32'h0e1bc2e4;
assign table1[239] = 32'h0d53db92;
assign table1[240] = 32'h0c8bd35e;
assign table1[241] = 32'h0bc3ac35;
assign table1[242] = 32'h0afb6805;
assign table1[243] = 32'h0a3308bc;
assign table1[244] = 32'h096a9049;
assign table1[245] = 32'h08a2009a;
assign table1[246] = 32'h07d95b9e;
assign table1[247] = 32'h0710a345;
assign table1[248] = 32'h0647d97c;
assign table1[249] = 32'h057f0035;
assign table1[250] = 32'h04b6195d;
assign table1[251] = 32'h03ed26e6;
assign table1[252] = 32'h03242abf;
assign table1[253] = 32'h025b26d7;
assign table1[254] = 32'h01921d20;
assign table1[255] = 32'h00c90f88;
