* NGSPICE file created from cust_rom.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

.subckt cust_rom addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] clk0
+ cs0 dout0[0] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[1]
+ dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] vccd1 vssd1
XFILLER_0_27_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_432_ net57 net65 _085_ _142_ vssd1 vssd1 vccd1 vccd1 _005_ sky130_fd_sc_hd__a22o_1
X_363_ _194_ net30 net28 _195_ vssd1 vssd1 vccd1 vccd1 _079_ sky130_fd_sc_hd__a22o_1
X_294_ _233_ _234_ vssd1 vssd1 vccd1 vccd1 _235_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_15_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_501_ clknet_1_1__leaf_clk0 _012_ vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_415_ _191_ _228_ vssd1 vssd1 vccd1 vccd1 _127_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_346_ _204_ net29 net27 _206_ vssd1 vssd1 vccd1 vccd1 _062_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_277_ _200_ net40 net37 _199_ _217_ vssd1 vssd1 vccd1 vccd1 _218_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_329_ addr0_reg\[6\] net36 net47 vssd1 vssd1 vccd1 vccd1 _045_ sky130_fd_sc_hd__and3b_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_78 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 dout0[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_18_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_68 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_500_ clknet_1_1__leaf_clk0 _011_ vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__dfxtp_1
X_431_ _137_ _141_ vssd1 vssd1 vccd1 vccd1 _142_ sky130_fd_sc_hd__or2_1
X_362_ _215_ net29 net27 _216_ vssd1 vssd1 vccd1 vccd1 _078_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_15_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_293_ net40 net37 _192_ vssd1 vssd1 vccd1 vccd1 _234_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_13_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_414_ _202_ _053_ _054_ vssd1 vssd1 vccd1 vccd1 _126_ sky130_fd_sc_hd__or3_1
X_345_ _059_ _060_ vssd1 vssd1 vccd1 vccd1 _061_ sky130_fd_sc_hd__or2_1
X_276_ net40 _215_ _216_ net37 vssd1 vssd1 vccd1 vccd1 _217_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_259_ net52 net54 net50 net48 vssd1 vssd1 vccd1 vccd1 _200_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_10_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_328_ _215_ net33 net31 _216_ vssd1 vssd1 vccd1 vccd1 _044_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Left_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput10 net10 vssd1 vssd1 vccd1 vccd1 dout0[10] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_18_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 dout0[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_69 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_430_ _197_ _101_ _139_ _140_ vssd1 vssd1 vccd1 vccd1 _141_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_15_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_292_ _189_ net40 net37 _190_ vssd1 vssd1 vccd1 vccd1 _233_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_361_ _222_ net29 net27 _223_ vssd1 vssd1 vccd1 vccd1 _077_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_20_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_413_ _072_ _075_ _124_ vssd1 vssd1 vccd1 vccd1 _125_ sky130_fd_sc_hd__or3_1
X_344_ _216_ net29 net27 _215_ vssd1 vssd1 vccd1 vccd1 _060_ sky130_fd_sc_hd__a22o_1
X_275_ net50 net48 net52 net54 vssd1 vssd1 vccd1 vccd1 _216_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Left_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_258_ net48 net52 net54 net50 vssd1 vssd1 vccd1 vccd1 _199_ sky130_fd_sc_hd__nor4b_2
X_327_ _222_ net33 net31 _223_ vssd1 vssd1 vccd1 vccd1 _043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold10 net23 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_11_Left_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput11 net11 vssd1 vssd1 vccd1 vccd1 dout0[11] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_18_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput9 net9 vssd1 vssd1 vccd1 vccd1 dout0[0] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 dout0[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_23_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_291_ net38 _222_ net35 net41 _231_ vssd1 vssd1 vccd1 vccd1 _232_ sky130_fd_sc_hd__a221o_1
X_360_ _072_ _075_ vssd1 vssd1 vccd1 vccd1 _076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_489_ clknet_1_0__leaf_clk0 _000_ vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_20_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_412_ _043_ _050_ _080_ vssd1 vssd1 vccd1 vccd1 _124_ sky130_fd_sc_hd__or3_1
X_343_ net42 net30 net28 _200_ vssd1 vssd1 vccd1 vccd1 _059_ sky130_fd_sc_hd__a22o_1
X_274_ net52 net54 net50 net48 vssd1 vssd1 vccd1 vccd1 _215_ sky130_fd_sc_hd__and4b_2
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_257_ net43 _194_ _195_ net45 vssd1 vssd1 vccd1 vccd1 _198_ sky130_fd_sc_hd__a22o_1
X_326_ _035_ _041_ vssd1 vssd1 vccd1 vccd1 _042_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_9_90 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_309_ addr0_reg\[4\] addr0_reg\[6\] net36 vssd1 vssd1 vccd1 vccd1 _025_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold11 net12 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_80 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 dout0[8] sky130_fd_sc_hd__buf_2
Xoutput12 net12 vssd1 vssd1 vccd1 vccd1 dout0[12] sky130_fd_sc_hd__buf_2
XFILLER_0_7_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_290_ _195_ net41 net38 _194_ vssd1 vssd1 vccd1 vccd1 _231_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_488_ clknet_1_0__leaf_clk0 net7 vssd1 vssd1 vccd1 vccd1 addr0_reg\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_70 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_411_ net56 net61 net25 _123_ vssd1 vssd1 vccd1 vccd1 _003_ sky130_fd_sc_hd__a22o_1
X_342_ net47 addr0_reg\[5\] addr0_reg\[6\] vssd1 vssd1 vccd1 vccd1 _058_ sky130_fd_sc_hd__nor3_1
X_273_ _200_ net40 net37 _199_ vssd1 vssd1 vccd1 vccd1 _214_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_256_ _188_ _191_ _196_ vssd1 vssd1 vccd1 vccd1 _197_ sky130_fd_sc_hd__or3_1
X_325_ _036_ _037_ _038_ _039_ vssd1 vssd1 vccd1 vccd1 _041_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_0_60 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload0 clknet_1_1__leaf_clk0 vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_24_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_308_ net46 _204_ _206_ net44 vssd1 vssd1 vccd1 vccd1 _024_ sky130_fd_sc_hd__a22o_1
Xhold12 net24 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_10_91 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_81 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput13 net13 vssd1 vssd1 vccd1 vccd1 dout0[13] sky130_fd_sc_hd__buf_2
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 dout0[9] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_487_ clknet_1_0__leaf_clk0 net6 vssd1 vssd1 vccd1 vccd1 addr0_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_71 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_410_ _097_ _120_ _121_ _122_ vssd1 vssd1 vccd1 vccd1 _123_ sky130_fd_sc_hd__or4_1
X_341_ addr0_reg\[6\] addr0_reg\[5\] net47 vssd1 vssd1 vccd1 vccd1 _057_ sky130_fd_sc_hd__and3b_1
X_272_ _211_ _212_ vssd1 vssd1 vccd1 vccd1 _213_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_324_ _036_ _038_ vssd1 vssd1 vccd1 vccd1 _040_ sky130_fd_sc_hd__or2_1
X_255_ net45 _194_ _195_ net43 vssd1 vssd1 vccd1 vccd1 _196_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_61 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_28_Left_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_307_ _021_ _022_ vssd1 vssd1 vccd1 vccd1 _023_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold13 net16 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_10_92 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput14 net14 vssd1 vssd1 vccd1 vccd1 dout0[14] sky130_fd_sc_hd__buf_2
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_486_ clknet_1_0__leaf_clk0 net5 vssd1 vssd1 vccd1 vccd1 addr0_reg\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_72 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_271_ _184_ net44 _187_ net46 vssd1 vssd1 vccd1 vccd1 _212_ sky130_fd_sc_hd__a22o_1
X_340_ _035_ _041_ _049_ _055_ vssd1 vssd1 vccd1 vccd1 _056_ sky130_fd_sc_hd__nor4_1
X_469_ _126_ _171_ _172_ _173_ vssd1 vssd1 vccd1 vccd1 _174_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_323_ _190_ net34 net32 _189_ vssd1 vssd1 vccd1 vccd1 _039_ sky130_fd_sc_hd__a22o_1
X_254_ net49 net53 net55 net51 vssd1 vssd1 vccd1 vccd1 _195_ sky130_fd_sc_hd__and4bb_2
XTAP_TAPCELL_ROW_0_62 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_306_ net43 _215_ _216_ net45 vssd1 vssd1 vccd1 vccd1 _022_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_3_Left_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold14 net13 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_93 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput15 net15 vssd1 vssd1 vccd1 vccd1 dout0[15] sky130_fd_sc_hd__buf_2
XFILLER_0_7_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_485_ clknet_1_0__leaf_clk0 net4 vssd1 vssd1 vccd1 vccd1 addr0_reg\[3\] sky130_fd_sc_hd__dfxtp_1
X_270_ net44 _189_ _190_ net46 vssd1 vssd1 vccd1 vccd1 _211_ sky130_fd_sc_hd__a22o_1
X_468_ _224_ _019_ _022_ _078_ vssd1 vssd1 vccd1 vccd1 _173_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_399_ _030_ _067_ vssd1 vssd1 vccd1 vccd1 _113_ sky130_fd_sc_hd__or2_1
X_322_ _195_ net34 net32 _194_ vssd1 vssd1 vccd1 vccd1 _038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_253_ net51 net49 net53 net55 vssd1 vssd1 vccd1 vccd1 _194_ sky130_fd_sc_hd__and4b_2
XTAP_TAPCELL_ROW_0_63 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout50 addr0_reg\[2\] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_2
XFILLER_0_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_305_ net43 _222_ net35 net45 vssd1 vssd1 vccd1 vccd1 _021_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold15 net9 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput16 net16 vssd1 vssd1 vccd1 vccd1 dout0[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_484_ clknet_1_0__leaf_clk0 net3 vssd1 vssd1 vccd1 vccd1 addr0_reg\[2\] sky130_fd_sc_hd__dfxtp_1
X_398_ _229_ _235_ _040_ _052_ vssd1 vssd1 vccd1 vccd1 _112_ sky130_fd_sc_hd__or4_1
X_467_ _188_ _016_ _127_ vssd1 vssd1 vccd1 vccd1 _172_ sky130_fd_sc_hd__or3_1
Xclkbuf_1_0__f_clk0 clknet_0_clk0 vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout40 _203_ vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_2
X_321_ net33 net31 _192_ vssd1 vssd1 vccd1 vccd1 _037_ sky130_fd_sc_hd__o21ba_1
X_252_ net46 net44 _192_ vssd1 vssd1 vccd1 vccd1 _193_ sky130_fd_sc_hd__o21ba_1
Xfanout51 addr0_reg\[2\] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_1
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_304_ _240_ _016_ _018_ _019_ vssd1 vssd1 vccd1 vccd1 _020_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold16 net19 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput17 net17 vssd1 vssd1 vccd1 vccd1 dout0[2] sky130_fd_sc_hd__buf_2
XFILLER_0_27_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_483_ clknet_1_0__leaf_clk0 net2 vssd1 vssd1 vccd1 vccd1 addr0_reg\[1\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_19_Left_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_466_ _047_ _064_ vssd1 vssd1 vccd1 vccd1 _171_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_397_ _082_ _108_ _110_ vssd1 vssd1 vccd1 vccd1 _111_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout41 _203_ vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_2
X_320_ _187_ net34 net32 _184_ vssd1 vssd1 vccd1 vccd1 _036_ sky130_fd_sc_hd__a22o_1
Xfanout30 _057_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_2
X_251_ net50 net52 net54 net48 vssd1 vssd1 vccd1 vccd1 _192_ sky130_fd_sc_hd__or4b_1
Xfanout52 addr0_reg\[1\] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_2
X_449_ _212_ _031_ _045_ _070_ vssd1 vssd1 vccd1 vccd1 _157_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_303_ net45 _222_ net35 net43 vssd1 vssd1 vccd1 vccd1 _019_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput18 net18 vssd1 vssd1 vccd1 vccd1 dout0[3] sky130_fd_sc_hd__buf_2
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_482_ clknet_1_0__leaf_clk0 net1 vssd1 vssd1 vccd1 vccd1 addr0_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_465_ net57 net60 _085_ _170_ vssd1 vssd1 vccd1 vccd1 _010_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_20_Left_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_396_ _226_ _102_ _109_ vssd1 vssd1 vccd1 vccd1 _110_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_250_ net46 _189_ _190_ net44 vssd1 vssd1 vccd1 vccd1 _191_ sky130_fd_sc_hd__a22o_1
Xfanout53 addr0_reg\[1\] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_1
Xfanout31 _029_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_2
XFILLER_0_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_448_ _188_ _193_ _074_ vssd1 vssd1 vccd1 vccd1 _156_ sky130_fd_sc_hd__or3_1
X_379_ _059_ _064_ vssd1 vssd1 vccd1 vccd1 _094_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_302_ net43 net42 _200_ net45 vssd1 vssd1 vccd1 vccd1 _018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput19 net19 vssd1 vssd1 vccd1 vccd1 dout0[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_481_ net56 net59 _027_ vssd1 vssd1 vccd1 vccd1 _015_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_464_ _156_ _167_ _169_ vssd1 vssd1 vccd1 vccd1 _170_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_395_ _207_ _220_ _046_ vssd1 vssd1 vccd1 vccd1 _109_ sky130_fd_sc_hd__or3_1
Xfanout43 net44 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_2
Xfanout32 _029_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout54 addr0_reg\[0\] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_447_ _089_ _098_ _115_ vssd1 vssd1 vccd1 vccd1 _155_ sky130_fd_sc_hd__or3_1
X_378_ net72 net56 net25 _093_ vssd1 vssd1 vccd1 vccd1 _000_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_301_ _240_ _016_ vssd1 vssd1 vccd1 vccd1 _017_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_480_ net8 net58 _084_ vssd1 vssd1 vccd1 vccd1 _014_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_7_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_463_ _035_ _066_ _112_ _168_ vssd1 vssd1 vccd1 vccd1 _169_ sky130_fd_sc_hd__or4_1
X_394_ _240_ _018_ _069_ _073_ vssd1 vssd1 vccd1 vccd1 _108_ sky130_fd_sc_hd__or4_1
Xfanout55 addr0_reg\[0\] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__buf_1
Xfanout44 _186_ vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_2
Xfanout33 _028_ vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_2
X_446_ net56 net66 net25 _154_ vssd1 vssd1 vccd1 vccd1 _007_ sky130_fd_sc_hd__a22o_1
X_377_ _239_ _087_ _088_ _092_ vssd1 vssd1 vccd1 vccd1 _093_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_9_88 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_300_ net43 net39 _206_ net45 vssd1 vssd1 vccd1 vccd1 _016_ sky130_fd_sc_hd__a22o_1
X_429_ _233_ _019_ _053_ _060_ vssd1 vssd1 vccd1 vccd1 _140_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput1 addr0[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_393_ net56 net70 net25 _107_ vssd1 vssd1 vccd1 vccd1 _001_ sky130_fd_sc_hd__a22o_1
X_462_ _017_ _047_ _081_ _099_ vssd1 vssd1 vccd1 vccd1 _168_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout45 net46 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_2
Xfanout34 _028_ vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_0_58 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout56 _182_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_89 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_376_ _040_ _068_ _089_ _091_ vssd1 vssd1 vccd1 vccd1 _092_ sky130_fd_sc_hd__or4_1
X_445_ _227_ _152_ _153_ vssd1 vssd1 vccd1 vccd1 _154_ sky130_fd_sc_hd__or3_1
X_428_ _052_ _103_ _129_ _138_ vssd1 vssd1 vccd1 vccd1 _139_ sky130_fd_sc_hd__or4_1
X_359_ _073_ _074_ vssd1 vssd1 vccd1 vccd1 _075_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 addr0[1] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_27_Left_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_79 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap42 _199_ vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_461_ _202_ _211_ _224_ _166_ vssd1 vssd1 vccd1 vccd1 _167_ sky130_fd_sc_hd__or4_1
X_392_ _097_ _104_ _106_ vssd1 vssd1 vccd1 vccd1 _107_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout57 _182_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_0_59 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout46 _183_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_2
X_375_ _213_ _030_ _031_ _090_ vssd1 vssd1 vccd1 vccd1 _091_ sky130_fd_sc_hd__or4_1
X_444_ _075_ _113_ _129_ _149_ vssd1 vssd1 vccd1 vccd1 _153_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_427_ net39 net29 net27 _206_ _080_ vssd1 vssd1 vccd1 vccd1 _138_ sky130_fd_sc_hd__a221o_1
X_358_ _189_ net30 net28 _190_ vssd1 vssd1 vccd1 vccd1 _074_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_289_ _228_ _229_ vssd1 vssd1 vccd1 vccd1 _230_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput3 addr0[2] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_391_ _101_ _102_ _105_ vssd1 vssd1 vccd1 vccd1 _106_ sky130_fd_sc_hd__or3_1
X_460_ _217_ _021_ _024_ _060_ vssd1 vssd1 vccd1 vccd1 _166_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout47 addr0_reg\[4\] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_2
Xfanout25 _085_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_2
X_443_ _020_ _094_ _151_ vssd1 vssd1 vccd1 vccd1 _152_ sky130_fd_sc_hd__or3_1
X_374_ addr0_reg\[4\] net36 _219_ _024_ _196_ vssd1 vssd1 vccd1 vccd1 _090_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_18_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_288_ _184_ net41 net38 _187_ vssd1 vssd1 vccd1 vccd1 _229_ sky130_fd_sc_hd__a22o_1
X_426_ _048_ _135_ _136_ vssd1 vssd1 vccd1 vccd1 _137_ sky130_fd_sc_hd__or3_1
X_357_ _184_ net30 net28 _187_ vssd1 vssd1 vccd1 vccd1 _073_ sky130_fd_sc_hd__a22o_1
Xinput4 addr0[3] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_409_ _025_ _033_ _048_ _054_ vssd1 vssd1 vccd1 vccd1 _122_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_390_ _193_ _196_ _224_ _100_ vssd1 vssd1 vccd1 vccd1 _105_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout37 _205_ vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_2
Xfanout48 addr0_reg\[3\] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_2
X_373_ _198_ _079_ vssd1 vssd1 vccd1 vccd1 _089_ sky130_fd_sc_hd__or2_1
X_442_ _193_ _022_ _034_ _150_ vssd1 vssd1 vccd1 vccd1 _151_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_287_ _194_ net41 net38 _195_ vssd1 vssd1 vccd1 vccd1 _228_ sky130_fd_sc_hd__a22o_1
X_425_ _231_ _023_ vssd1 vssd1 vccd1 vccd1 _136_ sky130_fd_sc_hd__or2_1
Xinput5 addr0[4] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_356_ _070_ _071_ vssd1 vssd1 vccd1 vccd1 _072_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_408_ _188_ _198_ _017_ _100_ vssd1 vssd1 vccd1 vccd1 _121_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_339_ _050_ _051_ _053_ _054_ vssd1 vssd1 vccd1 vccd1 _055_ sky130_fd_sc_hd__or4_2
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_18_Left_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout38 _205_ vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_2
Xfanout27 _058_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_2
Xfanout49 addr0_reg\[3\] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_1
X_441_ _231_ _234_ _054_ _079_ vssd1 vssd1 vccd1 vccd1 _150_ sky130_fd_sc_hd__or4_1
X_372_ _032_ _037_ _043_ _055_ vssd1 vssd1 vccd1 vccd1 _088_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_424_ _034_ _095_ _134_ vssd1 vssd1 vccd1 vccd1 _135_ sky130_fd_sc_hd__or3_1
X_355_ net29 net27 _192_ vssd1 vssd1 vccd1 vccd1 _071_ sky130_fd_sc_hd__o21ba_1
X_286_ _213_ _218_ _221_ _226_ vssd1 vssd1 vccd1 vccd1 _227_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput6 addr0[5] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_407_ _218_ _081_ _119_ vssd1 vssd1 vccd1 vccd1 _120_ sky130_fd_sc_hd__or3_1
X_338_ _189_ net33 net31 _190_ vssd1 vssd1 vccd1 vccd1 _054_ sky130_fd_sc_hd__a22o_1
X_269_ _193_ _197_ _202_ _209_ vssd1 vssd1 vccd1 vccd1 _210_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_6_Left_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap35 _223_ vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_16_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_82 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_440_ _229_ _051_ vssd1 vssd1 vccd1 vccd1 _149_ sky130_fd_sc_hd__or2_1
Xfanout28 _058_ vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_371_ _224_ _070_ _086_ vssd1 vssd1 vccd1 vccd1 _087_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_423_ _036_ _037_ _069_ _078_ vssd1 vssd1 vccd1 vccd1 _134_ sky130_fd_sc_hd__or4_1
X_354_ _190_ net29 net27 _189_ vssd1 vssd1 vccd1 vccd1 _070_ sky130_fd_sc_hd__a22o_1
X_285_ _224_ _225_ vssd1 vssd1 vccd1 vccd1 _226_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput7 addr0[6] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_406_ _066_ _072_ vssd1 vssd1 vccd1 vccd1 _119_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_22_Left_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_337_ _184_ net33 net31 _187_ vssd1 vssd1 vccd1 vccd1 _053_ sky130_fd_sc_hd__a22o_1
X_268_ net40 _208_ _207_ vssd1 vssd1 vccd1 vccd1 _209_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap36 _208_ vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_16_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_83 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_73 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout29 _057_ vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_2
XFILLER_0_25_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_370_ _214_ _062_ vssd1 vssd1 vccd1 vccd1 _086_ sky130_fd_sc_hd__nand2_1
X_499_ clknet_1_1__leaf_clk0 _010_ vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__dfxtp_1
X_422_ net57 net73 net25 _133_ vssd1 vssd1 vccd1 vccd1 _004_ sky130_fd_sc_hd__a22o_1
X_353_ _206_ net29 net27 _204_ vssd1 vssd1 vccd1 vccd1 _069_ sky130_fd_sc_hd__a22o_1
X_284_ net39 net37 _206_ net40 vssd1 vssd1 vccd1 vccd1 _225_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput8 cs0 vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_1
XFILLER_0_9_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_336_ _050_ _051_ vssd1 vssd1 vccd1 vccd1 _052_ sky130_fd_sc_hd__or2_1
X_405_ net57 net62 net25 _118_ vssd1 vssd1 vccd1 vccd1 _002_ sky130_fd_sc_hd__a22o_1
X_267_ net50 net48 net52 net54 vssd1 vssd1 vccd1 vccd1 _208_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_19_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_319_ _030_ _031_ _032_ _033_ vssd1 vssd1 vccd1 vccd1 _035_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_7_84 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_74 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_498_ clknet_1_0__leaf_clk0 _009_ vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__dfxtp_1
X_421_ _096_ _125_ _126_ _132_ vssd1 vssd1 vccd1 vccd1 _133_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_64 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_352_ _066_ _067_ vssd1 vssd1 vccd1 vccd1 _068_ sky130_fd_sc_hd__or2_1
X_283_ net40 _222_ _223_ net37 vssd1 vssd1 vccd1 vccd1 _224_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_335_ _194_ net34 net32 _195_ vssd1 vssd1 vccd1 vccd1 _051_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_404_ _111_ _112_ _114_ _117_ vssd1 vssd1 vccd1 vccd1 _118_ sky130_fd_sc_hd__or4_1
X_266_ net40 net39 net37 _206_ vssd1 vssd1 vccd1 vccd1 _207_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_318_ _032_ _033_ vssd1 vssd1 vccd1 vccd1 _034_ sky130_fd_sc_hd__or2_1
X_249_ net49 net53 net55 net51 vssd1 vssd1 vccd1 vccd1 _190_ sky130_fd_sc_hd__and4b_2
XTAP_TAPCELL_ROW_22_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1 net14 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_75 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_497_ clknet_1_1__leaf_clk0 _008_ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_420_ _017_ _064_ _130_ _131_ vssd1 vssd1 vccd1 vccd1 _132_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_1_65 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_282_ net50 net48 net54 net52 vssd1 vssd1 vccd1 vccd1 _223_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_351_ _195_ net29 net27 _194_ vssd1 vssd1 vccd1 vccd1 _067_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_334_ _200_ net34 net32 net42 vssd1 vssd1 vccd1 vccd1 _050_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_403_ _188_ _016_ _115_ _116_ vssd1 vssd1 vccd1 vccd1 _117_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_265_ net50 net48 net52 net54 vssd1 vssd1 vccd1 vccd1 _206_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_25_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap39 _204_ vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Left_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_317_ net39 net33 net31 _206_ vssd1 vssd1 vccd1 vccd1 _033_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_10_Left_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_248_ net51 net53 net55 net49 vssd1 vssd1 vccd1 vccd1 _189_ sky130_fd_sc_hd__and4bb_2
XTAP_TAPCELL_ROW_22_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold2 net15 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_13_Left_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_496_ clknet_1_0__leaf_clk0 _007_ vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_350_ _187_ net30 net28 _184_ vssd1 vssd1 vccd1 vccd1 _066_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_66 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_281_ net54 net52 net48 net50 vssd1 vssd1 vccd1 vccd1 _222_ sky130_fd_sc_hd__and4b_2
X_479_ net56 net71 net25 _181_ vssd1 vssd1 vccd1 vccd1 _013_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_28_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_402_ net38 _222_ net35 net41 _212_ vssd1 vssd1 vccd1 vccd1 _116_ sky130_fd_sc_hd__a221o_1
X_264_ addr0_reg\[5\] addr0_reg\[6\] net47 vssd1 vssd1 vccd1 vccd1 _205_ sky130_fd_sc_hd__and3b_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_333_ _043_ _044_ _045_ _046_ vssd1 vssd1 vccd1 vccd1 _049_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_25_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_247_ net45 _184_ net43 _187_ vssd1 vssd1 vccd1 vccd1 _188_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_1_Left_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_316_ _223_ net33 net31 _222_ vssd1 vssd1 vccd1 vccd1 _032_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3 net10 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_495_ clknet_1_1__leaf_clk0 _006_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_280_ _219_ _220_ vssd1 vssd1 vccd1 vccd1 _221_ sky130_fd_sc_hd__or2_1
X_478_ _056_ _065_ _180_ vssd1 vssd1 vccd1 vccd1 _181_ sky130_fd_sc_hd__nand3_1
XFILLER_0_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_401_ _024_ _059_ vssd1 vssd1 vccd1 vccd1 _115_ sky130_fd_sc_hd__or2_1
X_263_ net50 net48 net52 net54 vssd1 vssd1 vccd1 vccd1 _204_ sky130_fd_sc_hd__nor4b_2
X_332_ _043_ _044_ _046_ vssd1 vssd1 vccd1 vccd1 _048_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_25_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_315_ _216_ net33 net31 _215_ vssd1 vssd1 vccd1 vccd1 _031_ sky130_fd_sc_hd__a22o_1
X_246_ net49 net55 net53 net51 vssd1 vssd1 vccd1 vccd1 _187_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4 net18 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_494_ clknet_1_1__leaf_clk0 _005_ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_477_ _213_ _020_ _179_ vssd1 vssd1 vccd1 vccd1 _180_ sky130_fd_sc_hd__nor3_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_262_ net47 addr0_reg\[5\] addr0_reg\[6\] vssd1 vssd1 vccd1 vccd1 _203_ sky130_fd_sc_hd__and3b_1
X_331_ _045_ _046_ vssd1 vssd1 vccd1 vccd1 _047_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_400_ _031_ _033_ _072_ _113_ vssd1 vssd1 vccd1 vccd1 _114_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_245_ net47 addr0_reg\[5\] addr0_reg\[6\] vssd1 vssd1 vccd1 vccd1 _186_ sky130_fd_sc_hd__nor3b_1
X_314_ _199_ net33 net31 _200_ vssd1 vssd1 vccd1 vccd1 _030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5 net17 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_493_ clknet_1_1__leaf_clk0 _004_ vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Left_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_476_ _193_ _197_ _067_ vssd1 vssd1 vccd1 vccd1 _179_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_261_ _198_ _201_ vssd1 vssd1 vccd1 vccd1 _202_ sky130_fd_sc_hd__or2_1
X_330_ _206_ net33 net31 _204_ vssd1 vssd1 vccd1 vccd1 _046_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_459_ net56 net69 net25 _165_ vssd1 vssd1 vccd1 vccd1 _009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_313_ addr0_reg\[5\] addr0_reg\[6\] net47 vssd1 vssd1 vccd1 vccd1 _029_ sky130_fd_sc_hd__nor3b_1
X_244_ net47 addr0_reg\[5\] vssd1 vssd1 vccd1 vccd1 _185_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6 net21 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_492_ clknet_1_1__leaf_clk0 _003_ vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_475_ net56 net68 net25 _178_ vssd1 vssd1 vccd1 vccd1 _012_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_28_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_260_ net45 net42 _200_ net43 vssd1 vssd1 vccd1 vccd1 _201_ sky130_fd_sc_hd__a22o_1
X_389_ _098_ _099_ _103_ vssd1 vssd1 vccd1 vccd1 _104_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_458_ _161_ _164_ vssd1 vssd1 vccd1 vccd1 _165_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_312_ net47 addr0_reg\[6\] addr0_reg\[5\] vssd1 vssd1 vccd1 vccd1 _028_ sky130_fd_sc_hd__nor3b_1
X_243_ net51 net55 net53 net49 vssd1 vssd1 vccd1 vccd1 _184_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_23_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Left_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7 net11 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_491_ clknet_1_1__leaf_clk0 _002_ vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0_clk0 clk0 vssd1 vssd1 vccd1 vccd1 clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_474_ _026_ _042_ _177_ vssd1 vssd1 vccd1 vccd1 _178_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_388_ _201_ _211_ vssd1 vssd1 vccd1 vccd1 _103_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_457_ _087_ _108_ _162_ _163_ vssd1 vssd1 vccd1 vccd1 _164_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_16_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_242_ net47 addr0_reg\[5\] addr0_reg\[6\] vssd1 vssd1 vccd1 vccd1 _183_ sky130_fd_sc_hd__and3_1
X_311_ _210_ _227_ _239_ _026_ net8 vssd1 vssd1 vccd1 vccd1 _027_ sky130_fd_sc_hd__o41a_1
XFILLER_0_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold8 net20 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dlygate4sd3_1
X_490_ clknet_1_1__leaf_clk0 _001_ vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_473_ _055_ _119_ _128_ _176_ vssd1 vssd1 vccd1 vccd1 _177_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_387_ _021_ _025_ vssd1 vssd1 vccd1 vccd1 _102_ sky130_fd_sc_hd__or2_1
X_456_ _035_ _044_ _066_ _077_ vssd1 vssd1 vccd1 vccd1 _163_ sky130_fd_sc_hd__or4_1
X_310_ _020_ _023_ _024_ _025_ vssd1 vssd1 vccd1 vccd1 _026_ sky130_fd_sc_hd__or4_1
X_439_ net56 net63 _085_ _148_ vssd1 vssd1 vccd1 vccd1 _006_ sky130_fd_sc_hd__a22o_1
X_241_ net8 vssd1 vssd1 vccd1 vccd1 _182_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold9 net22 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Left_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_472_ _202_ _043_ _044_ _075_ vssd1 vssd1 vccd1 vccd1 _176_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_386_ _068_ _071_ vssd1 vssd1 vccd1 vccd1 _101_ sky130_fd_sc_hd__or2_1
X_455_ _061_ _089_ _102_ _149_ vssd1 vssd1 vccd1 vccd1 _162_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_438_ _114_ _143_ _147_ vssd1 vssd1 vccd1 vccd1 _148_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_369_ _027_ _084_ vssd1 vssd1 vccd1 vccd1 _085_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_21_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Left_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_471_ net57 net64 net25 _175_ vssd1 vssd1 vccd1 vccd1 _011_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_12_Left_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_385_ _031_ _036_ vssd1 vssd1 vccd1 vccd1 _100_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_454_ _191_ _193_ _221_ _160_ vssd1 vssd1 vccd1 vccd1 _161_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_437_ _086_ _116_ _144_ _146_ vssd1 vssd1 vccd1 vccd1 _147_ sky130_fd_sc_hd__or4_1
X_299_ net45 _215_ _216_ net43 vssd1 vssd1 vccd1 vccd1 _240_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_368_ _056_ _065_ _076_ net26 net56 vssd1 vssd1 vccd1 vccd1 _084_ sky130_fd_sc_hd__a41oi_1
XTAP_TAPCELL_ROW_21_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_470_ _042_ _120_ _174_ vssd1 vssd1 vccd1 vccd1 _175_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_384_ _039_ _077_ vssd1 vssd1 vccd1 vccd1 _099_ sky130_fd_sc_hd__or2_1
X_453_ _233_ _037_ _038_ _046_ vssd1 vssd1 vccd1 vccd1 _160_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_24_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_436_ _039_ _051_ _080_ _145_ vssd1 vssd1 vccd1 vccd1 _146_ sky130_fd_sc_hd__or4_1
X_298_ _230_ _232_ _235_ _238_ vssd1 vssd1 vccd1 vccd1 _239_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_367_ _185_ net36 _068_ _069_ _082_ vssd1 vssd1 vccd1 vccd1 _083_ sky130_fd_sc_hd__a2111oi_1
X_419_ _207_ _212_ _217_ _032_ vssd1 vssd1 vccd1 vccd1 _131_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_452_ net57 net67 _085_ _159_ vssd1 vssd1 vccd1 vccd1 _008_ sky130_fd_sc_hd__a22o_1
X_383_ _050_ _054_ vssd1 vssd1 vccd1 vccd1 _098_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_366_ _077_ _078_ _079_ _080_ vssd1 vssd1 vccd1 vccd1 _082_ sky130_fd_sc_hd__or4_2
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_435_ _201_ _219_ _234_ _016_ vssd1 vssd1 vccd1 vccd1 _145_ sky130_fd_sc_hd__or4_1
X_297_ _236_ _237_ vssd1 vssd1 vccd1 vccd1 _238_ sky130_fd_sc_hd__or2_1
X_504_ clknet_1_0__leaf_clk0 _015_ vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__dfxtp_1
Xwire26 _083_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_418_ _040_ _127_ _128_ _129_ vssd1 vssd1 vccd1 vccd1 _130_ sky130_fd_sc_hd__or4_1
X_349_ _061_ _064_ vssd1 vssd1 vccd1 vccd1 _065_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_8_85 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Left_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_451_ _137_ _155_ _156_ _158_ vssd1 vssd1 vccd1 vccd1 _159_ sky130_fd_sc_hd__or4_1
X_382_ _230_ _232_ _094_ _096_ vssd1 vssd1 vccd1 vccd1 _097_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_365_ _079_ _080_ vssd1 vssd1 vccd1 vccd1 _081_ sky130_fd_sc_hd__or2_1
X_434_ _053_ _054_ _077_ _078_ vssd1 vssd1 vccd1 vccd1 _144_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_296_ net37 _215_ _216_ net41 vssd1 vssd1 vccd1 vccd1 _237_ sky130_fd_sc_hd__a22o_1
X_503_ clknet_1_0__leaf_clk0 _014_ vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_417_ _237_ _025_ vssd1 vssd1 vccd1 vccd1 _129_ sky130_fd_sc_hd__or2_1
X_348_ _062_ _063_ vssd1 vssd1 vccd1 vccd1 _064_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_8_86 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_279_ _190_ net40 net37 _189_ vssd1 vssd1 vccd1 vccd1 _220_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Left_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_76 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_381_ _234_ _019_ _095_ vssd1 vssd1 vccd1 vccd1 _096_ sky130_fd_sc_hd__or3_1
X_450_ _230_ _018_ _019_ _157_ vssd1 vssd1 vccd1 vccd1 _158_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_433_ _197_ _049_ _136_ vssd1 vssd1 vccd1 vccd1 _143_ sky130_fd_sc_hd__or3_1
X_502_ clknet_1_0__leaf_clk0 _013_ vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_364_ _200_ net30 net28 net42 vssd1 vssd1 vccd1 vccd1 _080_ sky130_fd_sc_hd__a22o_1
Xclkbuf_1_1__f_clk0 clknet_0_clk0 vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
X_295_ net42 net41 net38 _200_ vssd1 vssd1 vccd1 vccd1 _236_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_278_ _187_ net41 net38 _184_ vssd1 vssd1 vccd1 vccd1 _219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_347_ _223_ net29 net27 _222_ vssd1 vssd1 vccd1 vccd1 _063_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_8_87 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_416_ _196_ _225_ vssd1 vssd1 vccd1 vccd1 _128_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_77 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_380_ _220_ _236_ vssd1 vssd1 vccd1 vccd1 _095_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_2_67 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
.ends

