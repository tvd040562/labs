module cust_rom0 (clk0,
    cs0,
    addr0,
    dout0);
 input clk0;
 input cs0;
 input [7:0] addr0;
 output [31:0] dout0;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire \addr0_reg[0] ;
 wire \addr0_reg[1] ;
 wire \addr0_reg[2] ;
 wire \addr0_reg[3] ;
 wire \addr0_reg[4] ;
 wire \addr0_reg[5] ;
 wire \addr0_reg[6] ;
 wire \addr0_reg[7] ;
 wire cs0_reg;
 wire clknet_0_clk0;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire clknet_2_0__leaf_clk0;
 wire clknet_2_1__leaf_clk0;
 wire clknet_2_2__leaf_clk0;
 wire clknet_2_3__leaf_clk0;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;

 sky130_fd_sc_hd__inv_2 _0716_ (.A(cs0_reg),
    .Y(_0629_));
 sky130_fd_sc_hd__and4bb_1 _0717_ (.A_N(net592),
    .B_N(net577),
    .C(net585),
    .D(net601),
    .X(_0639_));
 sky130_fd_sc_hd__and4bb_1 _0718_ (.A_N(net614),
    .B_N(net620),
    .C(net626),
    .D(net607),
    .X(_0649_));
 sky130_fd_sc_hd__and4bb_1 _0719_ (.A_N(net600),
    .B_N(net585),
    .C(net578),
    .D(net592),
    .X(_0660_));
 sky130_fd_sc_hd__and4b_1 _0720_ (.A_N(net606),
    .B(net612),
    .C(net624),
    .D(net618),
    .X(_0670_));
 sky130_fd_sc_hd__a22o_1 _0721_ (.A1(net555),
    .A2(net548),
    .B1(net542),
    .B2(net535),
    .X(_0680_));
 sky130_fd_sc_hd__and4bb_1 _0722_ (.A_N(net614),
    .B_N(net627),
    .C(net619),
    .D(net607),
    .X(_0690_));
 sky130_fd_sc_hd__and4bb_1 _0723_ (.A_N(net608),
    .B_N(net626),
    .C(net619),
    .D(net614),
    .X(_0695_));
 sky130_fd_sc_hd__a22o_1 _0724_ (.A1(net554),
    .A2(net531),
    .B1(net521),
    .B2(net542),
    .X(_0696_));
 sky130_fd_sc_hd__or2_1 _0725_ (.A(net336),
    .B(net334),
    .X(_0697_));
 sky130_fd_sc_hd__or4_1 _0726_ (.A(net609),
    .B(net612),
    .C(net623),
    .D(net617),
    .X(_0698_));
 sky130_fd_sc_hd__and4bb_1 _0727_ (.A_N(net602),
    .B_N(net577),
    .C(net587),
    .D(net594),
    .X(_0699_));
 sky130_fd_sc_hd__o21ba_1 _0728_ (.A1(net540),
    .A2(net508),
    .B1_N(net515),
    .X(_0700_));
 sky130_fd_sc_hd__and4b_1 _0729_ (.A_N(net617),
    .B(net623),
    .C(net611),
    .D(net605),
    .X(_0701_));
 sky130_fd_sc_hd__and4bb_1 _0730_ (.A_N(net605),
    .B_N(net611),
    .C(net624),
    .D(net621),
    .X(_0702_));
 sky130_fd_sc_hd__a22o_1 _0731_ (.A1(net557),
    .A2(net503),
    .B1(net495),
    .B2(net544),
    .X(_0703_));
 sky130_fd_sc_hd__or2_1 _0732_ (.A(net332),
    .B(net329),
    .X(_0704_));
 sky130_fd_sc_hd__and4_1 _0733_ (.A(net605),
    .B(net611),
    .C(net623),
    .D(net617),
    .X(_0705_));
 sky130_fd_sc_hd__nor4b_1 _0734_ (.A(net605),
    .B(net611),
    .C(net617),
    .D_N(net623),
    .Y(_0706_));
 sky130_fd_sc_hd__a22o_1 _0735_ (.A1(net557),
    .A2(net486),
    .B1(net478),
    .B2(net544),
    .X(_0707_));
 sky130_fd_sc_hd__or3_2 _0736_ (.A(net333),
    .B(net330),
    .C(net327),
    .X(_0708_));
 sky130_fd_sc_hd__and4b_1 _0737_ (.A_N(net625),
    .B(net618),
    .C(net606),
    .D(net612),
    .X(_0709_));
 sky130_fd_sc_hd__nor4b_1 _0738_ (.A(net606),
    .B(net613),
    .C(net624),
    .D_N(net618),
    .Y(_0710_));
 sky130_fd_sc_hd__a22o_1 _0739_ (.A1(net553),
    .A2(net470),
    .B1(net460),
    .B2(net540),
    .X(_0711_));
 sky130_fd_sc_hd__and4b_1 _0740_ (.A_N(net615),
    .B(net628),
    .C(net621),
    .D(net609),
    .X(_0712_));
 sky130_fd_sc_hd__and4bb_1 _0741_ (.A_N(net607),
    .B_N(net619),
    .C(net626),
    .D(net615),
    .X(_0713_));
 sky130_fd_sc_hd__a22o_1 _0742_ (.A1(net553),
    .A2(net453),
    .B1(net445),
    .B2(net540),
    .X(_0714_));
 sky130_fd_sc_hd__and4bb_1 _0743_ (.A_N(net626),
    .B_N(net619),
    .C(net608),
    .D(net615),
    .X(_0715_));
 sky130_fd_sc_hd__nor4b_1 _0744_ (.A(net607),
    .B(net627),
    .C(net620),
    .D_N(net614),
    .Y(_0031_));
 sky130_fd_sc_hd__a22o_1 _0745_ (.A1(net554),
    .A2(net436),
    .B1(net429),
    .B2(net541),
    .X(_0032_));
 sky130_fd_sc_hd__or2_1 _0746_ (.A(_0714_),
    .B(net323),
    .X(_0033_));
 sky130_fd_sc_hd__or3_1 _0747_ (.A(net330),
    .B(net328),
    .C(net325),
    .X(_0034_));
 sky130_fd_sc_hd__or4_1 _0748_ (.A(net333),
    .B(net329),
    .C(net327),
    .D(net324),
    .X(_0035_));
 sky130_fd_sc_hd__or2_1 _0749_ (.A(net68),
    .B(_0035_),
    .X(_0036_));
 sky130_fd_sc_hd__or3_1 _0750_ (.A(net335),
    .B(net334),
    .C(net323),
    .X(_0037_));
 sky130_fd_sc_hd__or4_2 _0751_ (.A(net335),
    .B(net334),
    .C(_0714_),
    .D(_0032_),
    .X(_0038_));
 sky130_fd_sc_hd__nor4b_1 _0752_ (.A(net594),
    .B(net602),
    .C(net577),
    .D_N(net587),
    .Y(_0039_));
 sky130_fd_sc_hd__and4b_1 _0753_ (.A_N(net585),
    .B(net577),
    .C(net600),
    .D(net592),
    .X(_0040_));
 sky130_fd_sc_hd__a22o_1 _0754_ (.A1(net529),
    .A2(net423),
    .B1(net416),
    .B2(net522),
    .X(_0041_));
 sky130_fd_sc_hd__a22o_1 _0755_ (.A1(net549),
    .A2(net423),
    .B1(net416),
    .B2(net536),
    .X(_0042_));
 sky130_fd_sc_hd__a22o_1 _0756_ (.A1(net437),
    .A2(net423),
    .B1(net416),
    .B2(net430),
    .X(_0043_));
 sky130_fd_sc_hd__or2_1 _0757_ (.A(net318),
    .B(net316),
    .X(_0044_));
 sky130_fd_sc_hd__a22o_1 _0758_ (.A1(net452),
    .A2(net421),
    .B1(net414),
    .B2(net443),
    .X(_0045_));
 sky130_fd_sc_hd__or2_1 _0759_ (.A(net318),
    .B(net315),
    .X(_0046_));
 sky130_fd_sc_hd__or3_1 _0760_ (.A(net318),
    .B(net317),
    .C(net313),
    .X(_0047_));
 sky130_fd_sc_hd__or2_1 _0761_ (.A(net320),
    .B(net313),
    .X(_0048_));
 sky130_fd_sc_hd__or4_1 _0762_ (.A(net320),
    .B(_0042_),
    .C(net316),
    .D(net312),
    .X(_0049_));
 sky130_fd_sc_hd__or4b_1 _0763_ (.A(net613),
    .B(net625),
    .C(net618),
    .D_N(net606),
    .X(_0050_));
 sky130_fd_sc_hd__o21ba_1 _0764_ (.A1(net421),
    .A2(net415),
    .B1_N(net410),
    .X(_0051_));
 sky130_fd_sc_hd__a22o_1 _0765_ (.A1(net523),
    .A2(net422),
    .B1(net414),
    .B2(net530),
    .X(_0052_));
 sky130_fd_sc_hd__a22o_1 _0766_ (.A1(net536),
    .A2(net422),
    .B1(net415),
    .B2(net549),
    .X(_0053_));
 sky130_fd_sc_hd__or2_1 _0767_ (.A(net309),
    .B(net308),
    .X(_0054_));
 sky130_fd_sc_hd__or2_1 _0768_ (.A(net311),
    .B(net308),
    .X(_0055_));
 sky130_fd_sc_hd__or3_1 _0769_ (.A(_0051_),
    .B(net309),
    .C(_0053_),
    .X(_0056_));
 sky130_fd_sc_hd__a22o_1 _0770_ (.A1(net548),
    .A2(net542),
    .B1(net535),
    .B2(net555),
    .X(_0057_));
 sky130_fd_sc_hd__o21ba_1 _0771_ (.A1(net555),
    .A2(net541),
    .B1_N(net410),
    .X(_0058_));
 sky130_fd_sc_hd__or2_1 _0772_ (.A(net307),
    .B(net305),
    .X(_0059_));
 sky130_fd_sc_hd__a22o_1 _0773_ (.A1(net541),
    .A2(net529),
    .B1(net522),
    .B2(net554),
    .X(_0060_));
 sky130_fd_sc_hd__a22o_1 _0774_ (.A1(net543),
    .A2(net451),
    .B1(net443),
    .B2(net556),
    .X(_0061_));
 sky130_fd_sc_hd__or4_2 _0775_ (.A(net307),
    .B(net305),
    .C(net304),
    .D(net300),
    .X(_0062_));
 sky130_fd_sc_hd__a22o_1 _0776_ (.A1(net544),
    .A2(net486),
    .B1(net478),
    .B2(net557),
    .X(_0063_));
 sky130_fd_sc_hd__a22o_1 _0777_ (.A1(net541),
    .A2(net436),
    .B1(net429),
    .B2(net554),
    .X(_0064_));
 sky130_fd_sc_hd__or2_1 _0778_ (.A(net297),
    .B(net296),
    .X(_0065_));
 sky130_fd_sc_hd__a22o_1 _0779_ (.A1(net540),
    .A2(net470),
    .B1(net460),
    .B2(net553),
    .X(_0066_));
 sky130_fd_sc_hd__a22o_1 _0780_ (.A1(net544),
    .A2(net505),
    .B1(net497),
    .B2(net557),
    .X(_0067_));
 sky130_fd_sc_hd__or2_1 _0781_ (.A(net293),
    .B(net292),
    .X(_0068_));
 sky130_fd_sc_hd__or4_1 _0782_ (.A(net297),
    .B(net294),
    .C(net293),
    .D(net291),
    .X(_0069_));
 sky130_fd_sc_hd__a22o_1 _0783_ (.A1(net470),
    .A2(net420),
    .B1(net412),
    .B2(net460),
    .X(_0070_));
 sky130_fd_sc_hd__a22o_1 _0784_ (.A1(net487),
    .A2(net419),
    .B1(net411),
    .B2(net479),
    .X(_0071_));
 sky130_fd_sc_hd__a22o_1 _0785_ (.A1(net504),
    .A2(net419),
    .B1(net411),
    .B2(net496),
    .X(_0072_));
 sky130_fd_sc_hd__o21ba_1 _0786_ (.A1(net553),
    .A2(net412),
    .B1_N(net515),
    .X(_0073_));
 sky130_fd_sc_hd__or2_2 _0787_ (.A(net287),
    .B(net283),
    .X(_0074_));
 sky130_fd_sc_hd__or3_1 _0788_ (.A(net287),
    .B(net285),
    .C(_0073_),
    .X(_0075_));
 sky130_fd_sc_hd__or2_1 _0789_ (.A(net289),
    .B(net282),
    .X(_0076_));
 sky130_fd_sc_hd__or4_1 _0790_ (.A(net290),
    .B(net288),
    .C(net286),
    .D(net281),
    .X(_0077_));
 sky130_fd_sc_hd__and4bb_1 _0791_ (.A_N(net574),
    .B_N(net581),
    .C(net590),
    .D(net598),
    .X(_0078_));
 sky130_fd_sc_hd__and4bb_1 _0792_ (.A_N(net590),
    .B_N(net597),
    .C(net574),
    .D(net581),
    .X(_0079_));
 sky130_fd_sc_hd__a22o_1 _0793_ (.A1(net501),
    .A2(net402),
    .B1(net395),
    .B2(net491),
    .X(_0080_));
 sky130_fd_sc_hd__a22o_1 _0794_ (.A1(net484),
    .A2(net406),
    .B1(net398),
    .B2(net475),
    .X(_0081_));
 sky130_fd_sc_hd__or2_1 _0795_ (.A(net277),
    .B(net275),
    .X(_0082_));
 sky130_fd_sc_hd__nor4b_1 _0796_ (.A(net593),
    .B(net516),
    .C(net600),
    .D_N(net586),
    .Y(_0083_));
 sky130_fd_sc_hd__a22o_1 _0797_ (.A1(net469),
    .A2(net407),
    .B1(net399),
    .B2(net459),
    .X(_0084_));
 sky130_fd_sc_hd__or2_1 _0798_ (.A(net279),
    .B(net273),
    .X(_0085_));
 sky130_fd_sc_hd__or4_2 _0799_ (.A(net278),
    .B(net275),
    .C(net272),
    .D(net269),
    .X(_0086_));
 sky130_fd_sc_hd__a22o_1 _0800_ (.A1(net525),
    .A2(net407),
    .B1(net399),
    .B2(net518),
    .X(_0087_));
 sky130_fd_sc_hd__a22o_1 _0801_ (.A1(net433),
    .A2(net401),
    .B1(net394),
    .B2(net426),
    .X(_0088_));
 sky130_fd_sc_hd__a22o_1 _0802_ (.A1(net449),
    .A2(net401),
    .B1(net394),
    .B2(net441),
    .X(_0089_));
 sky130_fd_sc_hd__or2_1 _0803_ (.A(net263),
    .B(net261),
    .X(_0090_));
 sky130_fd_sc_hd__a22o_1 _0804_ (.A1(net545),
    .A2(net402),
    .B1(net397),
    .B2(net532),
    .X(_0091_));
 sky130_fd_sc_hd__or3_1 _0805_ (.A(net263),
    .B(net261),
    .C(net259),
    .X(_0092_));
 sky130_fd_sc_hd__or4_1 _0806_ (.A(net266),
    .B(net263),
    .C(net262),
    .D(net259),
    .X(_0093_));
 sky130_fd_sc_hd__o21ba_1 _0807_ (.A1(net406),
    .A2(net398),
    .B1_N(net409),
    .X(_0094_));
 sky130_fd_sc_hd__a22o_1 _0808_ (.A1(net440),
    .A2(net401),
    .B1(net394),
    .B2(net448),
    .X(_0095_));
 sky130_fd_sc_hd__a22o_1 _0809_ (.A1(net518),
    .A2(net406),
    .B1(net398),
    .B2(net525),
    .X(_0096_));
 sky130_fd_sc_hd__a22o_1 _0810_ (.A1(net533),
    .A2(net403),
    .B1(net396),
    .B2(net546),
    .X(_0097_));
 sky130_fd_sc_hd__or3_1 _0811_ (.A(net256),
    .B(net254),
    .C(net251),
    .X(_0098_));
 sky130_fd_sc_hd__or2_1 _0812_ (.A(net258),
    .B(net252),
    .X(_0099_));
 sky130_fd_sc_hd__or4_1 _0813_ (.A(net257),
    .B(_0095_),
    .C(net253),
    .D(net251),
    .X(_0100_));
 sky130_fd_sc_hd__a22o_1 _0814_ (.A1(net426),
    .A2(net401),
    .B1(net394),
    .B2(net433),
    .X(_0101_));
 sky130_fd_sc_hd__a22o_1 _0815_ (.A1(net456),
    .A2(net404),
    .B1(net397),
    .B2(net466),
    .X(_0102_));
 sky130_fd_sc_hd__a22o_1 _0816_ (.A1(net475),
    .A2(net406),
    .B1(net398),
    .B2(net483),
    .X(_0103_));
 sky130_fd_sc_hd__a22o_1 _0817_ (.A1(net491),
    .A2(net404),
    .B1(net397),
    .B2(net500),
    .X(_0104_));
 sky130_fd_sc_hd__or2_1 _0818_ (.A(net245),
    .B(net242),
    .X(_0105_));
 sky130_fd_sc_hd__or2_1 _0819_ (.A(net250),
    .B(net245),
    .X(_0106_));
 sky130_fd_sc_hd__or2_1 _0820_ (.A(net247),
    .B(net244),
    .X(_0107_));
 sky130_fd_sc_hd__or4_1 _0821_ (.A(net248),
    .B(net246),
    .C(net245),
    .D(net242),
    .X(_0108_));
 sky130_fd_sc_hd__a22o_1 _0822_ (.A1(net429),
    .A2(net421),
    .B1(net414),
    .B2(net436),
    .X(_0109_));
 sky130_fd_sc_hd__a22o_1 _0823_ (.A1(net478),
    .A2(net419),
    .B1(net411),
    .B2(net486),
    .X(_0110_));
 sky130_fd_sc_hd__a22o_1 _0824_ (.A1(net495),
    .A2(net419),
    .B1(net411),
    .B2(net503),
    .X(_0111_));
 sky130_fd_sc_hd__or2_1 _0825_ (.A(net237),
    .B(net235),
    .X(_0112_));
 sky130_fd_sc_hd__or2_1 _0826_ (.A(net241),
    .B(net236),
    .X(_0113_));
 sky130_fd_sc_hd__a22o_1 _0827_ (.A1(net460),
    .A2(net423),
    .B1(net416),
    .B2(net470),
    .X(_0114_));
 sky130_fd_sc_hd__a22o_1 _0828_ (.A1(net443),
    .A2(net421),
    .B1(net414),
    .B2(net451),
    .X(_0115_));
 sky130_fd_sc_hd__or2_1 _0829_ (.A(net238),
    .B(net233),
    .X(_0116_));
 sky130_fd_sc_hd__or4_2 _0830_ (.A(net240),
    .B(net238),
    .C(net236),
    .D(net234),
    .X(_0117_));
 sky130_fd_sc_hd__nor4b_1 _0831_ (.A(net595),
    .B(net579),
    .C(net588),
    .D_N(net603),
    .Y(_0118_));
 sky130_fd_sc_hd__and4b_1 _0832_ (.A_N(net603),
    .B(net579),
    .C(net588),
    .D(net595),
    .X(_0119_));
 sky130_fd_sc_hd__a22o_1 _0833_ (.A1(net506),
    .A2(net390),
    .B1(net385),
    .B2(net498),
    .X(_0120_));
 sky130_fd_sc_hd__nor4b_1 _0834_ (.A(net597),
    .B(net574),
    .C(net581),
    .D_N(net590),
    .Y(_0121_));
 sky130_fd_sc_hd__o21ba_1 _0835_ (.A1(net387),
    .A2(net380),
    .B1_N(net515),
    .X(_0122_));
 sky130_fd_sc_hd__or2_1 _0836_ (.A(net227),
    .B(net224),
    .X(_0123_));
 sky130_fd_sc_hd__a22o_1 _0837_ (.A1(net551),
    .A2(net392),
    .B1(net386),
    .B2(net538),
    .X(_0124_));
 sky130_fd_sc_hd__a22o_1 _0838_ (.A1(net527),
    .A2(net391),
    .B1(net387),
    .B2(net520),
    .X(_0125_));
 sky130_fd_sc_hd__or2_1 _0839_ (.A(net222),
    .B(_0125_),
    .X(_0126_));
 sky130_fd_sc_hd__or4_1 _0840_ (.A(net228),
    .B(net226),
    .C(net221),
    .D(net220),
    .X(_0127_));
 sky130_fd_sc_hd__a22o_1 _0841_ (.A1(net454),
    .A2(net388),
    .B1(net383),
    .B2(net446),
    .X(_0128_));
 sky130_fd_sc_hd__a22o_1 _0842_ (.A1(net438),
    .A2(net392),
    .B1(net386),
    .B2(net431),
    .X(_0129_));
 sky130_fd_sc_hd__or2_1 _0843_ (.A(_0128_),
    .B(net217),
    .X(_0130_));
 sky130_fd_sc_hd__a22o_1 _0844_ (.A1(net473),
    .A2(net390),
    .B1(net385),
    .B2(net463),
    .X(_0131_));
 sky130_fd_sc_hd__a22o_1 _0845_ (.A1(net483),
    .A2(net388),
    .B1(net383),
    .B2(net475),
    .X(_0132_));
 sky130_fd_sc_hd__or4_1 _0846_ (.A(_0127_),
    .B(_0130_),
    .C(net214),
    .D(net212),
    .X(_0133_));
 sky130_fd_sc_hd__a22o_1 _0847_ (.A1(net431),
    .A2(net389),
    .B1(net384),
    .B2(net438),
    .X(_0134_));
 sky130_fd_sc_hd__a22o_1 _0848_ (.A1(net459),
    .A2(net389),
    .B1(net384),
    .B2(net469),
    .X(_0135_));
 sky130_fd_sc_hd__a22o_1 _0849_ (.A1(net494),
    .A2(net388),
    .B1(net383),
    .B2(net502),
    .X(_0136_));
 sky130_fd_sc_hd__a22o_1 _0850_ (.A1(net476),
    .A2(net388),
    .B1(net383),
    .B2(net483),
    .X(_0137_));
 sky130_fd_sc_hd__or3_1 _0851_ (.A(net207),
    .B(net205),
    .C(net204),
    .X(_0138_));
 sky130_fd_sc_hd__or2_1 _0852_ (.A(net210),
    .B(net204),
    .X(_0139_));
 sky130_fd_sc_hd__or4_2 _0853_ (.A(net209),
    .B(net207),
    .C(net205),
    .D(net204),
    .X(_0140_));
 sky130_fd_sc_hd__and4b_1 _0854_ (.A_N(net579),
    .B(net588),
    .C(net595),
    .D(net603),
    .X(_0141_));
 sky130_fd_sc_hd__nor4b_1 _0855_ (.A(net591),
    .B(net599),
    .C(net584),
    .D_N(net576),
    .Y(_0142_));
 sky130_fd_sc_hd__a22o_1 _0856_ (.A1(net492),
    .A2(net371),
    .B1(net364),
    .B2(net501),
    .X(_0143_));
 sky130_fd_sc_hd__a22o_1 _0857_ (.A1(net476),
    .A2(net375),
    .B1(net367),
    .B2(net484),
    .X(_0144_));
 sky130_fd_sc_hd__or2_1 _0858_ (.A(_0143_),
    .B(net200),
    .X(_0145_));
 sky130_fd_sc_hd__a22o_1 _0859_ (.A1(net458),
    .A2(net373),
    .B1(net366),
    .B2(net468),
    .X(_0146_));
 sky130_fd_sc_hd__a22o_1 _0860_ (.A1(net427),
    .A2(net370),
    .B1(net363),
    .B2(net434),
    .X(_0147_));
 sky130_fd_sc_hd__or2_1 _0861_ (.A(net198),
    .B(net196),
    .X(_0148_));
 sky130_fd_sc_hd__or3_1 _0862_ (.A(net202),
    .B(net199),
    .C(net196),
    .X(_0149_));
 sky130_fd_sc_hd__or4_2 _0863_ (.A(net203),
    .B(net199),
    .C(net198),
    .D(net196),
    .X(_0150_));
 sky130_fd_sc_hd__o21ba_1 _0864_ (.A1(net374),
    .A2(net367),
    .B1_N(net410),
    .X(_0151_));
 sky130_fd_sc_hd__a22o_1 _0865_ (.A1(net533),
    .A2(net369),
    .B1(net362),
    .B2(net546),
    .X(_0152_));
 sky130_fd_sc_hd__or2_1 _0866_ (.A(_0151_),
    .B(net193),
    .X(_0153_));
 sky130_fd_sc_hd__a22o_1 _0867_ (.A1(net441),
    .A2(net369),
    .B1(net362),
    .B2(net449),
    .X(_0154_));
 sky130_fd_sc_hd__a22o_1 _0868_ (.A1(net519),
    .A2(net375),
    .B1(net367),
    .B2(net526),
    .X(_0155_));
 sky130_fd_sc_hd__or2_2 _0869_ (.A(net191),
    .B(_0155_),
    .X(_0156_));
 sky130_fd_sc_hd__or4_2 _0870_ (.A(net195),
    .B(net192),
    .C(net189),
    .D(_0155_),
    .X(_0157_));
 sky130_fd_sc_hd__or2_1 _0871_ (.A(_0150_),
    .B(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__nor4_1 _0872_ (.A(net591),
    .B(net598),
    .C(net575),
    .D(net582),
    .Y(_0159_));
 sky130_fd_sc_hd__and4_1 _0873_ (.A(net591),
    .B(net597),
    .C(net575),
    .D(net582),
    .X(_0160_));
 sky130_fd_sc_hd__a22o_1 _0874_ (.A1(net449),
    .A2(net356),
    .B1(net349),
    .B2(net441),
    .X(_0161_));
 sky130_fd_sc_hd__a22o_1 _0875_ (.A1(net545),
    .A2(net356),
    .B1(net349),
    .B2(net532),
    .X(_0162_));
 sky130_fd_sc_hd__or2_1 _0876_ (.A(net187),
    .B(net185),
    .X(_0163_));
 sky130_fd_sc_hd__a22o_1 _0877_ (.A1(net434),
    .A2(net357),
    .B1(net350),
    .B2(net427),
    .X(_0164_));
 sky130_fd_sc_hd__a22o_1 _0878_ (.A1(net528),
    .A2(net360),
    .B1(net353),
    .B2(net519),
    .X(_0165_));
 sky130_fd_sc_hd__or2_1 _0879_ (.A(net188),
    .B(net184),
    .X(_0166_));
 sky130_fd_sc_hd__or2_1 _0880_ (.A(net186),
    .B(net183),
    .X(_0167_));
 sky130_fd_sc_hd__a22o_1 _0881_ (.A1(net521),
    .A2(net360),
    .B1(net353),
    .B2(net528),
    .X(_0168_));
 sky130_fd_sc_hd__o21ba_1 _0882_ (.A1(net361),
    .A2(net354),
    .B1_N(net409),
    .X(_0169_));
 sky130_fd_sc_hd__or2_1 _0883_ (.A(net181),
    .B(net180),
    .X(_0170_));
 sky130_fd_sc_hd__a22o_1 _0884_ (.A1(net442),
    .A2(net358),
    .B1(net351),
    .B2(net450),
    .X(_0171_));
 sky130_fd_sc_hd__a22o_1 _0885_ (.A1(net533),
    .A2(net357),
    .B1(net350),
    .B2(net546),
    .X(_0172_));
 sky130_fd_sc_hd__or2_1 _0886_ (.A(net179),
    .B(net177),
    .X(_0173_));
 sky130_fd_sc_hd__nor4_1 _0887_ (.A(net65),
    .B(_0167_),
    .C(_0170_),
    .D(_0173_),
    .Y(_0174_));
 sky130_fd_sc_hd__a22o_1 _0888_ (.A1(net547),
    .A2(net369),
    .B1(net362),
    .B2(net534),
    .X(_0175_));
 sky130_fd_sc_hd__a22o_1 _0889_ (.A1(net434),
    .A2(net369),
    .B1(net362),
    .B2(net427),
    .X(_0176_));
 sky130_fd_sc_hd__a22o_1 _0890_ (.A1(net448),
    .A2(net370),
    .B1(net363),
    .B2(net440),
    .X(_0177_));
 sky130_fd_sc_hd__a22o_1 _0891_ (.A1(net528),
    .A2(net374),
    .B1(net367),
    .B2(net521),
    .X(_0178_));
 sky130_fd_sc_hd__or2_1 _0892_ (.A(net172),
    .B(net170),
    .X(_0179_));
 sky130_fd_sc_hd__or2_1 _0893_ (.A(net174),
    .B(net169),
    .X(_0180_));
 sky130_fd_sc_hd__or4_1 _0894_ (.A(net174),
    .B(net173),
    .C(net170),
    .D(net168),
    .X(_0181_));
 sky130_fd_sc_hd__and4b_1 _0895_ (.A_N(net590),
    .B(net597),
    .C(net574),
    .D(net581),
    .X(_0182_));
 sky130_fd_sc_hd__a22o_1 _0896_ (.A1(net448),
    .A2(net377),
    .B1(net344),
    .B2(net440),
    .X(_0183_));
 sky130_fd_sc_hd__a22o_1 _0897_ (.A1(net433),
    .A2(net377),
    .B1(net344),
    .B2(net426),
    .X(_0184_));
 sky130_fd_sc_hd__a22o_1 _0898_ (.A1(net500),
    .A2(net379),
    .B1(net346),
    .B2(net493),
    .X(_0185_));
 sky130_fd_sc_hd__o21ba_1 _0899_ (.A1(net405),
    .A2(net346),
    .B1_N(net517),
    .X(_0186_));
 sky130_fd_sc_hd__or2_1 _0900_ (.A(_0185_),
    .B(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__a22o_1 _0901_ (.A1(net466),
    .A2(net379),
    .B1(net346),
    .B2(net456),
    .X(_0188_));
 sky130_fd_sc_hd__a22o_1 _0902_ (.A1(net485),
    .A2(net380),
    .B1(net347),
    .B2(net477),
    .X(_0189_));
 sky130_fd_sc_hd__or2_1 _0903_ (.A(net160),
    .B(net157),
    .X(_0190_));
 sky130_fd_sc_hd__or4_1 _0904_ (.A(net167),
    .B(net165),
    .C(net63),
    .D(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__a22o_1 _0905_ (.A1(net475),
    .A2(net380),
    .B1(net347),
    .B2(net483),
    .X(_0192_));
 sky130_fd_sc_hd__a22o_1 _0906_ (.A1(net456),
    .A2(net379),
    .B1(net348),
    .B2(net466),
    .X(_0193_));
 sky130_fd_sc_hd__or2_1 _0907_ (.A(_0192_),
    .B(net155),
    .X(_0194_));
 sky130_fd_sc_hd__a22o_1 _0908_ (.A1(net426),
    .A2(net378),
    .B1(net345),
    .B2(net433),
    .X(_0195_));
 sky130_fd_sc_hd__a22o_1 _0909_ (.A1(net491),
    .A2(net378),
    .B1(net345),
    .B2(net500),
    .X(_0196_));
 sky130_fd_sc_hd__or2_1 _0910_ (.A(net153),
    .B(net152),
    .X(_0197_));
 sky130_fd_sc_hd__or2_1 _0911_ (.A(net155),
    .B(net151),
    .X(_0198_));
 sky130_fd_sc_hd__or4_4 _0912_ (.A(_0192_),
    .B(net155),
    .C(net154),
    .D(net151),
    .X(_0199_));
 sky130_fd_sc_hd__a22o_1 _0913_ (.A1(net519),
    .A2(net381),
    .B1(net347),
    .B2(net526),
    .X(_0200_));
 sky130_fd_sc_hd__a22o_1 _0914_ (.A1(net440),
    .A2(net377),
    .B1(net344),
    .B2(net448),
    .X(_0201_));
 sky130_fd_sc_hd__or2_1 _0915_ (.A(net149),
    .B(net148),
    .X(_0202_));
 sky130_fd_sc_hd__a22o_1 _0916_ (.A1(net532),
    .A2(net378),
    .B1(net345),
    .B2(net545),
    .X(_0203_));
 sky130_fd_sc_hd__o21ba_1 _0917_ (.A1(net380),
    .A2(net347),
    .B1_N(net409),
    .X(_0204_));
 sky130_fd_sc_hd__or2_2 _0918_ (.A(net146),
    .B(net144),
    .X(_0205_));
 sky130_fd_sc_hd__or4_2 _0919_ (.A(net149),
    .B(net148),
    .C(net146),
    .D(net144),
    .X(_0206_));
 sky130_fd_sc_hd__nor2_1 _0920_ (.A(_0199_),
    .B(net61),
    .Y(_0207_));
 sky130_fd_sc_hd__a22o_1 _0921_ (.A1(net445),
    .A2(net391),
    .B1(net385),
    .B2(net453),
    .X(_0208_));
 sky130_fd_sc_hd__a22o_1 _0922_ (.A1(net518),
    .A2(net392),
    .B1(net386),
    .B2(net525),
    .X(_0209_));
 sky130_fd_sc_hd__a22o_1 _0923_ (.A1(net538),
    .A2(net390),
    .B1(net385),
    .B2(net551),
    .X(_0210_));
 sky130_fd_sc_hd__o21ba_1 _0924_ (.A1(net389),
    .A2(net384),
    .B1_N(net409),
    .X(_0211_));
 sky130_fd_sc_hd__or3_1 _0925_ (.A(net140),
    .B(net138),
    .C(net135),
    .X(_0212_));
 sky130_fd_sc_hd__or2_1 _0926_ (.A(net142),
    .B(net138),
    .X(_0213_));
 sky130_fd_sc_hd__or3_1 _0927_ (.A(net143),
    .B(net137),
    .C(net136),
    .X(_0214_));
 sky130_fd_sc_hd__or4_2 _0928_ (.A(net142),
    .B(net140),
    .C(net138),
    .D(net135),
    .X(_0215_));
 sky130_fd_sc_hd__and4bb_1 _0929_ (.A_N(net592),
    .B_N(net585),
    .C(net578),
    .D(net600),
    .X(_0216_));
 sky130_fd_sc_hd__a22o_1 _0930_ (.A1(net509),
    .A2(net437),
    .B1(net430),
    .B2(net337),
    .X(_0217_));
 sky130_fd_sc_hd__a22o_1 _0931_ (.A1(net548),
    .A2(net510),
    .B1(net339),
    .B2(net535),
    .X(_0218_));
 sky130_fd_sc_hd__a22o_1 _0932_ (.A1(net508),
    .A2(net486),
    .B1(net478),
    .B2(net338),
    .X(_0219_));
 sky130_fd_sc_hd__a22o_1 _0933_ (.A1(net511),
    .A2(net471),
    .B1(net461),
    .B2(net341),
    .X(_0220_));
 sky130_fd_sc_hd__or2_1 _0934_ (.A(net130),
    .B(net127),
    .X(_0221_));
 sky130_fd_sc_hd__or4_1 _0935_ (.A(net133),
    .B(net132),
    .C(net128),
    .D(net125),
    .X(_0222_));
 sky130_fd_sc_hd__a22o_1 _0936_ (.A1(net529),
    .A2(net510),
    .B1(net339),
    .B2(net522),
    .X(_0223_));
 sky130_fd_sc_hd__a22o_1 _0937_ (.A1(net511),
    .A2(net451),
    .B1(net444),
    .B2(net341),
    .X(_0224_));
 sky130_fd_sc_hd__or2_1 _0938_ (.A(net124),
    .B(net122),
    .X(_0225_));
 sky130_fd_sc_hd__a22o_1 _0939_ (.A1(net509),
    .A2(net503),
    .B1(net495),
    .B2(net337),
    .X(_0226_));
 sky130_fd_sc_hd__o21ba_1 _0940_ (.A1(net374),
    .A2(net338),
    .B1_N(net516),
    .X(_0227_));
 sky130_fd_sc_hd__or2_1 _0941_ (.A(net118),
    .B(net116),
    .X(_0228_));
 sky130_fd_sc_hd__or4_2 _0942_ (.A(_0217_),
    .B(net132),
    .C(net124),
    .D(_0224_),
    .X(_0229_));
 sky130_fd_sc_hd__or2_1 _0943_ (.A(net127),
    .B(net116),
    .X(_0230_));
 sky130_fd_sc_hd__or4_1 _0944_ (.A(net128),
    .B(net125),
    .C(net119),
    .D(net116),
    .X(_0231_));
 sky130_fd_sc_hd__a22o_1 _0945_ (.A1(net511),
    .A2(net461),
    .B1(net341),
    .B2(net471),
    .X(_0232_));
 sky130_fd_sc_hd__a22o_1 _0946_ (.A1(net535),
    .A2(net510),
    .B1(net340),
    .B2(net548),
    .X(_0233_));
 sky130_fd_sc_hd__a22o_1 _0947_ (.A1(net512),
    .A2(net429),
    .B1(net339),
    .B2(net436),
    .X(_0234_));
 sky130_fd_sc_hd__o21ba_1 _0948_ (.A1(net508),
    .A2(net338),
    .B1_N(net410),
    .X(_0235_));
 sky130_fd_sc_hd__or4_1 _0949_ (.A(net114),
    .B(net113),
    .C(net111),
    .D(net108),
    .X(_0236_));
 sky130_fd_sc_hd__a22o_1 _0950_ (.A1(net511),
    .A2(net443),
    .B1(net341),
    .B2(net451),
    .X(_0237_));
 sky130_fd_sc_hd__a22o_1 _0951_ (.A1(net522),
    .A2(net510),
    .B1(net339),
    .B2(net529),
    .X(_0238_));
 sky130_fd_sc_hd__or2_1 _0952_ (.A(_0237_),
    .B(net106),
    .X(_0239_));
 sky130_fd_sc_hd__a22o_1 _0953_ (.A1(net508),
    .A2(net479),
    .B1(net337),
    .B2(net487),
    .X(_0240_));
 sky130_fd_sc_hd__a22o_1 _0954_ (.A1(net509),
    .A2(net495),
    .B1(net337),
    .B2(net503),
    .X(_0241_));
 sky130_fd_sc_hd__or2_1 _0955_ (.A(net103),
    .B(net102),
    .X(_0242_));
 sky130_fd_sc_hd__or4_1 _0956_ (.A(_0237_),
    .B(net106),
    .C(net104),
    .D(net101),
    .X(_0243_));
 sky130_fd_sc_hd__or4_2 _0957_ (.A(_0229_),
    .B(_0231_),
    .C(_0236_),
    .D(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__a22o_1 _0958_ (.A1(net492),
    .A2(net356),
    .B1(net349),
    .B2(net501),
    .X(_0245_));
 sky130_fd_sc_hd__a22o_1 _0959_ (.A1(net427),
    .A2(net356),
    .B1(net349),
    .B2(net434),
    .X(_0246_));
 sky130_fd_sc_hd__or2_1 _0960_ (.A(net100),
    .B(net99),
    .X(_0247_));
 sky130_fd_sc_hd__a22o_1 _0961_ (.A1(net456),
    .A2(net359),
    .B1(net352),
    .B2(net467),
    .X(_0248_));
 sky130_fd_sc_hd__a22o_1 _0962_ (.A1(net476),
    .A2(net360),
    .B1(net353),
    .B2(net484),
    .X(_0249_));
 sky130_fd_sc_hd__or2_1 _0963_ (.A(net97),
    .B(net94),
    .X(_0250_));
 sky130_fd_sc_hd__a22o_1 _0964_ (.A1(net489),
    .A2(net374),
    .B1(net368),
    .B2(net481),
    .X(_0251_));
 sky130_fd_sc_hd__and2b_1 _0965_ (.A_N(net517),
    .B(net366),
    .X(_0252_));
 sky130_fd_sc_hd__or4_1 _0966_ (.A(net96),
    .B(net93),
    .C(net90),
    .D(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__a22o_1 _0967_ (.A1(net466),
    .A2(net372),
    .B1(net365),
    .B2(net457),
    .X(_0254_));
 sky130_fd_sc_hd__a22o_1 _0968_ (.A1(net501),
    .A2(net371),
    .B1(net364),
    .B2(net492),
    .X(_0255_));
 sky130_fd_sc_hd__a22o_1 _0969_ (.A1(net545),
    .A2(net377),
    .B1(net344),
    .B2(net532),
    .X(_0256_));
 sky130_fd_sc_hd__a22o_1 _0970_ (.A1(net525),
    .A2(net381),
    .B1(net348),
    .B2(net518),
    .X(_0257_));
 sky130_fd_sc_hd__or2_1 _0971_ (.A(net83),
    .B(net81),
    .X(_0258_));
 sky130_fd_sc_hd__or4_1 _0972_ (.A(net88),
    .B(net84),
    .C(net82),
    .D(net81),
    .X(_0259_));
 sky130_fd_sc_hd__a22o_1 _0973_ (.A1(net485),
    .A2(net360),
    .B1(net353),
    .B2(net477),
    .X(_0260_));
 sky130_fd_sc_hd__o21ba_1 _0974_ (.A1(net390),
    .A2(net354),
    .B1_N(net515),
    .X(_0261_));
 sky130_fd_sc_hd__or2_1 _0975_ (.A(net79),
    .B(net74),
    .X(_0262_));
 sky130_fd_sc_hd__a22o_1 _0976_ (.A1(net467),
    .A2(net359),
    .B1(net352),
    .B2(net457),
    .X(_0263_));
 sky130_fd_sc_hd__a22o_1 _0977_ (.A1(net500),
    .A2(net359),
    .B1(net352),
    .B2(net491),
    .X(_0264_));
 sky130_fd_sc_hd__or2_1 _0978_ (.A(net72),
    .B(net69),
    .X(_0265_));
 sky130_fd_sc_hd__or2_1 _0979_ (.A(net77),
    .B(net72),
    .X(_0266_));
 sky130_fd_sc_hd__or2_1 _0980_ (.A(net74),
    .B(net71),
    .X(_0267_));
 sky130_fd_sc_hd__or4_2 _0981_ (.A(net76),
    .B(net74),
    .C(net73),
    .D(net70),
    .X(_0268_));
 sky130_fd_sc_hd__or4_1 _0982_ (.A(_0035_),
    .B(_0038_),
    .C(_0062_),
    .D(_0069_),
    .X(_0269_));
 sky130_fd_sc_hd__or2_1 _0983_ (.A(_0077_),
    .B(_0117_),
    .X(_0270_));
 sky130_fd_sc_hd__or2_1 _0984_ (.A(net309),
    .B(net232),
    .X(_0271_));
 sky130_fd_sc_hd__or2_2 _0985_ (.A(net311),
    .B(net229),
    .X(_0272_));
 sky130_fd_sc_hd__or3_1 _0986_ (.A(_0049_),
    .B(_0054_),
    .C(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__or3_1 _0987_ (.A(_0269_),
    .B(_0270_),
    .C(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__or4_1 _0988_ (.A(_0086_),
    .B(_0093_),
    .C(_0100_),
    .D(_0108_),
    .X(_0275_));
 sky130_fd_sc_hd__or4bb_1 _0989_ (.A(_0133_),
    .B(_0158_),
    .C_N(net57),
    .D_N(_0207_),
    .X(_0276_));
 sky130_fd_sc_hd__or4_1 _0990_ (.A(_0140_),
    .B(_0215_),
    .C(_0259_),
    .D(_0268_),
    .X(_0277_));
 sky130_fd_sc_hd__or4_1 _0991_ (.A(net167),
    .B(net163),
    .C(_0247_),
    .D(_0253_),
    .X(_0278_));
 sky130_fd_sc_hd__or3_1 _0992_ (.A(_0181_),
    .B(net63),
    .C(_0190_),
    .X(_0279_));
 sky130_fd_sc_hd__or4_1 _0993_ (.A(_0275_),
    .B(_0277_),
    .C(_0278_),
    .D(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__o41a_1 _0994_ (.A1(_0244_),
    .A2(_0274_),
    .A3(_0276_),
    .A4(_0280_),
    .B1(cs0_reg),
    .X(_0281_));
 sky130_fd_sc_hd__or2_1 _0995_ (.A(net166),
    .B(net83),
    .X(_0282_));
 sky130_fd_sc_hd__or4_1 _0996_ (.A(_0212_),
    .B(_0245_),
    .C(net96),
    .D(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__or2_1 _0997_ (.A(net325),
    .B(net302),
    .X(_0284_));
 sky130_fd_sc_hd__or2_1 _0998_ (.A(net125),
    .B(net118),
    .X(_0285_));
 sky130_fd_sc_hd__or4_1 _0999_ (.A(_0097_),
    .B(net222),
    .C(_0284_),
    .D(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__or4_1 _1000_ (.A(net276),
    .B(net271),
    .C(net162),
    .D(_0186_),
    .X(_0287_));
 sky130_fd_sc_hd__or4_1 _1001_ (.A(net227),
    .B(net225),
    .C(net181),
    .D(net180),
    .X(_0288_));
 sky130_fd_sc_hd__or4_1 _1002_ (.A(net308),
    .B(net232),
    .C(net79),
    .D(net71),
    .X(_0289_));
 sky130_fd_sc_hd__or2_1 _1003_ (.A(net112),
    .B(net105),
    .X(_0290_));
 sky130_fd_sc_hd__or4_1 _1004_ (.A(net199),
    .B(net198),
    .C(net112),
    .D(net105),
    .X(_0291_));
 sky130_fd_sc_hd__or4_1 _1005_ (.A(net214),
    .B(net212),
    .C(net178),
    .D(net176),
    .X(_0292_));
 sky130_fd_sc_hd__or4_1 _1006_ (.A(net188),
    .B(net184),
    .C(net133),
    .D(net123),
    .X(_0293_));
 sky130_fd_sc_hd__or4_1 _1007_ (.A(net192),
    .B(net189),
    .C(net90),
    .D(net88),
    .X(_0294_));
 sky130_fd_sc_hd__or3_1 _1008_ (.A(net174),
    .B(net172),
    .C(net170),
    .X(_0295_));
 sky130_fd_sc_hd__or4_1 _1009_ (.A(net336),
    .B(net307),
    .C(net305),
    .D(net239),
    .X(_0296_));
 sky130_fd_sc_hd__or4_1 _1010_ (.A(net322),
    .B(net289),
    .C(net152),
    .D(net150),
    .X(_0297_));
 sky130_fd_sc_hd__or4_1 _1011_ (.A(_0289_),
    .B(_0293_),
    .C(_0296_),
    .D(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__or4_1 _1012_ (.A(_0138_),
    .B(_0288_),
    .C(_0291_),
    .D(_0292_),
    .X(_0299_));
 sky130_fd_sc_hd__nor2_1 _1013_ (.A(_0287_),
    .B(_0294_),
    .Y(_0300_));
 sky130_fd_sc_hd__or4b_1 _1014_ (.A(_0283_),
    .B(_0298_),
    .C(_0299_),
    .D_N(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__or4_1 _1015_ (.A(_0092_),
    .B(_0286_),
    .C(_0295_),
    .D(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__a22o_1 _1016_ (.A1(net631),
    .A2(net558),
    .B1(net41),
    .B2(_0302_),
    .X(_0000_));
 sky130_fd_sc_hd__or3_2 _1017_ (.A(net100),
    .B(net98),
    .C(net96),
    .X(_0303_));
 sky130_fd_sc_hd__or4_1 _1018_ (.A(net237),
    .B(net236),
    .C(net115),
    .D(net111),
    .X(_0304_));
 sky130_fd_sc_hd__or2_1 _1019_ (.A(net163),
    .B(net82),
    .X(_0305_));
 sky130_fd_sc_hd__or3_2 _1020_ (.A(net166),
    .B(net164),
    .C(net82),
    .X(_0306_));
 sky130_fd_sc_hd__or3_1 _1021_ (.A(net221),
    .B(net218),
    .C(net217),
    .X(_0307_));
 sky130_fd_sc_hd__or3_1 _1022_ (.A(net249),
    .B(net246),
    .C(net245),
    .X(_0308_));
 sky130_fd_sc_hd__or3_1 _1023_ (.A(net76),
    .B(net74),
    .C(net73),
    .X(_0309_));
 sky130_fd_sc_hd__or2_1 _1024_ (.A(net180),
    .B(net178),
    .X(_0310_));
 sky130_fd_sc_hd__or3_1 _1025_ (.A(_0169_),
    .B(net178),
    .C(net176),
    .X(_0311_));
 sky130_fd_sc_hd__or3_2 _1026_ (.A(_0149_),
    .B(net168),
    .C(_0179_),
    .X(_0312_));
 sky130_fd_sc_hd__or3_1 _1027_ (.A(net113),
    .B(net107),
    .C(_0237_),
    .X(_0313_));
 sky130_fd_sc_hd__or3_1 _1028_ (.A(_0055_),
    .B(net231),
    .C(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__or2_2 _1029_ (.A(net305),
    .B(net299),
    .X(_0315_));
 sky130_fd_sc_hd__or2_1 _1030_ (.A(net294),
    .B(net292),
    .X(_0316_));
 sky130_fd_sc_hd__or3_1 _1031_ (.A(net133),
    .B(net132),
    .C(net124),
    .X(_0317_));
 sky130_fd_sc_hd__nor2_1 _1032_ (.A(_0075_),
    .B(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__or4_1 _1033_ (.A(_0075_),
    .B(_0315_),
    .C(_0316_),
    .D(_0317_),
    .X(_0319_));
 sky130_fd_sc_hd__or3_1 _1034_ (.A(_0312_),
    .B(_0314_),
    .C(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__or2_1 _1035_ (.A(_0100_),
    .B(_0215_),
    .X(_0321_));
 sky130_fd_sc_hd__or2_1 _1036_ (.A(net209),
    .B(net205),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _1037_ (.A(_0696_),
    .B(_0084_),
    .X(_0323_));
 sky130_fd_sc_hd__or4_1 _1038_ (.A(net333),
    .B(net324),
    .C(net319),
    .D(net312),
    .X(_0324_));
 sky130_fd_sc_hd__or4_1 _1039_ (.A(net64),
    .B(net129),
    .C(net120),
    .D(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__or4_1 _1040_ (.A(net259),
    .B(net225),
    .C(_0322_),
    .D(_0323_),
    .X(_0326_));
 sky130_fd_sc_hd__or4_1 _1041_ (.A(_0137_),
    .B(net65),
    .C(_0167_),
    .D(_0197_),
    .X(_0327_));
 sky130_fd_sc_hd__or4_1 _1042_ (.A(_0321_),
    .B(_0325_),
    .C(_0326_),
    .D(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__or4_1 _1043_ (.A(net60),
    .B(_0304_),
    .C(_0306_),
    .D(_0308_),
    .X(_0329_));
 sky130_fd_sc_hd__or3_1 _1044_ (.A(_0307_),
    .B(_0309_),
    .C(_0311_),
    .X(_0330_));
 sky130_fd_sc_hd__or4_1 _1045_ (.A(net194),
    .B(_0156_),
    .C(_0329_),
    .D(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__or3_1 _1046_ (.A(_0320_),
    .B(_0328_),
    .C(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__a22o_1 _1047_ (.A1(net570),
    .A2(net639),
    .B1(net53),
    .B2(_0332_),
    .X(_0001_));
 sky130_fd_sc_hd__or2_1 _1048_ (.A(net114),
    .B(net102),
    .X(_0333_));
 sky130_fd_sc_hd__or3_1 _1049_ (.A(net115),
    .B(net104),
    .C(net101),
    .X(_0334_));
 sky130_fd_sc_hd__or2_1 _1050_ (.A(net307),
    .B(net291),
    .X(_0335_));
 sky130_fd_sc_hd__or2_1 _1051_ (.A(net181),
    .B(net179),
    .X(_0336_));
 sky130_fd_sc_hd__or4_1 _1052_ (.A(net297),
    .B(net181),
    .C(_0310_),
    .D(_0335_),
    .X(_0337_));
 sky130_fd_sc_hd__or4_1 _1053_ (.A(net239),
    .B(net235),
    .C(net79),
    .D(net75),
    .X(_0338_));
 sky130_fd_sc_hd__or2_2 _1054_ (.A(net166),
    .B(net80),
    .X(_0339_));
 sky130_fd_sc_hd__or4_1 _1055_ (.A(net201),
    .B(net198),
    .C(net130),
    .D(net121),
    .X(_0340_));
 sky130_fd_sc_hd__or2_1 _1056_ (.A(net260),
    .B(net210),
    .X(_0341_));
 sky130_fd_sc_hd__or2_1 _1057_ (.A(net332),
    .B(net299),
    .X(_0342_));
 sky130_fd_sc_hd__or2_1 _1058_ (.A(net252),
    .B(net183),
    .X(_0343_));
 sky130_fd_sc_hd__or2_1 _1059_ (.A(net220),
    .B(net216),
    .X(_0344_));
 sky130_fd_sc_hd__or4_1 _1060_ (.A(net60),
    .B(_0314_),
    .C(net59),
    .D(_0337_),
    .X(_0345_));
 sky130_fd_sc_hd__or4_1 _1061_ (.A(net261),
    .B(net207),
    .C(net173),
    .D(net90),
    .X(_0346_));
 sky130_fd_sc_hd__or3_1 _1062_ (.A(_0214_),
    .B(_0293_),
    .C(_0338_),
    .X(_0347_));
 sky130_fd_sc_hd__or4_1 _1063_ (.A(_0341_),
    .B(_0342_),
    .C(_0343_),
    .D(net58),
    .X(_0348_));
 sky130_fd_sc_hd__or4_1 _1064_ (.A(net244),
    .B(net62),
    .C(net146),
    .D(_0339_),
    .X(_0349_));
 sky130_fd_sc_hd__or3_1 _1065_ (.A(_0074_),
    .B(_0082_),
    .C(_0340_),
    .X(_0350_));
 sky130_fd_sc_hd__or4_1 _1066_ (.A(net271),
    .B(_0123_),
    .C(net196),
    .D(_0346_),
    .X(_0351_));
 sky130_fd_sc_hd__or4_1 _1067_ (.A(_0348_),
    .B(_0349_),
    .C(_0350_),
    .D(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__or3_1 _1068_ (.A(_0345_),
    .B(_0347_),
    .C(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__a22o_1 _1069_ (.A1(net572),
    .A2(net661),
    .B1(net55),
    .B2(_0353_),
    .X(_0002_));
 sky130_fd_sc_hd__or4_1 _1070_ (.A(net301),
    .B(net299),
    .C(net267),
    .D(net264),
    .X(_0354_));
 sky130_fd_sc_hd__or3_1 _1071_ (.A(net249),
    .B(_0107_),
    .C(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__or4_1 _1072_ (.A(_0680_),
    .B(net68),
    .C(_0046_),
    .D(_0225_),
    .X(_0356_));
 sky130_fd_sc_hd__or3_1 _1073_ (.A(net174),
    .B(net171),
    .C(net168),
    .X(_0357_));
 sky130_fd_sc_hd__or3_1 _1074_ (.A(net162),
    .B(net160),
    .C(net159),
    .X(_0358_));
 sky130_fd_sc_hd__or3_1 _1075_ (.A(net298),
    .B(net294),
    .C(net292),
    .X(_0359_));
 sky130_fd_sc_hd__or4_1 _1076_ (.A(_0708_),
    .B(_0357_),
    .C(_0358_),
    .D(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__or4_1 _1077_ (.A(_0086_),
    .B(_0214_),
    .C(net60),
    .D(_0304_),
    .X(_0361_));
 sky130_fd_sc_hd__or4_1 _1078_ (.A(net209),
    .B(net202),
    .C(net91),
    .D(net69),
    .X(_0362_));
 sky130_fd_sc_hd__or4_2 _1079_ (.A(net227),
    .B(net197),
    .C(_0197_),
    .D(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__or4_1 _1080_ (.A(_0057_),
    .B(net257),
    .C(net61),
    .D(net106),
    .X(_0364_));
 sky130_fd_sc_hd__or4_1 _1081_ (.A(_0360_),
    .B(_0361_),
    .C(_0363_),
    .D(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__or4_1 _1082_ (.A(_0054_),
    .B(_0153_),
    .C(_0262_),
    .D(_0285_),
    .X(_0366_));
 sky130_fd_sc_hd__or4_1 _1083_ (.A(net283),
    .B(net110),
    .C(_0310_),
    .D(_0339_),
    .X(_0367_));
 sky130_fd_sc_hd__or4_1 _1084_ (.A(_0355_),
    .B(_0356_),
    .C(_0366_),
    .D(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__or2_1 _1085_ (.A(_0365_),
    .B(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__a22o_1 _1086_ (.A1(net568),
    .A2(net658),
    .B1(net51),
    .B2(_0369_),
    .X(_0003_));
 sky130_fd_sc_hd__or3_1 _1087_ (.A(net298),
    .B(net293),
    .C(net291),
    .X(_0370_));
 sky130_fd_sc_hd__or3_2 _1088_ (.A(net113),
    .B(_0239_),
    .C(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__or2_1 _1089_ (.A(net332),
    .B(net98),
    .X(_0372_));
 sky130_fd_sc_hd__or2_1 _1090_ (.A(_0140_),
    .B(net61),
    .X(_0373_));
 sky130_fd_sc_hd__or3_2 _1091_ (.A(net228),
    .B(net214),
    .C(net211),
    .X(_0374_));
 sky130_fd_sc_hd__or4_1 _1092_ (.A(net267),
    .B(_0091_),
    .C(net175),
    .D(net168),
    .X(_0375_));
 sky130_fd_sc_hd__or3_1 _1093_ (.A(net163),
    .B(net82),
    .C(net81),
    .X(_0376_));
 sky130_fd_sc_hd__or3_2 _1094_ (.A(net185),
    .B(net184),
    .C(net182),
    .X(_0377_));
 sky130_fd_sc_hd__or4_1 _1095_ (.A(_0056_),
    .B(_0222_),
    .C(_0376_),
    .D(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__or4_1 _1096_ (.A(_0075_),
    .B(_0308_),
    .C(_0374_),
    .D(_0375_),
    .X(_0379_));
 sky130_fd_sc_hd__or4_1 _1097_ (.A(net255),
    .B(net236),
    .C(net234),
    .D(net139),
    .X(_0380_));
 sky130_fd_sc_hd__or4_1 _1098_ (.A(net319),
    .B(net316),
    .C(net194),
    .D(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__or4_1 _1099_ (.A(_0148_),
    .B(net64),
    .C(_0250_),
    .D(_0267_),
    .X(_0382_));
 sky130_fd_sc_hd__or4_1 _1100_ (.A(_0378_),
    .B(_0379_),
    .C(_0381_),
    .D(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__or4_1 _1101_ (.A(net301),
    .B(net277),
    .C(_0344_),
    .D(_0372_),
    .X(_0384_));
 sky130_fd_sc_hd__or4_1 _1102_ (.A(_0371_),
    .B(_0373_),
    .C(_0383_),
    .D(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__a22o_1 _1103_ (.A1(net571),
    .A2(net638),
    .B1(net54),
    .B2(_0385_),
    .X(_0004_));
 sky130_fd_sc_hd__or3_1 _1104_ (.A(net210),
    .B(net208),
    .C(net206),
    .X(_0386_));
 sky130_fd_sc_hd__or2_1 _1105_ (.A(net224),
    .B(net211),
    .X(_0387_));
 sky130_fd_sc_hd__or3_1 _1106_ (.A(net214),
    .B(_0386_),
    .C(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__or3_1 _1107_ (.A(net66),
    .B(_0152_),
    .C(_0156_),
    .X(_0389_));
 sky130_fd_sc_hd__or2_1 _1108_ (.A(net256),
    .B(net114),
    .X(_0390_));
 sky130_fd_sc_hd__or2_1 _1109_ (.A(net312),
    .B(net306),
    .X(_0391_));
 sky130_fd_sc_hd__or2_1 _1110_ (.A(_0186_),
    .B(net161),
    .X(_0392_));
 sky130_fd_sc_hd__or4_1 _1111_ (.A(_0116_),
    .B(_0390_),
    .C(_0391_),
    .D(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__or4_1 _1112_ (.A(_0093_),
    .B(_0388_),
    .C(_0389_),
    .D(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__or3_1 _1113_ (.A(net128),
    .B(net118),
    .C(net116),
    .X(_0395_));
 sky130_fd_sc_hd__or3_1 _1114_ (.A(net175),
    .B(net92),
    .C(net87),
    .X(_0396_));
 sky130_fd_sc_hd__or4_1 _1115_ (.A(_0034_),
    .B(_0370_),
    .C(_0395_),
    .D(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__or4_1 _1116_ (.A(net164),
    .B(_0192_),
    .C(net134),
    .D(net110),
    .X(_0398_));
 sky130_fd_sc_hd__or4_1 _1117_ (.A(net252),
    .B(net235),
    .C(net185),
    .D(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__or3_1 _1118_ (.A(net336),
    .B(net68),
    .C(_0212_),
    .X(_0400_));
 sky130_fd_sc_hd__or4_1 _1119_ (.A(net287),
    .B(net276),
    .C(net270),
    .D(net216),
    .X(_0401_));
 sky130_fd_sc_hd__or4_1 _1120_ (.A(_0106_),
    .B(net152),
    .C(net145),
    .D(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__or4_1 _1121_ (.A(net65),
    .B(_0170_),
    .C(_0247_),
    .D(_0266_),
    .X(_0403_));
 sky130_fd_sc_hd__or4_2 _1122_ (.A(_0399_),
    .B(_0400_),
    .C(_0402_),
    .D(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__or3_1 _1123_ (.A(_0394_),
    .B(_0397_),
    .C(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__a22o_1 _1124_ (.A1(net572),
    .A2(net656),
    .B1(net55),
    .B2(_0405_),
    .X(_0005_));
 sky130_fd_sc_hd__or3_1 _1125_ (.A(net129),
    .B(net126),
    .C(net119),
    .X(_0406_));
 sky130_fd_sc_hd__or2_1 _1126_ (.A(net59),
    .B(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__or4_1 _1127_ (.A(net276),
    .B(net275),
    .C(net268),
    .D(net265),
    .X(_0408_));
 sky130_fd_sc_hd__or2_1 _1128_ (.A(net271),
    .B(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__or4_1 _1129_ (.A(net227),
    .B(_0201_),
    .C(net147),
    .D(net95),
    .X(_0410_));
 sky130_fd_sc_hd__or2_1 _1130_ (.A(net206),
    .B(net140),
    .X(_0411_));
 sky130_fd_sc_hd__or2_1 _1131_ (.A(net329),
    .B(net291),
    .X(_0412_));
 sky130_fd_sc_hd__or2_1 _1132_ (.A(net133),
    .B(net122),
    .X(_0413_));
 sky130_fd_sc_hd__or4_1 _1133_ (.A(net187),
    .B(net186),
    .C(net76),
    .D(net70),
    .X(_0414_));
 sky130_fd_sc_hd__or4_1 _1134_ (.A(net241),
    .B(net233),
    .C(_0186_),
    .D(net157),
    .X(_0415_));
 sky130_fd_sc_hd__or3_2 _1135_ (.A(net290),
    .B(net286),
    .C(net281),
    .X(_0416_));
 sky130_fd_sc_hd__or3_1 _1136_ (.A(_0414_),
    .B(_0415_),
    .C(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__or4_1 _1137_ (.A(net327),
    .B(net257),
    .C(net179),
    .D(net123),
    .X(_0418_));
 sky130_fd_sc_hd__or4_1 _1138_ (.A(_0181_),
    .B(_0307_),
    .C(_0407_),
    .D(_0417_),
    .X(_0419_));
 sky130_fd_sc_hd__or4_1 _1139_ (.A(_0038_),
    .B(_0062_),
    .C(_0259_),
    .D(_0418_),
    .X(_0420_));
 sky130_fd_sc_hd__or4_1 _1140_ (.A(net256),
    .B(net253),
    .C(net62),
    .D(_0272_),
    .X(_0421_));
 sky130_fd_sc_hd__or4_1 _1141_ (.A(net67),
    .B(_0411_),
    .C(_0412_),
    .D(_0413_),
    .X(_0422_));
 sky130_fd_sc_hd__or4_1 _1142_ (.A(_0290_),
    .B(_0420_),
    .C(_0421_),
    .D(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__or4_1 _1143_ (.A(net248),
    .B(net242),
    .C(_0158_),
    .D(_0410_),
    .X(_0424_));
 sky130_fd_sc_hd__or4_1 _1144_ (.A(_0409_),
    .B(_0419_),
    .C(_0423_),
    .D(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__a22o_1 _1145_ (.A1(net562),
    .A2(net651),
    .B1(net45),
    .B2(_0425_),
    .X(_0006_));
 sky130_fd_sc_hd__or3_1 _1146_ (.A(net295),
    .B(net293),
    .C(_0315_),
    .X(_0426_));
 sky130_fd_sc_hd__or4_1 _1147_ (.A(net311),
    .B(net229),
    .C(net80),
    .D(net76),
    .X(_0427_));
 sky130_fd_sc_hd__or4_1 _1148_ (.A(net271),
    .B(net270),
    .C(net250),
    .D(net247),
    .X(_0428_));
 sky130_fd_sc_hd__or3_1 _1149_ (.A(net322),
    .B(net316),
    .C(net315),
    .X(_0429_));
 sky130_fd_sc_hd__or4_1 _1150_ (.A(net319),
    .B(net317),
    .C(net312),
    .D(net285),
    .X(_0430_));
 sky130_fd_sc_hd__or2_1 _1151_ (.A(net108),
    .B(_0239_),
    .X(_0431_));
 sky130_fd_sc_hd__or2_1 _1152_ (.A(net100),
    .B(net93),
    .X(_0432_));
 sky130_fd_sc_hd__or3_2 _1153_ (.A(net100),
    .B(net98),
    .C(net93),
    .X(_0433_));
 sky130_fd_sc_hd__or4_1 _1154_ (.A(_0427_),
    .B(_0428_),
    .C(_0431_),
    .D(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__or4_1 _1155_ (.A(_0127_),
    .B(_0295_),
    .C(_0317_),
    .D(_0358_),
    .X(_0435_));
 sky130_fd_sc_hd__or4_1 _1156_ (.A(_0112_),
    .B(_0228_),
    .C(_0310_),
    .D(_0343_),
    .X(_0436_));
 sky130_fd_sc_hd__or4_1 _1157_ (.A(_0202_),
    .B(_0242_),
    .C(net88),
    .D(net84),
    .X(_0437_));
 sky130_fd_sc_hd__or4_1 _1158_ (.A(_0322_),
    .B(_0435_),
    .C(_0436_),
    .D(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__or4_1 _1159_ (.A(_0036_),
    .B(_0389_),
    .C(_0426_),
    .D(_0430_),
    .X(_0439_));
 sky130_fd_sc_hd__or3_1 _1160_ (.A(_0434_),
    .B(_0438_),
    .C(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__a22o_1 _1161_ (.A1(net572),
    .A2(net659),
    .B1(net55),
    .B2(_0440_),
    .X(_0007_));
 sky130_fd_sc_hd__or4_1 _1162_ (.A(net173),
    .B(net95),
    .C(net86),
    .D(net69),
    .X(_0441_));
 sky130_fd_sc_hd__or4_1 _1163_ (.A(net195),
    .B(net193),
    .C(net180),
    .D(net178),
    .X(_0442_));
 sky130_fd_sc_hd__or3_1 _1164_ (.A(net332),
    .B(net289),
    .C(net283),
    .X(_0443_));
 sky130_fd_sc_hd__or4_1 _1165_ (.A(net208),
    .B(net206),
    .C(net155),
    .D(net148),
    .X(_0444_));
 sky130_fd_sc_hd__or4_1 _1166_ (.A(_0441_),
    .B(_0442_),
    .C(_0443_),
    .D(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__or3_2 _1167_ (.A(net125),
    .B(net118),
    .C(_0227_),
    .X(_0446_));
 sky130_fd_sc_hd__or3_1 _1168_ (.A(net324),
    .B(_0033_),
    .C(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__or2_1 _1169_ (.A(net298),
    .B(net230),
    .X(_0448_));
 sky130_fd_sc_hd__or2_1 _1170_ (.A(net306),
    .B(net304),
    .X(_0449_));
 sky130_fd_sc_hd__or4_1 _1171_ (.A(_0106_),
    .B(_0390_),
    .C(_0448_),
    .D(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__or4_1 _1172_ (.A(net278),
    .B(net266),
    .C(net261),
    .D(net259),
    .X(_0451_));
 sky130_fd_sc_hd__or4_2 _1173_ (.A(net185),
    .B(net182),
    .C(net146),
    .D(net144),
    .X(_0452_));
 sky130_fd_sc_hd__or3_1 _1174_ (.A(net67),
    .B(_0180_),
    .C(_0451_),
    .X(_0453_));
 sky130_fd_sc_hd__or3_1 _1175_ (.A(_0291_),
    .B(_0306_),
    .C(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__or4_1 _1176_ (.A(_0445_),
    .B(_0447_),
    .C(_0450_),
    .D(_0452_),
    .X(_0455_));
 sky130_fd_sc_hd__or4_1 _1177_ (.A(_0229_),
    .B(_0374_),
    .C(_0454_),
    .D(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__a22o_1 _1178_ (.A1(net570),
    .A2(net657),
    .B1(net53),
    .B2(_0456_),
    .X(_0008_));
 sky130_fd_sc_hd__or2_1 _1179_ (.A(net275),
    .B(_0192_),
    .X(_0457_));
 sky130_fd_sc_hd__or2_1 _1180_ (.A(net149),
    .B(net147),
    .X(_0458_));
 sky130_fd_sc_hd__or3_1 _1181_ (.A(net279),
    .B(net269),
    .C(net263),
    .X(_0459_));
 sky130_fd_sc_hd__or2_1 _1182_ (.A(net157),
    .B(_0392_),
    .X(_0460_));
 sky130_fd_sc_hd__or2_1 _1183_ (.A(net290),
    .B(_0074_),
    .X(_0461_));
 sky130_fd_sc_hd__or4_1 _1184_ (.A(_0265_),
    .B(_0411_),
    .C(_0457_),
    .D(_0458_),
    .X(_0462_));
 sky130_fd_sc_hd__or4_1 _1185_ (.A(_0697_),
    .B(_0099_),
    .C(_0153_),
    .D(_0230_),
    .X(_0463_));
 sky130_fd_sc_hd__or4_1 _1186_ (.A(net191),
    .B(net164),
    .C(net136),
    .D(net94),
    .X(_0464_));
 sky130_fd_sc_hd__or4_1 _1187_ (.A(net224),
    .B(_0130_),
    .C(net183),
    .D(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__or4_1 _1188_ (.A(_0312_),
    .B(_0462_),
    .C(_0463_),
    .D(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__or4_1 _1189_ (.A(_0708_),
    .B(_0108_),
    .C(_0236_),
    .D(_0459_),
    .X(_0467_));
 sky130_fd_sc_hd__or4_1 _1190_ (.A(_0113_),
    .B(_0316_),
    .C(_0460_),
    .D(_0461_),
    .X(_0468_));
 sky130_fd_sc_hd__or3_1 _1191_ (.A(_0466_),
    .B(_0467_),
    .C(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__a22o_1 _1192_ (.A1(net567),
    .A2(net642),
    .B1(net50),
    .B2(_0469_),
    .X(_0009_));
 sky130_fd_sc_hd__or3_1 _1193_ (.A(_0037_),
    .B(_0173_),
    .C(_0392_),
    .X(_0470_));
 sky130_fd_sc_hd__or4_1 _1194_ (.A(_0303_),
    .B(_0334_),
    .C(_0426_),
    .D(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__or3_1 _1195_ (.A(net137),
    .B(net135),
    .C(_0322_),
    .X(_0472_));
 sky130_fd_sc_hd__or4_1 _1196_ (.A(net266),
    .B(net262),
    .C(net248),
    .D(net242),
    .X(_0473_));
 sky130_fd_sc_hd__or4_1 _1197_ (.A(net258),
    .B(net255),
    .C(net113),
    .D(_0237_),
    .X(_0474_));
 sky130_fd_sc_hd__or4_1 _1198_ (.A(_0446_),
    .B(_0472_),
    .C(_0473_),
    .D(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__or2_1 _1199_ (.A(net228),
    .B(net134),
    .X(_0476_));
 sky130_fd_sc_hd__or2_1 _1200_ (.A(net164),
    .B(net80),
    .X(_0477_));
 sky130_fd_sc_hd__or4_1 _1201_ (.A(net269),
    .B(net220),
    .C(net215),
    .D(net94),
    .X(_0478_));
 sky130_fd_sc_hd__or4_1 _1202_ (.A(_0338_),
    .B(_0396_),
    .C(_0416_),
    .D(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__or4_1 _1203_ (.A(net309),
    .B(net150),
    .C(_0476_),
    .D(_0477_),
    .X(_0480_));
 sky130_fd_sc_hd__or4_1 _1204_ (.A(_0704_),
    .B(_0048_),
    .C(_0085_),
    .D(_0205_),
    .X(_0481_));
 sky130_fd_sc_hd__or3_1 _1205_ (.A(_0479_),
    .B(_0480_),
    .C(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__or3_1 _1206_ (.A(_0471_),
    .B(_0475_),
    .C(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__a22o_1 _1207_ (.A1(net570),
    .A2(net654),
    .B1(net53),
    .B2(_0483_),
    .X(_0010_));
 sky130_fd_sc_hd__or2_1 _1208_ (.A(net65),
    .B(_0268_),
    .X(_0484_));
 sky130_fd_sc_hd__or4_1 _1209_ (.A(net62),
    .B(net151),
    .C(_0202_),
    .D(net144),
    .X(_0485_));
 sky130_fd_sc_hd__or2_1 _1210_ (.A(_0337_),
    .B(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__or2_1 _1211_ (.A(_0153_),
    .B(_0155_),
    .X(_0487_));
 sky130_fd_sc_hd__or4_1 _1212_ (.A(net213),
    .B(net171),
    .C(net169),
    .D(net142),
    .X(_0488_));
 sky130_fd_sc_hd__or4_1 _1213_ (.A(net331),
    .B(net326),
    .C(_0076_),
    .D(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__or4_1 _1214_ (.A(net67),
    .B(_0271_),
    .C(_0341_),
    .D(_0476_),
    .X(_0490_));
 sky130_fd_sc_hd__or4_1 _1215_ (.A(net159),
    .B(net117),
    .C(net101),
    .D(_0306_),
    .X(_0491_));
 sky130_fd_sc_hd__or3_1 _1216_ (.A(net66),
    .B(net58),
    .C(_0433_),
    .X(_0492_));
 sky130_fd_sc_hd__or4_1 _1217_ (.A(_0489_),
    .B(_0490_),
    .C(_0491_),
    .D(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__or4_1 _1218_ (.A(net239),
    .B(_0112_),
    .C(_0428_),
    .D(_0487_),
    .X(_0494_));
 sky130_fd_sc_hd__or4_1 _1219_ (.A(_0484_),
    .B(_0486_),
    .C(_0493_),
    .D(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__a22o_1 _1220_ (.A1(net568),
    .A2(net643),
    .B1(net51),
    .B2(_0495_),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _1221_ (.A(net143),
    .B(net140),
    .X(_0496_));
 sky130_fd_sc_hd__or2_1 _1222_ (.A(net102),
    .B(net89),
    .X(_0497_));
 sky130_fd_sc_hd__or2_1 _1223_ (.A(net131),
    .B(_0413_),
    .X(_0498_));
 sky130_fd_sc_hd__or4_1 _1224_ (.A(net202),
    .B(net199),
    .C(net195),
    .D(net190),
    .X(_0499_));
 sky130_fd_sc_hd__or3_1 _1225_ (.A(net156),
    .B(net153),
    .C(_0205_),
    .X(_0500_));
 sky130_fd_sc_hd__or4_1 _1226_ (.A(net287),
    .B(net228),
    .C(net216),
    .D(net95),
    .X(_0501_));
 sky130_fd_sc_hd__or2_1 _1227_ (.A(net187),
    .B(net182),
    .X(_0502_));
 sky130_fd_sc_hd__or4_1 _1228_ (.A(_0098_),
    .B(_0498_),
    .C(_0499_),
    .D(_0500_),
    .X(_0503_));
 sky130_fd_sc_hd__or3_1 _1229_ (.A(_0105_),
    .B(_0497_),
    .C(_0502_),
    .X(_0504_));
 sky130_fd_sc_hd__or3_1 _1230_ (.A(_0371_),
    .B(_0409_),
    .C(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__or4_1 _1231_ (.A(_0267_),
    .B(_0271_),
    .C(_0342_),
    .D(_0496_),
    .X(_0506_));
 sky130_fd_sc_hd__or4_1 _1232_ (.A(_0139_),
    .B(_0282_),
    .C(_0501_),
    .D(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__or3_1 _1233_ (.A(_0037_),
    .B(net67),
    .C(_0180_),
    .X(_0508_));
 sky130_fd_sc_hd__or4_1 _1234_ (.A(_0126_),
    .B(net177),
    .C(_0415_),
    .D(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__or4_1 _1235_ (.A(_0503_),
    .B(_0505_),
    .C(_0507_),
    .D(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__a22o_1 _1236_ (.A1(net558),
    .A2(net648),
    .B1(net41),
    .B2(_0510_),
    .X(_0012_));
 sky130_fd_sc_hd__or3_1 _1237_ (.A(net248),
    .B(_0103_),
    .C(net243),
    .X(_0511_));
 sky130_fd_sc_hd__or4_2 _1238_ (.A(_0100_),
    .B(net99),
    .C(_0311_),
    .D(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__or2_1 _1239_ (.A(net297),
    .B(net241),
    .X(_0513_));
 sky130_fd_sc_hd__or2_1 _1240_ (.A(_0123_),
    .B(net211),
    .X(_0514_));
 sky130_fd_sc_hd__or2_1 _1241_ (.A(net63),
    .B(net161),
    .X(_0515_));
 sky130_fd_sc_hd__or2_1 _1242_ (.A(net142),
    .B(_0322_),
    .X(_0516_));
 sky130_fd_sc_hd__or4_1 _1243_ (.A(_0498_),
    .B(_0514_),
    .C(_0515_),
    .D(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__or4_1 _1244_ (.A(net218),
    .B(net170),
    .C(net103),
    .D(net84),
    .X(_0518_));
 sky130_fd_sc_hd__or4_1 _1245_ (.A(net192),
    .B(net189),
    .C(net114),
    .D(net112),
    .X(_0519_));
 sky130_fd_sc_hd__or4_1 _1246_ (.A(_0086_),
    .B(_0149_),
    .C(_0414_),
    .D(_0518_),
    .X(_0520_));
 sky130_fd_sc_hd__or3_1 _1247_ (.A(_0391_),
    .B(_0458_),
    .C(_0513_),
    .X(_0521_));
 sky130_fd_sc_hd__or3_1 _1248_ (.A(net62),
    .B(_0339_),
    .C(_0519_),
    .X(_0522_));
 sky130_fd_sc_hd__or4_1 _1249_ (.A(_0447_),
    .B(_0512_),
    .C(_0521_),
    .D(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__or3_1 _1250_ (.A(_0517_),
    .B(_0520_),
    .C(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__a22o_1 _1251_ (.A1(net561),
    .A2(net634),
    .B1(net44),
    .B2(_0524_),
    .X(_0013_));
 sky130_fd_sc_hd__or3_1 _1252_ (.A(net172),
    .B(net91),
    .C(net85),
    .X(_0525_));
 sky130_fd_sc_hd__or4_1 _1253_ (.A(_0459_),
    .B(_0474_),
    .C(_0515_),
    .D(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__or4_1 _1254_ (.A(_0076_),
    .B(_0139_),
    .C(net141),
    .D(net137),
    .X(_0527_));
 sky130_fd_sc_hd__or4_1 _1255_ (.A(net220),
    .B(net219),
    .C(net203),
    .D(_0146_),
    .X(_0528_));
 sky130_fd_sc_hd__or3_1 _1256_ (.A(_0106_),
    .B(_0156_),
    .C(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__or4_1 _1257_ (.A(net235),
    .B(net208),
    .C(net166),
    .D(net98),
    .X(_0530_));
 sky130_fd_sc_hd__or4_1 _1258_ (.A(net61),
    .B(_0288_),
    .C(_0429_),
    .D(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__or4_1 _1259_ (.A(_0221_),
    .B(_0527_),
    .C(_0529_),
    .D(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__or4_1 _1260_ (.A(_0163_),
    .B(_0262_),
    .C(_0315_),
    .D(_0413_),
    .X(_0533_));
 sky130_fd_sc_hd__or4_1 _1261_ (.A(_0198_),
    .B(net111),
    .C(_0241_),
    .D(_0448_),
    .X(_0534_));
 sky130_fd_sc_hd__or3_1 _1262_ (.A(_0036_),
    .B(_0533_),
    .C(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__or3_1 _1263_ (.A(_0526_),
    .B(_0532_),
    .C(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__a22o_1 _1264_ (.A1(net570),
    .A2(net641),
    .B1(net53),
    .B2(_0536_),
    .X(_0014_));
 sky130_fd_sc_hd__or4_1 _1265_ (.A(net334),
    .B(net68),
    .C(net203),
    .D(net66),
    .X(_0537_));
 sky130_fd_sc_hd__or4_1 _1266_ (.A(net283),
    .B(net282),
    .C(net92),
    .D(net87),
    .X(_0538_));
 sky130_fd_sc_hd__or4_1 _1267_ (.A(net301),
    .B(net276),
    .C(net159),
    .D(net103),
    .X(_0539_));
 sky130_fd_sc_hd__or4_1 _1268_ (.A(_0388_),
    .B(_0537_),
    .C(_0538_),
    .D(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__or4_1 _1269_ (.A(_0156_),
    .B(_0335_),
    .C(_0339_),
    .D(_0496_),
    .X(_0541_));
 sky130_fd_sc_hd__or4_1 _1270_ (.A(net265),
    .B(net187),
    .C(net162),
    .D(net151),
    .X(_0542_));
 sky130_fd_sc_hd__or4_1 _1271_ (.A(_0130_),
    .B(_0167_),
    .C(_0541_),
    .D(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__or4_1 _1272_ (.A(_0708_),
    .B(_0229_),
    .C(_0289_),
    .D(_0313_),
    .X(_0544_));
 sky130_fd_sc_hd__or4_1 _1273_ (.A(_0047_),
    .B(net240),
    .C(_0112_),
    .D(_0375_),
    .X(_0545_));
 sky130_fd_sc_hd__or4_1 _1274_ (.A(_0406_),
    .B(_0512_),
    .C(_0544_),
    .D(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__or3_1 _1275_ (.A(_0540_),
    .B(_0543_),
    .C(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__a22o_1 _1276_ (.A1(net572),
    .A2(net660),
    .B1(net55),
    .B2(_0547_),
    .X(_0015_));
 sky130_fd_sc_hd__or4_1 _1277_ (.A(net218),
    .B(_0170_),
    .C(net176),
    .D(net58),
    .X(_0548_));
 sky130_fd_sc_hd__or2_1 _1278_ (.A(net335),
    .B(net329),
    .X(_0549_));
 sky130_fd_sc_hd__or4_1 _1279_ (.A(net131),
    .B(net105),
    .C(_0497_),
    .D(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__or4_1 _1280_ (.A(_0044_),
    .B(_0230_),
    .C(_0272_),
    .D(_0387_),
    .X(_0551_));
 sky130_fd_sc_hd__or4_1 _1281_ (.A(_0065_),
    .B(net272),
    .C(net270),
    .D(_0496_),
    .X(_0552_));
 sky130_fd_sc_hd__or4_1 _1282_ (.A(_0145_),
    .B(_0548_),
    .C(_0551_),
    .D(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__or2_1 _1283_ (.A(_0194_),
    .B(net153),
    .X(_0554_));
 sky130_fd_sc_hd__or2_1 _1284_ (.A(net254),
    .B(_0099_),
    .X(_0555_));
 sky130_fd_sc_hd__or3_1 _1285_ (.A(_0113_),
    .B(net167),
    .C(net163),
    .X(_0556_));
 sky130_fd_sc_hd__or3_1 _1286_ (.A(_0554_),
    .B(_0555_),
    .C(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__or4_1 _1287_ (.A(_0357_),
    .B(_0433_),
    .C(_0452_),
    .D(_0473_),
    .X(_0558_));
 sky130_fd_sc_hd__or4_1 _1288_ (.A(_0714_),
    .B(net195),
    .C(net138),
    .D(net72),
    .X(_0559_));
 sky130_fd_sc_hd__or4_1 _1289_ (.A(net289),
    .B(net160),
    .C(net80),
    .D(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__or4_1 _1290_ (.A(_0062_),
    .B(_0138_),
    .C(_0558_),
    .D(_0560_),
    .X(_0561_));
 sky130_fd_sc_hd__or4_1 _1291_ (.A(_0550_),
    .B(_0553_),
    .C(_0557_),
    .D(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__a22o_1 _1292_ (.A1(net559),
    .A2(net653),
    .B1(net42),
    .B2(_0562_),
    .X(_0016_));
 sky130_fd_sc_hd__or4_1 _1293_ (.A(net250),
    .B(net246),
    .C(net90),
    .D(net88),
    .X(_0563_));
 sky130_fd_sc_hd__or3_1 _1294_ (.A(net131),
    .B(net123),
    .C(net122),
    .X(_0564_));
 sky130_fd_sc_hd__or3_1 _1295_ (.A(net303),
    .B(net300),
    .C(_0066_),
    .X(_0565_));
 sky130_fd_sc_hd__or4_1 _1296_ (.A(net63),
    .B(net157),
    .C(_0564_),
    .D(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__or4_1 _1297_ (.A(_0034_),
    .B(_0047_),
    .C(_0236_),
    .D(net60),
    .X(_0567_));
 sky130_fd_sc_hd__or2_1 _1298_ (.A(_0038_),
    .B(_0150_),
    .X(_0568_));
 sky130_fd_sc_hd__or4_1 _1299_ (.A(_0270_),
    .B(_0566_),
    .C(_0567_),
    .D(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__or3_1 _1300_ (.A(_0213_),
    .B(net58),
    .C(_0477_),
    .X(_0570_));
 sky130_fd_sc_hd__or4_1 _1301_ (.A(_0082_),
    .B(net78),
    .C(net69),
    .D(_0563_),
    .X(_0571_));
 sky130_fd_sc_hd__or3_1 _1302_ (.A(net310),
    .B(net211),
    .C(net189),
    .X(_0572_));
 sky130_fd_sc_hd__or4_1 _1303_ (.A(net265),
    .B(net253),
    .C(_0180_),
    .D(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__or4_1 _1304_ (.A(_0485_),
    .B(_0570_),
    .C(_0571_),
    .D(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__or2_1 _1305_ (.A(_0569_),
    .B(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__a22o_1 _1306_ (.A1(net560),
    .A2(net647),
    .B1(net43),
    .B2(_0575_),
    .X(_0017_));
 sky130_fd_sc_hd__or2_1 _1307_ (.A(net59),
    .B(_0359_),
    .X(_0576_));
 sky130_fd_sc_hd__or4_1 _1308_ (.A(net253),
    .B(net251),
    .C(net221),
    .D(net217),
    .X(_0577_));
 sky130_fd_sc_hd__or4_1 _1309_ (.A(net202),
    .B(net66),
    .C(_0525_),
    .D(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__nand2_1 _1310_ (.A(net57),
    .B(_0318_),
    .Y(_0579_));
 sky130_fd_sc_hd__or4_1 _1311_ (.A(_0431_),
    .B(_0451_),
    .C(_0460_),
    .D(_0511_),
    .X(_0580_));
 sky130_fd_sc_hd__or4_1 _1312_ (.A(net310),
    .B(net302),
    .C(net237),
    .D(net143),
    .X(_0581_));
 sky130_fd_sc_hd__or4_1 _1313_ (.A(_0049_),
    .B(_0199_),
    .C(_0395_),
    .D(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__or4_1 _1314_ (.A(net209),
    .B(net207),
    .C(_0305_),
    .D(_0549_),
    .X(_0583_));
 sky130_fd_sc_hd__or4_1 _1315_ (.A(net192),
    .B(_0155_),
    .C(net149),
    .D(net136),
    .X(_0584_));
 sky130_fd_sc_hd__or3_1 _1316_ (.A(_0123_),
    .B(_0262_),
    .C(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__or4_1 _1317_ (.A(_0578_),
    .B(_0582_),
    .C(_0583_),
    .D(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__or4_1 _1318_ (.A(_0576_),
    .B(_0579_),
    .C(_0580_),
    .D(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__a22o_1 _1319_ (.A1(net563),
    .A2(net646),
    .B1(net46),
    .B2(_0587_),
    .X(_0018_));
 sky130_fd_sc_hd__or3_1 _1320_ (.A(_0500_),
    .B(_0516_),
    .C(_0555_),
    .X(_0588_));
 sky130_fd_sc_hd__or2_1 _1321_ (.A(_0150_),
    .B(_0294_),
    .X(_0589_));
 sky130_fd_sc_hd__or4_1 _1322_ (.A(net314),
    .B(net239),
    .C(net128),
    .D(net107),
    .X(_0590_));
 sky130_fd_sc_hd__or4_1 _1323_ (.A(net284),
    .B(net217),
    .C(net215),
    .D(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__or4_1 _1324_ (.A(net278),
    .B(net172),
    .C(net167),
    .D(net123),
    .X(_0592_));
 sky130_fd_sc_hd__or3_1 _1325_ (.A(_0258_),
    .B(_0267_),
    .C(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__or4_1 _1326_ (.A(_0355_),
    .B(_0589_),
    .C(_0591_),
    .D(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__or4_1 _1327_ (.A(_0055_),
    .B(_0116_),
    .C(_0123_),
    .D(_0242_),
    .X(_0595_));
 sky130_fd_sc_hd__or4_1 _1328_ (.A(_0163_),
    .B(_0412_),
    .C(_0432_),
    .D(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__or4_1 _1329_ (.A(_0470_),
    .B(_0588_),
    .C(_0594_),
    .D(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__a22o_1 _1330_ (.A1(net563),
    .A2(net655),
    .B1(net46),
    .B2(_0597_),
    .X(_0019_));
 sky130_fd_sc_hd__or4_1 _1331_ (.A(net328),
    .B(net323),
    .C(net219),
    .D(net176),
    .X(_0598_));
 sky130_fd_sc_hd__or4_1 _1332_ (.A(net162),
    .B(net160),
    .C(_0457_),
    .D(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__or4_1 _1333_ (.A(net311),
    .B(net229),
    .C(net148),
    .D(net147),
    .X(_0600_));
 sky130_fd_sc_hd__or4_1 _1334_ (.A(_0059_),
    .B(net260),
    .C(net224),
    .D(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__or3_1 _1335_ (.A(_0283_),
    .B(_0599_),
    .C(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__or3_1 _1336_ (.A(net91),
    .B(net89),
    .C(net84),
    .X(_0603_));
 sky130_fd_sc_hd__or4_1 _1337_ (.A(_0333_),
    .B(_0502_),
    .C(_0555_),
    .D(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__or4_1 _1338_ (.A(_0108_),
    .B(_0222_),
    .C(_0309_),
    .D(_0416_),
    .X(_0605_));
 sky130_fd_sc_hd__or4_1 _1339_ (.A(net319),
    .B(net318),
    .C(net169),
    .D(net107),
    .X(_0606_));
 sky130_fd_sc_hd__or4_1 _1340_ (.A(net264),
    .B(net233),
    .C(_0168_),
    .D(net154),
    .X(_0607_));
 sky130_fd_sc_hd__or4_1 _1341_ (.A(_0054_),
    .B(_0068_),
    .C(_0126_),
    .D(_0153_),
    .X(_0608_));
 sky130_fd_sc_hd__or4_1 _1342_ (.A(_0605_),
    .B(_0606_),
    .C(_0607_),
    .D(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__or3_1 _1343_ (.A(_0602_),
    .B(_0604_),
    .C(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__a22o_1 _1344_ (.A1(net558),
    .A2(net652),
    .B1(net41),
    .B2(_0610_),
    .X(_0020_));
 sky130_fd_sc_hd__or4_1 _1345_ (.A(_0704_),
    .B(_0105_),
    .C(_0179_),
    .D(_0205_),
    .X(_0611_));
 sky130_fd_sc_hd__or4_1 _1346_ (.A(_0164_),
    .B(net177),
    .C(net127),
    .D(net109),
    .X(_0612_));
 sky130_fd_sc_hd__or3_1 _1347_ (.A(_0190_),
    .B(_0457_),
    .C(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__or4_1 _1348_ (.A(_0198_),
    .B(_0323_),
    .C(_0336_),
    .D(_0449_),
    .X(_0614_));
 sky130_fd_sc_hd__or4_1 _1349_ (.A(_0576_),
    .B(_0611_),
    .C(_0613_),
    .D(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__or4_1 _1350_ (.A(net281),
    .B(net251),
    .C(net225),
    .D(net99),
    .X(_0616_));
 sky130_fd_sc_hd__or4_1 _1351_ (.A(_0092_),
    .B(_0268_),
    .C(_0499_),
    .D(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__or4_1 _1352_ (.A(_0556_),
    .B(_0564_),
    .C(_0603_),
    .D(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__or3_1 _1353_ (.A(_0273_),
    .B(_0615_),
    .C(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__a22o_1 _1354_ (.A1(net560),
    .A2(net644),
    .B1(net43),
    .B2(_0619_),
    .X(_0021_));
 sky130_fd_sc_hd__or3_1 _1355_ (.A(net335),
    .B(net266),
    .C(net218),
    .X(_0620_));
 sky130_fd_sc_hd__or4_1 _1356_ (.A(net221),
    .B(net191),
    .C(net122),
    .D(net72),
    .X(_0621_));
 sky130_fd_sc_hd__or4_1 _1357_ (.A(_0098_),
    .B(_0311_),
    .C(_0620_),
    .D(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__or4_1 _1358_ (.A(_0107_),
    .B(_0213_),
    .C(_0305_),
    .D(_0432_),
    .X(_0623_));
 sky130_fd_sc_hd__or4_1 _1359_ (.A(net205),
    .B(net204),
    .C(net184),
    .D(net182),
    .X(_0624_));
 sky130_fd_sc_hd__or4_1 _1360_ (.A(_0090_),
    .B(net200),
    .C(net197),
    .D(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__or3_1 _1361_ (.A(_0622_),
    .B(_0623_),
    .C(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__or2_1 _1362_ (.A(_0181_),
    .B(_0603_),
    .X(_0627_));
 sky130_fd_sc_hd__or4_1 _1363_ (.A(_0446_),
    .B(_0461_),
    .C(_0514_),
    .D(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__or4_1 _1364_ (.A(net327),
    .B(net323),
    .C(net131),
    .D(net105),
    .X(_0630_));
 sky130_fd_sc_hd__or3_1 _1365_ (.A(net272),
    .B(net75),
    .C(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__or4_1 _1366_ (.A(net158),
    .B(net111),
    .C(net103),
    .D(net101),
    .X(_0632_));
 sky130_fd_sc_hd__or4_1 _1367_ (.A(net156),
    .B(net153),
    .C(_0458_),
    .D(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__or3_1 _1368_ (.A(_0117_),
    .B(_0315_),
    .C(_0316_),
    .X(_0634_));
 sky130_fd_sc_hd__or4_1 _1369_ (.A(_0273_),
    .B(_0631_),
    .C(_0633_),
    .D(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__or3_1 _1370_ (.A(_0626_),
    .B(_0628_),
    .C(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__a22o_1 _1371_ (.A1(net560),
    .A2(net632),
    .B1(net43),
    .B2(_0636_),
    .X(_0022_));
 sky130_fd_sc_hd__or4_1 _1372_ (.A(_0198_),
    .B(_0333_),
    .C(_0336_),
    .D(_0502_),
    .X(_0637_));
 sky130_fd_sc_hd__or3_1 _1373_ (.A(_0356_),
    .B(_0627_),
    .C(_0637_),
    .X(_0638_));
 sky130_fd_sc_hd__or4_1 _1374_ (.A(net64),
    .B(net158),
    .C(_0376_),
    .D(_0487_),
    .X(_0640_));
 sky130_fd_sc_hd__or4_1 _1375_ (.A(net246),
    .B(net213),
    .C(net201),
    .D(net150),
    .X(_0641_));
 sky130_fd_sc_hd__or4_1 _1376_ (.A(net328),
    .B(net256),
    .C(net130),
    .D(net117),
    .X(_0642_));
 sky130_fd_sc_hd__or4_1 _1377_ (.A(net219),
    .B(net216),
    .C(net95),
    .D(net93),
    .X(_0643_));
 sky130_fd_sc_hd__or4_1 _1378_ (.A(_0408_),
    .B(_0641_),
    .C(_0642_),
    .D(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__or4_1 _1379_ (.A(net308),
    .B(net231),
    .C(_0239_),
    .D(_0284_),
    .X(_0645_));
 sky130_fd_sc_hd__or4_1 _1380_ (.A(_0065_),
    .B(_0074_),
    .C(_0099_),
    .D(_0266_),
    .X(_0646_));
 sky130_fd_sc_hd__or4_1 _1381_ (.A(_0112_),
    .B(_0644_),
    .C(_0645_),
    .D(_0646_),
    .X(_0647_));
 sky130_fd_sc_hd__or4_1 _1382_ (.A(_0472_),
    .B(_0638_),
    .C(_0640_),
    .D(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__a22o_1 _1383_ (.A1(net567),
    .A2(net637),
    .B1(net50),
    .B2(_0648_),
    .X(_0023_));
 sky130_fd_sc_hd__or4_1 _1384_ (.A(_0139_),
    .B(net141),
    .C(net137),
    .D(_0513_),
    .X(_0650_));
 sky130_fd_sc_hd__or4_1 _1385_ (.A(net244),
    .B(net147),
    .C(net112),
    .D(net110),
    .X(_0651_));
 sky130_fd_sc_hd__or4_1 _1386_ (.A(net268),
    .B(net260),
    .C(_0372_),
    .D(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__or3_1 _1387_ (.A(_0537_),
    .B(_0650_),
    .C(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__or4_1 _1388_ (.A(_0287_),
    .B(net59),
    .C(_0377_),
    .D(_0427_),
    .X(_0654_));
 sky130_fd_sc_hd__or4_1 _1389_ (.A(net301),
    .B(net299),
    .C(net284),
    .D(net282),
    .X(_0655_));
 sky130_fd_sc_hd__or4_1 _1390_ (.A(_0044_),
    .B(net237),
    .C(net97),
    .D(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__or4_1 _1391_ (.A(_0157_),
    .B(_0292_),
    .C(_0654_),
    .D(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__or4_1 _1392_ (.A(_0554_),
    .B(_0564_),
    .C(_0577_),
    .D(_0627_),
    .X(_0658_));
 sky130_fd_sc_hd__or3_1 _1393_ (.A(_0653_),
    .B(_0657_),
    .C(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__a22o_1 _1394_ (.A1(net560),
    .A2(net650),
    .B1(net43),
    .B2(_0659_),
    .X(_0024_));
 sky130_fd_sc_hd__or4_1 _1395_ (.A(_0113_),
    .B(_0316_),
    .C(_0460_),
    .D(_0565_),
    .X(_0661_));
 sky130_fd_sc_hd__or3_1 _1396_ (.A(_0197_),
    .B(_0310_),
    .C(_0374_),
    .X(_0662_));
 sky130_fd_sc_hd__or2_1 _1397_ (.A(_0386_),
    .B(_0430_),
    .X(_0663_));
 sky130_fd_sc_hd__or4_1 _1398_ (.A(net223),
    .B(net135),
    .C(net134),
    .D(net117),
    .X(_0664_));
 sky130_fd_sc_hd__or4_1 _1399_ (.A(net145),
    .B(net78),
    .C(_0265_),
    .D(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__or4_1 _1400_ (.A(_0708_),
    .B(net324),
    .C(net278),
    .D(net249),
    .X(_0666_));
 sky130_fd_sc_hd__or4_1 _1401_ (.A(_0662_),
    .B(_0663_),
    .C(_0665_),
    .D(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__or4_1 _1402_ (.A(_0150_),
    .B(_0157_),
    .C(_0181_),
    .D(_0603_),
    .X(_0668_));
 sky130_fd_sc_hd__or3_1 _1403_ (.A(_0098_),
    .B(_0167_),
    .C(_0258_),
    .X(_0669_));
 sky130_fd_sc_hd__or4_1 _1404_ (.A(_0090_),
    .B(net233),
    .C(net229),
    .D(_0247_),
    .X(_0671_));
 sky130_fd_sc_hd__or4_1 _1405_ (.A(_0407_),
    .B(_0668_),
    .C(_0669_),
    .D(_0671_),
    .X(_0672_));
 sky130_fd_sc_hd__or3_1 _1406_ (.A(_0661_),
    .B(_0667_),
    .C(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__a22o_1 _1407_ (.A1(net564),
    .A2(net633),
    .B1(net47),
    .B2(_0673_),
    .X(_0025_));
 sky130_fd_sc_hd__or4_1 _1408_ (.A(net303),
    .B(net300),
    .C(_0234_),
    .D(net107),
    .X(_0674_));
 sky130_fd_sc_hd__or4_1 _1409_ (.A(net290),
    .B(net281),
    .C(net273),
    .D(net75),
    .X(_0675_));
 sky130_fd_sc_hd__or4_1 _1410_ (.A(_0229_),
    .B(_0231_),
    .C(_0674_),
    .D(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__or4_1 _1411_ (.A(net294),
    .B(net288),
    .C(_0081_),
    .D(net269),
    .X(_0677_));
 sky130_fd_sc_hd__or4_1 _1412_ (.A(net230),
    .B(_0117_),
    .C(_0548_),
    .D(_0669_),
    .X(_0678_));
 sky130_fd_sc_hd__or3_1 _1413_ (.A(_0371_),
    .B(_0373_),
    .C(_0676_),
    .X(_0679_));
 sky130_fd_sc_hd__or4_1 _1414_ (.A(_0108_),
    .B(_0374_),
    .C(_0668_),
    .D(_0677_),
    .X(_0681_));
 sky130_fd_sc_hd__or3_1 _1415_ (.A(_0678_),
    .B(_0679_),
    .C(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__a22o_1 _1416_ (.A1(net567),
    .A2(net640),
    .B1(net50),
    .B2(_0682_),
    .X(_0026_));
 sky130_fd_sc_hd__or2_1 _1417_ (.A(_0244_),
    .B(_0668_),
    .X(_0683_));
 sky130_fd_sc_hd__or4_1 _1418_ (.A(net230),
    .B(_0117_),
    .C(_0166_),
    .D(_0268_),
    .X(_0684_));
 sky130_fd_sc_hd__or4_1 _1419_ (.A(_0059_),
    .B(net257),
    .C(net226),
    .D(_0140_),
    .X(_0685_));
 sky130_fd_sc_hd__or2_1 _1420_ (.A(_0684_),
    .B(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__or3_1 _1421_ (.A(_0199_),
    .B(_0206_),
    .C(_0258_),
    .X(_0687_));
 sky130_fd_sc_hd__or4_1 _1422_ (.A(_0035_),
    .B(_0038_),
    .C(_0086_),
    .D(_0093_),
    .X(_0688_));
 sky130_fd_sc_hd__or4_1 _1423_ (.A(_0683_),
    .B(_0686_),
    .C(_0687_),
    .D(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__a22o_1 _1424_ (.A1(net567),
    .A2(net645),
    .B1(net50),
    .B2(_0689_),
    .X(_0027_));
 sky130_fd_sc_hd__or4_1 _1425_ (.A(_0049_),
    .B(_0056_),
    .C(_0077_),
    .D(_0215_),
    .X(_0691_));
 sky130_fd_sc_hd__or4_1 _1426_ (.A(_0133_),
    .B(_0269_),
    .C(_0687_),
    .D(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__or2_1 _1427_ (.A(_0683_),
    .B(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__a22o_1 _1428_ (.A1(net563),
    .A2(net636),
    .B1(net46),
    .B2(_0693_),
    .X(_0028_));
 sky130_fd_sc_hd__or4_1 _1429_ (.A(_0191_),
    .B(_0274_),
    .C(_0275_),
    .D(_0683_),
    .X(_0694_));
 sky130_fd_sc_hd__a22o_1 _1430_ (.A1(net563),
    .A2(net635),
    .B1(net46),
    .B2(_0694_),
    .X(_0029_));
 sky130_fd_sc_hd__a22o_1 _1431_ (.A1(net558),
    .A2(net649),
    .B1(_0252_),
    .B2(net41),
    .X(_0030_));
 sky130_fd_sc_hd__dfxtp_1 _1432_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net1),
    .Q(\addr0_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1433_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net2),
    .Q(\addr0_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1434_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net3),
    .Q(\addr0_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1435_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net4),
    .Q(\addr0_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1436_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net5),
    .Q(\addr0_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1437_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net6),
    .Q(\addr0_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1438_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net7),
    .Q(\addr0_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1439_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net8),
    .Q(\addr0_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1440_ (.CLK(clknet_2_2__leaf_clk0),
    .D(net9),
    .Q(cs0_reg));
 sky130_fd_sc_hd__dfxtp_1 _1441_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0000_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_1 _1442_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0001_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_1 _1443_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0002_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _1444_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0003_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _1445_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0004_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _1446_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0005_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _1447_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0006_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _1448_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0007_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _1449_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0008_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _1450_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0009_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _1451_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0010_),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_1 _1452_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0011_),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_1 _1453_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0012_),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_1 _1454_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0013_),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_1 _1455_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0014_),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_1 _1456_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0015_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_1 _1457_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0016_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_1 _1458_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0017_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_1 _1459_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0018_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_1 _1460_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0019_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_1 _1461_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0020_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_1 _1462_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0021_),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_1 _1463_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0022_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_1 _1464_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0023_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_1 _1465_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0024_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_1 _1466_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0025_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_1 _1467_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0026_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _1468_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0027_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_1 _1469_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0028_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _1470_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0029_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _1471_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0030_),
    .Q(net33));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk0 (.A(clk0),
    .X(clknet_0_clk0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_443 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(addr0[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(addr0[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(addr0[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(addr0[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(addr0[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(addr0[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(addr0[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(addr0[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(cs0),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(dout0[0]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(dout0[10]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(dout0[11]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(dout0[12]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(dout0[13]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(dout0[14]));
 sky130_fd_sc_hd__clkbuf_4 output16 (.A(net16),
    .X(dout0[15]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(dout0[16]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(dout0[17]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(dout0[18]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(dout0[19]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(dout0[1]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(dout0[20]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(dout0[21]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(dout0[22]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(dout0[23]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(dout0[24]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(dout0[25]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(dout0[26]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(dout0[27]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(dout0[28]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(dout0[29]));
 sky130_fd_sc_hd__clkbuf_4 output32 (.A(net32),
    .X(dout0[2]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(dout0[30]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(dout0[3]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(dout0[4]));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net36),
    .X(dout0[5]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(dout0[6]));
 sky130_fd_sc_hd__clkbuf_4 output38 (.A(net38),
    .X(dout0[7]));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net39),
    .X(dout0[8]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(dout0[9]));
 sky130_fd_sc_hd__buf_1 fanout41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 fanout42 (.A(net49),
    .X(net42));
 sky130_fd_sc_hd__buf_1 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__buf_1 fanout45 (.A(net48),
    .X(net45));
 sky130_fd_sc_hd__buf_1 fanout46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 fanout47 (.A(net48),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__buf_1 fanout49 (.A(net56),
    .X(net49));
 sky130_fd_sc_hd__buf_1 fanout50 (.A(net52),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 fanout52 (.A(net54),
    .X(net52));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__buf_1 fanout54 (.A(net56),
    .X(net54));
 sky130_fd_sc_hd__buf_1 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout56 (.A(_0281_),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 wire57 (.A(_0174_),
    .X(net57));
 sky130_fd_sc_hd__buf_1 fanout58 (.A(_0344_),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 fanout59 (.A(_0334_),
    .X(net59));
 sky130_fd_sc_hd__buf_1 fanout60 (.A(_0303_),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 fanout61 (.A(_0206_),
    .X(net61));
 sky130_fd_sc_hd__buf_1 fanout62 (.A(_0194_),
    .X(net62));
 sky130_fd_sc_hd__buf_1 fanout63 (.A(_0187_),
    .X(net63));
 sky130_fd_sc_hd__buf_1 fanout64 (.A(_0187_),
    .X(net64));
 sky130_fd_sc_hd__buf_1 fanout65 (.A(_0166_),
    .X(net65));
 sky130_fd_sc_hd__buf_1 fanout66 (.A(_0148_),
    .X(net66));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout67 (.A(_0046_),
    .X(net67));
 sky130_fd_sc_hd__buf_1 fanout68 (.A(_0033_),
    .X(net68));
 sky130_fd_sc_hd__buf_1 fanout69 (.A(net71),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 fanout71 (.A(_0264_),
    .X(net71));
 sky130_fd_sc_hd__buf_1 fanout72 (.A(_0263_),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 fanout73 (.A(_0263_),
    .X(net73));
 sky130_fd_sc_hd__buf_1 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 fanout75 (.A(_0261_),
    .X(net75));
 sky130_fd_sc_hd__buf_1 fanout76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 fanout77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__buf_1 fanout78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 fanout79 (.A(_0260_),
    .X(net79));
 sky130_fd_sc_hd__buf_1 fanout80 (.A(_0257_),
    .X(net80));
 sky130_fd_sc_hd__buf_1 fanout81 (.A(_0257_),
    .X(net81));
 sky130_fd_sc_hd__buf_1 fanout82 (.A(_0256_),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 fanout83 (.A(_0256_),
    .X(net83));
 sky130_fd_sc_hd__buf_1 fanout84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 fanout85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__buf_1 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__buf_1 fanout87 (.A(_0255_),
    .X(net87));
 sky130_fd_sc_hd__buf_1 fanout88 (.A(_0254_),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 fanout89 (.A(_0254_),
    .X(net89));
 sky130_fd_sc_hd__buf_1 fanout90 (.A(net92),
    .X(net90));
 sky130_fd_sc_hd__buf_1 fanout91 (.A(net92),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 fanout92 (.A(_0251_),
    .X(net92));
 sky130_fd_sc_hd__buf_1 fanout93 (.A(_0249_),
    .X(net93));
 sky130_fd_sc_hd__buf_1 fanout94 (.A(_0249_),
    .X(net94));
 sky130_fd_sc_hd__buf_1 fanout95 (.A(net97),
    .X(net95));
 sky130_fd_sc_hd__buf_1 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout97 (.A(_0248_),
    .X(net97));
 sky130_fd_sc_hd__buf_1 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout99 (.A(_0246_),
    .X(net99));
 sky130_fd_sc_hd__buf_1 fanout100 (.A(_0245_),
    .X(net100));
 sky130_fd_sc_hd__buf_1 fanout101 (.A(net102),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 fanout102 (.A(_0241_),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 fanout103 (.A(_0240_),
    .X(net103));
 sky130_fd_sc_hd__buf_1 fanout104 (.A(_0240_),
    .X(net104));
 sky130_fd_sc_hd__buf_1 fanout105 (.A(_0238_),
    .X(net105));
 sky130_fd_sc_hd__buf_1 fanout106 (.A(_0238_),
    .X(net106));
 sky130_fd_sc_hd__buf_1 fanout107 (.A(net109),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__buf_1 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout110 (.A(_0235_),
    .X(net110));
 sky130_fd_sc_hd__buf_1 fanout111 (.A(_0234_),
    .X(net111));
 sky130_fd_sc_hd__buf_1 fanout112 (.A(_0233_),
    .X(net112));
 sky130_fd_sc_hd__buf_1 fanout113 (.A(_0233_),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 fanout114 (.A(_0232_),
    .X(net114));
 sky130_fd_sc_hd__buf_1 fanout115 (.A(_0232_),
    .X(net115));
 sky130_fd_sc_hd__buf_1 fanout116 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__buf_1 fanout117 (.A(_0227_),
    .X(net117));
 sky130_fd_sc_hd__buf_1 fanout118 (.A(net120),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 fanout119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__buf_1 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__buf_1 fanout121 (.A(_0226_),
    .X(net121));
 sky130_fd_sc_hd__buf_1 fanout122 (.A(_0224_),
    .X(net122));
 sky130_fd_sc_hd__buf_1 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout124 (.A(_0223_),
    .X(net124));
 sky130_fd_sc_hd__buf_1 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 fanout126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 fanout127 (.A(_0220_),
    .X(net127));
 sky130_fd_sc_hd__buf_1 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__buf_1 fanout129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 fanout130 (.A(_0219_),
    .X(net130));
 sky130_fd_sc_hd__buf_1 fanout131 (.A(_0218_),
    .X(net131));
 sky130_fd_sc_hd__buf_1 fanout132 (.A(_0218_),
    .X(net132));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 fanout134 (.A(_0217_),
    .X(net134));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout135 (.A(_0211_),
    .X(net135));
 sky130_fd_sc_hd__buf_1 fanout136 (.A(_0211_),
    .X(net136));
 sky130_fd_sc_hd__buf_1 fanout137 (.A(net139),
    .X(net137));
 sky130_fd_sc_hd__buf_1 fanout138 (.A(_0210_),
    .X(net138));
 sky130_fd_sc_hd__buf_1 fanout139 (.A(_0210_),
    .X(net139));
 sky130_fd_sc_hd__buf_1 fanout140 (.A(_0209_),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 fanout141 (.A(_0209_),
    .X(net141));
 sky130_fd_sc_hd__buf_1 fanout142 (.A(_0208_),
    .X(net142));
 sky130_fd_sc_hd__buf_1 fanout143 (.A(_0208_),
    .X(net143));
 sky130_fd_sc_hd__buf_1 fanout144 (.A(_0204_),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 fanout145 (.A(_0204_),
    .X(net145));
 sky130_fd_sc_hd__buf_1 fanout146 (.A(_0203_),
    .X(net146));
 sky130_fd_sc_hd__buf_1 fanout147 (.A(_0203_),
    .X(net147));
 sky130_fd_sc_hd__buf_1 fanout148 (.A(_0201_),
    .X(net148));
 sky130_fd_sc_hd__buf_1 fanout149 (.A(_0200_),
    .X(net149));
 sky130_fd_sc_hd__buf_1 fanout150 (.A(_0200_),
    .X(net150));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout151 (.A(net152),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 fanout152 (.A(_0196_),
    .X(net152));
 sky130_fd_sc_hd__buf_1 fanout153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout154 (.A(_0195_),
    .X(net154));
 sky130_fd_sc_hd__buf_1 fanout155 (.A(_0193_),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 fanout156 (.A(_0193_),
    .X(net156));
 sky130_fd_sc_hd__buf_1 fanout157 (.A(_0189_),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout159 (.A(_0189_),
    .X(net159));
 sky130_fd_sc_hd__buf_1 fanout160 (.A(_0188_),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 fanout161 (.A(_0188_),
    .X(net161));
 sky130_fd_sc_hd__buf_1 fanout162 (.A(_0185_),
    .X(net162));
 sky130_fd_sc_hd__buf_1 fanout163 (.A(net165),
    .X(net163));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout164 (.A(_0184_),
    .X(net164));
 sky130_fd_sc_hd__buf_1 fanout165 (.A(_0184_),
    .X(net165));
 sky130_fd_sc_hd__buf_1 fanout166 (.A(_0183_),
    .X(net166));
 sky130_fd_sc_hd__buf_1 fanout167 (.A(_0183_),
    .X(net167));
 sky130_fd_sc_hd__buf_1 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 fanout169 (.A(_0178_),
    .X(net169));
 sky130_fd_sc_hd__buf_1 fanout170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__buf_1 fanout171 (.A(_0177_),
    .X(net171));
 sky130_fd_sc_hd__buf_1 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout173 (.A(_0176_),
    .X(net173));
 sky130_fd_sc_hd__buf_1 fanout174 (.A(_0175_),
    .X(net174));
 sky130_fd_sc_hd__buf_1 fanout175 (.A(_0175_),
    .X(net175));
 sky130_fd_sc_hd__buf_1 fanout176 (.A(_0172_),
    .X(net176));
 sky130_fd_sc_hd__buf_1 fanout177 (.A(_0172_),
    .X(net177));
 sky130_fd_sc_hd__buf_1 fanout178 (.A(_0171_),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 fanout179 (.A(_0171_),
    .X(net179));
 sky130_fd_sc_hd__buf_1 fanout180 (.A(_0169_),
    .X(net180));
 sky130_fd_sc_hd__buf_1 fanout181 (.A(_0168_),
    .X(net181));
 sky130_fd_sc_hd__buf_1 fanout182 (.A(_0165_),
    .X(net182));
 sky130_fd_sc_hd__buf_1 fanout183 (.A(_0165_),
    .X(net183));
 sky130_fd_sc_hd__buf_1 fanout184 (.A(_0164_),
    .X(net184));
 sky130_fd_sc_hd__buf_1 fanout185 (.A(_0162_),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 fanout186 (.A(_0162_),
    .X(net186));
 sky130_fd_sc_hd__buf_1 fanout187 (.A(_0161_),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 fanout188 (.A(_0161_),
    .X(net188));
 sky130_fd_sc_hd__buf_1 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 fanout190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__buf_1 fanout191 (.A(_0154_),
    .X(net191));
 sky130_fd_sc_hd__buf_1 fanout192 (.A(net194),
    .X(net192));
 sky130_fd_sc_hd__buf_1 fanout193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 fanout194 (.A(_0152_),
    .X(net194));
 sky130_fd_sc_hd__buf_1 fanout195 (.A(_0151_),
    .X(net195));
 sky130_fd_sc_hd__buf_1 fanout196 (.A(_0147_),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 fanout197 (.A(_0147_),
    .X(net197));
 sky130_fd_sc_hd__buf_1 fanout198 (.A(_0146_),
    .X(net198));
 sky130_fd_sc_hd__buf_1 fanout199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__buf_1 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__buf_1 fanout201 (.A(_0144_),
    .X(net201));
 sky130_fd_sc_hd__buf_1 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__buf_1 fanout203 (.A(_0143_),
    .X(net203));
 sky130_fd_sc_hd__buf_1 fanout204 (.A(_0137_),
    .X(net204));
 sky130_fd_sc_hd__buf_1 fanout205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout206 (.A(_0136_),
    .X(net206));
 sky130_fd_sc_hd__buf_1 fanout207 (.A(_0135_),
    .X(net207));
 sky130_fd_sc_hd__buf_1 fanout208 (.A(_0135_),
    .X(net208));
 sky130_fd_sc_hd__buf_1 fanout209 (.A(_0134_),
    .X(net209));
 sky130_fd_sc_hd__buf_1 fanout210 (.A(_0134_),
    .X(net210));
 sky130_fd_sc_hd__buf_1 fanout211 (.A(net213),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout213 (.A(_0132_),
    .X(net213));
 sky130_fd_sc_hd__buf_1 fanout214 (.A(_0131_),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 fanout215 (.A(_0131_),
    .X(net215));
 sky130_fd_sc_hd__buf_1 fanout216 (.A(_0129_),
    .X(net216));
 sky130_fd_sc_hd__buf_1 fanout217 (.A(_0129_),
    .X(net217));
 sky130_fd_sc_hd__buf_1 fanout218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__buf_1 fanout219 (.A(_0128_),
    .X(net219));
 sky130_fd_sc_hd__buf_1 fanout220 (.A(_0125_),
    .X(net220));
 sky130_fd_sc_hd__buf_1 fanout221 (.A(net223),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_1 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__buf_1 fanout223 (.A(_0124_),
    .X(net223));
 sky130_fd_sc_hd__buf_1 fanout224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 fanout225 (.A(_0122_),
    .X(net225));
 sky130_fd_sc_hd__buf_1 fanout226 (.A(_0122_),
    .X(net226));
 sky130_fd_sc_hd__buf_1 fanout227 (.A(_0120_),
    .X(net227));
 sky130_fd_sc_hd__buf_1 fanout228 (.A(_0120_),
    .X(net228));
 sky130_fd_sc_hd__buf_1 fanout229 (.A(net231),
    .X(net229));
 sky130_fd_sc_hd__buf_1 fanout230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 fanout231 (.A(_0115_),
    .X(net231));
 sky130_fd_sc_hd__buf_1 fanout232 (.A(_0115_),
    .X(net232));
 sky130_fd_sc_hd__buf_1 fanout233 (.A(_0114_),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 fanout234 (.A(_0114_),
    .X(net234));
 sky130_fd_sc_hd__buf_1 fanout235 (.A(_0111_),
    .X(net235));
 sky130_fd_sc_hd__buf_1 fanout236 (.A(_0111_),
    .X(net236));
 sky130_fd_sc_hd__buf_1 fanout237 (.A(_0110_),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 fanout238 (.A(_0110_),
    .X(net238));
 sky130_fd_sc_hd__buf_1 fanout239 (.A(_0109_),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 fanout240 (.A(net241),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 fanout241 (.A(_0109_),
    .X(net241));
 sky130_fd_sc_hd__buf_1 fanout242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__buf_1 fanout243 (.A(net244),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_2 fanout244 (.A(_0104_),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_2 fanout245 (.A(_0103_),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_2 fanout246 (.A(_0102_),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_1 fanout247 (.A(_0102_),
    .X(net247));
 sky130_fd_sc_hd__buf_1 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout249 (.A(net250),
    .X(net249));
 sky130_fd_sc_hd__buf_1 fanout250 (.A(_0101_),
    .X(net250));
 sky130_fd_sc_hd__buf_1 fanout251 (.A(net252),
    .X(net251));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout252 (.A(_0097_),
    .X(net252));
 sky130_fd_sc_hd__buf_1 fanout253 (.A(net255),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 fanout254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__buf_1 fanout255 (.A(_0096_),
    .X(net255));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout256 (.A(_0095_),
    .X(net256));
 sky130_fd_sc_hd__buf_1 fanout257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__buf_1 fanout258 (.A(_0094_),
    .X(net258));
 sky130_fd_sc_hd__buf_1 fanout259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_2 fanout260 (.A(_0091_),
    .X(net260));
 sky130_fd_sc_hd__buf_1 fanout261 (.A(_0089_),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 fanout262 (.A(_0089_),
    .X(net262));
 sky130_fd_sc_hd__buf_1 fanout263 (.A(_0088_),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_1 fanout264 (.A(net265),
    .X(net264));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout265 (.A(_0088_),
    .X(net265));
 sky130_fd_sc_hd__buf_1 fanout266 (.A(net268),
    .X(net266));
 sky130_fd_sc_hd__buf_1 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout268 (.A(_0087_),
    .X(net268));
 sky130_fd_sc_hd__buf_1 fanout269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__buf_1 fanout270 (.A(_0084_),
    .X(net270));
 sky130_fd_sc_hd__buf_1 fanout271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_2 fanout272 (.A(net274),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 fanout273 (.A(net274),
    .X(net273));
 sky130_fd_sc_hd__buf_1 wire274 (.A(_0083_),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_2 fanout275 (.A(_0081_),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_2 fanout276 (.A(net280),
    .X(net276));
 sky130_fd_sc_hd__buf_1 fanout277 (.A(net280),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_2 fanout278 (.A(net280),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 fanout279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_2 fanout280 (.A(_0080_),
    .X(net280));
 sky130_fd_sc_hd__buf_1 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_2 fanout282 (.A(_0073_),
    .X(net282));
 sky130_fd_sc_hd__buf_1 fanout283 (.A(net285),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 fanout284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_2 fanout285 (.A(_0072_),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_1 fanout286 (.A(_0072_),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_2 fanout287 (.A(_0071_),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_1 fanout288 (.A(_0071_),
    .X(net288));
 sky130_fd_sc_hd__buf_1 fanout289 (.A(_0070_),
    .X(net289));
 sky130_fd_sc_hd__buf_1 fanout290 (.A(_0070_),
    .X(net290));
 sky130_fd_sc_hd__buf_1 fanout291 (.A(_0067_),
    .X(net291));
 sky130_fd_sc_hd__buf_1 fanout292 (.A(_0067_),
    .X(net292));
 sky130_fd_sc_hd__buf_1 fanout293 (.A(_0066_),
    .X(net293));
 sky130_fd_sc_hd__buf_1 fanout294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 fanout295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__buf_1 fanout296 (.A(_0064_),
    .X(net296));
 sky130_fd_sc_hd__buf_1 fanout297 (.A(_0063_),
    .X(net297));
 sky130_fd_sc_hd__buf_1 fanout298 (.A(_0063_),
    .X(net298));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout299 (.A(_0061_),
    .X(net299));
 sky130_fd_sc_hd__buf_1 fanout300 (.A(_0061_),
    .X(net300));
 sky130_fd_sc_hd__buf_1 fanout301 (.A(net303),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_1 fanout302 (.A(net303),
    .X(net302));
 sky130_fd_sc_hd__buf_1 fanout303 (.A(_0060_),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 fanout304 (.A(_0060_),
    .X(net304));
 sky130_fd_sc_hd__buf_1 fanout305 (.A(_0058_),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 fanout306 (.A(_0058_),
    .X(net306));
 sky130_fd_sc_hd__buf_1 fanout307 (.A(_0057_),
    .X(net307));
 sky130_fd_sc_hd__buf_1 fanout308 (.A(_0053_),
    .X(net308));
 sky130_fd_sc_hd__buf_1 fanout309 (.A(net310),
    .X(net309));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout310 (.A(_0052_),
    .X(net310));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout311 (.A(_0051_),
    .X(net311));
 sky130_fd_sc_hd__buf_1 fanout312 (.A(net314),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_1 fanout313 (.A(net314),
    .X(net313));
 sky130_fd_sc_hd__buf_1 fanout314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__buf_1 fanout315 (.A(_0045_),
    .X(net315));
 sky130_fd_sc_hd__buf_1 fanout316 (.A(_0043_),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_1 fanout317 (.A(_0043_),
    .X(net317));
 sky130_fd_sc_hd__buf_1 fanout318 (.A(_0042_),
    .X(net318));
 sky130_fd_sc_hd__buf_1 fanout319 (.A(net321),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 fanout320 (.A(net321),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_1 fanout321 (.A(net322),
    .X(net321));
 sky130_fd_sc_hd__buf_1 fanout322 (.A(_0041_),
    .X(net322));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout323 (.A(_0032_),
    .X(net323));
 sky130_fd_sc_hd__buf_1 fanout324 (.A(net326),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_1 fanout325 (.A(net326),
    .X(net325));
 sky130_fd_sc_hd__buf_1 fanout326 (.A(_0711_),
    .X(net326));
 sky130_fd_sc_hd__buf_1 fanout327 (.A(net328),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_2 fanout328 (.A(_0707_),
    .X(net328));
 sky130_fd_sc_hd__buf_1 fanout329 (.A(net331),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_1 fanout330 (.A(net331),
    .X(net330));
 sky130_fd_sc_hd__buf_1 fanout331 (.A(_0703_),
    .X(net331));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout332 (.A(_0700_),
    .X(net332));
 sky130_fd_sc_hd__buf_1 fanout333 (.A(_0700_),
    .X(net333));
 sky130_fd_sc_hd__buf_1 fanout334 (.A(_0696_),
    .X(net334));
 sky130_fd_sc_hd__buf_1 fanout335 (.A(net336),
    .X(net335));
 sky130_fd_sc_hd__buf_1 fanout336 (.A(_0680_),
    .X(net336));
 sky130_fd_sc_hd__buf_1 fanout337 (.A(net338),
    .X(net337));
 sky130_fd_sc_hd__buf_1 fanout338 (.A(net343),
    .X(net338));
 sky130_fd_sc_hd__buf_1 fanout339 (.A(net340),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_1 fanout340 (.A(net342),
    .X(net340));
 sky130_fd_sc_hd__buf_1 fanout341 (.A(net342),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_1 fanout342 (.A(net343),
    .X(net342));
 sky130_fd_sc_hd__buf_1 fanout343 (.A(_0216_),
    .X(net343));
 sky130_fd_sc_hd__buf_1 fanout344 (.A(net345),
    .X(net344));
 sky130_fd_sc_hd__buf_1 fanout345 (.A(net346),
    .X(net345));
 sky130_fd_sc_hd__buf_1 fanout346 (.A(net348),
    .X(net346));
 sky130_fd_sc_hd__buf_1 fanout347 (.A(net348),
    .X(net347));
 sky130_fd_sc_hd__buf_1 fanout348 (.A(_0182_),
    .X(net348));
 sky130_fd_sc_hd__buf_1 fanout349 (.A(net351),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_1 fanout350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__buf_1 fanout351 (.A(net352),
    .X(net351));
 sky130_fd_sc_hd__buf_1 fanout352 (.A(net355),
    .X(net352));
 sky130_fd_sc_hd__buf_1 fanout353 (.A(net355),
    .X(net353));
 sky130_fd_sc_hd__buf_1 fanout354 (.A(net355),
    .X(net354));
 sky130_fd_sc_hd__buf_1 fanout355 (.A(_0160_),
    .X(net355));
 sky130_fd_sc_hd__buf_1 fanout356 (.A(net358),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_1 fanout357 (.A(net358),
    .X(net357));
 sky130_fd_sc_hd__buf_1 fanout358 (.A(net359),
    .X(net358));
 sky130_fd_sc_hd__buf_1 fanout359 (.A(net361),
    .X(net359));
 sky130_fd_sc_hd__buf_1 fanout360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__buf_1 fanout361 (.A(_0159_),
    .X(net361));
 sky130_fd_sc_hd__buf_1 fanout362 (.A(net363),
    .X(net362));
 sky130_fd_sc_hd__buf_1 fanout363 (.A(net364),
    .X(net363));
 sky130_fd_sc_hd__buf_1 fanout364 (.A(net365),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_1 fanout365 (.A(net366),
    .X(net365));
 sky130_fd_sc_hd__buf_1 fanout366 (.A(net368),
    .X(net366));
 sky130_fd_sc_hd__buf_1 fanout367 (.A(net368),
    .X(net367));
 sky130_fd_sc_hd__buf_1 fanout368 (.A(_0142_),
    .X(net368));
 sky130_fd_sc_hd__buf_1 fanout369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__buf_1 fanout370 (.A(net371),
    .X(net370));
 sky130_fd_sc_hd__buf_1 fanout371 (.A(net372),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_1 fanout372 (.A(net373),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_1 fanout373 (.A(net376),
    .X(net373));
 sky130_fd_sc_hd__buf_1 fanout374 (.A(net375),
    .X(net374));
 sky130_fd_sc_hd__buf_1 fanout375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__buf_1 fanout376 (.A(_0141_),
    .X(net376));
 sky130_fd_sc_hd__buf_1 fanout377 (.A(net378),
    .X(net377));
 sky130_fd_sc_hd__buf_1 fanout378 (.A(net379),
    .X(net378));
 sky130_fd_sc_hd__buf_1 fanout379 (.A(net382),
    .X(net379));
 sky130_fd_sc_hd__buf_1 fanout380 (.A(net382),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_1 fanout381 (.A(net382),
    .X(net381));
 sky130_fd_sc_hd__buf_1 fanout382 (.A(_0121_),
    .X(net382));
 sky130_fd_sc_hd__buf_1 fanout383 (.A(net384),
    .X(net383));
 sky130_fd_sc_hd__buf_1 fanout384 (.A(net387),
    .X(net384));
 sky130_fd_sc_hd__buf_1 fanout385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__buf_1 fanout386 (.A(net387),
    .X(net386));
 sky130_fd_sc_hd__buf_1 fanout387 (.A(_0119_),
    .X(net387));
 sky130_fd_sc_hd__buf_1 fanout388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__buf_1 fanout389 (.A(net393),
    .X(net389));
 sky130_fd_sc_hd__buf_1 fanout390 (.A(net393),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_1 fanout391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__buf_1 fanout392 (.A(net393),
    .X(net392));
 sky130_fd_sc_hd__buf_1 fanout393 (.A(_0118_),
    .X(net393));
 sky130_fd_sc_hd__buf_1 fanout394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_1 fanout395 (.A(net396),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_1 fanout396 (.A(net397),
    .X(net396));
 sky130_fd_sc_hd__buf_1 fanout397 (.A(net400),
    .X(net397));
 sky130_fd_sc_hd__buf_1 fanout398 (.A(net400),
    .X(net398));
 sky130_fd_sc_hd__buf_1 fanout399 (.A(net400),
    .X(net399));
 sky130_fd_sc_hd__buf_1 fanout400 (.A(_0079_),
    .X(net400));
 sky130_fd_sc_hd__buf_1 fanout401 (.A(net402),
    .X(net401));
 sky130_fd_sc_hd__buf_1 fanout402 (.A(net403),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_1 fanout403 (.A(net404),
    .X(net403));
 sky130_fd_sc_hd__buf_1 fanout404 (.A(net405),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_1 fanout405 (.A(net408),
    .X(net405));
 sky130_fd_sc_hd__buf_1 fanout406 (.A(net408),
    .X(net406));
 sky130_fd_sc_hd__buf_1 fanout407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__buf_1 fanout408 (.A(_0078_),
    .X(net408));
 sky130_fd_sc_hd__buf_1 fanout409 (.A(_0050_),
    .X(net409));
 sky130_fd_sc_hd__buf_1 fanout410 (.A(_0050_),
    .X(net410));
 sky130_fd_sc_hd__buf_1 fanout411 (.A(net413),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_1 fanout412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_1 fanout413 (.A(net418),
    .X(net413));
 sky130_fd_sc_hd__buf_1 fanout414 (.A(net417),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_1 fanout415 (.A(net417),
    .X(net415));
 sky130_fd_sc_hd__buf_1 fanout416 (.A(net418),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_1 fanout417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__buf_1 fanout418 (.A(_0040_),
    .X(net418));
 sky130_fd_sc_hd__buf_1 fanout419 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_1 fanout420 (.A(net425),
    .X(net420));
 sky130_fd_sc_hd__buf_1 fanout421 (.A(net424),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_1 fanout422 (.A(net424),
    .X(net422));
 sky130_fd_sc_hd__buf_1 fanout423 (.A(net425),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_1 fanout424 (.A(net425),
    .X(net424));
 sky130_fd_sc_hd__buf_1 fanout425 (.A(_0039_),
    .X(net425));
 sky130_fd_sc_hd__buf_1 fanout426 (.A(net428),
    .X(net426));
 sky130_fd_sc_hd__buf_1 fanout427 (.A(net428),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_1 fanout428 (.A(net432),
    .X(net428));
 sky130_fd_sc_hd__buf_1 fanout429 (.A(net430),
    .X(net429));
 sky130_fd_sc_hd__buf_1 fanout430 (.A(net431),
    .X(net430));
 sky130_fd_sc_hd__buf_1 fanout431 (.A(net432),
    .X(net431));
 sky130_fd_sc_hd__buf_1 fanout432 (.A(_0031_),
    .X(net432));
 sky130_fd_sc_hd__buf_1 fanout433 (.A(net435),
    .X(net433));
 sky130_fd_sc_hd__buf_1 fanout434 (.A(net435),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_1 fanout435 (.A(net439),
    .X(net435));
 sky130_fd_sc_hd__buf_1 fanout436 (.A(net437),
    .X(net436));
 sky130_fd_sc_hd__buf_1 fanout437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__buf_1 fanout438 (.A(net439),
    .X(net438));
 sky130_fd_sc_hd__buf_1 fanout439 (.A(_0715_),
    .X(net439));
 sky130_fd_sc_hd__buf_1 fanout440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__buf_1 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__buf_1 fanout442 (.A(net447),
    .X(net442));
 sky130_fd_sc_hd__buf_1 fanout443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_1 fanout444 (.A(net445),
    .X(net444));
 sky130_fd_sc_hd__buf_1 fanout445 (.A(net446),
    .X(net445));
 sky130_fd_sc_hd__buf_1 fanout446 (.A(net447),
    .X(net446));
 sky130_fd_sc_hd__buf_1 fanout447 (.A(_0713_),
    .X(net447));
 sky130_fd_sc_hd__buf_1 fanout448 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__buf_1 fanout449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__buf_1 fanout450 (.A(net455),
    .X(net450));
 sky130_fd_sc_hd__buf_1 fanout451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_1 fanout452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__buf_1 fanout453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__buf_1 fanout454 (.A(net455),
    .X(net454));
 sky130_fd_sc_hd__buf_1 fanout455 (.A(_0712_),
    .X(net455));
 sky130_fd_sc_hd__buf_1 fanout456 (.A(net457),
    .X(net456));
 sky130_fd_sc_hd__buf_1 fanout457 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__buf_1 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__buf_1 fanout459 (.A(net464),
    .X(net459));
 sky130_fd_sc_hd__buf_1 fanout460 (.A(net462),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_1 fanout461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_1 fanout462 (.A(net463),
    .X(net462));
 sky130_fd_sc_hd__buf_1 fanout463 (.A(net464),
    .X(net463));
 sky130_fd_sc_hd__buf_1 fanout464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_1 wire465 (.A(_0710_),
    .X(net465));
 sky130_fd_sc_hd__buf_1 fanout466 (.A(net467),
    .X(net466));
 sky130_fd_sc_hd__buf_1 fanout467 (.A(net468),
    .X(net467));
 sky130_fd_sc_hd__buf_1 fanout468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__buf_1 fanout469 (.A(net474),
    .X(net469));
 sky130_fd_sc_hd__buf_1 fanout470 (.A(net472),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_1 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_1 fanout472 (.A(net473),
    .X(net472));
 sky130_fd_sc_hd__buf_1 fanout473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__buf_1 fanout474 (.A(_0709_),
    .X(net474));
 sky130_fd_sc_hd__buf_1 fanout475 (.A(net477),
    .X(net475));
 sky130_fd_sc_hd__buf_1 fanout476 (.A(net477),
    .X(net476));
 sky130_fd_sc_hd__buf_1 fanout477 (.A(net482),
    .X(net477));
 sky130_fd_sc_hd__buf_1 fanout478 (.A(net480),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_1 fanout479 (.A(net480),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_1 fanout480 (.A(net481),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_1 fanout481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__buf_1 fanout482 (.A(_0706_),
    .X(net482));
 sky130_fd_sc_hd__buf_1 fanout483 (.A(net484),
    .X(net483));
 sky130_fd_sc_hd__buf_1 fanout484 (.A(net485),
    .X(net484));
 sky130_fd_sc_hd__buf_1 fanout485 (.A(net490),
    .X(net485));
 sky130_fd_sc_hd__buf_1 fanout486 (.A(net488),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_1 fanout487 (.A(net488),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_1 fanout488 (.A(net489),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_1 fanout489 (.A(net490),
    .X(net489));
 sky130_fd_sc_hd__buf_1 fanout490 (.A(_0705_),
    .X(net490));
 sky130_fd_sc_hd__buf_1 fanout491 (.A(net493),
    .X(net491));
 sky130_fd_sc_hd__buf_1 fanout492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__buf_1 fanout493 (.A(net494),
    .X(net493));
 sky130_fd_sc_hd__buf_1 fanout494 (.A(net499),
    .X(net494));
 sky130_fd_sc_hd__buf_1 fanout495 (.A(net496),
    .X(net495));
 sky130_fd_sc_hd__clkbuf_1 fanout496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_1 fanout497 (.A(net498),
    .X(net497));
 sky130_fd_sc_hd__buf_1 fanout498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__buf_1 fanout499 (.A(_0702_),
    .X(net499));
 sky130_fd_sc_hd__buf_1 fanout500 (.A(net502),
    .X(net500));
 sky130_fd_sc_hd__buf_1 fanout501 (.A(net502),
    .X(net501));
 sky130_fd_sc_hd__buf_1 fanout502 (.A(net507),
    .X(net502));
 sky130_fd_sc_hd__buf_1 fanout503 (.A(net504),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_1 fanout504 (.A(net505),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_1 fanout505 (.A(net506),
    .X(net505));
 sky130_fd_sc_hd__buf_1 fanout506 (.A(net507),
    .X(net506));
 sky130_fd_sc_hd__buf_1 fanout507 (.A(_0701_),
    .X(net507));
 sky130_fd_sc_hd__buf_1 fanout508 (.A(net514),
    .X(net508));
 sky130_fd_sc_hd__buf_1 fanout509 (.A(net514),
    .X(net509));
 sky130_fd_sc_hd__buf_1 fanout510 (.A(net512),
    .X(net510));
 sky130_fd_sc_hd__buf_1 fanout511 (.A(net513),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_1 fanout512 (.A(net513),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_1 fanout513 (.A(net514),
    .X(net513));
 sky130_fd_sc_hd__buf_1 fanout514 (.A(_0699_),
    .X(net514));
 sky130_fd_sc_hd__buf_1 fanout515 (.A(net517),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_1 fanout516 (.A(net517),
    .X(net516));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout517 (.A(_0698_),
    .X(net517));
 sky130_fd_sc_hd__buf_1 fanout518 (.A(net519),
    .X(net518));
 sky130_fd_sc_hd__buf_1 fanout519 (.A(net520),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_1 fanout520 (.A(net521),
    .X(net520));
 sky130_fd_sc_hd__buf_1 fanout521 (.A(net524),
    .X(net521));
 sky130_fd_sc_hd__buf_1 fanout522 (.A(net523),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_1 fanout523 (.A(net524),
    .X(net523));
 sky130_fd_sc_hd__buf_1 fanout524 (.A(_0695_),
    .X(net524));
 sky130_fd_sc_hd__buf_1 fanout525 (.A(net526),
    .X(net525));
 sky130_fd_sc_hd__buf_1 fanout526 (.A(net527),
    .X(net526));
 sky130_fd_sc_hd__clkbuf_1 fanout527 (.A(net528),
    .X(net527));
 sky130_fd_sc_hd__buf_1 fanout528 (.A(net531),
    .X(net528));
 sky130_fd_sc_hd__buf_1 fanout529 (.A(net530),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_1 fanout530 (.A(net531),
    .X(net530));
 sky130_fd_sc_hd__buf_1 fanout531 (.A(_0690_),
    .X(net531));
 sky130_fd_sc_hd__buf_1 fanout532 (.A(net533),
    .X(net532));
 sky130_fd_sc_hd__buf_1 fanout533 (.A(net534),
    .X(net533));
 sky130_fd_sc_hd__buf_1 fanout534 (.A(net539),
    .X(net534));
 sky130_fd_sc_hd__buf_1 fanout535 (.A(net537),
    .X(net535));
 sky130_fd_sc_hd__clkbuf_1 fanout536 (.A(net537),
    .X(net536));
 sky130_fd_sc_hd__clkbuf_1 fanout537 (.A(net538),
    .X(net537));
 sky130_fd_sc_hd__buf_1 fanout538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__buf_1 fanout539 (.A(_0670_),
    .X(net539));
 sky130_fd_sc_hd__buf_1 fanout540 (.A(net543),
    .X(net540));
 sky130_fd_sc_hd__buf_1 fanout541 (.A(net543),
    .X(net541));
 sky130_fd_sc_hd__buf_1 fanout542 (.A(net543),
    .X(net542));
 sky130_fd_sc_hd__buf_1 fanout543 (.A(_0660_),
    .X(net543));
 sky130_fd_sc_hd__buf_1 fanout544 (.A(_0660_),
    .X(net544));
 sky130_fd_sc_hd__buf_1 fanout545 (.A(net546),
    .X(net545));
 sky130_fd_sc_hd__buf_1 fanout546 (.A(net547),
    .X(net546));
 sky130_fd_sc_hd__buf_1 fanout547 (.A(net552),
    .X(net547));
 sky130_fd_sc_hd__buf_1 fanout548 (.A(net550),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_1 fanout549 (.A(net550),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_1 fanout550 (.A(net551),
    .X(net550));
 sky130_fd_sc_hd__buf_1 fanout551 (.A(net552),
    .X(net551));
 sky130_fd_sc_hd__buf_1 fanout552 (.A(_0649_),
    .X(net552));
 sky130_fd_sc_hd__buf_1 fanout553 (.A(net556),
    .X(net553));
 sky130_fd_sc_hd__buf_1 fanout554 (.A(net556),
    .X(net554));
 sky130_fd_sc_hd__buf_1 fanout555 (.A(net556),
    .X(net555));
 sky130_fd_sc_hd__buf_1 fanout556 (.A(_0639_),
    .X(net556));
 sky130_fd_sc_hd__buf_1 fanout557 (.A(_0639_),
    .X(net557));
 sky130_fd_sc_hd__buf_1 fanout558 (.A(net559),
    .X(net558));
 sky130_fd_sc_hd__clkbuf_1 fanout559 (.A(net566),
    .X(net559));
 sky130_fd_sc_hd__buf_1 fanout560 (.A(net561),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_1 fanout561 (.A(net562),
    .X(net561));
 sky130_fd_sc_hd__buf_1 fanout562 (.A(net565),
    .X(net562));
 sky130_fd_sc_hd__buf_1 fanout563 (.A(net564),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_1 fanout564 (.A(net565),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_1 fanout565 (.A(net566),
    .X(net565));
 sky130_fd_sc_hd__buf_1 fanout566 (.A(net573),
    .X(net566));
 sky130_fd_sc_hd__buf_1 fanout567 (.A(net569),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_1 fanout568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_1 fanout569 (.A(net571),
    .X(net569));
 sky130_fd_sc_hd__buf_1 fanout570 (.A(net571),
    .X(net570));
 sky130_fd_sc_hd__buf_1 fanout571 (.A(net573),
    .X(net571));
 sky130_fd_sc_hd__buf_1 fanout572 (.A(net573),
    .X(net572));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout573 (.A(_0629_),
    .X(net573));
 sky130_fd_sc_hd__buf_1 fanout574 (.A(net575),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_1 fanout575 (.A(net576),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_1 fanout576 (.A(net580),
    .X(net576));
 sky130_fd_sc_hd__buf_1 fanout577 (.A(net580),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_1 fanout578 (.A(net579),
    .X(net578));
 sky130_fd_sc_hd__buf_1 fanout579 (.A(net580),
    .X(net579));
 sky130_fd_sc_hd__buf_1 fanout580 (.A(\addr0_reg[7] ),
    .X(net580));
 sky130_fd_sc_hd__buf_1 fanout581 (.A(net583),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_1 fanout582 (.A(net583),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_1 fanout583 (.A(net584),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_1 fanout584 (.A(net589),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_1 fanout585 (.A(net586),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_1 fanout586 (.A(net587),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_1 fanout587 (.A(net588),
    .X(net587));
 sky130_fd_sc_hd__buf_1 fanout588 (.A(net589),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_1 fanout589 (.A(\addr0_reg[6] ),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_1 fanout590 (.A(net591),
    .X(net590));
 sky130_fd_sc_hd__buf_1 fanout591 (.A(net596),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_1 fanout592 (.A(net593),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_1 fanout593 (.A(net594),
    .X(net593));
 sky130_fd_sc_hd__buf_1 fanout594 (.A(net595),
    .X(net594));
 sky130_fd_sc_hd__buf_1 fanout595 (.A(net596),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_1 fanout596 (.A(\addr0_reg[5] ),
    .X(net596));
 sky130_fd_sc_hd__buf_1 fanout597 (.A(net599),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_1 fanout598 (.A(net599),
    .X(net598));
 sky130_fd_sc_hd__buf_1 fanout599 (.A(net604),
    .X(net599));
 sky130_fd_sc_hd__buf_1 fanout600 (.A(net601),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_1 fanout601 (.A(net602),
    .X(net601));
 sky130_fd_sc_hd__buf_1 fanout602 (.A(net603),
    .X(net602));
 sky130_fd_sc_hd__buf_1 fanout603 (.A(net604),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_1 fanout604 (.A(\addr0_reg[4] ),
    .X(net604));
 sky130_fd_sc_hd__buf_1 fanout605 (.A(net610),
    .X(net605));
 sky130_fd_sc_hd__buf_1 fanout606 (.A(net610),
    .X(net606));
 sky130_fd_sc_hd__buf_1 fanout607 (.A(net608),
    .X(net607));
 sky130_fd_sc_hd__clkbuf_1 fanout608 (.A(net609),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_1 fanout609 (.A(net610),
    .X(net609));
 sky130_fd_sc_hd__buf_1 fanout610 (.A(\addr0_reg[3] ),
    .X(net610));
 sky130_fd_sc_hd__buf_1 fanout611 (.A(net612),
    .X(net611));
 sky130_fd_sc_hd__buf_1 fanout612 (.A(net616),
    .X(net612));
 sky130_fd_sc_hd__clkbuf_1 fanout613 (.A(net616),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_1 fanout614 (.A(net615),
    .X(net614));
 sky130_fd_sc_hd__buf_1 fanout615 (.A(net616),
    .X(net615));
 sky130_fd_sc_hd__buf_1 fanout616 (.A(\addr0_reg[2] ),
    .X(net616));
 sky130_fd_sc_hd__buf_1 fanout617 (.A(net622),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_1 fanout618 (.A(net622),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_1 fanout619 (.A(net620),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_1 fanout620 (.A(net621),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_1 fanout621 (.A(net622),
    .X(net621));
 sky130_fd_sc_hd__buf_1 fanout622 (.A(\addr0_reg[1] ),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_1 fanout623 (.A(net624),
    .X(net623));
 sky130_fd_sc_hd__buf_1 fanout624 (.A(net629),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_1 fanout625 (.A(net629),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_1 fanout626 (.A(net627),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_1 fanout627 (.A(net628),
    .X(net627));
 sky130_fd_sc_hd__clkbuf_1 fanout628 (.A(net629),
    .X(net628));
 sky130_fd_sc_hd__buf_1 fanout629 (.A(\addr0_reg[0] ),
    .X(net629));
 sky130_fd_sc_hd__conb_1 cust_rom0_630 (.LO(net630));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_0__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_1__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_2__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_3__leaf_clk0));
 sky130_fd_sc_hd__clkinv_4 clkload0 (.A(clknet_2_0__leaf_clk0));
 sky130_fd_sc_hd__clkinv_4 clkload1 (.A(clknet_2_1__leaf_clk0));
 sky130_fd_sc_hd__bufinv_16 clkload2 (.A(clknet_2_3__leaf_clk0));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net10),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net24),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net27),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net14),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net31),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net30),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net25),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net35),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net21),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net28),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net15),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net40),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net12),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net23),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net29),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net19),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net18),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net13),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net33),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net26),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net37),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net22),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net17),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net11),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net20),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net36),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net39),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net34),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net38),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net16),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net32),
    .X(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0033_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0033_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0055_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0059_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0071_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_0097_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0103_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_0164_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0238_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_0272_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_0272_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_0312_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_0312_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_0352_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_0553_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_0560_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_0586_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_0644_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_0272_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_0512_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(clknet_2_1__leaf_clk0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_341 ();
 assign dout0[31] = net630;
endmodule
