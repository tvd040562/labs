VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cust_rom
  CLASS BLOCK ;
  FOREIGN cust_rom ;
  ORIGIN 0.000 0.000 ;
  SIZE 142.465 BY 153.185 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 141.680 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 141.680 ;
    END
  END VPWR
  PIN addr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END addr0[7]
  PIN clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END clk0
  PIN cs0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 149.185 113.070 153.185 ;
    END
  END cs0
  PIN dout0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 64.640 142.465 65.240 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 91.840 142.465 92.440 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 27.240 142.465 27.840 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 71.440 142.465 72.040 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 88.440 142.465 89.040 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 149.185 74.430 153.185 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 74.840 142.465 75.440 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 85.040 142.465 85.640 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 34.040 142.465 34.640 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 149.185 93.750 153.185 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 44.240 142.465 44.840 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 61.240 142.465 61.840 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 47.640 142.465 48.240 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 40.840 142.465 41.440 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 95.240 142.465 95.840 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 30.640 142.465 31.240 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 51.040 142.465 51.640 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 98.640 142.465 99.240 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 108.840 142.465 109.440 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 105.440 142.465 106.040 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 102.040 142.465 102.640 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 115.640 142.465 116.240 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 81.640 142.465 82.240 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 149.185 106.630 153.185 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 149.185 109.850 153.185 ;
    END
  END dout0[31]
  PIN dout0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 54.440 142.465 55.040 ;
    END
  END dout0[3]
  PIN dout0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 37.440 142.465 38.040 ;
    END
  END dout0[4]
  PIN dout0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 149.185 90.530 153.185 ;
    END
  END dout0[5]
  PIN dout0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 68.040 142.465 68.640 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 138.465 78.240 142.465 78.840 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 149.185 80.870 153.185 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 149.185 77.650 153.185 ;
    END
  END dout0[9]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 136.810 141.525 ;
      LAYER li1 ;
        RECT 5.520 10.795 136.620 141.525 ;
      LAYER met1 ;
        RECT 4.210 10.640 136.620 141.680 ;
      LAYER met2 ;
        RECT 4.230 148.905 73.870 149.185 ;
        RECT 74.710 148.905 77.090 149.185 ;
        RECT 77.930 148.905 80.310 149.185 ;
        RECT 81.150 148.905 89.970 149.185 ;
        RECT 90.810 148.905 93.190 149.185 ;
        RECT 94.030 148.905 106.070 149.185 ;
        RECT 106.910 148.905 109.290 149.185 ;
        RECT 110.130 148.905 112.510 149.185 ;
        RECT 113.350 148.905 136.060 149.185 ;
        RECT 4.230 10.695 136.060 148.905 ;
      LAYER met3 ;
        RECT 2.110 133.640 138.465 141.605 ;
        RECT 4.400 132.240 138.465 133.640 ;
        RECT 2.110 130.240 138.465 132.240 ;
        RECT 4.400 128.840 138.465 130.240 ;
        RECT 2.110 126.840 138.465 128.840 ;
        RECT 4.400 125.440 138.465 126.840 ;
        RECT 2.110 123.440 138.465 125.440 ;
        RECT 4.400 122.040 138.465 123.440 ;
        RECT 2.110 116.640 138.465 122.040 ;
        RECT 2.110 115.240 138.065 116.640 ;
        RECT 2.110 113.240 138.465 115.240 ;
        RECT 4.400 111.840 138.465 113.240 ;
        RECT 2.110 109.840 138.465 111.840 ;
        RECT 2.110 108.440 138.065 109.840 ;
        RECT 2.110 106.440 138.465 108.440 ;
        RECT 2.110 105.040 138.065 106.440 ;
        RECT 2.110 103.040 138.465 105.040 ;
        RECT 2.110 101.640 138.065 103.040 ;
        RECT 2.110 99.640 138.465 101.640 ;
        RECT 4.400 98.240 138.065 99.640 ;
        RECT 2.110 96.240 138.465 98.240 ;
        RECT 2.110 94.840 138.065 96.240 ;
        RECT 2.110 92.840 138.465 94.840 ;
        RECT 2.110 91.440 138.065 92.840 ;
        RECT 2.110 89.440 138.465 91.440 ;
        RECT 2.110 88.040 138.065 89.440 ;
        RECT 2.110 86.040 138.465 88.040 ;
        RECT 4.400 84.640 138.065 86.040 ;
        RECT 2.110 82.640 138.465 84.640 ;
        RECT 2.110 81.240 138.065 82.640 ;
        RECT 2.110 79.240 138.465 81.240 ;
        RECT 2.110 77.840 138.065 79.240 ;
        RECT 2.110 75.840 138.465 77.840 ;
        RECT 2.110 74.440 138.065 75.840 ;
        RECT 2.110 72.440 138.465 74.440 ;
        RECT 2.110 71.040 138.065 72.440 ;
        RECT 2.110 69.040 138.465 71.040 ;
        RECT 2.110 67.640 138.065 69.040 ;
        RECT 2.110 65.640 138.465 67.640 ;
        RECT 4.400 64.240 138.065 65.640 ;
        RECT 2.110 62.240 138.465 64.240 ;
        RECT 2.110 60.840 138.065 62.240 ;
        RECT 2.110 55.440 138.465 60.840 ;
        RECT 2.110 54.040 138.065 55.440 ;
        RECT 2.110 52.040 138.465 54.040 ;
        RECT 2.110 50.640 138.065 52.040 ;
        RECT 2.110 48.640 138.465 50.640 ;
        RECT 2.110 47.240 138.065 48.640 ;
        RECT 2.110 45.240 138.465 47.240 ;
        RECT 2.110 43.840 138.065 45.240 ;
        RECT 2.110 41.840 138.465 43.840 ;
        RECT 2.110 40.440 138.065 41.840 ;
        RECT 2.110 38.440 138.465 40.440 ;
        RECT 4.400 37.040 138.065 38.440 ;
        RECT 2.110 35.040 138.465 37.040 ;
        RECT 2.110 33.640 138.065 35.040 ;
        RECT 2.110 31.640 138.465 33.640 ;
        RECT 2.110 30.240 138.065 31.640 ;
        RECT 2.110 28.240 138.465 30.240 ;
        RECT 2.110 26.840 138.065 28.240 ;
        RECT 2.110 10.715 138.465 26.840 ;
      LAYER met4 ;
        RECT 2.135 17.175 20.640 139.905 ;
        RECT 23.040 17.175 23.940 139.905 ;
        RECT 26.340 17.175 127.585 139.905 ;
      LAYER met5 ;
        RECT 14.380 65.500 125.460 97.700 ;
  END
END cust_rom
END LIBRARY

