logic [0:(ROM_DEPTH/2)-1] [DATA_WIDTH-1:0] table2 = {
32'h00000000,
32'hff36f170,
32'hfe6deaa1,
32'hfda4f351,
32'hfcdc1342,
32'hfc135231,
32'hfb4ab7db,
32'hfa824bfd,
32'hf9ba1651,
32'hf8f21e8e,
32'hf82a6c6a,
32'hf7630799,
32'hf69bf7c9,
32'hf5d544a7,
32'hf50ef5de,
32'hf4491311,
32'hf383a3e2,
32'hf2beafed,
32'hf1fa3ecb,
32'hf136580d,
32'hf0730342,
32'hefb047f2,
32'heeee2d9d,
32'hee2cbbc1,
32'hed6bf9d1,
32'hecabef3d,
32'hebeca36c,
32'heb2e1dbe,
32'hea70658a,
32'he9b38223,
32'he8f77acf,
32'he83c56cf,
32'he7821d59,
32'he6c8d59c,
32'he61086bc,
32'he55937d5,
32'he4a2eff6,
32'he3edb628,
32'he3399167,
32'he28688a4,
32'he1d4a2c8,
32'he123e6ad,
32'he0745b24,
32'hdfc606f1,
32'hdf18f0ce,
32'hde6d1f65,
32'hddc29958,
32'hdd196538,
32'hdc71898d,
32'hdbcb0cce,
32'hdb25f566,
32'hda8249b4,
32'hd9e01006,
32'hd93f4e9e,
32'hd8a00bae,
32'hd8024d59,
32'hd76619b6,
32'hd6cb76c9,
32'hd6326a88,
32'hd59afadb,
32'hd5052d97,
32'hd4710883,
32'hd3de9156,
32'hd34dcdb4,
32'hd2bec333,
32'hd2317756,
32'hd1a5ef90,
32'hd11c3142,
32'hd09441bb,
32'hd00e2639,
32'hcf89e3e8,
32'hcf077fe1,
32'hce86ff2a,
32'hce0866b8,
32'hcd8bbb6d,
32'hcd110216,
32'hcc983f70,
32'hcc217822,
32'hcbacb0bf,
32'hcb39edca,
32'hcac933ae,
32'hca5a86c4,
32'hc9edeb50,
32'hc9836582,
32'hc91af976,
32'hc8b4ab32,
32'hc8507ea7,
32'hc7ee77b3,
32'hc78e9a1d,
32'hc730e997,
32'hc6d569be,
32'hc67c1e18,
32'hc6250a18,
32'hc5d03118,
32'hc57d965d,
32'hc52d3d18,
32'hc4df2862,
32'hc4935b3c,
32'hc449d892,
32'hc402a33c,
32'hc3bdbdf6,
32'hc37b2b6a,
32'hc33aee27,
32'hc2fd08a9,
32'hc2c17d52,
32'hc2884e6e,
32'hc2517e31,
32'hc21d0eb8,
32'hc1eb0209,
32'hc1bb5a11,
32'hc18e18a7,
32'hc1633f8a,
32'hc13ad060,
32'hc114ccb9,
32'hc0f1360b,
32'hc0d00db6,
32'hc0b15502,
32'hc0950d1d,
32'hc07b371e,
32'hc063d405,
32'hc04ee4b8,
32'hc03c6a07,
32'hc02c64a6,
32'hc01ed535,
32'hc013bc39,
32'hc00b1a20,
32'hc004ef3f,
32'hc0013bd3,
32'hc0000000,
32'hc0013bd3,
32'hc004ef3f,
32'hc00b1a20,
32'hc013bc39,
32'hc01ed535,
32'hc02c64a6,
32'hc03c6a07,
32'hc04ee4b8,
32'hc063d405,
32'hc07b371e,
32'hc0950d1d,
32'hc0b15502,
32'hc0d00db6,
32'hc0f1360b,
32'hc114ccb9,
32'hc13ad060,
32'hc1633f8a,
32'hc18e18a7,
32'hc1bb5a11,
32'hc1eb0209,
32'hc21d0eb8,
32'hc2517e31,
32'hc2884e6e,
32'hc2c17d52,
32'hc2fd08a9,
32'hc33aee27,
32'hc37b2b6a,
32'hc3bdbdf6,
32'hc402a33c,
32'hc449d892,
32'hc4935b3c,
32'hc4df2862,
32'hc52d3d18,
32'hc57d965d,
32'hc5d03118,
32'hc6250a18,
32'hc67c1e18,
32'hc6d569be,
32'hc730e997,
32'hc78e9a1d,
32'hc7ee77b3,
32'hc8507ea7,
32'hc8b4ab32,
32'hc91af976,
32'hc9836582,
32'hc9edeb50,
32'hca5a86c4,
32'hcac933ae,
32'hcb39edca,
32'hcbacb0bf,
32'hcc217822,
32'hcc983f70,
32'hcd110216,
32'hcd8bbb6d,
32'hce0866b8,
32'hce86ff2a,
32'hcf077fe1,
32'hcf89e3e8,
32'hd00e2639,
32'hd09441bb,
32'hd11c3142,
32'hd1a5ef90,
32'hd2317756,
32'hd2bec333,
32'hd34dcdb4,
32'hd3de9156,
32'hd4710883,
32'hd5052d97,
32'hd59afadb,
32'hd6326a88,
32'hd6cb76c9,
32'hd76619b6,
32'hd8024d59,
32'hd8a00bae,
32'hd93f4e9e,
32'hd9e01006,
32'hda8249b4,
32'hdb25f566,
32'hdbcb0cce,
32'hdc71898d,
32'hdd196538,
32'hddc29958,
32'hde6d1f65,
32'hdf18f0ce,
32'hdfc606f1,
32'he0745b24,
32'he123e6ad,
32'he1d4a2c8,
32'he28688a4,
32'he3399167,
32'he3edb628,
32'he4a2eff6,
32'he55937d5,
32'he61086bc,
32'he6c8d59c,
32'he7821d59,
32'he83c56cf,
32'he8f77acf,
32'he9b38223,
32'hea70658a,
32'heb2e1dbe,
32'hebeca36c,
32'hecabef3d,
32'hed6bf9d1,
32'hee2cbbc1,
32'heeee2d9d,
32'hefb047f2,
32'hf0730342,
32'hf136580d,
32'hf1fa3ecb,
32'hf2beafed,
32'hf383a3e2,
32'hf4491311,
32'hf50ef5de,
32'hf5d544a7,
32'hf69bf7c9,
32'hf7630799,
32'hf82a6c6a,
32'hf8f21e8e,
32'hf9ba1651,
32'hfa824bfd,
32'hfb4ab7db,
32'hfc135231,
32'hfcdc1342,
32'hfda4f351,
32'hfe6deaa1,
32'hff36f170
};
