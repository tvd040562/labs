assign table_[0] = 16'h0000;
assign table_[1] = 16'h0324;
assign table_[2] = 16'h0646;
assign table_[3] = 16'h0964;
assign table_[4] = 16'h0c7c;
assign table_[5] = 16'h0f8d;
assign table_[6] = 16'h1294;
assign table_[7] = 16'h1590;
assign table_[8] = 16'h187e;
assign table_[9] = 16'h1b5d;
assign table_[10] = 16'h1e2b;
assign table_[11] = 16'h20e7;
assign table_[12] = 16'h238e;
assign table_[13] = 16'h2620;
assign table_[14] = 16'h289a;
assign table_[15] = 16'h2afb;
assign table_[16] = 16'h2d41;
assign table_[17] = 16'h2f6c;
assign table_[18] = 16'h3179;
assign table_[19] = 16'h3368;
assign table_[20] = 16'h3537;
assign table_[21] = 16'h36e5;
assign table_[22] = 16'h3871;
assign table_[23] = 16'h39db;
assign table_[24] = 16'h3b21;
assign table_[25] = 16'h3c42;
assign table_[26] = 16'h3d3f;
assign table_[27] = 16'h3e15;
assign table_[28] = 16'h3ec5;
assign table_[29] = 16'h3f4f;
assign table_[30] = 16'h3fb1;
assign table_[31] = 16'h3fec;
assign table_[32] = 16'h4000;
assign table_[33] = 16'h3fec;
assign table_[34] = 16'h3fb1;
assign table_[35] = 16'h3f4f;
assign table_[36] = 16'h3ec5;
assign table_[37] = 16'h3e15;
assign table_[38] = 16'h3d3f;
assign table_[39] = 16'h3c42;
assign table_[40] = 16'h3b21;
assign table_[41] = 16'h39db;
assign table_[42] = 16'h3871;
assign table_[43] = 16'h36e5;
assign table_[44] = 16'h3537;
assign table_[45] = 16'h3368;
assign table_[46] = 16'h3179;
assign table_[47] = 16'h2f6c;
assign table_[48] = 16'h2d41;
assign table_[49] = 16'h2afb;
assign table_[50] = 16'h289a;
assign table_[51] = 16'h2620;
assign table_[52] = 16'h238e;
assign table_[53] = 16'h20e7;
assign table_[54] = 16'h1e2b;
assign table_[55] = 16'h1b5d;
assign table_[56] = 16'h187e;
assign table_[57] = 16'h1590;
assign table_[58] = 16'h1294;
assign table_[59] = 16'h0f8d;
assign table_[60] = 16'h0c7c;
assign table_[61] = 16'h0964;
assign table_[62] = 16'h0646;
assign table_[63] = 16'h0324;
assign table_[64] = 16'h0000;
assign table_[65] = 16'hfcdc;
assign table_[66] = 16'hf9ba;
assign table_[67] = 16'hf69c;
assign table_[68] = 16'hf384;
assign table_[69] = 16'hf073;
assign table_[70] = 16'hed6c;
assign table_[71] = 16'hea70;
assign table_[72] = 16'he782;
assign table_[73] = 16'he4a3;
assign table_[74] = 16'he1d5;
assign table_[75] = 16'hdf19;
assign table_[76] = 16'hdc72;
assign table_[77] = 16'hd9e0;
assign table_[78] = 16'hd766;
assign table_[79] = 16'hd505;
assign table_[80] = 16'hd2bf;
assign table_[81] = 16'hd094;
assign table_[82] = 16'hce87;
assign table_[83] = 16'hcc98;
assign table_[84] = 16'hcac9;
assign table_[85] = 16'hc91b;
assign table_[86] = 16'hc78f;
assign table_[87] = 16'hc625;
assign table_[88] = 16'hc4df;
assign table_[89] = 16'hc3be;
assign table_[90] = 16'hc2c1;
assign table_[91] = 16'hc1eb;
assign table_[92] = 16'hc13b;
assign table_[93] = 16'hc0b1;
assign table_[94] = 16'hc04f;
assign table_[95] = 16'hc014;
assign table_[96] = 16'hc000;
assign table_[97] = 16'hc014;
assign table_[98] = 16'hc04f;
assign table_[99] = 16'hc0b1;
assign table_[100] = 16'hc13b;
assign table_[101] = 16'hc1eb;
assign table_[102] = 16'hc2c1;
assign table_[103] = 16'hc3be;
assign table_[104] = 16'hc4df;
assign table_[105] = 16'hc625;
assign table_[106] = 16'hc78f;
assign table_[107] = 16'hc91b;
assign table_[108] = 16'hcac9;
assign table_[109] = 16'hcc98;
assign table_[110] = 16'hce87;
assign table_[111] = 16'hd094;
assign table_[112] = 16'hd2bf;
assign table_[113] = 16'hd505;
assign table_[114] = 16'hd766;
assign table_[115] = 16'hd9e0;
assign table_[116] = 16'hdc72;
assign table_[117] = 16'hdf19;
assign table_[118] = 16'he1d5;
assign table_[119] = 16'he4a3;
assign table_[120] = 16'he782;
assign table_[121] = 16'hea70;
assign table_[122] = 16'hed6c;
assign table_[123] = 16'hf073;
assign table_[124] = 16'hf384;
assign table_[125] = 16'hf69c;
assign table_[126] = 16'hf9ba;
assign table_[127] = 16'hfcdc;
