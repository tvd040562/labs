logic [0:ROM_DEPTH-1] [DATA_WIDTH-1:0] table_ = {
32'h00000000,
32'h001921fb,
32'h003243f1,
32'h004b65e1,
32'h006487c4,
32'h007da998,
32'h0096cb58,
32'h00afed02,
32'h00c90e90,
32'h00e22fff,
32'h00fb514b,
32'h01147271,
32'h012d936c,
32'h0146b438,
32'h015fd4d2,
32'h0178f536,
32'h0192155f,
32'h01ab354b,
32'h01c454f5,
32'h01dd7459,
32'h01f69373,
32'h020fb240,
32'h0228d0bb,
32'h0241eee2,
32'h025b0caf,
32'h02742a1f,
32'h028d472e,
32'h02a663d8,
32'h02bf801a,
32'h02d89bf0,
32'h02f1b755,
32'h030ad245,
32'h0323ecbe,
32'h033d06bb,
32'h03562038,
32'h036f3931,
32'h038851a2,
32'h03a16988,
32'h03ba80df,
32'h03d397a3,
32'h03ecadcf,
32'h0405c361,
32'h041ed854,
32'h0437eca4,
32'h0451004d,
32'h046a134c,
32'h0483259d,
32'h049c373c,
32'h04b54825,
32'h04ce5854,
32'h04e767c5,
32'h05007674,
32'h0519845e,
32'h0532917f,
32'h054b9dd3,
32'h0564a955,
32'h057db403,
32'h0596bdd7,
32'h05afc6d0,
32'h05c8cee7,
32'h05e1d61b,
32'h05fadc66,
32'h0613e1c5,
32'h062ce634,
32'h0645e9af,
32'h065eec33,
32'h0677edbb,
32'h0690ee44,
32'h06a9edc9,
32'h06c2ec48,
32'h06dbe9bb,
32'h06f4e620,
32'h070de172,
32'h0726dbae,
32'h073fd4cf,
32'h0758ccd2,
32'h0771c3b3,
32'h078ab96e,
32'h07a3adff,
32'h07bca163,
32'h07d59396,
32'h07ee8493,
32'h08077457,
32'h082062de,
32'h08395024,
32'h08523c25,
32'h086b26de,
32'h0884104b,
32'h089cf867,
32'h08b5df30,
32'h08cec4a0,
32'h08e7a8b5,
32'h09008b6a,
32'h09196cbc,
32'h09324ca7,
32'h094b2b27,
32'h09640837,
32'h097ce3d5,
32'h0995bdfd,
32'h09ae96aa,
32'h09c76dd8,
32'h09e04385,
32'h09f917ac,
32'h0a11ea49,
32'h0a2abb59,
32'h0a438ad7,
32'h0a5c58c0,
32'h0a752510,
32'h0a8defc3,
32'h0aa6b8d5,
32'h0abf8043,
32'h0ad84609,
32'h0af10a22,
32'h0b09cc8c,
32'h0b228d42,
32'h0b3b4c40,
32'h0b540982,
32'h0b6cc506,
32'h0b857ec7,
32'h0b9e36c0,
32'h0bb6ecef,
32'h0bcfa150,
32'h0be853de,
32'h0c010496,
32'h0c19b374,
32'h0c326075,
32'h0c4b0b94,
32'h0c63b4ce,
32'h0c7c5c1e,
32'h0c950182,
32'h0cada4f5,
32'h0cc64673,
32'h0cdee5f9,
32'h0cf78383,
32'h0d101f0e,
32'h0d28b894,
32'h0d415013,
32'h0d59e586,
32'h0d7278eb,
32'h0d8b0a3d,
32'h0da39978,
32'h0dbc2698,
32'h0dd4b19a,
32'h0ded3a7b,
32'h0e05c135,
32'h0e1e45c6,
32'h0e36c82a,
32'h0e4f485c,
32'h0e67c65a,
32'h0e80421e,
32'h0e98bba7,
32'h0eb132ef,
32'h0ec9a7f3,
32'h0ee21aaf,
32'h0efa8b20,
32'h0f12f941,
32'h0f2b650f,
32'h0f43ce86,
32'h0f5c35a3,
32'h0f749a61,
32'h0f8cfcbe,
32'h0fa55cb4,
32'h0fbdba40,
32'h0fd6155f,
32'h0fee6e0d,
32'h1006c446,
32'h101f1807,
32'h1037694b,
32'h104fb80e,
32'h1068044e,
32'h10804e06,
32'h10989532,
32'h10b0d9d0,
32'h10c91bda,
32'h10e15b4e,
32'h10f99827,
32'h1111d263,
32'h112a09fc,
32'h11423ef0,
32'h115a713a,
32'h1172a0d7,
32'h118acdc4,
32'h11a2f7fc,
32'h11bb1f7c,
32'h11d3443f,
32'h11eb6643,
32'h12038584,
32'h121ba1fd,
32'h1233bbac,
32'h124bd28c,
32'h1263e699,
32'h127bf7d1,
32'h1294062f,
32'h12ac11af,
32'h12c41a4f,
32'h12dc2009,
32'h12f422db,
32'h130c22c1,
32'h13241fb6,
32'h133c19b8,
32'h135410c3,
32'h136c04d2,
32'h1383f5e3,
32'h139be3f2,
32'h13b3cefa,
32'h13cbb6f8,
32'h13e39be9,
32'h13fb7dc9,
32'h14135c94,
32'h142b3846,
32'h144310dd,
32'h145ae653,
32'h1472b8a5,
32'h148a87d1,
32'h14a253d1,
32'h14ba1ca3,
32'h14d1e242,
32'h14e9a4ac,
32'h150163dc,
32'h15191fcf,
32'h1530d881,
32'h15488dee,
32'h15604013,
32'h1577eeec,
32'h158f9a76,
32'h15a742ac,
32'h15bee78c,
32'h15d68911,
32'h15ee2738,
32'h1605c1fd,
32'h161d595d,
32'h1634ed53,
32'h164c7ddd,
32'h16640af7,
32'h167b949d,
32'h16931acb,
32'h16aa9d7e,
32'h16c21cb2,
32'h16d99864,
32'h16f1108f,
32'h17088531,
32'h171ff646,
32'h173763c9,
32'h174ecdb8,
32'h1766340f,
32'h177d96ca,
32'h1794f5e6,
32'h17ac515f,
32'h17c3a931,
32'h17dafd59,
32'h17f24dd3,
32'h18099a9c,
32'h1820e3b0,
32'h1838290c,
32'h184f6aab,
32'h1866a88a,
32'h187de2a7,
32'h189518fc,
32'h18ac4b87,
32'h18c37a44,
32'h18daa52f,
32'h18f1cc45,
32'h1908ef82,
32'h19200ee3,
32'h19372a64,
32'h194e4201,
32'h196555b8,
32'h197c6584,
32'h19937161,
32'h19aa794d,
32'h19c17d44,
32'h19d87d42,
32'h19ef7944,
32'h1a067145,
32'h1a1d6544,
32'h1a34553b,
32'h1a4b4128,
32'h1a622907,
32'h1a790cd4,
32'h1a8fec8c,
32'h1aa6c82b,
32'h1abd9faf,
32'h1ad47312,
32'h1aeb4253,
32'h1b020d6c,
32'h1b18d45c,
32'h1b2f971e,
32'h1b4655ae,
32'h1b5d100a,
32'h1b73c62d,
32'h1b8a7815,
32'h1ba125bd,
32'h1bb7cf23,
32'h1bce7442,
32'h1be51518,
32'h1bfbb1a0,
32'h1c1249d8,
32'h1c28ddbb,
32'h1c3f6d47,
32'h1c55f878,
32'h1c6c7f4a,
32'h1c8301b9,
32'h1c997fc4,
32'h1caff965,
32'h1cc66e99,
32'h1cdcdf5e,
32'h1cf34baf,
32'h1d09b389,
32'h1d2016e9,
32'h1d3675cb,
32'h1d4cd02c,
32'h1d632608,
32'h1d79775c,
32'h1d8fc424,
32'h1da60c5d,
32'h1dbc5004,
32'h1dd28f15,
32'h1de8c98c,
32'h1dfeff67,
32'h1e1530a1,
32'h1e2b5d38,
32'h1e418528,
32'h1e57a86d,
32'h1e6dc705,
32'h1e83e0eb,
32'h1e99f61d,
32'h1eb00696,
32'h1ec61254,
32'h1edc1953,
32'h1ef21b90,
32'h1f081907,
32'h1f1e11b5,
32'h1f340596,
32'h1f49f4a8,
32'h1f5fdee6,
32'h1f75c44e,
32'h1f8ba4dc,
32'h1fa1808c,
32'h1fb7575c,
32'h1fcd2948,
32'h1fe2f64c,
32'h1ff8be65,
32'h200e8190,
32'h20243fca,
32'h2039f90f,
32'h204fad5b,
32'h20655cac,
32'h207b06fe,
32'h2090ac4d,
32'h20a64c97,
32'h20bbe7d8,
32'h20d17e0d,
32'h20e70f32,
32'h20fc9b44,
32'h21122240,
32'h2127a423,
32'h213d20e8,
32'h2152988d,
32'h21680b0f,
32'h217d786a,
32'h2192e09b,
32'h21a8439e,
32'h21bda171,
32'h21d2fa0f,
32'h21e84d76,
32'h21fd9ba3,
32'h2212e492,
32'h2228283f,
32'h223d66a8,
32'h22529fca,
32'h2267d3a0,
32'h227d0228,
32'h22922b5e,
32'h22a74f40,
32'h22bc6dca,
32'h22d186f8,
32'h22e69ac8,
32'h22fba936,
32'h2310b23e,
32'h2325b5df,
32'h233ab414,
32'h234facda,
32'h2364a02e,
32'h23798e0d,
32'h238e7673,
32'h23a3595e,
32'h23b836ca,
32'h23cd0eb3,
32'h23e1e117,
32'h23f6adf3,
32'h240b7543,
32'h24203704,
32'h2434f332,
32'h2449a9cc,
32'h245e5acc,
32'h24730631,
32'h2487abf7,
32'h249c4c1b,
32'h24b0e699,
32'h24c57b6f,
32'h24da0a9a,
32'h24ee9415,
32'h250317df,
32'h251795f3,
32'h252c0e4f,
32'h254080ef,
32'h2554edd1,
32'h256954f1,
32'h257db64c,
32'h259211df,
32'h25a667a7,
32'h25bab7a0,
32'h25cf01c8,
32'h25e3461b,
32'h25f78497,
32'h260bbd37,
32'h261feffa,
32'h26341cdb,
32'h264843d9,
32'h265c64ef,
32'h2670801a,
32'h26849558,
32'h2698a4a6,
32'h26acadff,
32'h26c0b162,
32'h26d4aecb,
32'h26e8a637,
32'h26fc97a3,
32'h2710830c,
32'h2724686e,
32'h273847c8,
32'h274c2115,
32'h275ff452,
32'h2773c17d,
32'h27878893,
32'h279b4990,
32'h27af0472,
32'h27c2b934,
32'h27d667d5,
32'h27ea1052,
32'h27fdb2a7,
32'h28114ed0,
32'h2824e4cc,
32'h28387498,
32'h284bfe2f,
32'h285f8190,
32'h2872feb6,
32'h288675a0,
32'h2899e64a,
32'h28ad50b1,
32'h28c0b4d2,
32'h28d412ab,
32'h28e76a37,
32'h28fabb75,
32'h290e0661,
32'h29214af8,
32'h29348937,
32'h2947c11c,
32'h295af2a3,
32'h296e1dc9,
32'h2981428c,
32'h299460e8,
32'h29a778db,
32'h29ba8a61,
32'h29cd9578,
32'h29e09a1c,
32'h29f3984c,
32'h2a069003,
32'h2a19813f,
32'h2a2c6bfd,
32'h2a3f503a,
32'h2a522df3,
32'h2a650525,
32'h2a77d5ce,
32'h2a8a9fea,
32'h2a9d6377,
32'h2ab02071,
32'h2ac2d6d6,
32'h2ad586a3,
32'h2ae82fd5,
32'h2afad269,
32'h2b0d6e5c,
32'h2b2003ac,
32'h2b329255,
32'h2b451a55,
32'h2b579ba8,
32'h2b6a164d,
32'h2b7c8a3f,
32'h2b8ef77d,
32'h2ba15e03,
32'h2bb3bdce,
32'h2bc616dd,
32'h2bd8692b,
32'h2beab4b6,
32'h2bfcf97c,
32'h2c0f3779,
32'h2c216eaa,
32'h2c339f0e,
32'h2c45c8a0,
32'h2c57eb5e,
32'h2c6a0746,
32'h2c7c1c55,
32'h2c8e2a87,
32'h2ca031da,
32'h2cb2324c,
32'h2cc42bd9,
32'h2cd61e7f,
32'h2ce80a3a,
32'h2cf9ef09,
32'h2d0bcce8,
32'h2d1da3d5,
32'h2d2f73cd
};
