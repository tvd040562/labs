* NGSPICE file created from cust_rom1.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

.subckt cust_rom1 addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7]
+ clk0 cs0 dout0[0] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[16]
+ dout0[17] dout0[18] dout0[19] dout0[1] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24]
+ dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[2] dout0[30] dout0[31] dout0[3]
+ dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] vccd1 vssd1
XTAP_TAPCELL_ROW_52_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1270_ net223 net220 net218 vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0985_ _0278_ _0284_ _0294_ _0296_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__or4_1
X_1399_ clknet_2_3__leaf_clk0 _0017_ vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__dfxtp_1
Xfanout127 _0211_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout105 net106 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__buf_1
Xfanout138 _0202_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
Xfanout116 net118 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__buf_1
Xfanout149 _0187_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0770_ net561 net567 net574 net581 vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__and4b_1
X_1322_ net217 net199 net153 net129 vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__or4_1
X_1253_ _0062_ net202 _0459_ _0540_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__or4_1
X_1184_ _0309_ _0481_ _0483_ _0484_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_19_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0968_ net195 net193 vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0899_ net471 net346 net339 net462 vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout480 net481 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout491 net492 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_16_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0822_ net440 net395 net387 net433 vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0753_ net524 net422 net415 net536 vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1236_ _0499_ _0519_ _0529_ _0532_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__or4_1
X_1305_ net309 _0206_ _0239_ _0596_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__or4_1
X_1167_ _0179_ _0192_ _0339_ _0347_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1098_ net300 net296 net215 net212 vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__or4_1
XFILLER_0_51_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1021_ _0073_ net89 net85 vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__or3_2
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0805_ net571 net578 net559 net564 vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__and4b_1
X_0736_ net304 net301 net296 vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1219_ _0040_ _0157_ _0514_ _0516_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold30 net36 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_5 _0123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1004_ _0299_ _0301_ _0314_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_32_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0719_ net322 net315 vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 dout0[29] sky130_fd_sc_hd__buf_2
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 dout0[19] sky130_fd_sc_hd__buf_2
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout309 _0038_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_1
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0984_ net246 net120 _0282_ _0295_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1398_ clknet_2_1__leaf_clk0 _0016_ vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__dfxtp_1
Xfanout128 _0210_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_1
Xfanout139 net140 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_1
Xfanout117 net118 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_1
Xfanout106 _0229_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_49_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_19_Left_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1252_ _0147_ net79 net78 _0547_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__or4_1
X_1321_ _0069_ net180 net67 vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__or3_1
X_1183_ _0075_ _0103_ _0113_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_19_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0967_ net285 net208 vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0898_ net454 net345 net338 net447 vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout470 net471 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_1
Xfanout481 _0680_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_1
Xfanout492 net493 vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_16_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0821_ net497 net394 net388 net503 vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__a22o_1
X_0752_ net287 net285 vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1166_ _0123_ _0171_ _0412_ _0467_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_39_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1235_ _0475_ _0520_ _0521_ _0531_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__or4_1
X_1304_ net232 net226 net222 net152 vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__or4_1
X_1097_ net88 net86 net83 vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1020_ _0190_ _0243_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0804_ net580 net560 net566 net573 vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__nor4b_1
X_0735_ net304 net298 vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__or2_1
X_1218_ net233 net113 _0246_ _0515_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1149_ _0240_ _0270_ _0445_ _0451_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold31 net18 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 net28 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_6 _0140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Left_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1003_ _0192_ _0199_ _0250_ net60 vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0718_ net531 net450 net443 net518 vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 dout0[1] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_33_Left_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput10 net10 vssd1 vssd1 vccd1 vccd1 dout0[0] sky130_fd_sc_hd__buf_2
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 dout0[2] sky130_fd_sc_hd__buf_2
XFILLER_0_41_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0983_ net187 net183 net173 net168 vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__or4_1
Xfanout129 net131 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_1
Xfanout118 _0223_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__buf_1
Xfanout107 net109 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__buf_1
X_1397_ clknet_2_2__leaf_clk0 _0015_ vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1320_ _0180_ _0199_ _0204_ _0304_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__or4_1
X_1251_ net137 net113 net110 net104 vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__or4_1
X_1182_ _0080_ net259 net199 _0482_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_20_Left_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0897_ net486 net344 net339 net479 vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0966_ _0164_ _0277_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout471 net472 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_1
Xfanout460 net461 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_1
Xfanout482 net483 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_1
Xfanout493 net494 vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_16_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0751_ net509 net426 net420 net516 vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0820_ net437 net367 net361 net429 vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1303_ _0299_ _0460_ _0593_ _0594_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__or4_1
X_1096_ net172 net167 net159 net155 vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__or4_1
X_1234_ net212 net204 _0181_ _0530_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__or4_1
X_1165_ net320 net223 net97 net73 vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__or4_1
X_0949_ net447 net427 net419 net454 vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout290 net291 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_1
X_0803_ _0107_ net63 _0113_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0734_ net521 net483 net476 net533 vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1217_ net265 net153 net145 vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__or3_1
X_1148_ net275 net107 net92 _0450_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__or4_1
X_1079_ net236 net120 net81 net80 vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold10 net30 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 net19 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 _0160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1002_ _0277_ _0309_ _0310_ _0312_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0717_ net589 net597 net603 net613 vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_50_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput11 net11 vssd1 vssd1 vccd1 vccd1 dout0[10] sky130_fd_sc_hd__clkbuf_4
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 dout0[20] sky130_fd_sc_hd__clkbuf_4
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 dout0[30] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0982_ _0180_ _0279_ _0280_ _0281_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout119 net120 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__buf_1
Xfanout108 net109 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1396_ clknet_2_3__leaf_clk0 _0014_ vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1250_ net286 net210 _0253_ _0536_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__or4_1
X_1181_ net210 net176 net129 net124 vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0965_ net130 net128 net126 vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__or3_2
X_0896_ net138 net136 net134 net133 vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__or4_2
XFILLER_0_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1379_ _0130_ net203 net201 _0218_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout472 net473 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_1
Xfanout483 net484 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__buf_1
Xfanout450 net452 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_1
Xfanout461 net466 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_1
Xfanout494 net496 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_16_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0750_ net491 net423 net416 net499 vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__a22o_1
Xfanout90 _0245_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_1
X_1302_ _0064_ _0148_ _0326_ _0348_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__or4_1
X_1233_ net251 net244 net237 net235 vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1164_ _0462_ _0463_ _0464_ _0465_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__or4_1
X_1095_ _0221_ _0237_ _0399_ _0400_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__or4_1
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0948_ net429 net425 net418 net436 vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0879_ net150 net148 net146 vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout280 net281 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_1
Xfanout291 _0056_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_2
X_0802_ net240 _0112_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__or2_2
XFILLER_0_8_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0733_ net520 net467 net459 net532 vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__a22o_1
X_1216_ _0364_ _0462_ _0513_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1078_ net167 net139 net133 net128 vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__or4_1
X_1147_ net315 net260 net252 net236 vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold22 net13 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 net40 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_8 _0181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ net228 net226 net190 _0311_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0716_ net602 net611 net588 net596 vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__and4b_1
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 dout0[21] sky130_fd_sc_hd__clkbuf_4
Xoutput34 net34 vssd1 vssd1 vccd1 vccd1 dout0[31] sky130_fd_sc_hd__buf_2
Xoutput12 net12 vssd1 vssd1 vccd1 vccd1 dout0[11] sky130_fd_sc_hd__buf_2
XFILLER_0_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0981_ _0088_ _0093_ _0291_ _0292_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__or4_1
XFILLER_0_13_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1395_ clknet_2_3__leaf_clk0 _0013_ vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout109 _0228_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_49_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout610 net611 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1180_ _0678_ _0365_ _0417_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__or3_1
X_0964_ _0218_ _0271_ _0275_ cs0_reg vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__o31a_1
XFILLER_0_27_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0895_ net136 net132 vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__or2_1
X_1378_ net553 net625 net53 _0665_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout440 net441 vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_1
Xfanout462 net463 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_1
Xfanout473 net474 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout451 net452 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_1
Xfanout484 net488 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_1
Xfanout495 net496 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_1
Xfanout80 _0256_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_24_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout91 _0245_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dlymetal6s2s_1
X_1301_ net74 net66 _0521_ _0536_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__or4_1
X_1232_ _0281_ _0525_ _0526_ _0528_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_47_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1094_ net311 net307 net138 net107 vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__or4_1
X_1163_ net300 net296 net121 net118 vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__or4_1
X_0947_ net79 net59 vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0878_ net151 net149 vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload0 clknet_2_0__leaf_clk0 vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_18_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout270 _0078_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_1
Xfanout281 _0069_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_1
Xfanout292 _0055_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__buf_1
X_0801_ net238 _0112_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0732_ net520 net436 net430 net532 vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1146_ net206 net186 net162 net156 vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__or4_1
X_1215_ net262 net257 net254 vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1077_ _0191_ _0328_ _0380_ _0381_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold23 net17 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 net39 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_9 _0186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1000_ net253 net250 net214 net103 vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0715_ net575 net457 net582 net568 vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_12_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1129_ _0397_ _0415_ _0431_ _0432_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 dout0[22] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput13 net13 vssd1 vssd1 vccd1 vccd1 dout0[12] sky130_fd_sc_hd__buf_2
Xoutput35 net35 vssd1 vssd1 vccd1 vccd1 dout0[3] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0980_ net294 net248 net231 net225 vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1394_ clknet_2_2__leaf_clk0 _0012_ vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__dfxtp_1
Xfanout611 net615 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_1
Xfanout600 net602 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0963_ _0051_ _0272_ _0273_ _0274_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_27_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0894_ net498 net343 net337 net495 vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1377_ _0051_ _0183_ _0651_ _0664_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout463 net464 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__clkbuf_1
Xfanout474 _0682_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_1
Xfanout441 net442 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_1
Xfanout430 net431 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_1
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_1
Xfanout485 net487 vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_1
Xfanout496 _0673_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__buf_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout70 net71 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__buf_1
Xfanout81 _0255_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_24_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout92 _0242_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_24_Left_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1231_ _0129_ _0513_ _0522_ _0527_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__or4_1
X_1300_ _0060_ _0491_ _0588_ _0591_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__or4_1
X_1162_ net251 net248 net247 vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1093_ net322 net134 net112 _0398_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0946_ net81 net77 vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0877_ net148 net147 vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_38_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload1 clknet_2_1__leaf_clk0 vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout293 _0055_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__buf_1
Xfanout282 net284 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_1
Xfanout271 _0077_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_1
Xfanout260 net261 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_44_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0800_ net503 net406 net398 net496 vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__a22o_1
X_0731_ net521 net450 net443 net533 vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1145_ net207 net186 vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__or2_1
X_1214_ _0378_ _0427_ _0510_ _0511_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1076_ _0107_ _0128_ _0379_ _0382_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0929_ net482 net379 net373 net475 vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__a22o_1
Xhold24 net22 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 net32 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0714_ net605 net614 net591 net598 vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_27_Left_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1128_ net173 net168 net162 net156 vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_11_Left_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1059_ _0164_ _0266_ _0341_ _0366_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__or4_1
XFILLER_0_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput14 net14 vssd1 vssd1 vccd1 vccd1 dout0[13] sky130_fd_sc_hd__buf_2
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 dout0[23] sky130_fd_sc_hd__buf_2
Xoutput36 net36 vssd1 vssd1 vccd1 vccd1 dout0[4] sky130_fd_sc_hd__buf_2
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1393_ clknet_2_1__leaf_clk0 _0011_ vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout612 net613 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_1
Xfanout601 net602 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0893_ net538 net342 net335 net526 vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__a22o_1
X_0962_ _0061_ _0149_ _0266_ _0270_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1376_ net247 _0201_ _0225_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout486 net487 vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__clkbuf_1
Xfanout464 net465 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_1
Xfanout420 net421 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout442 _0034_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_1
Xfanout497 _0673_ vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__clkbuf_1
Xfanout453 net456 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__buf_1
Xfanout431 net435 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_1
Xfanout475 net476 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__buf_1
Xfanout71 _0261_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__buf_1
Xfanout60 _0258_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout82 _0255_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_1
Xfanout93 _0242_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1092_ net189 net184 net182 vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__or3_1
X_1230_ net197 net71 net69 vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__or3_1
X_1161_ net143 net139 net136 net133 vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_47_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0945_ net473 net397 net391 net465 vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0876_ net493 net342 net336 net501 vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1359_ _0066_ _0644_ _0646_ _0647_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_41_Left_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout272 net274 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_1
Xfanout283 net284 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_1
Xfanout250 net251 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_1
Xfanout294 _0054_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_1
Xfanout261 _0087_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_44_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0730_ net312 net310 net309 net307 vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__or4_1
XFILLER_0_21_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1213_ _0058_ _0073_ _0170_ _0264_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__or4_1
X_1144_ net293 net289 net71 net64 vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1075_ net267 net262 net255 vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0859_ net172 net169 net167 net165 vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0928_ _0233_ net102 net99 net96 vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__or4_1
Xhold25 net11 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 net10 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0713_ net323 net318 vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1127_ net331 net271 net98 net96 vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__or4_1
X_1058_ _0032_ _0362_ _0364_ _0365_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput15 net15 vssd1 vssd1 vccd1 vccd1 dout0[14] sky130_fd_sc_hd__buf_2
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 dout0[24] sky130_fd_sc_hd__buf_2
Xoutput37 net37 vssd1 vssd1 vccd1 vccd1 dout0[5] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1392_ clknet_2_3__leaf_clk0 _0010_ vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout613 net614 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_1
Xfanout602 net606 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0961_ _0142_ _0225_ _0232_ _0254_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0892_ net137 _0203_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__or2_2
XFILLER_0_49_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1375_ net551 net620 net51 _0663_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout487 net488 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_1
Xfanout465 net466 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout454 net455 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_1
Xfanout432 net433 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__buf_1
Xfanout410 net411 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__buf_1
Xfanout421 _0053_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_1
Xfanout476 net477 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_1
Xfanout443 net445 vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_1
Xfanout498 net502 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_1
XFILLER_0_51_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout50 net52 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_1
Xfanout61 _0135_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_1
Xfanout72 net76 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_24_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout83 net84 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__buf_1
Xfanout94 _0241_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_1
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1091_ net293 net291 net231 net228 vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__or4_1
X_1160_ net334 net327 net149 net101 vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__or4_1
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0944_ net454 net393 net387 net447 vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0875_ net524 net343 net335 net536 vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__a22o_1
X_1358_ _0207_ net107 net72 _0429_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__or4_1
X_1289_ net280 net198 net126 net80 vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_38_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout240 _0109_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_1
Xfanout273 net274 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_1
Xfanout251 _0101_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout262 net263 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_1
Xfanout295 _0054_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_1
Xfanout284 _0065_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1212_ _0148_ _0304_ _0444_ _0509_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_35_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1143_ net224 net222 net85 net84 vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1074_ net217 net204 net200 vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0927_ net103 net96 vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__or2_1
X_0858_ net171 net167 vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0789_ net380 net374 net490 vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__o21ba_1
Xhold26 net34 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 net21 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0712_ net532 net467 net459 net520 vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1126_ _0133_ net199 net192 net161 vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__or4_1
X_1057_ net267 net263 net88 net83 vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput16 net16 vssd1 vssd1 vccd1 vccd1 dout0[15] sky130_fd_sc_hd__buf_2
Xoutput38 net38 vssd1 vssd1 vccd1 vccd1 dout0[6] sky130_fd_sc_hd__buf_2
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 dout0[25] sky130_fd_sc_hd__buf_2
Xclkbuf_2_3__f_clk0 clknet_0_clk0 vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1109_ _0042_ net62 vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1391_ clknet_2_1__leaf_clk0 _0009_ vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout603 net604 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__buf_1
Xfanout614 net615 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_5_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0960_ _0090_ _0097_ _0267_ _0268_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0891_ net515 net343 net337 net508 vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__a22o_1
X_1374_ _0652_ _0661_ _0662_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_2_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout411 net412 vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__clkbuf_1
Xfanout400 net401 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_1
Xfanout422 net423 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_1
Xfanout488 _0679_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_1
Xfanout466 _0683_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_1
Xfanout455 net456 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_1
Xfanout433 net434 vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_1
Xfanout444 net445 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_1
Xfanout499 net500 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_1
Xfanout477 net481 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_1
Xfanout51 net52 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout73 net76 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
Xfanout62 _0123_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout84 _0252_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout95 _0241_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1090_ net333 net197 net72 _0395_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__or4_2
X_0943_ net485 net393 net387 net478 vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0874_ net507 net342 net335 net514 vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1288_ _0096_ _0106_ _0161_ _0175_ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_38_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1357_ _0155_ net156 net122 _0645_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout241 _0109_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_1
Xfanout252 _0095_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__buf_1
Xfanout263 _0086_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout230 _0121_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
Xfanout274 net275 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_1
Xfanout296 net297 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_1
Xfanout285 net286 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__buf_1
XFILLER_0_12_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1211_ net137 net132 vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__or2_1
X_1142_ _0040_ _0200_ _0381_ _0416_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1073_ net94 net92 _0244_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__or3_1
X_0857_ _0167_ net165 vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0926_ net102 net98 net97 vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__or3_1
XFILLER_0_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold27 net24 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ clknet_2_3__leaf_clk0 _0027_ vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__dfxtp_1
Xhold16 net12 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__dlygate4sd3_1
X_0788_ net566 net560 net580 net573 vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__and4b_1
XFILLER_0_38_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0711_ net603 net589 net597 net612 vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__nor4b_1
X_1125_ net139 net125 vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1056_ net121 net119 net116 vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__or3_1
Xoutput17 net17 vssd1 vssd1 vccd1 vccd1 dout0[16] sky130_fd_sc_hd__clkbuf_4
Xoutput39 net39 vssd1 vssd1 vccd1 vccd1 dout0[7] sky130_fd_sc_hd__buf_2
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 dout0[26] sky130_fd_sc_hd__buf_2
X_0909_ net123 net122 vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Left_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1039_ net113 net104 vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__or2_1
X_1108_ net205 net186 net105 net78 vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1390_ clknet_2_2__leaf_clk0 _0008_ vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout604 net605 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_1
Xfanout615 addr0_reg\[0\] vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0890_ net342 net335 net489 vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__o21ba_1
X_1373_ _0247_ _0278_ _0660_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout434 net435 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_1
Xfanout456 _0688_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_1
Xfanout401 net402 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__clkbuf_1
Xfanout412 net413 vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_1
Xfanout423 net424 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_1
Xfanout445 net446 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_18_Left_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout478 net480 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_1
Xfanout489 _0675_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_1
Xfanout467 net468 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_1
Xfanout74 net76 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__buf_1
Xfanout52 net55 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout63 _0110_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_1
Xfanout85 _0251_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__buf_1
Xfanout96 _0236_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__buf_1
XFILLER_0_51_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0873_ net439 net344 net338 net432 vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__a22o_1
X_0942_ net88 net87 net85 net83 vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1287_ _0191_ _0488_ _0578_ _0579_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__or4_1
X_1356_ net310 net309 net152 net146 vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_46_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout253 _0095_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_1
Xfanout286 _0063_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_1
Xfanout264 _0085_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_1
Xfanout242 net243 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_1
Xfanout231 _0120_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_3_Left_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout220 net222 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_1
Xfanout275 _0076_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_1
Xfanout297 net298 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_1
XFILLER_0_49_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1210_ net550 net622 net50 _0508_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__a22o_1
X_1072_ net277 net268 net157 net154 vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__or4_1
X_1141_ net286 net283 vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0856_ net528 net355 net348 net540 vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0925_ net99 net96 vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0787_ net570 net577 net558 net565 vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__nor4b_1
Xhold28 net23 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_45_Left_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1408_ clknet_2_1__leaf_clk0 _0026_ vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__dfxtp_1
Xhold17 net16 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__dlygate4sd3_1
X_1339_ net304 net294 net290 net230 vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_49_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0710_ net603 net612 net589 net597 vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1055_ net122 net118 vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__or2_1
X_1124_ _0032_ _0036_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 dout0[27] sky130_fd_sc_hd__buf_2
Xoutput18 net18 vssd1 vssd1 vccd1 vccd1 dout0[17] sky130_fd_sc_hd__buf_2
X_0908_ net459 net379 net373 net467 vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__a22o_1
X_0839_ net574 net582 net562 net568 vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__and4_1
XFILLER_0_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Left_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1038_ net192 net81 vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__or2_1
X_1107_ net241 net239 net87 net85 vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Left_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout605 net606 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__buf_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1372_ _0050_ _0158_ net58 _0351_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout479 net480 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_1
Xfanout435 _0035_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__buf_1
Xfanout402 net403 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_1
Xfanout446 net449 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_1
Xfanout413 net414 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_1
Xfanout468 net469 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_1
Xfanout457 _0686_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_1
Xfanout424 net425 vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout64 net65 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_1
Xfanout75 net76 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_1
Xfanout53 net54 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_1
Xfanout86 _0251_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
Xfanout97 _0236_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__buf_1
Xfanout42 net46 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_51_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0941_ net87 net84 vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__or2_1
X_0872_ net580 net560 net566 net573 vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__and4b_1
X_1355_ net306 _0075_ net150 net134 vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_38_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1286_ net311 net307 net195 net193 vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_46_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout210 net211 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_1
Xfanout265 _0085_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_1
Xfanout254 _0094_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout276 net277 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__buf_1
Xfanout221 net222 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_1
Xfanout243 _0108_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_1
Xfanout298 net299 vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_1
Xfanout287 _0062_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_1
Xfanout232 _0120_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_1
XFILLER_0_49_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1140_ net151 net149 net121 net116 vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__or4_2
X_1071_ net319 net315 net230 _0377_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_43_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0924_ net436 net381 net375 net430 vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__a22o_1
X_0786_ _0090_ _0097_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__or2_1
X_0855_ net508 net355 net349 net515 vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold29 net41 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1338_ _0379_ _0431_ _0463_ _0555_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__or4_1
X_1407_ clknet_2_2__leaf_clk0 _0025_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__dfxtp_1
Xhold18 net27 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__dlygate4sd3_1
X_1269_ net553 net646 net53 _0563_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1123_ _0425_ _0426_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__or2_1
X_1054_ net333 net328 net324 vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0907_ net443 net383 net377 net450 vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0769_ _0075_ net272 net271 _0080_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput19 net19 vssd1 vssd1 vccd1 vccd1 dout0[18] sky130_fd_sc_hd__buf_2
X_0838_ net575 net582 net562 net568 vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__nor4_1
XFILLER_0_34_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1106_ net215 net213 net202 vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__or3_1
XFILLER_0_48_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1037_ _0171_ _0345_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout606 addr0_reg\[1\] vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1371_ _0113_ _0169_ _0254_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout447 net448 vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__buf_1
Xfanout458 _0686_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__buf_1
Xfanout403 net404 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_1
Xfanout436 net438 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_1
Xfanout425 net428 vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_1
Xfanout414 _0067_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_1
Xfanout469 net474 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout87 _0249_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_1
Xfanout65 net66 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
Xfanout54 net55 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__buf_1
XFILLER_0_36_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout76 _0260_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__buf_2
Xfanout43 net45 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_1
Xfanout98 net99 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__buf_1
XFILLER_0_35_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0940_ net477 net407 net398 net484 vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__a22o_1
X_0871_ _0158_ _0164_ _0171_ _0182_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1354_ _0409_ _0425_ _0553_ _0641_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__or4_1
X_1285_ net330 net303 net214 vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_46_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout211 _0134_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_1
XFILLER_0_41_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout200 net201 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_1
Xfanout222 _0126_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_2
Xfanout233 _0119_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_1
Xfanout277 _0072_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__buf_1
Xfanout266 _0084_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_1
Xfanout255 _0094_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout288 _0057_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__buf_1
Xfanout244 _0105_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_1
Xfanout299 _0046_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__buf_1
XFILLER_0_24_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1070_ net306 net297 net177 net175 vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_43_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0923_ net504 net382 net376 net511 vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__a22o_1
X_0854_ net494 net360 net354 net502 vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0785_ net258 net256 net254 net252 vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__or4_1
X_1268_ _0556_ _0560_ _0562_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__or3_1
X_1406_ clknet_2_3__leaf_clk0 _0024_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__dfxtp_1
Xhold19 net25 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__dlygate4sd3_1
X_1337_ _0565_ _0622_ _0623_ _0625_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__or4_1
X_1199_ net547 net637 net47 _0498_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1122_ net89 _0249_ _0252_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1053_ net242 _0114_ _0359_ _0360_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0906_ _0183_ _0193_ _0216_ _0217_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0837_ net197 net196 net193 net191 vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0768_ net270 net269 vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0699_ net530 net514 net507 net519 vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1105_ net295 net287 vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1036_ net211 net161 net142 net100 vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout607 net609 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1019_ _0327_ _0328_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1370_ net551 net635 net51 _0659_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout404 net405 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_1
Xfanout448 net449 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_1
Xfanout426 net428 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__buf_1
Xfanout459 net460 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout437 net438 vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_1
Xfanout415 net416 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_1
Xfanout55 net56 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout44 net45 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
Xfanout66 _0263_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__buf_1
Xfanout88 _0248_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__buf_1
Xfanout77 _0257_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__buf_1
Xfanout99 net100 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0870_ net163 net159 _0176_ net154 vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__or4_1
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1422_ net34 vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_50_Left_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1284_ _0337_ _0376_ _0519_ _0566_ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__or4_1
X_1353_ _0032_ _0128_ _0352_ _0404_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_46_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0999_ _0048_ _0089_ _0307_ _0308_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout256 _0092_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_2
Xfanout234 net235 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_1
Xfanout245 _0105_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_1
Xfanout212 _0132_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_1
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout223 _0125_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_1
Xfanout201 _0141_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
Xfanout289 _0057_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_1
Xfanout278 _0071_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_1
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout267 _0084_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_1
XFILLER_0_24_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0853_ net439 net358 net352 net433 vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__a22o_1
X_0922_ net523 net379 net373 net535 vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0784_ net254 net253 vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__or2_1
X_1405_ clknet_2_2__leaf_clk0 _0023_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__dfxtp_1
X_1267_ _0172_ _0473_ _0552_ _0561_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__or4_1
Xinput1 addr0[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
X_1198_ _0380_ _0401_ _0495_ _0497_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__or4_1
X_1336_ _0031_ _0224_ _0269_ _0624_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1052_ net61 _0175_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__or2_1
X_1121_ net250 net249 net244 vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_31_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0905_ _0201_ _0208_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__or2_1
X_0767_ net426 net402 net458 vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__o21ba_1
X_0836_ net198 net194 vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0698_ net607 net593 net587 net601 vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_11_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1319_ net554 net643 net54 _0609_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_50 _0255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1104_ net101 net95 net93 net91 vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__or4_1
X_1035_ _0088_ net243 net101 _0343_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__or4_2
XFILLER_0_17_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0819_ net495 net368 net362 net498 vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout608 net609 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1018_ net74 net71 net66 vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__or3_2
XFILLER_0_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout427 net428 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_1
Xfanout438 net442 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_1
Xfanout416 net417 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_1
Xfanout405 _0068_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__clkbuf_1
Xfanout449 _0689_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout67 net69 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__buf_1
Xfanout56 net57 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_1
Xfanout89 _0248_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__buf_1
Xfanout78 _0257_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
Xfanout45 net46 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_24_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1421_ clknet_2_3__leaf_clk0 net9 vssd1 vssd1 vccd1 vccd1 cs0_reg sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1352_ net325 net171 net169 vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__or3_1
X_1283_ net543 net636 net43 _0576_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_46_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0998_ _0041_ _0169_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout213 net214 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_1
Xfanout202 _0140_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_1
Xfanout257 _0092_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_1
Xfanout268 _0079_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_1
Xfanout279 _0070_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__buf_1
Xfanout224 _0125_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_1
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout235 _0119_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_1
Xfanout246 _0104_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_1
XFILLER_0_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_39_Left_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0921_ net492 net382 net378 net500 vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_23_Left_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0852_ net181 net179 net177 net175 vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__or4_2
X_0783_ net515 net396 net390 net508 vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__a22o_1
X_1404_ clknet_2_1__leaf_clk0 _0022_ vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__dfxtp_1
X_1335_ net258 net235 vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__or2_1
Xinput2 addr0[1] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_1266_ net185 _0181_ _0189_ net111 vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__or4_1
X_1197_ _0340_ _0360_ _0476_ _0496_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1051_ net185 net183 net114 net112 vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__or4_2
X_1120_ net553 net627 net53 _0424_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__a22o_1
X_0904_ _0214_ _0215_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0835_ net194 net191 vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__or2_1
X_0697_ net607 net585 net595 net601 vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__and4bb_1
X_0766_ net473 net410 net401 net465 vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1318_ _0601_ _0607_ _0608_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__or3_1
X_1249_ _0535_ _0538_ _0541_ _0544_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__or4_1
XANTENNA_51 _0504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_40 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1103_ net542 net616 net42 _0408_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__a22o_1
X_1034_ net294 net292 net246 net120 vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_26_Left_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0818_ net62 _0129_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__or2_1
X_0749_ net295 net292 net290 net288 vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_10_Left_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout609 net610 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1017_ net258 net256 net252 vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout439 net440 vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_1
Xfanout428 _0052_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__buf_1
Xfanout417 net418 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_1
Xfanout406 net408 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout68 net69 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
Xfanout57 _0276_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__buf_1
Xfanout79 net80 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__buf_1
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout46 net47 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_24_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1351_ net544 net617 net44 _0640_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__a22o_1
X_1420_ clknet_2_0__leaf_clk0 net8 vssd1 vssd1 vccd1 vccd1 addr0_reg\[7\] sky130_fd_sc_hd__dfxtp_1
X_1282_ _0428_ _0565_ _0566_ _0575_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_46_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0997_ net195 net191 net72 net67 vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_1
Xfanout269 _0079_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_1
Xfanout258 _0091_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout247 _0104_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_1
Xfanout225 net227 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout214 _0132_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_2
Xfanout236 _0118_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0920_ net114 net111 net109 net105 vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_43_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0851_ net540 net355 net348 net528 vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__a22o_1
X_0782_ net392 net386 net489 vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1403_ clknet_2_3__leaf_clk0 _0021_ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__dfxtp_1
X_1265_ _0135_ _0557_ _0558_ _0559_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__or4_1
X_1334_ _0358_ _0393_ _0579_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput3 addr0[2] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1196_ _0487_ _0490_ _0491_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_40_Left_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1050_ net305 net215 vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__or2_1
X_0834_ net470 net427 net420 net462 vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0903_ net128 net124 vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_47_Left_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0696_ net538 net531 net526 net518 vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__a22o_1
X_0765_ net453 net406 net398 net446 vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__a22o_1
X_1317_ net58 _0217_ _0277_ _0600_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__or4_1
X_1248_ _0327_ _0432_ _0542_ _0543_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1179_ _0230_ _0259_ _0476_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_41 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_30 _0676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1102_ _0401_ _0405_ _0407_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__or3_1
X_1033_ _0337_ _0338_ _0341_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__or3_1
X_0817_ net226 net224 net221 net219 vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__or4_1
X_0748_ net295 net292 net288 vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1016_ net259 net252 vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout407 net408 vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_1
Xfanout429 net431 vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_1
Xfanout418 net421 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout69 _0262_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__buf_1
Xfanout58 _0193_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_1
XFILLER_0_36_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout47 net57 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1350_ _0487_ _0634_ _0635_ _0639_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__or4_1
X_1281_ _0569_ _0570_ _0572_ _0574_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0996_ net282 net268 net180 net132 vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout204 _0140_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_2
Xfanout259 _0091_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout237 _0118_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_1
Xfanout248 _0102_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_1
Xfanout215 _0131_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_1
Xfanout226 net227 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_37_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0850_ net498 net360 net354 net495 vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__a22o_1
X_1402_ clknet_2_1__leaf_clk0 _0020_ vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__dfxtp_1
X_0781_ net258 net256 vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1333_ _0253_ net74 net66 _0621_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__or4_2
XFILLER_0_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 addr0[3] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_1264_ _0031_ _0049_ _0204_ _0282_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1195_ _0047_ _0149_ _0493_ _0494_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0979_ net311 net98 net94 _0290_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout590 net591 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_1
X_0902_ net131 net127 vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0833_ net451 net423 net416 net444 vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0695_ net570 net577 net558 net564 vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__and4bb_1
X_0764_ net484 net408 net399 net477 vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1247_ net279 net276 net90 vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__or3_1
X_1316_ _0474_ _0604_ _0605_ _0606_ vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1178_ _0066_ _0284_ _0477_ _0478_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__or4_1
XANTENNA_20 _0249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_31 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_53 _0467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_42 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1032_ net254 _0326_ _0340_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__or3_1
X_1101_ _0394_ _0396_ _0406_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0747_ net293 net289 vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__or2_1
X_0816_ net225 net224 net218 vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1015_ _0322_ _0323_ _0324_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__or3_1
XFILLER_0_48_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout419 net420 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_1
Xfanout408 net414 vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_1
Xfanout48 net49 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_1
XFILLER_0_44_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout59 _0258_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_29_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1280_ _0158_ _0323_ _0333_ _0573_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0995_ _0243_ _0246_ _0303_ _0305_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout216 net217 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__clkbuf_1
Xfanout205 _0139_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_1
Xfanout238 net239 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__buf_1
Xfanout227 _0124_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout249 _0102_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0780_ net539 net396 net390 net527 vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1401_ clknet_2_2__leaf_clk0 _0019_ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__dfxtp_1
X_1332_ net189 net182 net173 net164 vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__or4_1
X_1263_ net269 net100 _0250_ net79 vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__or4_1
X_1194_ _0103_ net234 _0488_ _0489_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__or4_1
Xinput5 addr0[4] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0978_ net333 net288 net148 net125 vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_40_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout591 net592 vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_1
Xfanout580 net583 vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_31_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0901_ net127 net124 vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__or2_1
X_0763_ net280 _0070_ net278 net276 vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__or4_2
X_0832_ net483 net425 net418 net476 vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__a22o_1
X_0694_ net600 net593 net584 net608 vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__and4bb_1
X_1315_ _0047_ _0148_ _0169_ _0363_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__or4_1
X_1246_ net209 net188 net158 net144 vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__or4_1
X_1177_ _0448_ _0473_ _0474_ _0475_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_43 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _0249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 _0189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1031_ net273 _0077_ net270 vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1100_ _0200_ _0307_ _0353_ _0404_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__or4_1
X_0746_ net291 net289 vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0815_ net537 net370 net364 net525 vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1229_ net61 _0190_ net138 net135 vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_2__f_clk0 clknet_0_clk0 vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1014_ net212 net202 net201 net82 vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_14_Left_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap385 _0099_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0729_ net312 net307 vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout409 net410 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__buf_1
Xfanout49 net56 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0994_ net240 net238 _0112_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout206 _0138_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_1
Xfanout228 net229 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_1
Xfanout239 _0111_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_2
Xfanout217 _0131_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_49_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_17_Left_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1331_ net548 net642 net48 _0620_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__a22o_1
X_1400_ clknet_2_2__leaf_clk0 _0018_ vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__dfxtp_1
X_1262_ _0040_ _0201_ _0362_ _0447_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__or4_1
X_1193_ net285 _0288_ _0353_ _0492_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__or4_1
Xinput6 addr0[5] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0977_ _0285_ _0286_ _0287_ _0288_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__or4_1
XFILLER_0_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Left_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout592 addr0_reg\[3\] vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_1
Xfanout570 net571 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__buf_1
Xfanout581 net583 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0900_ net368 net336 net457 vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__o21ba_1
X_0831_ net419 net393 net458 vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_36_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0762_ net281 net279 net276 vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__or3_2
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0693_ net558 net564 net570 net577 vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1314_ _0114_ net227 net224 _0339_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1245_ _0465_ _0476_ _0488_ _0539_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1176_ _0189_ _0237_ _0246_ _0280_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__or4_1
XANTENNA_22 _0252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_33 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_44_Left_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_11 _0192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1030_ net272 net270 vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__or2_1
X_0814_ net370 net364 net490 vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_24_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0745_ net512 net424 net417 net505 vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__a22o_1
X_1228_ _0523_ _0524_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1159_ _0098_ _0231_ _0459_ _0460_ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1013_ net159 net157 _0209_ net126 vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_29_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0728_ _0037_ net309 net308 vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__or3_2
XFILLER_0_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0993_ net240 net239 vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout207 _0138_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_1
Xfanout229 net230 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout218 _0127_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_1
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1330_ _0230_ _0588_ _0616_ _0619_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__or4_1
X_1261_ _0464_ _0553_ _0554_ _0555_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__or4_1
X_1192_ net291 net281 _0162_ net146 vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__or4_1
Xinput7 addr0[6] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0976_ net243 net240 net238 vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__or3_1
XFILLER_0_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout560 net563 vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_48_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout593 net594 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_1
Xfanout571 net572 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_1
Xfanout582 net583 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__buf_1
X_0830_ net206 net205 net202 net199 vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0761_ _0071_ net277 vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__or2_1
X_0692_ net584 net594 net600 net607 vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__and4b_1
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1244_ net265 net261 net129 _0210_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__or4_1
X_1313_ _0142_ _0287_ _0602_ _0603_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__or4_1
X_1175_ net75 net68 net64 vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__or3_1
XANTENNA_34 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _0281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0959_ _0081_ _0115_ _0130_ _0247_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__or4_1
XANTENNA_12 _0201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_45 clknet_2_1__leaf_clk0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout390 net391 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0813_ net499 net369 net363 net491 vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0744_ net422 net415 net490 vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__o21ba_1
X_1227_ net289 net111 net104 net100 vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__or4_1
X_1158_ net280 net91 vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1089_ net275 net150 net90 net77 vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Left_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1012_ _0133_ net206 net205 vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0727_ net521 net499 net491 net533 vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0992_ _0059_ _0073_ _0302_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout219 _0127_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_1
Xfanout208 _0137_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_1
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1260_ net131 _0215_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__or2_1
X_1191_ net213 net200 net171 net164 vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__or4_1
Xinput8 addr0[7] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0975_ net315 net313 net107 net106 vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__or4_1
X_1389_ clknet_2_3__leaf_clk0 _0007_ vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout550 net552 vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__buf_1
Xfanout583 addr0_reg\[4\] vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__buf_1
Xfanout572 net576 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_1
Xfanout561 net563 vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_1
Xfanout594 net595 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__clkbuf_1
X_0760_ net509 net411 net402 net516 vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0691_ cs0_reg vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1243_ net273 _0078_ net268 vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__or3_1
X_1312_ net281 net279 net228 net84 vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__or4_1
X_1174_ net243 net116 vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__or2_1
XANTENNA_13 _0201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_46 _0060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0889_ net145 net144 net141 net140 vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__or4_2
XFILLER_0_6_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_35 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_24 _0281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0958_ net287 net285 net282 net208 vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout391 _0083_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_1
Xfanout380 net381 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_1
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0743_ net499 net422 net415 net492 vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__a22o_1
X_0812_ net511 net369 net363 net505 vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__a22o_1
X_1226_ net229 net173 _0197_ net128 vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__or4_1
X_1157_ net312 net310 vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1088_ net227 net220 _0392_ _0393_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1011_ _0050_ _0318_ _0319_ _0320_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0726_ net521 net511 net504 net533 vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1209_ _0283_ _0306_ _0499_ _0507_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__or4_1
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0709_ net532 net482 net475 net520 vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_23_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0991_ _0056_ net206 net205 vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout209 _0137_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__buf_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput9 cs0 vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1190_ net264 net261 net256 net253 vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_42_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0974_ _0041_ net59 vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1388_ clknet_2_2__leaf_clk0 _0006_ vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__clkbuf_1
Xfanout551 net552 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_1
Xfanout540 net541 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_1
Xfanout584 net586 vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_1
Xfanout573 net576 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_1
Xfanout562 net563 vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1311_ net208 net178 net170 _0244_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__or4_1
X_1242_ net103 net99 _0392_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__or3_1
X_1173_ _0038_ net191 vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_36 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_14 _0201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 _0094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 _0329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0888_ net144 net141 net140 vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0957_ net282 net208 vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout392 net397 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_1
Xfanout381 net382 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_1
Xfanout370 net371 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_1
X_0811_ net236 net235 net231 net230 vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__or4_2
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0742_ net535 net422 net415 net523 vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__a22o_1
X_1156_ net549 net644 net49 _0458_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__a22o_1
X_1225_ net94 net91 net72 vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__or3_1
X_1087_ net178 net175 vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_50_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1010_ net242 net239 net218 net121 vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__or4_1
X_0725_ net531 net526 net518 net538 vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1208_ _0503_ _0504_ _0505_ _0506_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1139_ net543 net626 net43 _0442_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_9_Left_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1 net38 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0708_ net612 net589 net597 net604 vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__nor4b_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_35_Left_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0990_ _0677_ _0300_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0973_ net61 net207 vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__or2_1
X_1387_ clknet_2_2__leaf_clk0 _0005_ vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout552 net555 vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_1
Xfanout596 net599 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_1
Xfanout541 _0638_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_1
Xfanout585 net586 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_1
Xfanout574 net575 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_1
Xfanout530 net531 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__buf_1
Xfanout563 addr0_reg\[7\] vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__buf_1
XFILLER_0_28_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_38_Left_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1310_ _0677_ _0060_ _0157_ _0490_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__or4_1
X_1241_ net148 _0244_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_22_Left_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1172_ net229 net219 vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_37 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 _0344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 _0212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0956_ _0133_ net211 net81 net77 vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__or4_1
XANTENNA_48 _0108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0887_ _0195_ net141 vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout393 net394 vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_1
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout382 net383 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_1
Xfanout371 net372 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__buf_1
Xfanout360 _0150_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_1
X_0810_ net232 net228 vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0741_ net570 net564 net558 net577 vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__and4bb_1
X_1224_ net308 _0112_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_50_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1155_ _0452_ _0453_ _0457_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__or3_1
X_1086_ net248 net244 vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__or2_1
X_0939_ net465 net410 net403 net473 vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout190 _0152_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_1
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_47 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0724_ net534 net438 net431 net519 vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__a22o_1
X_1207_ _0080_ _0096_ _0122_ net60 vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1138_ _0427_ _0428_ _0440_ _0441_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__or4_1
X_1069_ _0060_ _0238_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 net26 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_17_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0707_ net612 net590 net599 net603 vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__and4b_1
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0972_ net145 _0198_ _0204_ net134 vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1386_ clknet_2_2__leaf_clk0 _0004_ vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout520 net522 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__buf_1
XFILLER_0_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout542 net546 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout531 net534 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__buf_1
Xfanout553 net554 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__buf_1
Xfanout597 net598 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__buf_1
Xfanout586 net587 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_1
Xfanout564 net565 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_1
Xfanout575 net576 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_1
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1171_ net548 net640 net48 _0472_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1240_ net330 net177 vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0955_ net217 net214 _0136_ net79 vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__or4_1
XANTENNA_49 _0142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 _0481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0886_ net141 net140 vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_16 _0220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1369_ _0081_ _0414_ _0652_ _0657_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout350 net351 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_1
Xfanout361 net366 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_1
Xfanout383 net385 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_1
Xfanout372 _0116_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_1
Xfanout394 net395 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_1
X_0740_ net579 net559 net565 net572 vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__and4bb_1
X_1154_ _0115_ _0278_ _0454_ _0456_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__or4_1
X_1223_ net296 net82 vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_50_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1085_ net544 net619 net44 _0391_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__a22o_1
X_0938_ net89 net87 vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__or2_1
X_0869_ net159 net154 vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout191 _0146_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__buf_1
Xfanout180 _0159_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_1
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0723_ net605 net614 net591 net598 vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1206_ net74 net70 _0501_ _0502_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__or4_1
X_1137_ net58 _0208_ _0225_ _0232_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1068_ _0064_ net283 net61 _0139_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__or4_2
XFILLER_0_7_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3 net20 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0706_ net334 net332 net327 net324 vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0971_ _0198_ _0204_ net135 vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1385_ clknet_2_2__leaf_clk0 _0003_ vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout554 net555 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_1
Xfanout510 _0670_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__buf_1
Xfanout543 net545 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_1
Xfanout532 net534 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_1
Xfanout565 net569 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_1
Xfanout521 net522 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__buf_1
Xfanout598 net599 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__buf_1
Xfanout587 net588 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_1
Xfanout576 addr0_reg\[5\] vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__buf_1
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1170_ _0375_ _0461_ _0471_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__or3_1
X_0954_ net75 net70 net67 net65 vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__or4_2
XANTENNA_28 _0506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0885_ net464 net345 net338 net472 vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__a22o_1
XANTENNA_39 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_17 _0220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1368_ _0641_ _0654_ _0655_ _0656_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__or4_1
X_1299_ _0090_ _0201_ _0589_ _0590_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_53_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout340 net341 vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__buf_1
Xfanout351 net352 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__buf_1
Xfanout395 net396 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_1
Xfanout373 net374 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_1
Xfanout362 net366 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__buf_1
X_1153_ net280 net279 _0122_ _0455_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__or4_1
X_1084_ _0383_ _0388_ _0390_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__or3_1
X_1222_ _0032_ _0403_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_50_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0868_ net162 net158 vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__or2_1
X_0937_ net448 net409 net400 net455 vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__a22o_1
X_0799_ net513 net406 net398 net506 vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout192 _0146_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_1
Xfanout181 _0159_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout170 _0166_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0722_ net605 net614 net591 net598 vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1136_ _0433_ _0435_ _0437_ _0439_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__or4_1
X_1067_ net542 net645 net42 _0374_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__a22o_1
X_1205_ _0042_ _0238_ _0354_ _0500_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4 net37 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0705_ net331 net327 net324 vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1119_ _0418_ _0420_ _0423_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_0_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Left_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0970_ net216 net203 vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1384_ clknet_2_2__leaf_clk0 _0002_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout555 net556 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_1
Xfanout599 addr0_reg\[2\] vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__buf_1
Xfanout588 net592 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_1
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_1
Xfanout566 net569 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_1
Xfanout533 net534 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_1
Xfanout577 net578 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__buf_1
Xfanout511 net512 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__buf_1
Xfanout500 net501 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_1
Xfanout522 _0666_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__buf_1
XFILLER_0_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_29 _0527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_18 _0228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0953_ net75 net68 vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__or2_1
X_0884_ net478 net345 net338 net485 vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1367_ _0158_ _0240_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1298_ net238 net236 net178 vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__or3_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout352 net353 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_1
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_1
Xfanout330 _0674_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout374 net375 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_1
Xfanout341 _0184_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_1
Xfanout363 net366 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_1
X_1221_ net550 net621 net50 _0518_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1083_ _0375_ _0376_ _0378_ _0389_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__or4_1
X_1152_ net331 net330 net135 net132 vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_50_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0936_ net434 net407 net399 net441 vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__a22o_1
X_0867_ net160 net157 vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__or2_1
X_0798_ net242 net241 vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1419_ clknet_2_0__leaf_clk0 net7 vssd1 vssd1 vccd1 vccd1 addr0_reg\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout182 net183 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_1
Xfanout160 net161 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__buf_1
Xfanout171 net174 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_1
Xfanout193 _0145_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0721_ net322 net318 net316 net314 vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1204_ _0107_ _0402_ _0426_ _0443_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1135_ net59 _0326_ _0438_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__or3_1
X_1066_ _0361_ _0367_ _0373_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0919_ net113 net110 vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 net29 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_29_Left_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0704_ net530 net518 net489 vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1118_ _0301_ _0414_ _0421_ _0422_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__or4_1
X_1049_ net542 net624 net42 _0357_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1383_ clknet_2_1__leaf_clk0 _0001_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout556 net557 vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_1
Xfanout589 net590 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__buf_1
Xfanout545 net546 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout523 net524 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_1
Xfanout578 net579 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_1
Xfanout501 net502 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_16_Left_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout534 _0648_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_1
Xfanout512 net513 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__buf_1
Xfanout567 net569 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_1
XFILLER_0_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0952_ net67 net64 vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_19 _0242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0883_ net432 net344 net339 net439 vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1366_ _0179_ _0264_ _0537_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1297_ net189 net184 net158 vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__or3_1
Xfanout331 _0671_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_2
Xfanout320 net321 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_1
Xfanout353 net354 vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_1
Xfanout397 _0082_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_1
Xfanout386 net391 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_1_Left_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout375 net376 vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_1
Xfanout342 net343 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__buf_1
Xfanout364 net365 vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_1
X_1151_ _0147_ net190 net182 _0449_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__or4_1
X_1220_ _0325_ _0512_ _0517_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_9_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1082_ net325 _0155_ _0231_ net89 vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_50_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0866_ net348 net344 net458 vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__o21ba_1
X_0935_ _0240_ _0243_ _0246_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0797_ net539 net409 net400 net527 vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Left_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1349_ _0359_ _0411_ _0426_ _0637_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1418_ clknet_2_0__leaf_clk0 net6 vssd1 vssd1 vccd1 vccd1 addr0_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout183 _0156_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_1
Xfanout172 net174 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
Xfanout161 _0174_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_1
Xfanout150 _0186_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout194 _0145_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0720_ net323 net318 net316 vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap317 _0687_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__buf_1
XFILLER_0_20_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1203_ net286 net210 net152 net129 vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__or4_1
X_1134_ net333 net326 net266 net264 vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1065_ _0368_ _0369_ _0372_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__or3_1
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0918_ net111 net109 net104 vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__or3_1
X_0849_ net181 net179 vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_1__f_clk0 clknet_0_clk0 vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
Xhold6 net15 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0703_ net600 net607 net593 net584 vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__or4b_1
XFILLER_0_29_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1117_ _0198_ _0392_ _0410_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_0_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1048_ _0342_ _0350_ _0356_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_30_Left_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1382_ clknet_2_1__leaf_clk0 _0000_ vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout502 net503 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__buf_1
Xfanout524 net525 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__buf_1
Xfanout513 net514 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_1
Xfanout557 _0628_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__buf_1
Xfanout546 net547 vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__buf_1
Xfanout535 net536 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__buf_1
Xfanout579 net583 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__clkbuf_1
Xfanout568 net569 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_1
X_0951_ net463 net426 net419 net470 vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0882_ net446 net347 net341 net453 vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1365_ net63 net177 net163 _0653_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__or4_1
X_1296_ net272 net271 net268 vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_53_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout321 _0684_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__buf_1
Xfanout343 net347 vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout365 net366 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__buf_1
Xfanout332 _0671_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_1
Xfanout354 _0151_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__buf_1
Xfanout310 net311 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_1
Xfanout387 net388 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_1
Xfanout376 net378 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_1
Xfanout398 net399 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_1
XFILLER_0_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1150_ _0259_ _0443_ _0446_ _0447_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_9_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1081_ _0384_ _0385_ _0386_ _0387_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__or4_2
XFILLER_0_23_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0865_ net573 net560 net566 net580 vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_15_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0934_ _0244_ net90 vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__or2_2
XFILLER_0_23_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0796_ net413 net404 net489 vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1417_ clknet_2_0__leaf_clk0 net5 vssd1 vssd1 vccd1 vccd1 addr0_reg\[4\] sky130_fd_sc_hd__dfxtp_1
X_1348_ _0048_ _0300_ _0340_ _0636_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__or4_1
X_1279_ net195 _0205_ net119 net95 vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout162 _0173_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__buf_1
Xfanout184 _0154_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_1
Xfanout173 _0165_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_1
Xfanout140 _0197_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout151 _0186_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__buf_1
Xfanout195 net196 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_29_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1202_ net261 net192 vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1064_ _0075_ net62 _0370_ _0371_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__or4_1
X_1133_ _0114_ _0429_ _0436_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0779_ _0672_ net394 net388 net497 vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0917_ net530 net362 net457 vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__o21ba_1
X_0848_ net360 net354 net490 vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_3_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7 net14 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0702_ net530 net498 net495 net519 vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__a22o_1
X_1116_ _0409_ _0411_ _0412_ _0415_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_0_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1047_ _0074_ _0351_ _0352_ _0355_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk0 clk0 vssd1 vssd1 vccd1 vccd1 clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1381_ net554 net641 net54 vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_33_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout503 _0672_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout547 net557 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout536 net537 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__buf_1
Xfanout525 net526 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout514 net517 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__buf_1
Xfanout558 net559 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__buf_1
Xfanout569 addr0_reg\[6\] vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__buf_1
XFILLER_0_36_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0950_ net478 net427 net419 net485 vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__a22o_1
X_0881_ _0190_ _0192_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1364_ net314 _0212_ net70 vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__or3_1
X_1295_ net546 net618 net46 _0587_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout344 net345 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_1
Xfanout388 net389 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_1
Xfanout355 net359 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_1
Xfanout377 _0100_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_1
Xfanout311 _0037_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__buf_1
Xfanout333 _0668_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_2
Xfanout322 _0681_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_1
Xfanout366 _0117_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__buf_1
Xfanout300 net302 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__buf_1
Xfanout399 net405 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_1
XFILLER_0_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1080_ net331 net197 net196 _0305_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0864_ net455 net356 net350 net447 vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__a22o_1
X_0795_ net250 net248 net246 net245 vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__or4_2
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0933_ net468 net383 net377 net460 vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1416_ clknet_2_0__leaf_clk0 net4 vssd1 vssd1 vccd1 vccd1 addr0_reg\[3\] sky130_fd_sc_hd__dfxtp_1
X_1347_ net262 net221 net170 vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1278_ net262 net255 _0410_ _0571_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__or4_1
Xfanout185 _0154_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_1
Xfanout152 _0185_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__buf_1
Xfanout163 _0173_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_1
Xfanout174 _0165_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_1
Xfanout130 net131 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_1
Xfanout141 net142 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_1
Xfanout196 _0144_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_6_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1201_ net297 net271 net123 net115 vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1063_ net170 net137 net101 net94 vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__or4_1
X_1132_ net306 net299 net92 net90 vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__or4_1
XFILLER_0_50_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0916_ net450 net368 net362 net443 vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__a22o_1
X_0847_ net515 net355 net348 net508 vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__a22o_1
X_0778_ net266 net264 net263 net260 vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__or4_1
XFILLER_0_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold8 net31 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0701_ net593 net585 net608 net601 vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__and4b_1
XFILLER_0_20_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1115_ _0208_ _0214_ _0413_ _0419_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_0_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1046_ _0040_ _0333_ _0353_ _0354_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1029_ net302 net251 net244 net112 vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1380_ net553 net623 net53 _0667_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout548 net549 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__buf_1
Xfanout515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__buf_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout526 net529 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout537 net538 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_1
Xfanout559 net563 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_1
Xfanout504 net505 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__buf_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0880_ net152 net146 vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__or2_2
X_1363_ _0208_ _0425_ _0651_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__or3_1
XFILLER_0_53_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1294_ _0577_ _0580_ _0586_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__or3_1
XFILLER_0_53_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Left_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout345 net346 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_1
Xfanout356 net357 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__buf_1
Xfanout389 net390 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__clkbuf_1
Xfanout367 net372 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_1
Xfanout334 _0668_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__buf_1
Xfanout378 _0100_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_1
Xfanout312 _0036_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_1
Xfanout323 _0681_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_1
Xfanout301 net302 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0932_ net451 net381 net375 net444 vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0863_ net162 net160 vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__or2_1
X_0794_ net247 net245 vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1415_ clknet_2_0__leaf_clk0 net3 vssd1 vssd1 vccd1 vccd1 addr0_reg\[2\] sky130_fd_sc_hd__dfxtp_1
X_1346_ _0488_ _0538_ _0568_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__or3_1
X_1277_ net259 net215 net201 net83 vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__or4_1
Xfanout131 _0209_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_1
Xfanout120 _0222_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_5_Left_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout186 net188 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_1
Xfanout142 net143 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_1
Xfanout197 _0143_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout153 _0185_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_1
Xfanout175 _0163_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__buf_1
Xfanout164 net166 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_6_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1200_ _0157_ net181 vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1131_ _0328_ _0398_ _0430_ _0434_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1062_ net290 net246 net193 net125 vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__or4_1
XFILLER_0_50_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0915_ net482 net371 net365 net475 vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__a22o_1
X_0846_ net189 net187 net184 net182 vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__or4_2
X_0777_ net266 net264 net260 vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1329_ _0446_ _0535_ _0554_ _0618_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_3_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold9 net35 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_17_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0700_ net600 net584 net595 net610 vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__and4bb_1
Xwire384 _0099_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1114_ net220 net218 _0192_ _0224_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_0_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1045_ net223 net220 net212 net204 vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0829_ net504 net369 net363 net511 vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1028_ net287 _0243_ net91 _0269_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout549 net556 vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_1
Xfanout527 net529 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__buf_1
Xfanout516 net517 vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_1
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout538 net541 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_1
Xfanout505 net506 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__buf_1
XFILLER_0_8_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1362_ net216 net213 _0232_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__or3_1
X_1293_ _0283_ _0581_ _0583_ _0585_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__buf_1
Xfanout313 net314 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_2
Xfanout357 net358 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_1
Xfanout346 net347 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_1
Xfanout379 net380 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_1
Xfanout335 net337 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_1
Xfanout368 net372 vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_1
Xfanout324 _0676_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_52_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Left_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0862_ net486 net357 net351 net479 vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__a22o_1
X_0931_ net95 net93 vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_21_Left_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0793_ net512 net382 net376 net504 vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1414_ clknet_2_0__leaf_clk0 net2 vssd1 vssd1 vccd1 vccd1 addr0_reg\[1\] sky130_fd_sc_hd__dfxtp_1
X_1345_ _0552_ _0600_ _0632_ _0633_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1276_ net108 net73 _0520_ _0567_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout143 _0196_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_1
Xfanout110 _0228_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_1
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_1
Xfanout165 net166 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_1
Xfanout121 net122 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__buf_1
Xfanout132 net133 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_1
Xfanout187 net188 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_1
Xfanout198 _0143_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_1
Xfanout176 _0163_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__buf_1
XFILLER_0_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1130_ net270 net233 net226 net144 vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__or4_1
X_1061_ _0041_ _0189_ _0358_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__or3_1
X_0845_ _0155_ net183 vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0914_ net468 net369 net363 net460 vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0776_ net263 net260 vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1259_ net257 _0096_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1328_ net322 net304 _0279_ _0617_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1044_ net130 net126 net124 vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__or3_2
X_1113_ _0308_ _0382_ _0416_ _0417_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_0_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0759_ net527 net409 net400 net539 vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0828_ net523 net371 net365 net535 vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1027_ net542 net628 net42 _0336_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout506 net507 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_1
Xfanout539 net541 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__buf_1
Xfanout528 net529 vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_1
Xfanout517 _0669_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1292_ _0170_ _0231_ _0265_ _0584_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1361_ net543 net633 net43 _0650_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout325 net326 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout347 _0177_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__buf_1
Xfanout336 net337 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_1
Xfanout303 _0045_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__buf_1
Xfanout314 _0690_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_2
Xfanout358 net359 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_1
Xfanout369 net372 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__buf_1
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0861_ net470 net356 net350 net462 vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__a22o_1
X_0792_ net500 net384 net376 net491 vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__a22o_1
X_0930_ net406 net377 net457 vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1413_ clknet_2_0__leaf_clk0 net1 vssd1 vssd1 vccd1 vccd1 addr0_reg\[0\] sky130_fd_sc_hd__dfxtp_1
X_1275_ _0074_ _0464_ _0568_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__or3_1
X_1344_ _0685_ _0509_ _0567_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__or3_1
Xfanout111 net112 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_1
Xfanout155 net156 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_1
Xfanout188 _0153_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_1
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_1
Xfanout166 _0168_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_1
Xfanout144 _0195_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_1
Xfanout133 _0206_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_1
Xfanout177 _0162_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_2
Xfanout100 _0235_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout122 _0220_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1060_ _0064_ _0207_ _0239_ net59 vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0844_ net448 net356 net350 net454 vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0775_ net477 net392 net386 net484 vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__a22o_1
X_0913_ net123 _0220_ _0222_ net117 vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1258_ net63 net86 vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__or2_1
X_1189_ net326 net88 net80 net77 vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__or4_1
X_1327_ net326 net310 net303 net266 vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_49_Left_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1043_ net237 net233 net181 net176 vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_0_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1112_ net318 net313 net305 net301 vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0827_ net509 net396 net390 net516 vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__a22o_1
X_0758_ net441 net412 net403 net434 vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1026_ _0321_ _0325_ _0335_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout529 _0658_ vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__buf_1
XFILLER_0_13_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout518 net522 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_1
Xfanout507 net510 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__buf_1
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1009_ net274 net196 net175 net166 vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1360_ _0642_ _0643_ _0649_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__or3_1
X_1291_ net190 net186 vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout348 net349 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_1
Xfanout359 net360 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_1
Xfanout326 _0676_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__clkbuf_2
Xfanout304 _0044_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__buf_1
Xfanout337 net341 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_1
Xfanout315 _0687_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_1
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0860_ _0164_ _0171_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__or2_1
X_0791_ net250 net249 vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1412_ clknet_2_3__leaf_clk0 _0030_ vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__dfxtp_1
X_1343_ _0041_ _0059_ net63 _0215_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__or4_1
X_1274_ net327 net324 net151 net147 vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0989_ net160 net157 net154 vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout156 _0178_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout189 net190 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__buf_1
Xfanout167 _0167_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_2
Xfanout145 _0194_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_1
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout123 _0219_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__buf_1
Xfanout112 _0227_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_2
Xfanout134 net135 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_1
Xfanout101 _0234_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__buf_1
Xfanout178 _0160_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_1
XFILLER_0_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0912_ net119 net116 vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__or2_1
X_0843_ net188 net184 vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__or2_2
XFILLER_0_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0774_ net461 net392 net386 net469 vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__a22o_1
X_1326_ _0610_ _0611_ _0613_ _0615_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__or4_1
X_1257_ net209 _0149_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__or2_1
X_1188_ net231 net225 net223 vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__or3_2
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1111_ net171 net168 net164 vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_0_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1042_ net334 net332 net328 vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0826_ net527 net394 net388 net539 vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__a22o_1
X_0757_ net496 net409 net400 net503 vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__a22o_1
X_1309_ net278 _0522_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1025_ _0329_ _0330_ _0331_ _0334_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__or4_1
X_0809_ net429 net367 net361 net437 vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_1 _0056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout508 net509 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__buf_1
Xfanout519 net522 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__buf_1
XFILLER_0_44_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1008_ _0685_ net108 net106 _0317_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1290_ _0110_ net234 _0219_ _0582_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout338 net340 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__buf_1
Xfanout349 net353 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_1
Xfanout305 net306 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__buf_1
Xfanout327 net329 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_1
Xfanout316 net317 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0790_ net535 net380 net374 net523 vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__a22o_1
X_1411_ clknet_2_3__leaf_clk0 _0029_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__dfxtp_1
X_1342_ net547 net634 net47 _0631_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__a22o_1
X_1273_ net123 net117 vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0988_ net313 _0031_ _0221_ net119 vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__or4_2
Xfanout113 net115 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__buf_1
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout102 _0234_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
Xfanout157 net158 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__buf_1
Xfanout124 net125 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_1
Xfanout179 _0160_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_1
Xfanout168 _0166_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout135 _0205_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_2
Xfanout146 _0188_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_1
XFILLER_0_49_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Left_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0842_ net462 net356 net350 net470 vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0911_ net475 net379 net373 net482 vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__a22o_1
X_0773_ net433 net393 net387 net440 vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1256_ net548 net638 net48 _0551_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__a22o_1
X_1325_ net233 net232 net150 _0614_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__or4_1
X_1187_ net180 net178 _0194_ net142 vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1110_ net278 net276 net180 net176 vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__or4_1
X_1041_ net58 _0344_ _0346_ _0349_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0825_ net439 net426 net420 net432 vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0756_ net581 net567 net561 net574 vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__and4bb_1
X_1308_ net548 net639 net48 _0599_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__a22o_1
X_1239_ net321 net313 net92 _0534_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1024_ _0677_ net62 _0332_ _0333_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_44_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Left_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0808_ net444 net367 net361 net451 vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_12_Left_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0739_ _0678_ _0033_ _0042_ _0050_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_2 _0057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout509 net510 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_1
X_1007_ net288 net225 net103 net98 vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout339 net340 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_1
Xfanout306 _0043_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_1
Xfanout328 net329 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1410_ clknet_2_3__leaf_clk0 _0028_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1272_ _0322_ _0539_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1341_ _0626_ _0627_ _0630_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__or3_1
X_0987_ net629 net547 net47 _0298_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__a22o_1
Xfanout114 net115 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_1
Xfanout136 _0203_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout147 _0188_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_1
Xfanout103 _0233_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__buf_1
Xfanout125 _0212_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout169 net170 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_1
Xfanout158 _0176_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_1
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0841_ net478 net357 net351 net485 vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0910_ net429 net383 net377 net436 vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__a22o_1
X_0772_ net446 net392 net386 net453 vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1255_ _0545_ _0550_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1186_ net550 net631 net50 _0486_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__a22o_1
X_1324_ net277 net168 net164 vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Left_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1040_ net70 net64 _0347_ _0348_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0824_ net458 net389 vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0755_ net574 net561 net567 net581 vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__and4bb_1
X_1169_ _0466_ _0468_ _0469_ _0470_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__or4_1
X_1307_ _0592_ _0595_ _0598_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__or3_1
X_1238_ net294 net292 net290 vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1023_ net145 net139 net136 vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__or3_2
XFILLER_0_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0807_ net459 net371 net365 net467 vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0738_ net305 _0044_ net300 net297 vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__or4_1
XFILLER_0_21_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_3 _0060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1006_ net550 net630 net50 _0316_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 dout0[8] sky130_fd_sc_hd__buf_2
XFILLER_0_53_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout307 net308 vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_1
Xfanout329 net330 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_1
Xfanout318 net319 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_1
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1340_ _0089_ _0330_ _0338_ _0629_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1271_ net242 _0114_ _0564_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0986_ _0289_ _0293_ _0297_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__or3_1
Xfanout159 net160 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_1
Xfanout104 net106 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__buf_1
Xfanout126 _0211_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_1
Xfanout137 net138 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout148 _0187_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_1
Xfanout115 _0226_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0840_ net432 net359 net349 net440 vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0771_ net575 net581 net567 net561 vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__nor4b_1
X_1323_ _0501_ _0584_ _0612_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__or3_1
X_1254_ _0537_ _0546_ _0548_ _0549_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__or4_1
X_1185_ _0479_ _0480_ _0485_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_19_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0969_ net278 net272 vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout490 _0675_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_1
XFILLER_0_28_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0823_ _0133_ net210 vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0754_ _0061_ _0064_ net282 vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1306_ _0277_ _0285_ _0331_ _0597_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__or4_1
X_1168_ _0058_ _0161_ _0213_ _0282_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__or4_1
X_1099_ _0397_ _0402_ _0403_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__or3_1
X_1237_ net543 net632 net43 _0533_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk0 clknet_0_clk0 vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_40_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1022_ net312 net284 net267 net147 vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_44_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0806_ net476 net367 net361 net483 vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0737_ net305 net300 vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _0105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1005_ _0306_ _0313_ _0315_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__or3_1
XFILLER_0_29_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 dout0[9] sky130_fd_sc_hd__clkbuf_4
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 dout0[28] sky130_fd_sc_hd__buf_2
XFILLER_0_53_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout308 _0039_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__buf_1
Xfanout319 net320 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_1
.ends

