assign table_[0] = 32'h00000000;
assign table_[1] = 32'h0192155f;
assign table_[2] = 32'h0323ecbe;
assign table_[3] = 32'h04b54825;
assign table_[4] = 32'h0645e9af;
assign table_[5] = 32'h07d59396;
assign table_[6] = 32'h09640837;
assign table_[7] = 32'h0af10a22;
assign table_[8] = 32'h0c7c5c1e;
assign table_[9] = 32'h0e05c135;
assign table_[10] = 32'h0f8cfcbe;
assign table_[11] = 32'h1111d263;
assign table_[12] = 32'h1294062f;
assign table_[13] = 32'h14135c94;
assign table_[14] = 32'h158f9a76;
assign table_[15] = 32'h17088531;
assign table_[16] = 32'h187de2a7;
assign table_[17] = 32'h19ef7944;
assign table_[18] = 32'h1b5d100a;
assign table_[19] = 32'h1cc66e99;
assign table_[20] = 32'h1e2b5d38;
assign table_[21] = 32'h1f8ba4dc;
assign table_[22] = 32'h20e70f32;
assign table_[23] = 32'h223d66a8;
assign table_[24] = 32'h238e7673;
assign table_[25] = 32'h24da0a9a;
assign table_[26] = 32'h261feffa;
assign table_[27] = 32'h275ff452;
assign table_[28] = 32'h2899e64a;
assign table_[29] = 32'h29cd9578;
assign table_[30] = 32'h2afad269;
assign table_[31] = 32'h2c216eaa;
assign table_[32] = 32'h2d413ccd;
assign table_[33] = 32'h2e5a1070;
assign table_[34] = 32'h2f6bbe45;
assign table_[35] = 32'h30761c18;
assign table_[36] = 32'h317900d6;
assign table_[37] = 32'h32744493;
assign table_[38] = 32'h3367c090;
assign table_[39] = 32'h34534f41;
assign table_[40] = 32'h3536cc52;
assign table_[41] = 32'h361214b0;
assign table_[42] = 32'h36e5068a;
assign table_[43] = 32'h37af8159;
assign table_[44] = 32'h387165e3;
assign table_[45] = 32'h392a9642;
assign table_[46] = 32'h39daf5e8;
assign table_[47] = 32'h3a8269a3;
assign table_[48] = 32'h3b20d79e;
assign table_[49] = 32'h3bb6276e;
assign table_[50] = 32'h3c42420a;
assign table_[51] = 32'h3cc511d9;
assign table_[52] = 32'h3d3e82ae;
assign table_[53] = 32'h3dae81cf;
assign table_[54] = 32'h3e14fdf7;
assign table_[55] = 32'h3e71e759;
assign table_[56] = 32'h3ec52fa0;
assign table_[57] = 32'h3f0ec9f5;
assign table_[58] = 32'h3f4eaafe;
assign table_[59] = 32'h3f84c8e2;
assign table_[60] = 32'h3fb11b48;
assign table_[61] = 32'h3fd39b5a;
assign table_[62] = 32'h3fec43c7;
assign table_[63] = 32'h3ffb10c1;
assign table_[64] = 32'h40000000;
assign table_[65] = 32'h3ffb10c1;
assign table_[66] = 32'h3fec43c7;
assign table_[67] = 32'h3fd39b5a;
assign table_[68] = 32'h3fb11b48;
assign table_[69] = 32'h3f84c8e2;
assign table_[70] = 32'h3f4eaafe;
assign table_[71] = 32'h3f0ec9f5;
assign table_[72] = 32'h3ec52fa0;
assign table_[73] = 32'h3e71e759;
assign table_[74] = 32'h3e14fdf7;
assign table_[75] = 32'h3dae81cf;
assign table_[76] = 32'h3d3e82ae;
assign table_[77] = 32'h3cc511d9;
assign table_[78] = 32'h3c42420a;
assign table_[79] = 32'h3bb6276e;
assign table_[80] = 32'h3b20d79e;
assign table_[81] = 32'h3a8269a3;
assign table_[82] = 32'h39daf5e8;
assign table_[83] = 32'h392a9642;
assign table_[84] = 32'h387165e3;
assign table_[85] = 32'h37af8159;
assign table_[86] = 32'h36e5068a;
assign table_[87] = 32'h361214b0;
assign table_[88] = 32'h3536cc52;
assign table_[89] = 32'h34534f41;
assign table_[90] = 32'h3367c090;
assign table_[91] = 32'h32744493;
assign table_[92] = 32'h317900d6;
assign table_[93] = 32'h30761c18;
assign table_[94] = 32'h2f6bbe45;
assign table_[95] = 32'h2e5a1070;
assign table_[96] = 32'h2d413ccd;
assign table_[97] = 32'h2c216eaa;
assign table_[98] = 32'h2afad269;
assign table_[99] = 32'h29cd9578;
assign table_[100] = 32'h2899e64a;
assign table_[101] = 32'h275ff452;
assign table_[102] = 32'h261feffa;
assign table_[103] = 32'h24da0a9a;
assign table_[104] = 32'h238e7673;
assign table_[105] = 32'h223d66a8;
assign table_[106] = 32'h20e70f32;
assign table_[107] = 32'h1f8ba4dc;
assign table_[108] = 32'h1e2b5d38;
assign table_[109] = 32'h1cc66e99;
assign table_[110] = 32'h1b5d100a;
assign table_[111] = 32'h19ef7944;
assign table_[112] = 32'h187de2a7;
assign table_[113] = 32'h17088531;
assign table_[114] = 32'h158f9a76;
assign table_[115] = 32'h14135c94;
assign table_[116] = 32'h1294062f;
assign table_[117] = 32'h1111d263;
assign table_[118] = 32'h0f8cfcbe;
assign table_[119] = 32'h0e05c135;
assign table_[120] = 32'h0c7c5c1e;
assign table_[121] = 32'h0af10a22;
assign table_[122] = 32'h09640837;
assign table_[123] = 32'h07d59396;
assign table_[124] = 32'h0645e9af;
assign table_[125] = 32'h04b54825;
assign table_[126] = 32'h0323ecbe;
assign table_[127] = 32'h0192155f;
assign table_[128] = 32'h00000000;
assign table_[129] = 32'hfe6deaa1;
assign table_[130] = 32'hfcdc1342;
assign table_[131] = 32'hfb4ab7db;
assign table_[132] = 32'hf9ba1651;
assign table_[133] = 32'hf82a6c6a;
assign table_[134] = 32'hf69bf7c9;
assign table_[135] = 32'hf50ef5de;
assign table_[136] = 32'hf383a3e2;
assign table_[137] = 32'hf1fa3ecb;
assign table_[138] = 32'hf0730342;
assign table_[139] = 32'heeee2d9d;
assign table_[140] = 32'hed6bf9d1;
assign table_[141] = 32'hebeca36c;
assign table_[142] = 32'hea70658a;
assign table_[143] = 32'he8f77acf;
assign table_[144] = 32'he7821d59;
assign table_[145] = 32'he61086bc;
assign table_[146] = 32'he4a2eff6;
assign table_[147] = 32'he3399167;
assign table_[148] = 32'he1d4a2c8;
assign table_[149] = 32'he0745b24;
assign table_[150] = 32'hdf18f0ce;
assign table_[151] = 32'hddc29958;
assign table_[152] = 32'hdc71898d;
assign table_[153] = 32'hdb25f566;
assign table_[154] = 32'hd9e01006;
assign table_[155] = 32'hd8a00bae;
assign table_[156] = 32'hd76619b6;
assign table_[157] = 32'hd6326a88;
assign table_[158] = 32'hd5052d97;
assign table_[159] = 32'hd3de9156;
assign table_[160] = 32'hd2bec333;
assign table_[161] = 32'hd1a5ef90;
assign table_[162] = 32'hd09441bb;
assign table_[163] = 32'hcf89e3e8;
assign table_[164] = 32'hce86ff2a;
assign table_[165] = 32'hcd8bbb6d;
assign table_[166] = 32'hcc983f70;
assign table_[167] = 32'hcbacb0bf;
assign table_[168] = 32'hcac933ae;
assign table_[169] = 32'hc9edeb50;
assign table_[170] = 32'hc91af976;
assign table_[171] = 32'hc8507ea7;
assign table_[172] = 32'hc78e9a1d;
assign table_[173] = 32'hc6d569be;
assign table_[174] = 32'hc6250a18;
assign table_[175] = 32'hc57d965d;
assign table_[176] = 32'hc4df2862;
assign table_[177] = 32'hc449d892;
assign table_[178] = 32'hc3bdbdf6;
assign table_[179] = 32'hc33aee27;
assign table_[180] = 32'hc2c17d52;
assign table_[181] = 32'hc2517e31;
assign table_[182] = 32'hc1eb0209;
assign table_[183] = 32'hc18e18a7;
assign table_[184] = 32'hc13ad060;
assign table_[185] = 32'hc0f1360b;
assign table_[186] = 32'hc0b15502;
assign table_[187] = 32'hc07b371e;
assign table_[188] = 32'hc04ee4b8;
assign table_[189] = 32'hc02c64a6;
assign table_[190] = 32'hc013bc39;
assign table_[191] = 32'hc004ef3f;
assign table_[192] = 32'hc0000000;
assign table_[193] = 32'hc004ef3f;
assign table_[194] = 32'hc013bc39;
assign table_[195] = 32'hc02c64a6;
assign table_[196] = 32'hc04ee4b8;
assign table_[197] = 32'hc07b371e;
assign table_[198] = 32'hc0b15502;
assign table_[199] = 32'hc0f1360b;
assign table_[200] = 32'hc13ad060;
assign table_[201] = 32'hc18e18a7;
assign table_[202] = 32'hc1eb0209;
assign table_[203] = 32'hc2517e31;
assign table_[204] = 32'hc2c17d52;
assign table_[205] = 32'hc33aee27;
assign table_[206] = 32'hc3bdbdf6;
assign table_[207] = 32'hc449d892;
assign table_[208] = 32'hc4df2862;
assign table_[209] = 32'hc57d965d;
assign table_[210] = 32'hc6250a18;
assign table_[211] = 32'hc6d569be;
assign table_[212] = 32'hc78e9a1d;
assign table_[213] = 32'hc8507ea7;
assign table_[214] = 32'hc91af976;
assign table_[215] = 32'hc9edeb50;
assign table_[216] = 32'hcac933ae;
assign table_[217] = 32'hcbacb0bf;
assign table_[218] = 32'hcc983f70;
assign table_[219] = 32'hcd8bbb6d;
assign table_[220] = 32'hce86ff2a;
assign table_[221] = 32'hcf89e3e8;
assign table_[222] = 32'hd09441bb;
assign table_[223] = 32'hd1a5ef90;
assign table_[224] = 32'hd2bec333;
assign table_[225] = 32'hd3de9156;
assign table_[226] = 32'hd5052d97;
assign table_[227] = 32'hd6326a88;
assign table_[228] = 32'hd76619b6;
assign table_[229] = 32'hd8a00bae;
assign table_[230] = 32'hd9e01006;
assign table_[231] = 32'hdb25f566;
assign table_[232] = 32'hdc71898d;
assign table_[233] = 32'hddc29958;
assign table_[234] = 32'hdf18f0ce;
assign table_[235] = 32'he0745b24;
assign table_[236] = 32'he1d4a2c8;
assign table_[237] = 32'he3399167;
assign table_[238] = 32'he4a2eff6;
assign table_[239] = 32'he61086bc;
assign table_[240] = 32'he7821d59;
assign table_[241] = 32'he8f77acf;
assign table_[242] = 32'hea70658a;
assign table_[243] = 32'hebeca36c;
assign table_[244] = 32'hed6bf9d1;
assign table_[245] = 32'heeee2d9d;
assign table_[246] = 32'hf0730342;
assign table_[247] = 32'hf1fa3ecb;
assign table_[248] = 32'hf383a3e2;
assign table_[249] = 32'hf50ef5de;
assign table_[250] = 32'hf69bf7c9;
assign table_[251] = 32'hf82a6c6a;
assign table_[252] = 32'hf9ba1651;
assign table_[253] = 32'hfb4ab7db;
assign table_[254] = 32'hfcdc1342;
assign table_[255] = 32'hfe6deaa1;
