module cust_rom (clk0,
    cs0,
    addr0,
    dout0);
 input clk0;
 input cs0;
 input [7:0] addr0;
 output [31:0] dout0;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire \addr0_reg[0] ;
 wire \addr0_reg[1] ;
 wire \addr0_reg[2] ;
 wire \addr0_reg[3] ;
 wire \addr0_reg[4] ;
 wire \addr0_reg[5] ;
 wire \addr0_reg[6] ;
 wire \addr0_reg[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire clknet_0_clk0;
 wire clknet_2_0__leaf_clk0;
 wire clknet_2_1__leaf_clk0;
 wire clknet_2_2__leaf_clk0;
 wire clknet_2_3__leaf_clk0;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;

 sky130_fd_sc_hd__inv_2 _0707_ (.A(net9),
    .Y(_0648_));
 sky130_fd_sc_hd__and4b_1 _0708_ (.A_N(net129),
    .B(net127),
    .C(net131),
    .D(net133),
    .X(_0658_));
 sky130_fd_sc_hd__and4_1 _0709_ (.A(net125),
    .B(net123),
    .C(net119),
    .D(net121),
    .X(_0668_));
 sky130_fd_sc_hd__and4bb_1 _0710_ (.A_N(net127),
    .B_N(net131),
    .C(net133),
    .D(net129),
    .X(_0677_));
 sky130_fd_sc_hd__nor4b_1 _0711_ (.A(net126),
    .B(net124),
    .C(net122),
    .D_N(net120),
    .Y(_0685_));
 sky130_fd_sc_hd__a22o_2 _0712_ (.A1(net118),
    .A2(net116),
    .B1(net114),
    .B2(net111),
    .X(_0686_));
 sky130_fd_sc_hd__or4b_4 _0713_ (.A(net129),
    .B(net131),
    .C(net133),
    .D_N(net127),
    .X(_0687_));
 sky130_fd_sc_hd__o21ba_2 _0714_ (.A1(net116),
    .A2(net111),
    .B1_N(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__and4b_1 _0715_ (.A_N(net127),
    .B(net131),
    .C(net133),
    .D(net129),
    .X(_0689_));
 sky130_fd_sc_hd__and4bb_1 _0716_ (.A_N(net129),
    .B_N(net131),
    .C(net133),
    .D(net127),
    .X(_0690_));
 sky130_fd_sc_hd__a22o_2 _0717_ (.A1(net111),
    .A2(net108),
    .B1(net106),
    .B2(net116),
    .X(_0691_));
 sky130_fd_sc_hd__and4bb_1 _0718_ (.A_N(net130),
    .B_N(net134),
    .C(net131),
    .D(net127),
    .X(_0692_));
 sky130_fd_sc_hd__and4bb_1 _0719_ (.A_N(net128),
    .B_N(net133),
    .C(net132),
    .D(net130),
    .X(_0693_));
 sky130_fd_sc_hd__a22o_2 _0720_ (.A1(net116),
    .A2(net105),
    .B1(net103),
    .B2(net111),
    .X(_0694_));
 sky130_fd_sc_hd__or2_1 _0721_ (.A(_0691_),
    .B(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__or2_1 _0722_ (.A(_0688_),
    .B(_0691_),
    .X(_0696_));
 sky130_fd_sc_hd__or3_1 _0723_ (.A(_0688_),
    .B(_0691_),
    .C(_0694_),
    .X(_0697_));
 sky130_fd_sc_hd__or4_2 _0724_ (.A(_0686_),
    .B(_0688_),
    .C(_0691_),
    .D(_0694_),
    .X(_0698_));
 sky130_fd_sc_hd__a22o_1 _0725_ (.A1(net116),
    .A2(net113),
    .B1(net110),
    .B2(net117),
    .X(_0699_));
 sky130_fd_sc_hd__nor4b_1 _0726_ (.A(net128),
    .B(net132),
    .C(net134),
    .D_N(net130),
    .Y(_0700_));
 sky130_fd_sc_hd__and4bb_1 _0727_ (.A_N(net132),
    .B_N(net133),
    .C(net130),
    .D(net128),
    .X(_0701_));
 sky130_fd_sc_hd__a22o_2 _0728_ (.A1(net115),
    .A2(net98),
    .B1(net96),
    .B2(net110),
    .X(_0702_));
 sky130_fd_sc_hd__or2_1 _0729_ (.A(_0699_),
    .B(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__a22o_1 _0730_ (.A1(net111),
    .A2(net105),
    .B1(net103),
    .B2(net116),
    .X(_0704_));
 sky130_fd_sc_hd__a22o_1 _0731_ (.A1(net115),
    .A2(net108),
    .B1(net106),
    .B2(net110),
    .X(_0705_));
 sky130_fd_sc_hd__or2_2 _0732_ (.A(_0704_),
    .B(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__or4_2 _0733_ (.A(_0699_),
    .B(_0702_),
    .C(_0704_),
    .D(_0705_),
    .X(_0032_));
 sky130_fd_sc_hd__or2_1 _0734_ (.A(_0698_),
    .B(_0032_),
    .X(_0033_));
 sky130_fd_sc_hd__and4b_1 _0735_ (.A_N(net131),
    .B(net133),
    .C(net129),
    .D(net127),
    .X(_0034_));
 sky130_fd_sc_hd__and4bb_1 _0736_ (.A_N(net129),
    .B_N(net127),
    .C(net131),
    .D(net133),
    .X(_0035_));
 sky130_fd_sc_hd__a22o_2 _0737_ (.A1(net115),
    .A2(net94),
    .B1(net92),
    .B2(net110),
    .X(_0036_));
 sky130_fd_sc_hd__nor4b_1 _0738_ (.A(net129),
    .B(net128),
    .C(net131),
    .D_N(net134),
    .Y(_0037_));
 sky130_fd_sc_hd__and4_1 _0739_ (.A(net130),
    .B(net127),
    .C(net132),
    .D(net134),
    .X(_0038_));
 sky130_fd_sc_hd__a22o_2 _0740_ (.A1(net110),
    .A2(net89),
    .B1(net87),
    .B2(net115),
    .X(_0039_));
 sky130_fd_sc_hd__or2_1 _0741_ (.A(_0036_),
    .B(_0039_),
    .X(_0040_));
 sky130_fd_sc_hd__a22o_1 _0742_ (.A1(net110),
    .A2(net98),
    .B1(net96),
    .B2(net115),
    .X(_0041_));
 sky130_fd_sc_hd__and4b_1 _0743_ (.A_N(net134),
    .B(net132),
    .C(net128),
    .D(net129),
    .X(_0042_));
 sky130_fd_sc_hd__nor4b_1 _0744_ (.A(net130),
    .B(net128),
    .C(net134),
    .D_N(net132),
    .Y(_0043_));
 sky130_fd_sc_hd__a22o_2 _0745_ (.A1(net115),
    .A2(net85),
    .B1(net81),
    .B2(net110),
    .X(_0044_));
 sky130_fd_sc_hd__or2_1 _0746_ (.A(_0041_),
    .B(_0044_),
    .X(_0045_));
 sky130_fd_sc_hd__or2_2 _0747_ (.A(_0036_),
    .B(_0041_),
    .X(_0046_));
 sky130_fd_sc_hd__or4_2 _0748_ (.A(_0036_),
    .B(_0039_),
    .C(_0041_),
    .D(_0044_),
    .X(_0047_));
 sky130_fd_sc_hd__a22o_1 _0749_ (.A1(net115),
    .A2(net89),
    .B1(net87),
    .B2(net110),
    .X(_0048_));
 sky130_fd_sc_hd__a22o_2 _0750_ (.A1(net110),
    .A2(net94),
    .B1(net92),
    .B2(net115),
    .X(_0049_));
 sky130_fd_sc_hd__or4_4 _0751_ (.A(net129),
    .B(net127),
    .C(net131),
    .D(net133),
    .X(_0050_));
 sky130_fd_sc_hd__and4bb_1 _0752_ (.A_N(net123),
    .B_N(net121),
    .C(net119),
    .D(net125),
    .X(_0051_));
 sky130_fd_sc_hd__o21ba_2 _0753_ (.A1(net115),
    .A2(net79),
    .B1_N(_0050_),
    .X(_0052_));
 sky130_fd_sc_hd__a22o_1 _0754_ (.A1(net110),
    .A2(net85),
    .B1(net81),
    .B2(net115),
    .X(_0053_));
 sky130_fd_sc_hd__or3_1 _0755_ (.A(_0049_),
    .B(_0052_),
    .C(_0053_),
    .X(_0054_));
 sky130_fd_sc_hd__or2_1 _0756_ (.A(_0048_),
    .B(_0049_),
    .X(_0055_));
 sky130_fd_sc_hd__or2_1 _0757_ (.A(_0048_),
    .B(_0053_),
    .X(_0056_));
 sky130_fd_sc_hd__or4_1 _0758_ (.A(_0048_),
    .B(_0049_),
    .C(_0052_),
    .D(_0053_),
    .X(_0057_));
 sky130_fd_sc_hd__or4_1 _0759_ (.A(_0698_),
    .B(_0032_),
    .C(_0047_),
    .D(_0057_),
    .X(_0058_));
 sky130_fd_sc_hd__and4b_1 _0760_ (.A_N(net123),
    .B(net119),
    .C(net121),
    .D(net125),
    .X(_0059_));
 sky130_fd_sc_hd__nand3b_1 _0761_ (.A_N(net126),
    .B(net124),
    .C(net120),
    .Y(_0060_));
 sky130_fd_sc_hd__and4bb_1 _0762_ (.A_N(net125),
    .B_N(net121),
    .C(net119),
    .D(net123),
    .X(_0061_));
 sky130_fd_sc_hd__a22o_1 _0763_ (.A1(net92),
    .A2(net77),
    .B1(net75),
    .B2(net94),
    .X(_0062_));
 sky130_fd_sc_hd__a22o_1 _0764_ (.A1(net81),
    .A2(net78),
    .B1(net76),
    .B2(net85),
    .X(_0063_));
 sky130_fd_sc_hd__or2_1 _0765_ (.A(_0062_),
    .B(_0063_),
    .X(_0064_));
 sky130_fd_sc_hd__and4b_1 _0766_ (.A_N(net121),
    .B(net119),
    .C(net123),
    .D(net125),
    .X(_0065_));
 sky130_fd_sc_hd__o21ba_1 _0767_ (.A1(net77),
    .A2(net74),
    .B1_N(_0050_),
    .X(_0066_));
 sky130_fd_sc_hd__a22o_2 _0768_ (.A1(net89),
    .A2(net77),
    .B1(net75),
    .B2(net87),
    .X(_0067_));
 sky130_fd_sc_hd__or2_2 _0769_ (.A(_0062_),
    .B(_0066_),
    .X(_0068_));
 sky130_fd_sc_hd__or4_2 _0770_ (.A(_0062_),
    .B(_0063_),
    .C(_0066_),
    .D(_0067_),
    .X(_0069_));
 sky130_fd_sc_hd__and4b_1 _0771_ (.A_N(net125),
    .B(net123),
    .C(net119),
    .D(net121),
    .X(_0070_));
 sky130_fd_sc_hd__a22o_2 _0772_ (.A1(net113),
    .A2(net79),
    .B1(net71),
    .B2(net117),
    .X(_0071_));
 sky130_fd_sc_hd__a22o_2 _0773_ (.A1(net102),
    .A2(net80),
    .B1(net72),
    .B2(net104),
    .X(_0072_));
 sky130_fd_sc_hd__and4bb_1 _0774_ (.A_N(net125),
    .B_N(net123),
    .C(net119),
    .D(net121),
    .X(_0073_));
 sky130_fd_sc_hd__a22o_1 _0775_ (.A1(net87),
    .A2(net74),
    .B1(net70),
    .B2(net89),
    .X(_0074_));
 sky130_fd_sc_hd__a22o_2 _0776_ (.A1(net94),
    .A2(net74),
    .B1(net70),
    .B2(net92),
    .X(_0075_));
 sky130_fd_sc_hd__or4_1 _0777_ (.A(_0071_),
    .B(_0072_),
    .C(_0074_),
    .D(_0075_),
    .X(_0076_));
 sky130_fd_sc_hd__a22o_2 _0778_ (.A1(net89),
    .A2(net79),
    .B1(net72),
    .B2(net88),
    .X(_0077_));
 sky130_fd_sc_hd__a22o_1 _0779_ (.A1(net81),
    .A2(net80),
    .B1(net72),
    .B2(net85),
    .X(_0078_));
 sky130_fd_sc_hd__or2_1 _0780_ (.A(_0077_),
    .B(net48),
    .X(_0079_));
 sky130_fd_sc_hd__a22o_2 _0781_ (.A1(net98),
    .A2(net80),
    .B1(net72),
    .B2(net96),
    .X(_0080_));
 sky130_fd_sc_hd__a22o_2 _0782_ (.A1(net92),
    .A2(net79),
    .B1(net71),
    .B2(net94),
    .X(_0081_));
 sky130_fd_sc_hd__or3_1 _0783_ (.A(_0077_),
    .B(net48),
    .C(_0081_),
    .X(_0082_));
 sky130_fd_sc_hd__or4_1 _0784_ (.A(_0077_),
    .B(net48),
    .C(_0080_),
    .D(_0081_),
    .X(_0083_));
 sky130_fd_sc_hd__a22o_2 _0785_ (.A1(net117),
    .A2(net74),
    .B1(net70),
    .B2(net113),
    .X(_0084_));
 sky130_fd_sc_hd__a22o_2 _0786_ (.A1(net96),
    .A2(net73),
    .B1(net69),
    .B2(net98),
    .X(_0085_));
 sky130_fd_sc_hd__a22o_2 _0787_ (.A1(net106),
    .A2(net73),
    .B1(net69),
    .B2(net108),
    .X(_0086_));
 sky130_fd_sc_hd__a22o_1 _0788_ (.A1(net104),
    .A2(net73),
    .B1(net70),
    .B2(net102),
    .X(_0087_));
 sky130_fd_sc_hd__or4_2 _0789_ (.A(_0084_),
    .B(_0085_),
    .C(_0086_),
    .D(_0087_),
    .X(_0088_));
 sky130_fd_sc_hd__or4_1 _0790_ (.A(_0069_),
    .B(_0076_),
    .C(_0083_),
    .D(_0088_),
    .X(_0089_));
 sky130_fd_sc_hd__a22o_2 _0791_ (.A1(net81),
    .A2(net73),
    .B1(net69),
    .B2(net85),
    .X(_0090_));
 sky130_fd_sc_hd__a22o_2 _0792_ (.A1(net92),
    .A2(net73),
    .B1(net69),
    .B2(net94),
    .X(_0091_));
 sky130_fd_sc_hd__a22o_2 _0793_ (.A1(net89),
    .A2(net73),
    .B1(net69),
    .B2(net87),
    .X(_0092_));
 sky130_fd_sc_hd__a22o_1 _0794_ (.A1(net98),
    .A2(net73),
    .B1(net69),
    .B2(net96),
    .X(_0093_));
 sky130_fd_sc_hd__or2_2 _0795_ (.A(_0090_),
    .B(_0093_),
    .X(_0094_));
 sky130_fd_sc_hd__or2_1 _0796_ (.A(_0090_),
    .B(_0092_),
    .X(_0095_));
 sky130_fd_sc_hd__or4_2 _0797_ (.A(_0090_),
    .B(_0091_),
    .C(_0092_),
    .D(_0093_),
    .X(_0096_));
 sky130_fd_sc_hd__a22o_1 _0798_ (.A1(net98),
    .A2(net78),
    .B1(net76),
    .B2(net96),
    .X(_0097_));
 sky130_fd_sc_hd__a22o_2 _0799_ (.A1(net108),
    .A2(net77),
    .B1(net75),
    .B2(net106),
    .X(_0098_));
 sky130_fd_sc_hd__a22o_2 _0800_ (.A1(net113),
    .A2(net77),
    .B1(net75),
    .B2(net117),
    .X(_0099_));
 sky130_fd_sc_hd__a22o_1 _0801_ (.A1(net102),
    .A2(net77),
    .B1(net75),
    .B2(net104),
    .X(_0100_));
 sky130_fd_sc_hd__or2_2 _0802_ (.A(_0098_),
    .B(_0100_),
    .X(_0101_));
 sky130_fd_sc_hd__or4_1 _0803_ (.A(net47),
    .B(_0098_),
    .C(_0099_),
    .D(_0100_),
    .X(_0102_));
 sky130_fd_sc_hd__a22o_2 _0804_ (.A1(net106),
    .A2(net79),
    .B1(net71),
    .B2(net108),
    .X(_0103_));
 sky130_fd_sc_hd__a22o_1 _0805_ (.A1(net96),
    .A2(net79),
    .B1(net72),
    .B2(net98),
    .X(_0104_));
 sky130_fd_sc_hd__or2_1 _0806_ (.A(_0103_),
    .B(_0104_),
    .X(_0105_));
 sky130_fd_sc_hd__a22o_1 _0807_ (.A1(net104),
    .A2(net79),
    .B1(net71),
    .B2(net102),
    .X(_0106_));
 sky130_fd_sc_hd__a22o_2 _0808_ (.A1(net117),
    .A2(net79),
    .B1(net71),
    .B2(net113),
    .X(_0107_));
 sky130_fd_sc_hd__or3_1 _0809_ (.A(_0103_),
    .B(_0104_),
    .C(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__or4_4 _0810_ (.A(_0103_),
    .B(_0104_),
    .C(_0106_),
    .D(_0107_),
    .X(_0109_));
 sky130_fd_sc_hd__nor2_2 _0811_ (.A(_0050_),
    .B(_0060_),
    .Y(_0110_));
 sky130_fd_sc_hd__a22o_2 _0812_ (.A1(net87),
    .A2(net80),
    .B1(net71),
    .B2(net89),
    .X(_0111_));
 sky130_fd_sc_hd__or2_1 _0813_ (.A(_0110_),
    .B(_0111_),
    .X(_0112_));
 sky130_fd_sc_hd__a22o_1 _0814_ (.A1(net95),
    .A2(net79),
    .B1(net71),
    .B2(net93),
    .X(_0113_));
 sky130_fd_sc_hd__a22o_2 _0815_ (.A1(net85),
    .A2(net80),
    .B1(net71),
    .B2(net81),
    .X(_0114_));
 sky130_fd_sc_hd__or3_2 _0816_ (.A(_0110_),
    .B(_0111_),
    .C(_0114_),
    .X(_0115_));
 sky130_fd_sc_hd__or4_1 _0817_ (.A(_0110_),
    .B(_0111_),
    .C(_0113_),
    .D(_0114_),
    .X(_0116_));
 sky130_fd_sc_hd__or4_1 _0818_ (.A(_0096_),
    .B(_0102_),
    .C(_0109_),
    .D(_0116_),
    .X(_0117_));
 sky130_fd_sc_hd__a22o_1 _0819_ (.A1(net94),
    .A2(net77),
    .B1(net75),
    .B2(net92),
    .X(_0118_));
 sky130_fd_sc_hd__a22o_2 _0820_ (.A1(net96),
    .A2(net77),
    .B1(net75),
    .B2(net98),
    .X(_0119_));
 sky130_fd_sc_hd__or2_2 _0821_ (.A(_0118_),
    .B(_0119_),
    .X(_0120_));
 sky130_fd_sc_hd__a22o_1 _0822_ (.A1(net87),
    .A2(net78),
    .B1(net76),
    .B2(net89),
    .X(_0121_));
 sky130_fd_sc_hd__a22o_2 _0823_ (.A1(net85),
    .A2(net78),
    .B1(net76),
    .B2(net81),
    .X(_0122_));
 sky130_fd_sc_hd__or2_1 _0824_ (.A(_0121_),
    .B(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__or4_2 _0825_ (.A(_0118_),
    .B(_0119_),
    .C(_0121_),
    .D(_0122_),
    .X(_0124_));
 sky130_fd_sc_hd__a22o_1 _0826_ (.A1(net117),
    .A2(net77),
    .B1(net75),
    .B2(net113),
    .X(_0125_));
 sky130_fd_sc_hd__a22o_1 _0827_ (.A1(net104),
    .A2(net78),
    .B1(net75),
    .B2(net102),
    .X(_0126_));
 sky130_fd_sc_hd__or2_2 _0828_ (.A(_0125_),
    .B(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__a22o_2 _0829_ (.A1(net106),
    .A2(net77),
    .B1(net75),
    .B2(net108),
    .X(_0128_));
 sky130_fd_sc_hd__o21ba_2 _0830_ (.A1(net78),
    .A2(net76),
    .B1_N(_0687_),
    .X(_0129_));
 sky130_fd_sc_hd__or4_4 _0831_ (.A(_0125_),
    .B(_0126_),
    .C(_0128_),
    .D(_0129_),
    .X(_0130_));
 sky130_fd_sc_hd__a22o_2 _0832_ (.A1(net113),
    .A2(net73),
    .B1(net69),
    .B2(net117),
    .X(_0131_));
 sky130_fd_sc_hd__a22o_2 _0833_ (.A1(net108),
    .A2(net73),
    .B1(net69),
    .B2(net106),
    .X(_0132_));
 sky130_fd_sc_hd__or2_1 _0834_ (.A(_0131_),
    .B(_0132_),
    .X(_0133_));
 sky130_fd_sc_hd__a22o_1 _0835_ (.A1(net85),
    .A2(net74),
    .B1(net70),
    .B2(net81),
    .X(_0134_));
 sky130_fd_sc_hd__and2b_1 _0836_ (.A_N(_0050_),
    .B(net70),
    .X(_0135_));
 sky130_fd_sc_hd__a22o_2 _0837_ (.A1(net102),
    .A2(net74),
    .B1(net69),
    .B2(net104),
    .X(_0136_));
 sky130_fd_sc_hd__o21ba_1 _0838_ (.A1(net73),
    .A2(net69),
    .B1_N(_0687_),
    .X(_0137_));
 sky130_fd_sc_hd__o21ba_2 _0839_ (.A1(net80),
    .A2(net71),
    .B1_N(_0687_),
    .X(_0138_));
 sky130_fd_sc_hd__a22o_2 _0840_ (.A1(net108),
    .A2(net79),
    .B1(net71),
    .B2(net106),
    .X(_0139_));
 sky130_fd_sc_hd__or2_1 _0841_ (.A(_0131_),
    .B(_0136_),
    .X(_0140_));
 sky130_fd_sc_hd__or4_1 _0842_ (.A(_0131_),
    .B(_0132_),
    .C(_0136_),
    .D(_0137_),
    .X(_0141_));
 sky130_fd_sc_hd__or4_1 _0843_ (.A(_0134_),
    .B(_0135_),
    .C(_0138_),
    .D(_0139_),
    .X(_0142_));
 sky130_fd_sc_hd__or4_1 _0844_ (.A(_0124_),
    .B(_0130_),
    .C(_0141_),
    .D(_0142_),
    .X(_0143_));
 sky130_fd_sc_hd__or4_1 _0845_ (.A(_0058_),
    .B(_0089_),
    .C(_0117_),
    .D(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__nor4b_1 _0846_ (.A(net126),
    .B(net124),
    .C(net120),
    .D_N(net121),
    .Y(_0145_));
 sky130_fd_sc_hd__and4bb_1 _0847_ (.A_N(net120),
    .B_N(net122),
    .C(net126),
    .D(net124),
    .X(_0146_));
 sky130_fd_sc_hd__o21ba_2 _0848_ (.A1(net67),
    .A2(net65),
    .B1_N(_0687_),
    .X(_0147_));
 sky130_fd_sc_hd__a22o_2 _0849_ (.A1(net99),
    .A2(net67),
    .B1(net65),
    .B2(net97),
    .X(_0148_));
 sky130_fd_sc_hd__a22o_2 _0850_ (.A1(net92),
    .A2(net66),
    .B1(net64),
    .B2(net94),
    .X(_0149_));
 sky130_fd_sc_hd__a22o_1 _0851_ (.A1(net90),
    .A2(net66),
    .B1(net64),
    .B2(net87),
    .X(_0150_));
 sky130_fd_sc_hd__a22o_1 _0852_ (.A1(net82),
    .A2(net66),
    .B1(net64),
    .B2(net86),
    .X(_0151_));
 sky130_fd_sc_hd__or2_2 _0853_ (.A(_0150_),
    .B(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__or4_2 _0854_ (.A(_0148_),
    .B(_0149_),
    .C(_0150_),
    .D(_0151_),
    .X(_0153_));
 sky130_fd_sc_hd__a22o_2 _0855_ (.A1(net102),
    .A2(net66),
    .B1(net64),
    .B2(net104),
    .X(_0154_));
 sky130_fd_sc_hd__a22o_1 _0856_ (.A1(net113),
    .A2(net66),
    .B1(net64),
    .B2(net117),
    .X(_0155_));
 sky130_fd_sc_hd__a22o_1 _0857_ (.A1(net109),
    .A2(net66),
    .B1(net64),
    .B2(net107),
    .X(_0156_));
 sky130_fd_sc_hd__or2_1 _0858_ (.A(_0154_),
    .B(_0155_),
    .X(_0157_));
 sky130_fd_sc_hd__or2_1 _0859_ (.A(_0154_),
    .B(_0156_),
    .X(_0158_));
 sky130_fd_sc_hd__or3_1 _0860_ (.A(_0154_),
    .B(_0155_),
    .C(_0156_),
    .X(_0159_));
 sky130_fd_sc_hd__or2_1 _0861_ (.A(_0153_),
    .B(_0159_),
    .X(_0160_));
 sky130_fd_sc_hd__or4_4 _0862_ (.A(_0147_),
    .B(_0154_),
    .C(_0155_),
    .D(_0156_),
    .X(_0161_));
 sky130_fd_sc_hd__or2_1 _0863_ (.A(_0153_),
    .B(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__a22o_2 _0864_ (.A1(net88),
    .A2(net67),
    .B1(net65),
    .B2(net90),
    .X(_0163_));
 sky130_fd_sc_hd__a22o_1 _0865_ (.A1(net95),
    .A2(net66),
    .B1(net64),
    .B2(net93),
    .X(_0164_));
 sky130_fd_sc_hd__or2_1 _0866_ (.A(_0163_),
    .B(_0164_),
    .X(_0165_));
 sky130_fd_sc_hd__a22o_1 _0867_ (.A1(net86),
    .A2(net66),
    .B1(net64),
    .B2(net82),
    .X(_0166_));
 sky130_fd_sc_hd__and4bb_1 _0868_ (.A_N(net123),
    .B_N(net119),
    .C(net121),
    .D(net125),
    .X(_0167_));
 sky130_fd_sc_hd__o21ba_2 _0869_ (.A1(net64),
    .A2(_0167_),
    .B1_N(_0050_),
    .X(_0168_));
 sky130_fd_sc_hd__or2_2 _0870_ (.A(_0163_),
    .B(_0168_),
    .X(_0169_));
 sky130_fd_sc_hd__or2_1 _0871_ (.A(_0163_),
    .B(_0166_),
    .X(_0170_));
 sky130_fd_sc_hd__or2_1 _0872_ (.A(_0164_),
    .B(_0168_),
    .X(_0171_));
 sky130_fd_sc_hd__or4_1 _0873_ (.A(_0163_),
    .B(_0164_),
    .C(_0166_),
    .D(_0168_),
    .X(_0172_));
 sky130_fd_sc_hd__a22o_2 _0874_ (.A1(net104),
    .A2(net67),
    .B1(net65),
    .B2(net102),
    .X(_0173_));
 sky130_fd_sc_hd__a22o_2 _0875_ (.A1(net107),
    .A2(net66),
    .B1(net65),
    .B2(net109),
    .X(_0174_));
 sky130_fd_sc_hd__a22o_1 _0876_ (.A1(net97),
    .A2(net67),
    .B1(net65),
    .B2(net99),
    .X(_0175_));
 sky130_fd_sc_hd__a22o_1 _0877_ (.A1(net118),
    .A2(net66),
    .B1(net64),
    .B2(net114),
    .X(_0176_));
 sky130_fd_sc_hd__or2_2 _0878_ (.A(_0175_),
    .B(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__or4_1 _0879_ (.A(_0173_),
    .B(_0174_),
    .C(_0175_),
    .D(_0176_),
    .X(_0178_));
 sky130_fd_sc_hd__or4_1 _0880_ (.A(_0153_),
    .B(_0161_),
    .C(_0172_),
    .D(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__nor4b_2 _0881_ (.A(net125),
    .B(net119),
    .C(_0050_),
    .D_N(net123),
    .Y(_0180_));
 sky130_fd_sc_hd__nor4b_1 _0882_ (.A(net125),
    .B(net119),
    .C(net121),
    .D_N(net123),
    .Y(_0181_));
 sky130_fd_sc_hd__a22o_2 _0883_ (.A1(net85),
    .A2(net62),
    .B1(net60),
    .B2(net81),
    .X(_0182_));
 sky130_fd_sc_hd__a22o_2 _0884_ (.A1(net87),
    .A2(net62),
    .B1(net60),
    .B2(net89),
    .X(_0183_));
 sky130_fd_sc_hd__a22o_1 _0885_ (.A1(net94),
    .A2(net63),
    .B1(net60),
    .B2(net92),
    .X(_0184_));
 sky130_fd_sc_hd__or4_1 _0886_ (.A(net46),
    .B(_0182_),
    .C(_0183_),
    .D(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__a22o_2 _0887_ (.A1(net117),
    .A2(net62),
    .B1(net60),
    .B2(net113),
    .X(_0186_));
 sky130_fd_sc_hd__a22o_1 _0888_ (.A1(net96),
    .A2(net62),
    .B1(net60),
    .B2(net98),
    .X(_0187_));
 sky130_fd_sc_hd__a22o_2 _0889_ (.A1(net106),
    .A2(net62),
    .B1(net61),
    .B2(net108),
    .X(_0188_));
 sky130_fd_sc_hd__a22o_2 _0890_ (.A1(net104),
    .A2(net63),
    .B1(net60),
    .B2(net102),
    .X(_0189_));
 sky130_fd_sc_hd__or2_1 _0891_ (.A(_0188_),
    .B(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__or4_1 _0892_ (.A(_0186_),
    .B(_0187_),
    .C(_0188_),
    .D(_0189_),
    .X(_0191_));
 sky130_fd_sc_hd__or2_1 _0893_ (.A(_0185_),
    .B(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__a22o_2 _0894_ (.A1(net108),
    .A2(net63),
    .B1(net61),
    .B2(net106),
    .X(_0193_));
 sky130_fd_sc_hd__a22o_2 _0895_ (.A1(net102),
    .A2(net63),
    .B1(net61),
    .B2(net104),
    .X(_0194_));
 sky130_fd_sc_hd__a22o_2 _0896_ (.A1(net113),
    .A2(net62),
    .B1(net61),
    .B2(net117),
    .X(_0195_));
 sky130_fd_sc_hd__o21ba_2 _0897_ (.A1(net62),
    .A2(net60),
    .B1_N(_0687_),
    .X(_0196_));
 sky130_fd_sc_hd__or2_1 _0898_ (.A(_0195_),
    .B(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__or2_1 _0899_ (.A(_0194_),
    .B(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__or4_1 _0900_ (.A(_0193_),
    .B(_0194_),
    .C(_0195_),
    .D(_0196_),
    .X(_0199_));
 sky130_fd_sc_hd__a22o_2 _0901_ (.A1(net92),
    .A2(net63),
    .B1(net61),
    .B2(net94),
    .X(_0200_));
 sky130_fd_sc_hd__a22o_1 _0902_ (.A1(net89),
    .A2(net62),
    .B1(net60),
    .B2(net87),
    .X(_0201_));
 sky130_fd_sc_hd__a22o_2 _0903_ (.A1(net98),
    .A2(net62),
    .B1(net60),
    .B2(net96),
    .X(_0202_));
 sky130_fd_sc_hd__a22o_2 _0904_ (.A1(net81),
    .A2(net62),
    .B1(net60),
    .B2(net85),
    .X(_0203_));
 sky130_fd_sc_hd__or2_1 _0905_ (.A(_0201_),
    .B(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__or3_2 _0906_ (.A(_0201_),
    .B(_0202_),
    .C(_0203_),
    .X(_0205_));
 sky130_fd_sc_hd__or2_1 _0907_ (.A(_0200_),
    .B(_0202_),
    .X(_0206_));
 sky130_fd_sc_hd__or3_1 _0908_ (.A(_0199_),
    .B(_0200_),
    .C(_0205_),
    .X(_0207_));
 sky130_fd_sc_hd__or3_1 _0909_ (.A(_0179_),
    .B(_0192_),
    .C(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__and4bb_1 _0910_ (.A_N(net126),
    .B_N(net120),
    .C(net122),
    .D(net124),
    .X(_0209_));
 sky130_fd_sc_hd__nor4b_1 _0911_ (.A(net124),
    .B(net120),
    .C(net122),
    .D_N(net126),
    .Y(_0210_));
 sky130_fd_sc_hd__o21ba_1 _0912_ (.A1(net58),
    .A2(net54),
    .B1_N(_0687_),
    .X(_0211_));
 sky130_fd_sc_hd__a22o_1 _0913_ (.A1(net103),
    .A2(net59),
    .B1(net55),
    .B2(net105),
    .X(_0212_));
 sky130_fd_sc_hd__a22o_1 _0914_ (.A1(net114),
    .A2(net58),
    .B1(net54),
    .B2(net118),
    .X(_0213_));
 sky130_fd_sc_hd__or2_1 _0915_ (.A(_0212_),
    .B(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__a22o_1 _0916_ (.A1(net109),
    .A2(net58),
    .B1(net54),
    .B2(net107),
    .X(_0215_));
 sky130_fd_sc_hd__or2_1 _0917_ (.A(_0212_),
    .B(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__or2_1 _0918_ (.A(_0214_),
    .B(_0215_),
    .X(_0217_));
 sky130_fd_sc_hd__or2_1 _0919_ (.A(_0211_),
    .B(_0213_),
    .X(_0218_));
 sky130_fd_sc_hd__or2_1 _0920_ (.A(_0211_),
    .B(_0215_),
    .X(_0219_));
 sky130_fd_sc_hd__or4_2 _0921_ (.A(_0211_),
    .B(_0212_),
    .C(_0213_),
    .D(_0215_),
    .X(_0220_));
 sky130_fd_sc_hd__a22o_1 _0922_ (.A1(net99),
    .A2(net59),
    .B1(net55),
    .B2(net97),
    .X(_0221_));
 sky130_fd_sc_hd__a22o_2 _0923_ (.A1(net90),
    .A2(net59),
    .B1(net54),
    .B2(net88),
    .X(_0222_));
 sky130_fd_sc_hd__or2_1 _0924_ (.A(_0221_),
    .B(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__a22o_2 _0925_ (.A1(net82),
    .A2(net58),
    .B1(net54),
    .B2(net86),
    .X(_0224_));
 sky130_fd_sc_hd__a22o_2 _0926_ (.A1(net93),
    .A2(net58),
    .B1(net54),
    .B2(net95),
    .X(_0225_));
 sky130_fd_sc_hd__or4_1 _0927_ (.A(_0221_),
    .B(_0222_),
    .C(_0224_),
    .D(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__or2_1 _0928_ (.A(_0220_),
    .B(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__and4b_1 _0929_ (.A_N(net120),
    .B(net122),
    .C(net126),
    .D(net124),
    .X(_0228_));
 sky130_fd_sc_hd__nor4_1 _0930_ (.A(net126),
    .B(net124),
    .C(net120),
    .D(net122),
    .Y(_0229_));
 sky130_fd_sc_hd__a22o_2 _0931_ (.A1(net97),
    .A2(net52),
    .B1(net50),
    .B2(net99),
    .X(_0230_));
 sky130_fd_sc_hd__a22o_1 _0932_ (.A1(net118),
    .A2(net52),
    .B1(net49),
    .B2(net114),
    .X(_0231_));
 sky130_fd_sc_hd__or2_2 _0933_ (.A(_0230_),
    .B(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__a22o_1 _0934_ (.A1(net105),
    .A2(net52),
    .B1(net49),
    .B2(net103),
    .X(_0233_));
 sky130_fd_sc_hd__a22o_1 _0935_ (.A1(net107),
    .A2(net52),
    .B1(net49),
    .B2(net109),
    .X(_0234_));
 sky130_fd_sc_hd__or2_2 _0936_ (.A(_0233_),
    .B(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__or2_1 _0937_ (.A(_0231_),
    .B(_0234_),
    .X(_0236_));
 sky130_fd_sc_hd__o21ba_2 _0938_ (.A1(net54),
    .A2(net53),
    .B1_N(_0050_),
    .X(_0237_));
 sky130_fd_sc_hd__a22o_2 _0939_ (.A1(net95),
    .A2(net58),
    .B1(net54),
    .B2(net93),
    .X(_0238_));
 sky130_fd_sc_hd__or2_1 _0940_ (.A(_0237_),
    .B(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__a22o_2 _0941_ (.A1(net86),
    .A2(net59),
    .B1(net55),
    .B2(net82),
    .X(_0240_));
 sky130_fd_sc_hd__a22o_2 _0942_ (.A1(net88),
    .A2(net59),
    .B1(net55),
    .B2(net90),
    .X(_0241_));
 sky130_fd_sc_hd__or2_1 _0943_ (.A(_0240_),
    .B(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__or2_1 _0944_ (.A(_0238_),
    .B(_0241_),
    .X(_0243_));
 sky130_fd_sc_hd__or4_1 _0945_ (.A(_0237_),
    .B(_0238_),
    .C(_0240_),
    .D(_0241_),
    .X(_0244_));
 sky130_fd_sc_hd__or3_1 _0946_ (.A(_0232_),
    .B(_0235_),
    .C(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__a22o_1 _0947_ (.A1(net109),
    .A2(net52),
    .B1(net49),
    .B2(net107),
    .X(_0246_));
 sky130_fd_sc_hd__a22o_2 _0948_ (.A1(net114),
    .A2(net52),
    .B1(net49),
    .B2(net118),
    .X(_0247_));
 sky130_fd_sc_hd__o21ba_2 _0949_ (.A1(net53),
    .A2(net49),
    .B1_N(_0687_),
    .X(_0248_));
 sky130_fd_sc_hd__a22o_2 _0950_ (.A1(net103),
    .A2(net53),
    .B1(net49),
    .B2(net105),
    .X(_0249_));
 sky130_fd_sc_hd__or2_1 _0951_ (.A(_0248_),
    .B(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__or4_1 _0952_ (.A(_0246_),
    .B(_0247_),
    .C(_0248_),
    .D(_0249_),
    .X(_0251_));
 sky130_fd_sc_hd__a22o_2 _0953_ (.A1(net95),
    .A2(net52),
    .B1(net49),
    .B2(net93),
    .X(_0252_));
 sky130_fd_sc_hd__a22o_2 _0954_ (.A1(net86),
    .A2(net53),
    .B1(net50),
    .B2(net82),
    .X(_0253_));
 sky130_fd_sc_hd__or2_1 _0955_ (.A(_0252_),
    .B(_0253_),
    .X(_0254_));
 sky130_fd_sc_hd__or4_1 _0956_ (.A(net126),
    .B(net124),
    .C(net122),
    .D(_0050_),
    .X(_0255_));
 sky130_fd_sc_hd__a22o_2 _0957_ (.A1(net88),
    .A2(net52),
    .B1(net49),
    .B2(net90),
    .X(_0256_));
 sky130_fd_sc_hd__or4b_1 _0958_ (.A(_0251_),
    .B(_0254_),
    .C(_0256_),
    .D_N(_0255_),
    .X(_0257_));
 sky130_fd_sc_hd__a22o_2 _0959_ (.A1(net99),
    .A2(net52),
    .B1(net50),
    .B2(net97),
    .X(_0258_));
 sky130_fd_sc_hd__a22o_2 _0960_ (.A1(net93),
    .A2(net53),
    .B1(net49),
    .B2(net95),
    .X(_0259_));
 sky130_fd_sc_hd__or2_1 _0961_ (.A(_0258_),
    .B(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__a22o_2 _0962_ (.A1(net90),
    .A2(net53),
    .B1(net50),
    .B2(net88),
    .X(_0261_));
 sky130_fd_sc_hd__a22o_1 _0963_ (.A1(net82),
    .A2(net52),
    .B1(net50),
    .B2(net86),
    .X(_0262_));
 sky130_fd_sc_hd__or2_1 _0964_ (.A(_0261_),
    .B(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__or2_1 _0965_ (.A(_0258_),
    .B(_0261_),
    .X(_0264_));
 sky130_fd_sc_hd__or2_1 _0966_ (.A(_0259_),
    .B(_0262_),
    .X(_0265_));
 sky130_fd_sc_hd__or4_1 _0967_ (.A(_0258_),
    .B(_0259_),
    .C(_0261_),
    .D(_0262_),
    .X(_0266_));
 sky130_fd_sc_hd__a22oi_4 _0968_ (.A1(net105),
    .A2(net59),
    .B1(net55),
    .B2(net103),
    .Y(_0267_));
 sky130_fd_sc_hd__a22oi_4 _0969_ (.A1(net97),
    .A2(net58),
    .B1(net55),
    .B2(net99),
    .Y(_0268_));
 sky130_fd_sc_hd__a22o_2 _0970_ (.A1(net97),
    .A2(net58),
    .B1(net55),
    .B2(net99),
    .X(_0269_));
 sky130_fd_sc_hd__nand2_1 _0971_ (.A(_0267_),
    .B(_0268_),
    .Y(_0270_));
 sky130_fd_sc_hd__a22oi_4 _0972_ (.A1(net107),
    .A2(net58),
    .B1(net54),
    .B2(net109),
    .Y(_0271_));
 sky130_fd_sc_hd__a22oi_4 _0973_ (.A1(net118),
    .A2(net58),
    .B1(net54),
    .B2(net114),
    .Y(_0272_));
 sky130_fd_sc_hd__nand2_1 _0974_ (.A(_0271_),
    .B(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__nand2_1 _0975_ (.A(_0267_),
    .B(_0271_),
    .Y(_0274_));
 sky130_fd_sc_hd__nand2_1 _0976_ (.A(_0268_),
    .B(_0272_),
    .Y(_0275_));
 sky130_fd_sc_hd__nand4_2 _0977_ (.A(_0267_),
    .B(_0268_),
    .C(_0271_),
    .D(_0272_),
    .Y(_0276_));
 sky130_fd_sc_hd__or2_1 _0978_ (.A(_0266_),
    .B(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__or2_1 _0979_ (.A(_0253_),
    .B(_0256_),
    .X(_0278_));
 sky130_fd_sc_hd__or4_1 _0980_ (.A(_0227_),
    .B(_0245_),
    .C(_0257_),
    .D(_0277_),
    .X(_0279_));
 sky130_fd_sc_hd__o21ai_1 _0981_ (.A1(_0208_),
    .A2(_0279_),
    .B1(net9),
    .Y(_0280_));
 sky130_fd_sc_hd__o31a_1 _0982_ (.A1(_0144_),
    .A2(_0208_),
    .A3(_0279_),
    .B1(net9),
    .X(_0281_));
 sky130_fd_sc_hd__or3_1 _0983_ (.A(_0091_),
    .B(net47),
    .C(_0099_),
    .X(_0282_));
 sky130_fd_sc_hd__or3_1 _0984_ (.A(_0140_),
    .B(_0239_),
    .C(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__or2_1 _0985_ (.A(_0699_),
    .B(_0705_),
    .X(_0284_));
 sky130_fd_sc_hd__or3_2 _0986_ (.A(_0699_),
    .B(_0702_),
    .C(_0705_),
    .X(_0285_));
 sky130_fd_sc_hd__or2_1 _0987_ (.A(_0048_),
    .B(_0052_),
    .X(_0286_));
 sky130_fd_sc_hd__or3_1 _0988_ (.A(_0283_),
    .B(_0285_),
    .C(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__or2_1 _0989_ (.A(_0150_),
    .B(_0224_),
    .X(_0288_));
 sky130_fd_sc_hd__or4_1 _0990_ (.A(_0252_),
    .B(_0256_),
    .C(_0264_),
    .D(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__or4_1 _0991_ (.A(_0694_),
    .B(_0039_),
    .C(_0086_),
    .D(_0114_),
    .X(_0290_));
 sky130_fd_sc_hd__or4_1 _0992_ (.A(_0067_),
    .B(_0110_),
    .C(_0180_),
    .D(_0182_),
    .X(_0291_));
 sky130_fd_sc_hd__or3_1 _0993_ (.A(_0289_),
    .B(_0290_),
    .C(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__or3_1 _0994_ (.A(_0046_),
    .B(_0186_),
    .C(_0188_),
    .X(_0293_));
 sky130_fd_sc_hd__or2_2 _0995_ (.A(_0074_),
    .B(_0134_),
    .X(_0294_));
 sky130_fd_sc_hd__or3_1 _0996_ (.A(_0125_),
    .B(_0128_),
    .C(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__or4_1 _0997_ (.A(_0081_),
    .B(_0138_),
    .C(_0246_),
    .D(_0247_),
    .X(_0296_));
 sky130_fd_sc_hd__or3_1 _0998_ (.A(_0211_),
    .B(_0230_),
    .C(_0233_),
    .X(_0297_));
 sky130_fd_sc_hd__or4_1 _0999_ (.A(_0156_),
    .B(_0164_),
    .C(_0195_),
    .D(_0202_),
    .X(_0298_));
 sky130_fd_sc_hd__or4_1 _1000_ (.A(_0122_),
    .B(_0132_),
    .C(_0151_),
    .D(_0201_),
    .X(_0299_));
 sky130_fd_sc_hd__or3_2 _1001_ (.A(_0173_),
    .B(_0174_),
    .C(_0176_),
    .X(_0300_));
 sky130_fd_sc_hd__or4_1 _1002_ (.A(_0297_),
    .B(_0298_),
    .C(_0299_),
    .D(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__or4_1 _1003_ (.A(_0293_),
    .B(_0295_),
    .C(_0296_),
    .D(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__or3_1 _1004_ (.A(_0287_),
    .B(_0292_),
    .C(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__a22o_1 _1005_ (.A1(net163),
    .A2(net138),
    .B1(net45),
    .B2(_0303_),
    .X(_0000_));
 sky130_fd_sc_hd__or4_1 _1006_ (.A(_0186_),
    .B(_0187_),
    .C(_0237_),
    .D(_0240_),
    .X(_0304_));
 sky130_fd_sc_hd__or3_1 _1007_ (.A(_0706_),
    .B(_0056_),
    .C(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__or3_1 _1008_ (.A(_0072_),
    .B(_0128_),
    .C(_0129_),
    .X(_0306_));
 sky130_fd_sc_hd__or2_1 _1009_ (.A(_0173_),
    .B(_0175_),
    .X(_0307_));
 sky130_fd_sc_hd__or3_1 _1010_ (.A(_0173_),
    .B(_0175_),
    .C(_0176_),
    .X(_0308_));
 sky130_fd_sc_hd__or3_1 _1011_ (.A(_0305_),
    .B(_0306_),
    .C(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__or2_1 _1012_ (.A(_0686_),
    .B(_0119_),
    .X(_0310_));
 sky130_fd_sc_hd__or2_1 _1013_ (.A(_0258_),
    .B(_0262_),
    .X(_0311_));
 sky130_fd_sc_hd__nand2b_1 _1014_ (.A_N(_0194_),
    .B(_0267_),
    .Y(_0312_));
 sky130_fd_sc_hd__or3_1 _1015_ (.A(_0068_),
    .B(_0099_),
    .C(_0100_),
    .X(_0313_));
 sky130_fd_sc_hd__or3_1 _1016_ (.A(_0163_),
    .B(_0166_),
    .C(_0168_),
    .X(_0314_));
 sky130_fd_sc_hd__or2_1 _1017_ (.A(_0247_),
    .B(_0250_),
    .X(_0315_));
 sky130_fd_sc_hd__or4_1 _1018_ (.A(_0036_),
    .B(_0044_),
    .C(net48),
    .D(_0081_),
    .X(_0316_));
 sky130_fd_sc_hd__or3_1 _1019_ (.A(_0084_),
    .B(_0086_),
    .C(_0087_),
    .X(_0317_));
 sky130_fd_sc_hd__or4_1 _1020_ (.A(_0313_),
    .B(_0314_),
    .C(_0315_),
    .D(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__or4_1 _1021_ (.A(_0223_),
    .B(_0310_),
    .C(_0311_),
    .D(_0312_),
    .X(_0319_));
 sky130_fd_sc_hd__or3_1 _1022_ (.A(_0115_),
    .B(_0316_),
    .C(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__or4_1 _1023_ (.A(_0109_),
    .B(_0220_),
    .C(_0232_),
    .D(_0235_),
    .X(_0321_));
 sky130_fd_sc_hd__or4_1 _1024_ (.A(_0074_),
    .B(_0075_),
    .C(_0149_),
    .D(_0196_),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _1025_ (.A(_0096_),
    .B(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__or4_1 _1026_ (.A(_0696_),
    .B(_0157_),
    .C(_0206_),
    .D(_0278_),
    .X(_0324_));
 sky130_fd_sc_hd__or4_1 _1027_ (.A(_0299_),
    .B(_0321_),
    .C(_0323_),
    .D(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__or4_1 _1028_ (.A(_0309_),
    .B(_0318_),
    .C(_0320_),
    .D(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__a22o_1 _1029_ (.A1(net136),
    .A2(net144),
    .B1(net43),
    .B2(_0326_),
    .X(_0001_));
 sky130_fd_sc_hd__or2_1 _1030_ (.A(_0067_),
    .B(_0256_),
    .X(_0327_));
 sky130_fd_sc_hd__or2_1 _1031_ (.A(_0062_),
    .B(_0084_),
    .X(_0328_));
 sky130_fd_sc_hd__or2_1 _1032_ (.A(_0327_),
    .B(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__nand2b_1 _1033_ (.A_N(_0262_),
    .B(_0272_),
    .Y(_0330_));
 sky130_fd_sc_hd__or4_1 _1034_ (.A(_0074_),
    .B(_0075_),
    .C(_0132_),
    .D(_0151_),
    .X(_0331_));
 sky130_fd_sc_hd__or3_1 _1035_ (.A(net46),
    .B(_0182_),
    .C(_0187_),
    .X(_0332_));
 sky130_fd_sc_hd__or4_1 _1036_ (.A(_0090_),
    .B(_0091_),
    .C(_0111_),
    .D(_0114_),
    .X(_0333_));
 sky130_fd_sc_hd__or2_1 _1037_ (.A(_0332_),
    .B(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__or4_1 _1038_ (.A(_0237_),
    .B(_0241_),
    .C(_0252_),
    .D(_0253_),
    .X(_0335_));
 sky130_fd_sc_hd__or3_1 _1039_ (.A(_0246_),
    .B(_0248_),
    .C(_0249_),
    .X(_0336_));
 sky130_fd_sc_hd__or4_1 _1040_ (.A(_0691_),
    .B(_0699_),
    .C(_0055_),
    .D(_0308_),
    .X(_0337_));
 sky130_fd_sc_hd__or4_2 _1041_ (.A(_0232_),
    .B(_0233_),
    .C(_0336_),
    .D(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__or3_1 _1042_ (.A(_0125_),
    .B(_0128_),
    .C(_0129_),
    .X(_0339_));
 sky130_fd_sc_hd__or3_1 _1043_ (.A(net47),
    .B(_0099_),
    .C(_0100_),
    .X(_0340_));
 sky130_fd_sc_hd__or3_1 _1044_ (.A(_0071_),
    .B(_0072_),
    .C(_0138_),
    .X(_0341_));
 sky130_fd_sc_hd__or4_1 _1045_ (.A(_0082_),
    .B(_0331_),
    .C(_0335_),
    .D(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__or3_1 _1046_ (.A(_0169_),
    .B(_0339_),
    .C(_0340_),
    .X(_0343_));
 sky130_fd_sc_hd__or4_1 _1047_ (.A(_0109_),
    .B(_0158_),
    .C(_0260_),
    .D(_0330_),
    .X(_0344_));
 sky130_fd_sc_hd__or4_1 _1048_ (.A(_0329_),
    .B(_0334_),
    .C(_0343_),
    .D(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__or3_1 _1049_ (.A(_0338_),
    .B(_0342_),
    .C(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__a22o_1 _1050_ (.A1(net136),
    .A2(net146),
    .B1(net43),
    .B2(_0346_),
    .X(_0002_));
 sky130_fd_sc_hd__or2_1 _1051_ (.A(_0240_),
    .B(_0253_),
    .X(_0347_));
 sky130_fd_sc_hd__or2_1 _1052_ (.A(_0080_),
    .B(_0184_),
    .X(_0348_));
 sky130_fd_sc_hd__nor3_1 _1053_ (.A(_0686_),
    .B(_0691_),
    .C(_0694_),
    .Y(_0349_));
 sky130_fd_sc_hd__or3b_1 _1054_ (.A(_0269_),
    .B(_0273_),
    .C_N(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__or3_1 _1055_ (.A(_0118_),
    .B(_0119_),
    .C(_0122_),
    .X(_0351_));
 sky130_fd_sc_hd__or2_1 _1056_ (.A(_0174_),
    .B(_0177_),
    .X(_0352_));
 sky130_fd_sc_hd__or2_1 _1057_ (.A(_0072_),
    .B(_0139_),
    .X(_0353_));
 sky130_fd_sc_hd__or3_2 _1058_ (.A(_0072_),
    .B(_0138_),
    .C(_0139_),
    .X(_0354_));
 sky130_fd_sc_hd__or3_2 _1059_ (.A(_0084_),
    .B(_0085_),
    .C(_0086_),
    .X(_0355_));
 sky130_fd_sc_hd__or3_1 _1060_ (.A(_0064_),
    .B(_0148_),
    .C(_0149_),
    .X(_0356_));
 sky130_fd_sc_hd__or4_1 _1061_ (.A(_0172_),
    .B(_0226_),
    .C(_0339_),
    .D(_0351_),
    .X(_0357_));
 sky130_fd_sc_hd__or4_1 _1062_ (.A(_0057_),
    .B(_0230_),
    .C(_0238_),
    .D(_0258_),
    .X(_0358_));
 sky130_fd_sc_hd__or4_1 _1063_ (.A(_0107_),
    .B(_0113_),
    .C(_0154_),
    .D(_0203_),
    .X(_0359_));
 sky130_fd_sc_hd__or4_1 _1064_ (.A(_0036_),
    .B(_0077_),
    .C(net47),
    .D(_0136_),
    .X(_0360_));
 sky130_fd_sc_hd__or4_1 _1065_ (.A(_0357_),
    .B(_0358_),
    .C(_0359_),
    .D(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__or4_1 _1066_ (.A(_0180_),
    .B(_0352_),
    .C(_0354_),
    .D(_0356_),
    .X(_0362_));
 sky130_fd_sc_hd__or4_1 _1067_ (.A(_0194_),
    .B(_0195_),
    .C(_0250_),
    .D(_0294_),
    .X(_0363_));
 sky130_fd_sc_hd__or4_1 _1068_ (.A(_0216_),
    .B(_0284_),
    .C(_0347_),
    .D(_0348_),
    .X(_0364_));
 sky130_fd_sc_hd__or4_1 _1069_ (.A(_0327_),
    .B(_0350_),
    .C(_0363_),
    .D(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__or4_1 _1070_ (.A(_0355_),
    .B(_0361_),
    .C(_0362_),
    .D(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__a22o_1 _1071_ (.A1(net136),
    .A2(net151),
    .B1(net43),
    .B2(_0366_),
    .X(_0003_));
 sky130_fd_sc_hd__or4_1 _1072_ (.A(_0084_),
    .B(_0085_),
    .C(_0158_),
    .D(_0220_),
    .X(_0367_));
 sky130_fd_sc_hd__nand2_1 _1073_ (.A(_0267_),
    .B(_0272_),
    .Y(_0368_));
 sky130_fd_sc_hd__or3_1 _1074_ (.A(_0193_),
    .B(_0197_),
    .C(_0269_),
    .X(_0369_));
 sky130_fd_sc_hd__or3_1 _1075_ (.A(_0367_),
    .B(_0368_),
    .C(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__or3_1 _1076_ (.A(_0259_),
    .B(_0263_),
    .C(_0336_),
    .X(_0371_));
 sky130_fd_sc_hd__or3_1 _1077_ (.A(_0067_),
    .B(net47),
    .C(_0101_),
    .X(_0372_));
 sky130_fd_sc_hd__or2_1 _1078_ (.A(_0126_),
    .B(_0238_),
    .X(_0373_));
 sky130_fd_sc_hd__or2_1 _1079_ (.A(_0104_),
    .B(_0139_),
    .X(_0374_));
 sky130_fd_sc_hd__or2_1 _1080_ (.A(_0121_),
    .B(_0128_),
    .X(_0375_));
 sky130_fd_sc_hd__or3_1 _1081_ (.A(_0699_),
    .B(_0702_),
    .C(_0052_),
    .X(_0376_));
 sky130_fd_sc_hd__or3_1 _1082_ (.A(_0186_),
    .B(_0187_),
    .C(_0189_),
    .X(_0377_));
 sky130_fd_sc_hd__or4_2 _1083_ (.A(_0231_),
    .B(_0233_),
    .C(_0253_),
    .D(_0256_),
    .X(_0378_));
 sky130_fd_sc_hd__or4_1 _1084_ (.A(_0173_),
    .B(_0174_),
    .C(_0183_),
    .D(_0184_),
    .X(_0379_));
 sky130_fd_sc_hd__or4_1 _1085_ (.A(_0092_),
    .B(_0094_),
    .C(_0376_),
    .D(_0377_),
    .X(_0380_));
 sky130_fd_sc_hd__or4_1 _1086_ (.A(_0046_),
    .B(_0171_),
    .C(_0294_),
    .D(_0373_),
    .X(_0381_));
 sky130_fd_sc_hd__or4_1 _1087_ (.A(_0691_),
    .B(_0225_),
    .C(_0374_),
    .D(_0375_),
    .X(_0382_));
 sky130_fd_sc_hd__or4_1 _1088_ (.A(_0371_),
    .B(_0372_),
    .C(_0381_),
    .D(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__or3_1 _1089_ (.A(_0122_),
    .B(_0131_),
    .C(_0149_),
    .X(_0384_));
 sky130_fd_sc_hd__or3_1 _1090_ (.A(_0064_),
    .B(_0079_),
    .C(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__or2_1 _1091_ (.A(_0115_),
    .B(_0378_),
    .X(_0386_));
 sky130_fd_sc_hd__or4_1 _1092_ (.A(_0379_),
    .B(_0380_),
    .C(_0385_),
    .D(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__or3_1 _1093_ (.A(_0370_),
    .B(_0383_),
    .C(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__a22o_1 _1094_ (.A1(net135),
    .A2(net159),
    .B1(net42),
    .B2(_0388_),
    .X(_0004_));
 sky130_fd_sc_hd__or3_1 _1095_ (.A(_0230_),
    .B(_0235_),
    .C(_0254_),
    .X(_0389_));
 sky130_fd_sc_hd__or4bb_1 _1096_ (.A(_0686_),
    .B(_0039_),
    .C_N(_0267_),
    .D_N(_0268_),
    .X(_0390_));
 sky130_fd_sc_hd__or3b_1 _1097_ (.A(_0090_),
    .B(_0091_),
    .C_N(_0271_),
    .X(_0391_));
 sky130_fd_sc_hd__or2_1 _1098_ (.A(_0390_),
    .B(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__or2_1 _1099_ (.A(_0212_),
    .B(_0225_),
    .X(_0393_));
 sky130_fd_sc_hd__or2_1 _1100_ (.A(_0222_),
    .B(_0224_),
    .X(_0394_));
 sky130_fd_sc_hd__or3_1 _1101_ (.A(_0246_),
    .B(_0247_),
    .C(_0249_),
    .X(_0395_));
 sky130_fd_sc_hd__or4_1 _1102_ (.A(_0130_),
    .B(_0211_),
    .C(_0237_),
    .D(_0261_),
    .X(_0396_));
 sky130_fd_sc_hd__or2_1 _1103_ (.A(_0075_),
    .B(_0294_),
    .X(_0397_));
 sky130_fd_sc_hd__or2_1 _1104_ (.A(_0131_),
    .B(_0137_),
    .X(_0398_));
 sky130_fd_sc_hd__or3_1 _1105_ (.A(_0131_),
    .B(_0132_),
    .C(_0137_),
    .X(_0399_));
 sky130_fd_sc_hd__or3_1 _1106_ (.A(_0205_),
    .B(_0395_),
    .C(_0397_),
    .X(_0400_));
 sky130_fd_sc_hd__or4_1 _1107_ (.A(_0307_),
    .B(_0311_),
    .C(_0393_),
    .D(_0394_),
    .X(_0401_));
 sky130_fd_sc_hd__or4_1 _1108_ (.A(_0082_),
    .B(_0108_),
    .C(_0351_),
    .D(_0399_),
    .X(_0402_));
 sky130_fd_sc_hd__or4_1 _1109_ (.A(_0161_),
    .B(_0313_),
    .C(_0396_),
    .D(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__or4_1 _1110_ (.A(_0049_),
    .B(_0163_),
    .C(_0183_),
    .D(_0193_),
    .X(_0404_));
 sky130_fd_sc_hd__or4_1 _1111_ (.A(_0688_),
    .B(_0071_),
    .C(_0085_),
    .D(_0110_),
    .X(_0405_));
 sky130_fd_sc_hd__or2_1 _1112_ (.A(_0404_),
    .B(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__or4_1 _1113_ (.A(_0389_),
    .B(_0392_),
    .C(_0401_),
    .D(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__or3_1 _1114_ (.A(_0400_),
    .B(_0403_),
    .C(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__a22o_1 _1115_ (.A1(net137),
    .A2(net157),
    .B1(net44),
    .B2(_0408_),
    .X(_0005_));
 sky130_fd_sc_hd__or3_1 _1116_ (.A(_0211_),
    .B(_0212_),
    .C(_0213_),
    .X(_0409_));
 sky130_fd_sc_hd__or2_1 _1117_ (.A(_0200_),
    .B(_0203_),
    .X(_0410_));
 sky130_fd_sc_hd__or3_1 _1118_ (.A(_0202_),
    .B(_0409_),
    .C(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__or3_2 _1119_ (.A(_0221_),
    .B(_0224_),
    .C(_0225_),
    .X(_0412_));
 sky130_fd_sc_hd__or3_1 _1120_ (.A(_0049_),
    .B(_0286_),
    .C(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__or2_1 _1121_ (.A(_0702_),
    .B(_0137_),
    .X(_0414_));
 sky130_fd_sc_hd__or2_2 _1122_ (.A(_0188_),
    .B(_0247_),
    .X(_0415_));
 sky130_fd_sc_hd__or2_1 _1123_ (.A(_0182_),
    .B(_0183_),
    .X(_0416_));
 sky130_fd_sc_hd__or2_1 _1124_ (.A(_0241_),
    .B(_0256_),
    .X(_0417_));
 sky130_fd_sc_hd__or2_1 _1125_ (.A(_0118_),
    .B(_0187_),
    .X(_0418_));
 sky130_fd_sc_hd__or4_1 _1126_ (.A(_0706_),
    .B(_0101_),
    .C(_0197_),
    .D(_0330_),
    .X(_0419_));
 sky130_fd_sc_hd__or4_1 _1127_ (.A(net48),
    .B(_0103_),
    .C(_0111_),
    .D(net46),
    .X(_0420_));
 sky130_fd_sc_hd__or4_1 _1128_ (.A(_0066_),
    .B(_0067_),
    .C(_0127_),
    .D(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__or4_1 _1129_ (.A(_0094_),
    .B(_0415_),
    .C(_0416_),
    .D(_0417_),
    .X(_0422_));
 sky130_fd_sc_hd__or3_1 _1130_ (.A(_0165_),
    .B(_0414_),
    .C(_0418_),
    .X(_0423_));
 sky130_fd_sc_hd__or4_1 _1131_ (.A(_0419_),
    .B(_0421_),
    .C(_0422_),
    .D(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__or3_1 _1132_ (.A(_0080_),
    .B(_0081_),
    .C(_0353_),
    .X(_0425_));
 sky130_fd_sc_hd__or2_1 _1133_ (.A(_0044_),
    .B(_0046_),
    .X(_0426_));
 sky130_fd_sc_hd__or4_1 _1134_ (.A(_0698_),
    .B(_0300_),
    .C(_0425_),
    .D(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__or3_1 _1135_ (.A(_0160_),
    .B(_0411_),
    .C(_0413_),
    .X(_0428_));
 sky130_fd_sc_hd__or3_1 _1136_ (.A(_0424_),
    .B(_0427_),
    .C(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__a22o_1 _1137_ (.A1(net135),
    .A2(net169),
    .B1(net42),
    .B2(_0429_),
    .X(_0006_));
 sky130_fd_sc_hd__or2_1 _1138_ (.A(_0697_),
    .B(_0040_),
    .X(_0430_));
 sky130_fd_sc_hd__or3_1 _1139_ (.A(_0113_),
    .B(_0114_),
    .C(_0222_),
    .X(_0431_));
 sky130_fd_sc_hd__or4_1 _1140_ (.A(_0104_),
    .B(_0107_),
    .C(_0216_),
    .D(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__or2_1 _1141_ (.A(_0193_),
    .B(_0249_),
    .X(_0433_));
 sky130_fd_sc_hd__or3_1 _1142_ (.A(_0077_),
    .B(net48),
    .C(_0080_),
    .X(_0434_));
 sky130_fd_sc_hd__or4_1 _1143_ (.A(_0205_),
    .B(_0232_),
    .C(_0253_),
    .D(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__or4_1 _1144_ (.A(_0285_),
    .B(_0306_),
    .C(_0308_),
    .D(_0377_),
    .X(_0436_));
 sky130_fd_sc_hd__or4_1 _1145_ (.A(_0095_),
    .B(_0123_),
    .C(_0152_),
    .D(_0171_),
    .X(_0437_));
 sky130_fd_sc_hd__or4_1 _1146_ (.A(_0056_),
    .B(_0239_),
    .C(_0273_),
    .D(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__or4_1 _1147_ (.A(_0193_),
    .B(_0194_),
    .C(_0249_),
    .D(_0259_),
    .X(_0439_));
 sky130_fd_sc_hd__or4_1 _1148_ (.A(_0099_),
    .B(_0118_),
    .C(_0132_),
    .D(_0138_),
    .X(_0440_));
 sky130_fd_sc_hd__or4_1 _1149_ (.A(_0062_),
    .B(_0075_),
    .C(_0085_),
    .D(_0180_),
    .X(_0441_));
 sky130_fd_sc_hd__or4_1 _1150_ (.A(_0161_),
    .B(_0439_),
    .C(_0440_),
    .D(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__or3_1 _1151_ (.A(_0435_),
    .B(_0436_),
    .C(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__or4_1 _1152_ (.A(_0430_),
    .B(_0432_),
    .C(_0438_),
    .D(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__a22o_1 _1153_ (.A1(net136),
    .A2(net158),
    .B1(net43),
    .B2(_0444_),
    .X(_0007_));
 sky130_fd_sc_hd__or4_1 _1154_ (.A(_0101_),
    .B(_0169_),
    .C(_0232_),
    .D(_0328_),
    .X(_0445_));
 sky130_fd_sc_hd__or2_1 _1155_ (.A(_0704_),
    .B(_0164_),
    .X(_0446_));
 sky130_fd_sc_hd__or3_1 _1156_ (.A(_0071_),
    .B(_0138_),
    .C(_0139_),
    .X(_0447_));
 sky130_fd_sc_hd__or3_1 _1157_ (.A(_0148_),
    .B(_0149_),
    .C(_0151_),
    .X(_0448_));
 sky130_fd_sc_hd__or4_1 _1158_ (.A(_0054_),
    .B(_0127_),
    .C(_0129_),
    .D(_0447_),
    .X(_0449_));
 sky130_fd_sc_hd__or4_1 _1159_ (.A(_0094_),
    .B(_0270_),
    .C(_0393_),
    .D(_0446_),
    .X(_0450_));
 sky130_fd_sc_hd__or4_1 _1160_ (.A(_0147_),
    .B(_0156_),
    .C(_0188_),
    .D(_0195_),
    .X(_0451_));
 sky130_fd_sc_hd__or4_1 _1161_ (.A(_0703_),
    .B(_0074_),
    .C(_0087_),
    .D(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__or4_1 _1162_ (.A(_0697_),
    .B(_0108_),
    .C(_0115_),
    .D(_0205_),
    .X(_0453_));
 sky130_fd_sc_hd__or4_1 _1163_ (.A(_0241_),
    .B(_0246_),
    .C(_0256_),
    .D(_0261_),
    .X(_0454_));
 sky130_fd_sc_hd__or4_1 _1164_ (.A(_0124_),
    .B(_0300_),
    .C(_0316_),
    .D(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__or4_1 _1165_ (.A(_0448_),
    .B(_0449_),
    .C(_0453_),
    .D(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__or4_1 _1166_ (.A(_0445_),
    .B(_0450_),
    .C(_0452_),
    .D(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__a22o_1 _1167_ (.A1(net137),
    .A2(net149),
    .B1(net44),
    .B2(_0457_),
    .X(_0008_));
 sky130_fd_sc_hd__or2_2 _1168_ (.A(_0110_),
    .B(_0113_),
    .X(_0458_));
 sky130_fd_sc_hd__or2_1 _1169_ (.A(_0147_),
    .B(_0154_),
    .X(_0459_));
 sky130_fd_sc_hd__or3_1 _1170_ (.A(_0221_),
    .B(_0222_),
    .C(_0224_),
    .X(_0460_));
 sky130_fd_sc_hd__or3_1 _1171_ (.A(_0063_),
    .B(_0067_),
    .C(_0098_),
    .X(_0461_));
 sky130_fd_sc_hd__or2_1 _1172_ (.A(_0119_),
    .B(_0121_),
    .X(_0462_));
 sky130_fd_sc_hd__or2_1 _1173_ (.A(_0118_),
    .B(_0121_),
    .X(_0463_));
 sky130_fd_sc_hd__or3_2 _1174_ (.A(_0118_),
    .B(_0119_),
    .C(_0121_),
    .X(_0464_));
 sky130_fd_sc_hd__or4_1 _1175_ (.A(_0448_),
    .B(_0460_),
    .C(_0461_),
    .D(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__or4_1 _1176_ (.A(_0174_),
    .B(_0175_),
    .C(_0182_),
    .D(_0200_),
    .X(_0466_));
 sky130_fd_sc_hd__or4_1 _1177_ (.A(_0706_),
    .B(_0055_),
    .C(_0074_),
    .D(_0311_),
    .X(_0467_));
 sky130_fd_sc_hd__or4_1 _1178_ (.A(_0434_),
    .B(_0465_),
    .C(_0466_),
    .D(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__or3_1 _1179_ (.A(_0047_),
    .B(_0127_),
    .C(_0129_),
    .X(_0469_));
 sky130_fd_sc_hd__or4_1 _1180_ (.A(_0688_),
    .B(_0694_),
    .C(_0236_),
    .D(_0458_),
    .X(_0470_));
 sky130_fd_sc_hd__or4_1 _1181_ (.A(_0283_),
    .B(_0459_),
    .C(_0469_),
    .D(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__or4_1 _1182_ (.A(_0107_),
    .B(_0194_),
    .C(_0212_),
    .D(_0314_),
    .X(_0472_));
 sky130_fd_sc_hd__or4_1 _1183_ (.A(_0071_),
    .B(_0084_),
    .C(_0086_),
    .D(_0219_),
    .X(_0473_));
 sky130_fd_sc_hd__or4_1 _1184_ (.A(_0274_),
    .B(_0415_),
    .C(_0472_),
    .D(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__or3_1 _1185_ (.A(_0468_),
    .B(_0471_),
    .C(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__a22o_1 _1186_ (.A1(net137),
    .A2(net161),
    .B1(net44),
    .B2(_0475_),
    .X(_0009_));
 sky130_fd_sc_hd__or3_1 _1187_ (.A(_0091_),
    .B(_0173_),
    .C(_0174_),
    .X(_0476_));
 sky130_fd_sc_hd__or4_1 _1188_ (.A(_0094_),
    .B(_0131_),
    .C(_0163_),
    .D(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__or2_1 _1189_ (.A(_0168_),
    .B(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__or4_1 _1190_ (.A(_0052_),
    .B(_0053_),
    .C(_0067_),
    .D(_0099_),
    .X(_0479_));
 sky130_fd_sc_hd__or4_1 _1191_ (.A(_0103_),
    .B(_0114_),
    .C(_0284_),
    .D(_0373_),
    .X(_0480_));
 sky130_fd_sc_hd__or3_1 _1192_ (.A(_0079_),
    .B(_0278_),
    .C(_0479_),
    .X(_0481_));
 sky130_fd_sc_hd__or2_1 _1193_ (.A(_0182_),
    .B(_0184_),
    .X(_0482_));
 sky130_fd_sc_hd__or4_1 _1194_ (.A(net46),
    .B(_0250_),
    .C(_0462_),
    .D(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__or4_1 _1195_ (.A(_0411_),
    .B(_0480_),
    .C(_0481_),
    .D(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__or4_1 _1196_ (.A(_0193_),
    .B(_0196_),
    .C(_0258_),
    .D(_0259_),
    .X(_0485_));
 sky130_fd_sc_hd__or3_1 _1197_ (.A(_0221_),
    .B(_0222_),
    .C(_0225_),
    .X(_0486_));
 sky130_fd_sc_hd__or4_1 _1198_ (.A(_0686_),
    .B(_0695_),
    .C(_0485_),
    .D(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__or4_1 _1199_ (.A(_0088_),
    .B(_0147_),
    .C(_0194_),
    .D(_0261_),
    .X(_0488_));
 sky130_fd_sc_hd__or4_1 _1200_ (.A(_0276_),
    .B(_0397_),
    .C(_0487_),
    .D(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__or4_1 _1201_ (.A(_0293_),
    .B(_0478_),
    .C(_0484_),
    .D(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__a22o_1 _1202_ (.A1(net137),
    .A2(net168),
    .B1(net44),
    .B2(_0490_),
    .X(_0010_));
 sky130_fd_sc_hd__or2_1 _1203_ (.A(_0243_),
    .B(_0265_),
    .X(_0491_));
 sky130_fd_sc_hd__or4_1 _1204_ (.A(_0096_),
    .B(_0102_),
    .C(_0285_),
    .D(_0286_),
    .X(_0492_));
 sky130_fd_sc_hd__or2_1 _1205_ (.A(_0066_),
    .B(net48),
    .X(_0493_));
 sky130_fd_sc_hd__or4_1 _1206_ (.A(_0127_),
    .B(_0133_),
    .C(_0294_),
    .D(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__or4_1 _1207_ (.A(_0173_),
    .B(_0188_),
    .C(_0196_),
    .D(_0201_),
    .X(_0495_));
 sky130_fd_sc_hd__or3_1 _1208_ (.A(_0389_),
    .B(_0432_),
    .C(_0483_),
    .X(_0496_));
 sky130_fd_sc_hd__or4_1 _1209_ (.A(_0356_),
    .B(_0390_),
    .C(_0447_),
    .D(_0491_),
    .X(_0497_));
 sky130_fd_sc_hd__or4_1 _1210_ (.A(_0161_),
    .B(_0492_),
    .C(_0494_),
    .D(_0495_),
    .X(_0498_));
 sky130_fd_sc_hd__or3_1 _1211_ (.A(_0496_),
    .B(_0497_),
    .C(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__a22o_1 _1212_ (.A1(net135),
    .A2(net164),
    .B1(net42),
    .B2(_0499_),
    .X(_0011_));
 sky130_fd_sc_hd__or3_1 _1213_ (.A(_0702_),
    .B(_0705_),
    .C(_0106_),
    .X(_0500_));
 sky130_fd_sc_hd__or3_1 _1214_ (.A(_0105_),
    .B(_0242_),
    .C(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__or2_1 _1215_ (.A(_0134_),
    .B(_0317_),
    .X(_0502_));
 sky130_fd_sc_hd__or3_2 _1216_ (.A(_0148_),
    .B(_0149_),
    .C(_0150_),
    .X(_0503_));
 sky130_fd_sc_hd__or3_1 _1217_ (.A(_0399_),
    .B(_0426_),
    .C(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__or4_1 _1218_ (.A(_0695_),
    .B(_0327_),
    .C(_0353_),
    .D(_0410_),
    .X(_0505_));
 sky130_fd_sc_hd__or4_1 _1219_ (.A(_0193_),
    .B(_0218_),
    .C(_0269_),
    .D(_0286_),
    .X(_0506_));
 sky130_fd_sc_hd__or4_1 _1220_ (.A(_0501_),
    .B(_0502_),
    .C(_0505_),
    .D(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__or3_1 _1221_ (.A(_0092_),
    .B(_0094_),
    .C(_0185_),
    .X(_0508_));
 sky130_fd_sc_hd__or3_1 _1222_ (.A(_0315_),
    .B(_0340_),
    .C(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__or4_1 _1223_ (.A(_0071_),
    .B(_0081_),
    .C(_0224_),
    .D(_0225_),
    .X(_0510_));
 sky130_fd_sc_hd__or4_1 _1224_ (.A(_0111_),
    .B(_0119_),
    .C(_0173_),
    .D(_0231_),
    .X(_0511_));
 sky130_fd_sc_hd__or2_1 _1225_ (.A(_0130_),
    .B(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__or4_1 _1226_ (.A(_0171_),
    .B(_0265_),
    .C(_0510_),
    .D(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__or4_1 _1227_ (.A(_0504_),
    .B(_0507_),
    .C(_0509_),
    .D(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__a22o_1 _1228_ (.A1(net135),
    .A2(net166),
    .B1(net42),
    .B2(_0514_),
    .X(_0012_));
 sky130_fd_sc_hd__or3_1 _1229_ (.A(_0048_),
    .B(_0049_),
    .C(_0053_),
    .X(_0515_));
 sky130_fd_sc_hd__or2_1 _1230_ (.A(_0103_),
    .B(_0182_),
    .X(_0516_));
 sky130_fd_sc_hd__or4_1 _1231_ (.A(_0205_),
    .B(_0237_),
    .C(_0238_),
    .D(_0241_),
    .X(_0517_));
 sky130_fd_sc_hd__or4_1 _1232_ (.A(_0099_),
    .B(_0101_),
    .C(_0409_),
    .D(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__or4_1 _1233_ (.A(_0072_),
    .B(_0113_),
    .C(_0114_),
    .D(_0180_),
    .X(_0519_));
 sky130_fd_sc_hd__or4_1 _1234_ (.A(_0230_),
    .B(_0249_),
    .C(_0253_),
    .D(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__or4_1 _1235_ (.A(_0040_),
    .B(_0068_),
    .C(_0223_),
    .D(_0273_),
    .X(_0521_));
 sky130_fd_sc_hd__or4_1 _1236_ (.A(net48),
    .B(_0080_),
    .C(_0459_),
    .D(_0516_),
    .X(_0522_));
 sky130_fd_sc_hd__or4_1 _1237_ (.A(_0477_),
    .B(_0520_),
    .C(_0521_),
    .D(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__or4_1 _1238_ (.A(_0698_),
    .B(_0130_),
    .C(_0285_),
    .D(_0355_),
    .X(_0524_));
 sky130_fd_sc_hd__or4_1 _1239_ (.A(_0397_),
    .B(_0464_),
    .C(_0515_),
    .D(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__or3_1 _1240_ (.A(_0518_),
    .B(_0523_),
    .C(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__a22o_1 _1241_ (.A1(net137),
    .A2(net170),
    .B1(net44),
    .B2(_0526_),
    .X(_0013_));
 sky130_fd_sc_hd__or3b_1 _1242_ (.A(_0230_),
    .B(_0254_),
    .C_N(_0349_),
    .X(_0527_));
 sky130_fd_sc_hd__or4_1 _1243_ (.A(_0093_),
    .B(_0460_),
    .C(_0476_),
    .D(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__or4b_1 _1244_ (.A(_0092_),
    .B(_0103_),
    .C(_0259_),
    .D_N(_0271_),
    .X(_0529_));
 sky130_fd_sc_hd__or3_1 _1245_ (.A(_0056_),
    .B(net48),
    .C(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__or4_1 _1246_ (.A(_0702_),
    .B(_0039_),
    .C(_0398_),
    .D(_0458_),
    .X(_0531_));
 sky130_fd_sc_hd__or4_1 _1247_ (.A(_0151_),
    .B(_0155_),
    .C(_0156_),
    .D(_0269_),
    .X(_0532_));
 sky130_fd_sc_hd__or4_1 _1248_ (.A(_0062_),
    .B(_0085_),
    .C(_0087_),
    .D(_0190_),
    .X(_0533_));
 sky130_fd_sc_hd__or4_1 _1249_ (.A(_0530_),
    .B(_0531_),
    .C(_0532_),
    .D(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__or4_1 _1250_ (.A(_0166_),
    .B(_0168_),
    .C(_0186_),
    .D(_0196_),
    .X(_0535_));
 sky130_fd_sc_hd__or4_1 _1251_ (.A(_0076_),
    .B(_0124_),
    .C(_0251_),
    .D(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__or4_1 _1252_ (.A(_0518_),
    .B(_0528_),
    .C(_0534_),
    .D(_0536_),
    .X(_0537_));
 sky130_fd_sc_hd__a22o_1 _1253_ (.A1(net137),
    .A2(net150),
    .B1(net44),
    .B2(_0537_),
    .X(_0014_));
 sky130_fd_sc_hd__nand2b_1 _1254_ (.A_N(_0189_),
    .B(_0272_),
    .Y(_0538_));
 sky130_fd_sc_hd__or3_1 _1255_ (.A(_0049_),
    .B(_0085_),
    .C(_0237_),
    .X(_0539_));
 sky130_fd_sc_hd__or3_1 _1256_ (.A(_0414_),
    .B(_0538_),
    .C(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__or4_1 _1257_ (.A(_0149_),
    .B(_0168_),
    .C(_0214_),
    .D(_0516_),
    .X(_0541_));
 sky130_fd_sc_hd__or4_1 _1258_ (.A(_0372_),
    .B(_0430_),
    .C(_0540_),
    .D(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__or2_1 _1259_ (.A(_0197_),
    .B(_0410_),
    .X(_0543_));
 sky130_fd_sc_hd__or4_1 _1260_ (.A(_0091_),
    .B(_0095_),
    .C(_0112_),
    .D(_0263_),
    .X(_0544_));
 sky130_fd_sc_hd__or4_1 _1261_ (.A(_0083_),
    .B(_0159_),
    .C(_0354_),
    .D(_0412_),
    .X(_0545_));
 sky130_fd_sc_hd__or4_1 _1262_ (.A(_0464_),
    .B(_0543_),
    .C(_0544_),
    .D(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__or3_1 _1263_ (.A(_0232_),
    .B(_0253_),
    .C(_0395_),
    .X(_0547_));
 sky130_fd_sc_hd__or3_1 _1264_ (.A(_0178_),
    .B(_0295_),
    .C(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__or3_1 _1265_ (.A(_0542_),
    .B(_0546_),
    .C(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__a22o_1 _1266_ (.A1(net136),
    .A2(net156),
    .B1(net43),
    .B2(_0549_),
    .X(_0015_));
 sky130_fd_sc_hd__or4_1 _1267_ (.A(_0688_),
    .B(_0694_),
    .C(_0194_),
    .D(_0195_),
    .X(_0550_));
 sky130_fd_sc_hd__or3_1 _1268_ (.A(_0232_),
    .B(_0234_),
    .C(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__or2_1 _1269_ (.A(_0048_),
    .B(_0125_),
    .X(_0552_));
 sky130_fd_sc_hd__or2_1 _1270_ (.A(_0463_),
    .B(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__or4_2 _1271_ (.A(_0093_),
    .B(_0098_),
    .C(_0129_),
    .D(_0174_),
    .X(_0554_));
 sky130_fd_sc_hd__or2_1 _1272_ (.A(_0237_),
    .B(_0242_),
    .X(_0555_));
 sky130_fd_sc_hd__or4_1 _1273_ (.A(_0069_),
    .B(_0276_),
    .C(_0296_),
    .D(_0332_),
    .X(_0556_));
 sky130_fd_sc_hd__or4_1 _1274_ (.A(_0702_),
    .B(_0039_),
    .C(_0103_),
    .D(_0114_),
    .X(_0557_));
 sky130_fd_sc_hd__or4_1 _1275_ (.A(_0502_),
    .B(_0551_),
    .C(_0553_),
    .D(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__or4_1 _1276_ (.A(_0486_),
    .B(_0503_),
    .C(_0554_),
    .D(_0555_),
    .X(_0559_));
 sky130_fd_sc_hd__or4_1 _1277_ (.A(_0095_),
    .B(_0140_),
    .C(_0147_),
    .D(_0202_),
    .X(_0560_));
 sky130_fd_sc_hd__or4_1 _1278_ (.A(_0214_),
    .B(_0254_),
    .C(_0265_),
    .D(_0446_),
    .X(_0561_));
 sky130_fd_sc_hd__or4_1 _1279_ (.A(_0190_),
    .B(_0556_),
    .C(_0560_),
    .D(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__or3_1 _1280_ (.A(_0558_),
    .B(_0559_),
    .C(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__a22o_1 _1281_ (.A1(net137),
    .A2(net145),
    .B1(net44),
    .B2(_0563_),
    .X(_0016_));
 sky130_fd_sc_hd__or2_1 _1282_ (.A(_0052_),
    .B(_0119_),
    .X(_0564_));
 sky130_fd_sc_hd__or4_1 _1283_ (.A(_0177_),
    .B(_0190_),
    .C(_0288_),
    .D(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__or4_1 _1284_ (.A(_0091_),
    .B(net47),
    .C(_0100_),
    .D(_0134_),
    .X(_0566_));
 sky130_fd_sc_hd__or4_1 _1285_ (.A(_0149_),
    .B(_0183_),
    .C(_0200_),
    .D(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__or4_1 _1286_ (.A(_0204_),
    .B(_0482_),
    .C(_0493_),
    .D(_0552_),
    .X(_0568_));
 sky130_fd_sc_hd__or4_1 _1287_ (.A(_0046_),
    .B(_0170_),
    .C(_0278_),
    .D(_0374_),
    .X(_0569_));
 sky130_fd_sc_hd__or4_1 _1288_ (.A(_0565_),
    .B(_0567_),
    .C(_0568_),
    .D(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__or3_1 _1289_ (.A(_0132_),
    .B(_0136_),
    .C(_0137_),
    .X(_0571_));
 sky130_fd_sc_hd__or4_1 _1290_ (.A(_0111_),
    .B(_0458_),
    .C(_0491_),
    .D(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__or4_1 _1291_ (.A(_0033_),
    .B(_0370_),
    .C(_0570_),
    .D(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__a22o_1 _1292_ (.A1(net135),
    .A2(net152),
    .B1(net42),
    .B2(_0573_),
    .X(_0017_));
 sky130_fd_sc_hd__or3_1 _1293_ (.A(net47),
    .B(_0098_),
    .C(_0348_),
    .X(_0574_));
 sky130_fd_sc_hd__or4_1 _1294_ (.A(_0090_),
    .B(_0128_),
    .C(_0225_),
    .D(_0252_),
    .X(_0575_));
 sky130_fd_sc_hd__or4_1 _1295_ (.A(_0039_),
    .B(_0044_),
    .C(_0085_),
    .D(_0122_),
    .X(_0576_));
 sky130_fd_sc_hd__or4_1 _1296_ (.A(_0462_),
    .B(_0574_),
    .C(_0575_),
    .D(_0576_),
    .X(_0577_));
 sky130_fd_sc_hd__or4_1 _1297_ (.A(_0105_),
    .B(_0186_),
    .C(_0189_),
    .D(_0409_),
    .X(_0578_));
 sky130_fd_sc_hd__or2_1 _1298_ (.A(_0071_),
    .B(_0274_),
    .X(_0579_));
 sky130_fd_sc_hd__or3_1 _1299_ (.A(_0165_),
    .B(_0311_),
    .C(_0331_),
    .X(_0580_));
 sky130_fd_sc_hd__or4_1 _1300_ (.A(_0069_),
    .B(_0115_),
    .C(_0161_),
    .D(_0244_),
    .X(_0581_));
 sky130_fd_sc_hd__or4_1 _1301_ (.A(_0198_),
    .B(_0579_),
    .C(_0580_),
    .D(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__or4_1 _1302_ (.A(_0338_),
    .B(_0577_),
    .C(_0578_),
    .D(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__a22o_1 _1303_ (.A1(net137),
    .A2(net162),
    .B1(net44),
    .B2(_0583_),
    .X(_0018_));
 sky130_fd_sc_hd__or4_1 _1304_ (.A(_0177_),
    .B(_0250_),
    .C(_0410_),
    .D(_0418_),
    .X(_0584_));
 sky130_fd_sc_hd__or3_1 _1305_ (.A(_0049_),
    .B(_0075_),
    .C(_0195_),
    .X(_0585_));
 sky130_fd_sc_hd__or4_1 _1306_ (.A(_0066_),
    .B(_0067_),
    .C(_0152_),
    .D(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__or4_1 _1307_ (.A(_0072_),
    .B(_0081_),
    .C(_0182_),
    .D(_0183_),
    .X(_0587_));
 sky130_fd_sc_hd__or3_1 _1308_ (.A(net47),
    .B(_0101_),
    .C(_0285_),
    .X(_0588_));
 sky130_fd_sc_hd__or4_1 _1309_ (.A(_0091_),
    .B(_0095_),
    .C(_0571_),
    .D(_0587_),
    .X(_0589_));
 sky130_fd_sc_hd__or3_1 _1310_ (.A(_0112_),
    .B(_0263_),
    .C(_0412_),
    .X(_0590_));
 sky130_fd_sc_hd__or4_1 _1311_ (.A(_0555_),
    .B(_0588_),
    .C(_0589_),
    .D(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__or2_1 _1312_ (.A(_0047_),
    .B(_0130_),
    .X(_0592_));
 sky130_fd_sc_hd__or4_1 _1313_ (.A(_0350_),
    .B(_0367_),
    .C(_0584_),
    .D(_0586_),
    .X(_0593_));
 sky130_fd_sc_hd__or3_1 _1314_ (.A(_0591_),
    .B(_0592_),
    .C(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__a22o_1 _1315_ (.A1(net135),
    .A2(net160),
    .B1(net42),
    .B2(_0594_),
    .X(_0019_));
 sky130_fd_sc_hd__or2_1 _1316_ (.A(_0077_),
    .B(_0224_),
    .X(_0595_));
 sky130_fd_sc_hd__or3_1 _1317_ (.A(_0398_),
    .B(_0415_),
    .C(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__or4_1 _1318_ (.A(_0099_),
    .B(_0100_),
    .C(_0202_),
    .D(_0203_),
    .X(_0597_));
 sky130_fd_sc_hd__or4_1 _1319_ (.A(_0045_),
    .B(_0080_),
    .C(_0081_),
    .D(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__or3_1 _1320_ (.A(_0236_),
    .B(_0252_),
    .C(_0256_),
    .X(_0599_));
 sky130_fd_sc_hd__or2_1 _1321_ (.A(_0067_),
    .B(_0068_),
    .X(_0600_));
 sky130_fd_sc_hd__or4_1 _1322_ (.A(_0694_),
    .B(_0163_),
    .C(_0175_),
    .D(_0221_),
    .X(_0601_));
 sky130_fd_sc_hd__or4_1 _1323_ (.A(_0341_),
    .B(_0485_),
    .C(_0503_),
    .D(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__or4_1 _1324_ (.A(_0217_),
    .B(_0599_),
    .C(_0600_),
    .D(_0602_),
    .X(_0603_));
 sky130_fd_sc_hd__or4_1 _1325_ (.A(_0305_),
    .B(_0502_),
    .C(_0596_),
    .D(_0598_),
    .X(_0604_));
 sky130_fd_sc_hd__or4_1 _1326_ (.A(_0122_),
    .B(_0126_),
    .C(_0248_),
    .D(_0379_),
    .X(_0605_));
 sky130_fd_sc_hd__or4_1 _1327_ (.A(_0111_),
    .B(_0391_),
    .C(_0458_),
    .D(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__or3_1 _1328_ (.A(_0603_),
    .B(_0604_),
    .C(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__a22o_1 _1329_ (.A1(net135),
    .A2(net143),
    .B1(net42),
    .B2(_0607_),
    .X(_0020_));
 sky130_fd_sc_hd__or2_1 _1330_ (.A(_0032_),
    .B(_0515_),
    .X(_0608_));
 sky130_fd_sc_hd__or4_1 _1331_ (.A(_0198_),
    .B(_0352_),
    .C(_0377_),
    .D(_0461_),
    .X(_0609_));
 sky130_fd_sc_hd__or4_1 _1332_ (.A(_0078_),
    .B(_0081_),
    .C(_0169_),
    .D(_0235_),
    .X(_0610_));
 sky130_fd_sc_hd__or3_1 _1333_ (.A(_0394_),
    .B(_0458_),
    .C(_0482_),
    .X(_0611_));
 sky130_fd_sc_hd__or3_1 _1334_ (.A(_0392_),
    .B(_0608_),
    .C(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__or4_1 _1335_ (.A(_0071_),
    .B(_0075_),
    .C(_0136_),
    .D(_0138_),
    .X(_0613_));
 sky130_fd_sc_hd__or3_1 _1336_ (.A(_0152_),
    .B(_0206_),
    .C(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__or4_1 _1337_ (.A(_0041_),
    .B(_0137_),
    .C(_0148_),
    .D(_0248_),
    .X(_0615_));
 sky130_fd_sc_hd__or4_1 _1338_ (.A(_0109_),
    .B(_0317_),
    .C(_0335_),
    .D(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__or4_1 _1339_ (.A(_0375_),
    .B(_0610_),
    .C(_0614_),
    .D(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__or3_1 _1340_ (.A(_0609_),
    .B(_0612_),
    .C(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__a22o_1 _1341_ (.A1(net135),
    .A2(net155),
    .B1(net42),
    .B2(_0618_),
    .X(_0021_));
 sky130_fd_sc_hd__or2_1 _1342_ (.A(_0092_),
    .B(_0104_),
    .X(_0619_));
 sky130_fd_sc_hd__or4_1 _1343_ (.A(_0140_),
    .B(_0312_),
    .C(_0459_),
    .D(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__or4_1 _1344_ (.A(_0202_),
    .B(_0203_),
    .C(_0224_),
    .D(_0225_),
    .X(_0621_));
 sky130_fd_sc_hd__or4_1 _1345_ (.A(_0036_),
    .B(_0080_),
    .C(_0152_),
    .D(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__or4_1 _1346_ (.A(_0192_),
    .B(_0245_),
    .C(_0620_),
    .D(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__or4_1 _1347_ (.A(_0039_),
    .B(_0044_),
    .C(_0164_),
    .D(_0166_),
    .X(_0624_));
 sky130_fd_sc_hd__or4_1 _1348_ (.A(_0099_),
    .B(_0106_),
    .C(_0111_),
    .D(_0149_),
    .X(_0625_));
 sky130_fd_sc_hd__or3_1 _1349_ (.A(_0213_),
    .B(_0215_),
    .C(_0248_),
    .X(_0626_));
 sky130_fd_sc_hd__or4_1 _1350_ (.A(_0355_),
    .B(_0447_),
    .C(_0625_),
    .D(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__or4_1 _1351_ (.A(_0554_),
    .B(_0600_),
    .C(_0624_),
    .D(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__or3_1 _1352_ (.A(_0608_),
    .B(_0623_),
    .C(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__a22o_1 _1353_ (.A1(net137),
    .A2(net141),
    .B1(net44),
    .B2(_0629_),
    .X(_0022_));
 sky130_fd_sc_hd__or4_1 _1354_ (.A(_0165_),
    .B(_0311_),
    .C(_0550_),
    .D(_0599_),
    .X(_0630_));
 sky130_fd_sc_hd__or4_1 _1355_ (.A(_0045_),
    .B(net48),
    .C(_0080_),
    .D(_0094_),
    .X(_0631_));
 sky130_fd_sc_hd__or4_1 _1356_ (.A(_0124_),
    .B(_0130_),
    .C(_0413_),
    .D(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__or3_1 _1357_ (.A(_0147_),
    .B(_0176_),
    .C(_0249_),
    .X(_0633_));
 sky130_fd_sc_hd__or4_1 _1358_ (.A(_0106_),
    .B(_0107_),
    .C(_0132_),
    .D(_0155_),
    .X(_0634_));
 sky130_fd_sc_hd__or4_1 _1359_ (.A(_0086_),
    .B(_0087_),
    .C(_0136_),
    .D(_0139_),
    .X(_0635_));
 sky130_fd_sc_hd__or4_1 _1360_ (.A(_0153_),
    .B(_0633_),
    .C(_0634_),
    .D(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__or4_1 _1361_ (.A(net47),
    .B(_0098_),
    .C(_0204_),
    .D(_0243_),
    .X(_0637_));
 sky130_fd_sc_hd__or4_1 _1362_ (.A(_0068_),
    .B(_0219_),
    .C(_0284_),
    .D(_0368_),
    .X(_0638_));
 sky130_fd_sc_hd__or4_1 _1363_ (.A(_0112_),
    .B(_0636_),
    .C(_0637_),
    .D(_0638_),
    .X(_0639_));
 sky130_fd_sc_hd__or3_1 _1364_ (.A(_0630_),
    .B(_0632_),
    .C(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__a22o_1 _1365_ (.A1(net135),
    .A2(net165),
    .B1(net42),
    .B2(_0640_),
    .X(_0023_));
 sky130_fd_sc_hd__or3_1 _1366_ (.A(_0334_),
    .B(_0372_),
    .C(_0501_),
    .X(_0641_));
 sky130_fd_sc_hd__or4_1 _1367_ (.A(_0378_),
    .B(_0425_),
    .C(_0543_),
    .D(_0571_),
    .X(_0642_));
 sky130_fd_sc_hd__or4_1 _1368_ (.A(_0036_),
    .B(_0041_),
    .C(_0125_),
    .D(_0128_),
    .X(_0643_));
 sky130_fd_sc_hd__or4_1 _1369_ (.A(_0696_),
    .B(_0247_),
    .C(_0249_),
    .D(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__or3_1 _1370_ (.A(_0049_),
    .B(_0052_),
    .C(_0225_),
    .X(_0645_));
 sky130_fd_sc_hd__or3_1 _1371_ (.A(_0177_),
    .B(_0263_),
    .C(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__or4_1 _1372_ (.A(_0169_),
    .B(_0218_),
    .C(_0463_),
    .D(_0538_),
    .X(_0647_));
 sky130_fd_sc_hd__or4_1 _1373_ (.A(_0160_),
    .B(_0644_),
    .C(_0646_),
    .D(_0647_),
    .X(_0649_));
 sky130_fd_sc_hd__or3_1 _1374_ (.A(_0641_),
    .B(_0642_),
    .C(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__a22o_1 _1375_ (.A1(net135),
    .A2(net142),
    .B1(net42),
    .B2(_0650_),
    .X(_0024_));
 sky130_fd_sc_hd__or4_1 _1376_ (.A(_0699_),
    .B(_0097_),
    .C(_0201_),
    .D(_0246_),
    .X(_0651_));
 sky130_fd_sc_hd__or4_1 _1377_ (.A(_0064_),
    .B(_0120_),
    .C(_0128_),
    .D(_0129_),
    .X(_0652_));
 sky130_fd_sc_hd__or4_1 _1378_ (.A(_0040_),
    .B(_0347_),
    .C(_0433_),
    .D(_0595_),
    .X(_0653_));
 sky130_fd_sc_hd__or4_1 _1379_ (.A(_0162_),
    .B(_0551_),
    .C(_0578_),
    .D(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__or3_1 _1380_ (.A(_0269_),
    .B(_0273_),
    .C(_0651_),
    .X(_0655_));
 sky130_fd_sc_hd__or4_1 _1381_ (.A(_0054_),
    .B(_0111_),
    .C(_0458_),
    .D(_0587_),
    .X(_0656_));
 sky130_fd_sc_hd__or4_1 _1382_ (.A(_0264_),
    .B(_0652_),
    .C(_0655_),
    .D(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__or3_1 _1383_ (.A(_0478_),
    .B(_0654_),
    .C(_0657_),
    .X(_0659_));
 sky130_fd_sc_hd__a22o_1 _1384_ (.A1(net138),
    .A2(net167),
    .B1(net45),
    .B2(_0659_),
    .X(_0025_));
 sky130_fd_sc_hd__or3_1 _1385_ (.A(net46),
    .B(_0354_),
    .C(_0416_),
    .X(_0660_));
 sky130_fd_sc_hd__or4_1 _1386_ (.A(_0079_),
    .B(_0120_),
    .C(_0127_),
    .D(_0232_),
    .X(_0661_));
 sky130_fd_sc_hd__or3_1 _1387_ (.A(_0695_),
    .B(_0275_),
    .C(_0619_),
    .X(_0662_));
 sky130_fd_sc_hd__or4_1 _1388_ (.A(_0162_),
    .B(_0371_),
    .C(_0661_),
    .D(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__or4_1 _1389_ (.A(_0217_),
    .B(_0376_),
    .C(_0431_),
    .D(_0624_),
    .X(_0664_));
 sky130_fd_sc_hd__or4_1 _1390_ (.A(net47),
    .B(_0188_),
    .C(_0238_),
    .D(_0252_),
    .X(_0665_));
 sky130_fd_sc_hd__or4_1 _1391_ (.A(_0069_),
    .B(_0178_),
    .C(_0199_),
    .D(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__or4_1 _1392_ (.A(_0660_),
    .B(_0663_),
    .C(_0664_),
    .D(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__a22o_1 _1393_ (.A1(net138),
    .A2(net153),
    .B1(net45),
    .B2(_0667_),
    .X(_0026_));
 sky130_fd_sc_hd__or2_1 _1394_ (.A(_0244_),
    .B(_0275_),
    .X(_0669_));
 sky130_fd_sc_hd__or2_1 _1395_ (.A(_0686_),
    .B(_0107_),
    .X(_0670_));
 sky130_fd_sc_hd__or4_1 _1396_ (.A(_0120_),
    .B(_0200_),
    .C(_0205_),
    .D(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__or4_1 _1397_ (.A(_0703_),
    .B(_0103_),
    .C(_0106_),
    .D(_0235_),
    .X(_0672_));
 sky130_fd_sc_hd__or4_1 _1398_ (.A(_0660_),
    .B(_0669_),
    .C(_0671_),
    .D(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__or4_1 _1399_ (.A(_0099_),
    .B(_0101_),
    .C(_0226_),
    .D(_0515_),
    .X(_0674_));
 sky130_fd_sc_hd__or4_1 _1400_ (.A(_0179_),
    .B(_0336_),
    .C(_0592_),
    .D(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__or2_1 _1401_ (.A(_0673_),
    .B(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__a22o_1 _1402_ (.A1(net138),
    .A2(net154),
    .B1(net45),
    .B2(_0676_),
    .X(_0027_));
 sky130_fd_sc_hd__or4_1 _1403_ (.A(_0706_),
    .B(_0123_),
    .C(_0184_),
    .D(_0247_),
    .X(_0678_));
 sky130_fd_sc_hd__or4_1 _1404_ (.A(_0109_),
    .B(_0116_),
    .C(_0207_),
    .D(_0669_),
    .X(_0679_));
 sky130_fd_sc_hd__or3_1 _1405_ (.A(_0191_),
    .B(_0266_),
    .C(_0354_),
    .X(_0680_));
 sky130_fd_sc_hd__or4_1 _1406_ (.A(_0698_),
    .B(_0047_),
    .C(_0678_),
    .D(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__or3_1 _1407_ (.A(_0179_),
    .B(_0679_),
    .C(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__a22o_1 _1408_ (.A1(net137),
    .A2(net147),
    .B1(net44),
    .B2(_0682_),
    .X(_0028_));
 sky130_fd_sc_hd__or4_1 _1409_ (.A(_0058_),
    .B(_0083_),
    .C(_0227_),
    .D(_0579_),
    .X(_0683_));
 sky130_fd_sc_hd__or2_1 _1410_ (.A(_0208_),
    .B(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__a22o_1 _1411_ (.A1(net138),
    .A2(net148),
    .B1(net45),
    .B2(_0684_),
    .X(_0029_));
 sky130_fd_sc_hd__o21a_1 _1412_ (.A1(net9),
    .A2(net139),
    .B1(_0280_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _1413_ (.A0(net140),
    .A1(_0144_),
    .S(net9),
    .X(_0031_));
 sky130_fd_sc_hd__dfxtp_1 _1414_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net1),
    .Q(\addr0_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1415_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net2),
    .Q(\addr0_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1416_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net3),
    .Q(\addr0_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1417_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net4),
    .Q(\addr0_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1418_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net5),
    .Q(\addr0_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1419_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net6),
    .Q(\addr0_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1420_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net7),
    .Q(\addr0_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1421_ (.CLK(clknet_2_0__leaf_clk0),
    .D(net8),
    .Q(\addr0_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1422_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0000_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_1 _1423_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0001_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_1 _1424_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0002_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _1425_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0003_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _1426_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0004_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _1427_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0005_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _1428_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0006_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _1429_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0007_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _1430_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0008_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _1431_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0009_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _1432_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0010_),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_1 _1433_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0011_),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_1 _1434_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0012_),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_1 _1435_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0013_),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_1 _1436_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0014_),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_1 _1437_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0015_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_1 _1438_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0016_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_1 _1439_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0017_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_1 _1440_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0018_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_1 _1441_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0019_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_1 _1442_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0020_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_1 _1443_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0021_),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_1 _1444_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0022_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_1 _1445_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0023_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_1 _1446_ (.CLK(clknet_2_2__leaf_clk0),
    .D(_0024_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_1 _1447_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0025_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_1 _1448_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0026_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _1449_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0027_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_1 _1450_ (.CLK(clknet_2_1__leaf_clk0),
    .D(_0028_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _1451_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0029_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _1452_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0030_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _1453_ (.CLK(clknet_2_3__leaf_clk0),
    .D(_0031_),
    .Q(net34));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_345 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(addr0[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(addr0[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(addr0[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(addr0[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(addr0[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(addr0[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(addr0[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(addr0[7]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(cs0),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(dout0[0]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(dout0[10]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(dout0[11]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(dout0[12]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(dout0[13]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(dout0[14]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(dout0[15]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(dout0[16]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(dout0[17]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(dout0[18]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(dout0[19]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(dout0[1]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(dout0[20]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(dout0[21]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(dout0[22]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(dout0[23]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(dout0[24]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(dout0[25]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(dout0[26]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(dout0[27]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(dout0[28]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(dout0[29]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(dout0[2]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(dout0[30]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(dout0[31]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(dout0[3]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(dout0[4]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(dout0[5]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(dout0[6]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(dout0[7]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(dout0[8]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(dout0[9]));
 sky130_fd_sc_hd__buf_2 fanout42 (.A(_0281_),
    .X(net42));
 sky130_fd_sc_hd__buf_1 fanout43 (.A(_0281_),
    .X(net43));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(_0281_),
    .X(net44));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout45 (.A(_0281_),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 max_cap46 (.A(_0180_),
    .X(net46));
 sky130_fd_sc_hd__buf_2 fanout47 (.A(_0097_),
    .X(net47));
 sky130_fd_sc_hd__buf_2 fanout48 (.A(_0078_),
    .X(net48));
 sky130_fd_sc_hd__buf_2 fanout49 (.A(_0229_),
    .X(net49));
 sky130_fd_sc_hd__buf_1 fanout50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 max_cap51 (.A(_0229_),
    .X(net51));
 sky130_fd_sc_hd__buf_2 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 fanout53 (.A(_0228_),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(net57),
    .X(net54));
 sky130_fd_sc_hd__buf_2 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 max_cap56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 wire57 (.A(_0210_),
    .X(net57));
 sky130_fd_sc_hd__buf_4 fanout58 (.A(_0209_),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 fanout59 (.A(_0209_),
    .X(net59));
 sky130_fd_sc_hd__buf_2 fanout60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout61 (.A(_0181_),
    .X(net61));
 sky130_fd_sc_hd__buf_2 fanout62 (.A(_0167_),
    .X(net62));
 sky130_fd_sc_hd__buf_1 fanout63 (.A(_0167_),
    .X(net63));
 sky130_fd_sc_hd__buf_2 fanout64 (.A(_0146_),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 fanout65 (.A(_0146_),
    .X(net65));
 sky130_fd_sc_hd__buf_2 fanout66 (.A(_0145_),
    .X(net66));
 sky130_fd_sc_hd__buf_1 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 max_cap68 (.A(_0145_),
    .X(net68));
 sky130_fd_sc_hd__buf_2 fanout69 (.A(_0073_),
    .X(net69));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout70 (.A(_0073_),
    .X(net70));
 sky130_fd_sc_hd__buf_2 fanout71 (.A(_0070_),
    .X(net71));
 sky130_fd_sc_hd__buf_1 fanout72 (.A(_0070_),
    .X(net72));
 sky130_fd_sc_hd__buf_2 fanout73 (.A(_0065_),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 fanout74 (.A(_0065_),
    .X(net74));
 sky130_fd_sc_hd__buf_2 fanout75 (.A(_0061_),
    .X(net75));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout76 (.A(_0061_),
    .X(net76));
 sky130_fd_sc_hd__buf_2 fanout77 (.A(_0059_),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 fanout78 (.A(_0059_),
    .X(net78));
 sky130_fd_sc_hd__buf_2 fanout79 (.A(_0051_),
    .X(net79));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout80 (.A(_0051_),
    .X(net80));
 sky130_fd_sc_hd__buf_2 fanout81 (.A(net83),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 fanout82 (.A(net84),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 max_cap83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 wire84 (.A(_0043_),
    .X(net84));
 sky130_fd_sc_hd__buf_2 fanout85 (.A(_0042_),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 fanout86 (.A(_0042_),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 fanout87 (.A(_0038_),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 fanout88 (.A(_0038_),
    .X(net88));
 sky130_fd_sc_hd__buf_2 fanout89 (.A(net91),
    .X(net89));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout90 (.A(_0037_),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 max_cap91 (.A(_0037_),
    .X(net91));
 sky130_fd_sc_hd__buf_2 fanout92 (.A(_0035_),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 fanout93 (.A(_0035_),
    .X(net93));
 sky130_fd_sc_hd__buf_2 fanout94 (.A(_0034_),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 fanout95 (.A(_0034_),
    .X(net95));
 sky130_fd_sc_hd__buf_2 fanout96 (.A(_0701_),
    .X(net96));
 sky130_fd_sc_hd__buf_2 fanout97 (.A(_0701_),
    .X(net97));
 sky130_fd_sc_hd__buf_2 fanout98 (.A(net100),
    .X(net98));
 sky130_fd_sc_hd__buf_2 fanout99 (.A(net101),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 wire100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 wire101 (.A(_0700_),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_4 fanout102 (.A(_0693_),
    .X(net102));
 sky130_fd_sc_hd__buf_2 fanout103 (.A(_0693_),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 fanout104 (.A(_0692_),
    .X(net104));
 sky130_fd_sc_hd__buf_2 fanout105 (.A(_0692_),
    .X(net105));
 sky130_fd_sc_hd__buf_2 fanout106 (.A(_0690_),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 fanout107 (.A(_0690_),
    .X(net107));
 sky130_fd_sc_hd__buf_2 fanout108 (.A(_0689_),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 fanout109 (.A(_0689_),
    .X(net109));
 sky130_fd_sc_hd__buf_2 fanout110 (.A(net112),
    .X(net110));
 sky130_fd_sc_hd__buf_1 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 wire112 (.A(_0685_),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 fanout113 (.A(_0677_),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 fanout114 (.A(_0677_),
    .X(net114));
 sky130_fd_sc_hd__buf_2 fanout115 (.A(_0668_),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 fanout116 (.A(_0668_),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_4 fanout117 (.A(_0658_),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 fanout118 (.A(_0658_),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 fanout119 (.A(\addr0_reg[7] ),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 fanout120 (.A(\addr0_reg[7] ),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 fanout121 (.A(\addr0_reg[6] ),
    .X(net121));
 sky130_fd_sc_hd__buf_1 fanout122 (.A(\addr0_reg[6] ),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 fanout123 (.A(\addr0_reg[5] ),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 fanout124 (.A(\addr0_reg[5] ),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 fanout125 (.A(\addr0_reg[4] ),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 fanout126 (.A(\addr0_reg[4] ),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 fanout127 (.A(\addr0_reg[3] ),
    .X(net127));
 sky130_fd_sc_hd__buf_1 fanout128 (.A(\addr0_reg[3] ),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 fanout129 (.A(\addr0_reg[2] ),
    .X(net129));
 sky130_fd_sc_hd__buf_1 fanout130 (.A(\addr0_reg[2] ),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 fanout131 (.A(\addr0_reg[1] ),
    .X(net131));
 sky130_fd_sc_hd__buf_1 fanout132 (.A(\addr0_reg[1] ),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 fanout133 (.A(\addr0_reg[0] ),
    .X(net133));
 sky130_fd_sc_hd__buf_1 fanout134 (.A(\addr0_reg[0] ),
    .X(net134));
 sky130_fd_sc_hd__buf_2 fanout135 (.A(_0648_),
    .X(net135));
 sky130_fd_sc_hd__buf_1 fanout136 (.A(_0648_),
    .X(net136));
 sky130_fd_sc_hd__buf_2 fanout137 (.A(_0648_),
    .X(net137));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout138 (.A(_0648_),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk0 (.A(clk0),
    .X(clknet_0_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_0__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_1__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_2__leaf_clk0));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk0 (.A(clknet_0_clk0),
    .X(clknet_2_3__leaf_clk0));
 sky130_fd_sc_hd__clkinv_4 clkload0 (.A(clknet_2_0__leaf_clk0));
 sky130_fd_sc_hd__clkinv_4 clkload1 (.A(clknet_2_1__leaf_clk0));
 sky130_fd_sc_hd__bufinv_16 clkload2 (.A(clknet_2_3__leaf_clk0));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net33),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net34),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net24),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net26),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net22),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net21),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net17),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net32),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net30),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net31),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net40),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net15),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net35),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net18),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net28),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net29),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net23),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net16),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net37),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net39),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net36),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net20),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net41),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net19),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net10),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net12),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net25),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net13),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net27),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net11),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net38),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net14),
    .X(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0044_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0044_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0093_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_0094_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_0149_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_0240_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_0300_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_0595_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_0644_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_0225_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_0240_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_0464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_0225_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_0464_));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_281 ();
endmodule
