* NGSPICE file created from cust_rom.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

.subckt cust_rom VGND VPWR addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6]
+ addr0[7] clk0 cs0 dout0[0] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15]
+ dout0[16] dout0[17] dout0[18] dout0[19] dout0[1] dout0[20] dout0[21] dout0[22] dout0[23]
+ dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[2] dout0[30] dout0[31]
+ dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9]
XTAP_TAPCELL_ROW_9_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1270_ _0463_ _0552_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0985_ _0699_ _0705_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__or2_1
Xfanout127 addr0_reg\[3\] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
Xfanout105 _0692_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_2
Xfanout138 _0648_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dlymetal6s2s_1
X_1399_ _0099_ _0101_ _0226_ _0515_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__or4_1
Xfanout116 _0668_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_37_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0770_ _0062_ _0063_ _0066_ _0067_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__or4_2
X_1253_ net137 net150 net44 _0537_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__a22o_1
X_1322_ _0694_ _0163_ _0175_ _0221_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__or4_1
X_1184_ _0274_ _0415_ _0472_ _0473_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__or4_1
X_0968_ net105 net59 net55 net103 VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__a22oi_4
X_0899_ _0194_ _0197_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0822_ net87 net78 net76 net89 VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0753_ net115 net79 _0050_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__o21ba_2
X_1236_ net48 _0080_ _0459_ _0516_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1305_ _0049_ _0075_ _0195_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__or3_1
X_1167_ net137 net149 net44 _0457_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a22o_1
X_1098_ _0390_ _0391_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_22_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire100 net101 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1021_ _0223_ _0310_ _0311_ _0312_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0805_ net96 net79 net72 net98 VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0736_ net129 net127 net131 net133 VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1219_ _0193_ _0218_ _0269_ _0286_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold30 net11 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_5 _0088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1004_ _0287_ _0292_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__or3_1
X_0719_ net128 net133 net132 net130 VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput31 net31 VGND VGND VPWR VPWR dout0[29] sky130_fd_sc_hd__buf_2
Xoutput20 net20 VGND VGND VPWR VPWR dout0[19] sky130_fd_sc_hd__buf_2
XFILLER_0_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0984_ _0140_ _0239_ _0282_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout128 addr0_reg\[3\] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_1
X_1398_ _0660_ _0669_ _0671_ _0672_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__or4_1
Xfanout106 _0690_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_2
Xfanout117 _0658_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_37_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1252_ _0518_ _0528_ _0534_ _0536_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__or4_1
X_1321_ _0067_ _0068_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1183_ _0071_ _0084_ _0086_ _0219_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__or4_1
X_0967_ _0258_ _0259_ _0261_ _0262_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0898_ _0195_ _0196_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0821_ _0118_ _0119_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__or2_2
X_0752_ net123 net121 net119 net125 VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_28_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1166_ _0445_ _0450_ _0452_ _0456_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__or4_1
X_1235_ _0040_ _0068_ _0223_ _0273_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__or4_1
X_1304_ _0177_ _0250_ _0410_ _0418_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__or4_1
X_1097_ _0090_ _0091_ _0271_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__or3b_1
XFILLER_0_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire101 _0700_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
Xwire112 _0685_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
X_1020_ _0313_ _0314_ _0315_ _0317_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__or4_1
X_0735_ net131 net133 net129 net127 VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__and4b_1
X_0804_ net106 net79 net71 net108 VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__a22o_2
XFILLER_0_24_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1218_ _0695_ _0327_ _0353_ _0410_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__or4_1
X_1149_ _0062_ _0075_ _0085_ _0180_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold31 net38 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 net39 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_6 _0093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1003_ _0293_ _0295_ _0296_ _0301_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0718_ net130 net134 net131 net127 VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput21 net21 VGND VGND VPWR VPWR dout0[1] sky130_fd_sc_hd__buf_2
Xoutput10 net10 VGND VGND VPWR VPWR dout0[0] sky130_fd_sc_hd__buf_2
Xoutput32 net32 VGND VGND VPWR VPWR dout0[2] sky130_fd_sc_hd__buf_2
XFILLER_0_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0983_ _0091_ net47 _0099_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__or3_1
Xfanout107 _0690_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_2
Xfanout129 addr0_reg\[2\] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
Xfanout118 _0658_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
X_1397_ _0703_ _0103_ _0106_ _0235_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_37_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1320_ _0236_ _0252_ _0256_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__or3_1
X_1182_ _0107_ _0194_ _0212_ _0314_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__or4_1
X_1251_ _0076_ _0124_ _0251_ _0535_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_19_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0966_ _0259_ _0262_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0897_ net62 net60 _0687_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__o21ba_2
X_1449_ clknet_2_1__leaf_clk0 _0027_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_2_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0751_ net129 net127 net131 net133 VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__or4_4
X_0820_ net96 net77 net75 net98 VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__a22o_2
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1303_ net137 net162 net44 _0583_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__a22o_1
X_1234_ _0230_ _0249_ _0253_ _0519_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__or4_1
X_1096_ _0686_ _0039_ _0267_ _0268_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__or4bb_1
X_1165_ _0448_ _0449_ _0453_ _0455_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0949_ net53 net49 _0687_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0803_ net47 _0098_ _0099_ _0100_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__or4_1
X_0734_ _0698_ _0032_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1217_ _0399_ _0426_ _0503_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__or3_1
X_1148_ _0099_ _0118_ _0132_ _0138_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__or4_1
X_1079_ _0104_ _0139_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold32 net14 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 net31 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 net36 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_7 _0094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1002_ _0297_ _0298_ _0299_ _0300_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0717_ net111 net108 net106 net116 VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__a22o_2
XFILLER_0_35_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput33 net33 VGND VGND VPWR VPWR dout0[30] sky130_fd_sc_hd__buf_2
Xoutput11 net11 VGND VGND VPWR VPWR dout0[10] sky130_fd_sc_hd__buf_2
Xoutput22 net22 VGND VGND VPWR VPWR dout0[20] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0982_ _0144_ _0208_ _0279_ net9 VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__o31a_1
XFILLER_0_14_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout108 _0689_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_2
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout119 addr0_reg\[7\] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1396_ _0120_ _0200_ _0205_ _0670_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_37_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1181_ _0283_ _0459_ _0469_ _0470_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__or4_1
X_1250_ _0166_ _0168_ _0186_ _0196_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0965_ _0258_ _0261_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__or2_1
X_0896_ net113 net62 net61 net117 VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__a22o_2
X_1448_ clknet_2_1__leaf_clk0 _0026_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1379_ _0162_ _0551_ _0578_ _0653_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_25_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout90 _0037_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0750_ net110 net94 net92 net115 VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__a22o_2
X_1302_ _0338_ _0577_ _0578_ _0582_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1233_ _0072_ _0113_ _0114_ _0180_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_47_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1164_ _0124_ _0300_ _0316_ _0454_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__or4_1
X_1095_ _0230_ _0235_ _0254_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__or3_1
X_0948_ net114 net52 net49 net118 VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_30_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0879_ _0173_ _0174_ _0175_ _0176_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0802_ _0098_ _0100_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__or2_2
X_0733_ _0699_ _0702_ _0704_ _0705_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__or4_2
XFILLER_0_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1216_ _0148_ _0149_ _0150_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__or3_2
X_1147_ _0193_ _0194_ _0249_ _0259_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__or4_1
X_1078_ _0126_ _0238_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold11 net40 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_45_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold22 net20 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_8 _0094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1001_ _0173_ _0174_ _0176_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__or3_2
XFILLER_0_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0716_ net129 net131 net133 net127 VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput34 net34 VGND VGND VPWR VPWR dout0[31] sky130_fd_sc_hd__buf_2
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput12 net12 VGND VGND VPWR VPWR dout0[11] sky130_fd_sc_hd__buf_2
Xoutput23 net23 VGND VGND VPWR VPWR dout0[21] sky130_fd_sc_hd__buf_2
XFILLER_0_27_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0981_ _0208_ _0279_ net9 VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_32_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1395_ _0686_ _0107_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__or2_1
Xfanout109 _0689_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1180_ _0688_ _0694_ _0236_ _0458_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0964_ _0261_ _0262_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0895_ net102 net63 net61 net104 VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__a22o_2
X_1447_ clknet_2_3__leaf_clk0 _0025_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfxtp_1
X_1378_ _0040_ _0347_ _0433_ _0595_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout80 _0051_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlymetal6s2s_1
X_1301_ _0198_ _0579_ _0580_ _0581_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__or4_1
X_1232_ _0099_ _0101_ _0409_ _0517_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_47_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1163_ _0241_ _0246_ _0256_ _0261_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__or4_1
X_1094_ net135 net159 net42 _0388_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0947_ net109 net52 net49 net107 VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0878_ _0175_ _0176_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__or2_2
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload0 clknet_2_0__leaf_clk0 VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0801_ net102 net77 net75 net104 VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__a22o_1
X_0732_ _0704_ _0705_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__or2_2
XFILLER_0_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1215_ _0134_ _0317_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__or2_1
X_1146_ _0056_ _0239_ _0273_ _0437_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__or4_1
X_1077_ _0067_ net47 _0101_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__or3_1
Xhold23 net41 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 net15 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_9 _0107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1000_ _0122_ _0132_ _0151_ _0201_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0715_ net127 net131 net133 net129 VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__and4b_1
XFILLER_0_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1129_ _0094_ _0415_ _0416_ _0417_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput24 net24 VGND VGND VPWR VPWR dout0[22] sky130_fd_sc_hd__buf_2
Xoutput35 net35 VGND VGND VPWR VPWR dout0[3] sky130_fd_sc_hd__buf_2
Xoutput13 net13 VGND VGND VPWR VPWR dout0[12] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0980_ _0227_ _0245_ _0257_ _0277_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__or4_1
XFILLER_0_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1394_ _0244_ _0275_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0963_ net82 net52 net50 net86 VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__a22o_1
X_0894_ net108 net63 net61 net106 VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__a22o_2
XFILLER_0_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1377_ _0064_ _0120_ _0128_ _0129_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__or4_1
X_1446_ clknet_2_2__leaf_clk0 _0024_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_25_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout92 _0035_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_2
Xfanout70 _0073_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout81 net83 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_2
X_1162_ _0697_ _0108_ _0115_ _0205_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__or4_1
X_1300_ _0069_ _0115_ _0161_ _0244_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__or4_1
X_1231_ _0205_ _0237_ _0238_ _0241_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1093_ _0370_ _0383_ _0387_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__or3_1
X_0946_ _0232_ _0235_ _0244_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__or3_1
X_0877_ net118 net66 net64 net114 VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1429_ clknet_2_2__leaf_clk0 _0007_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfxtp_1
Xclkload1 clknet_2_1__leaf_clk0 VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0800_ net113 net77 net75 net117 VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__a22o_2
X_0731_ net115 net108 net106 net110 VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1214_ _0105_ _0242_ _0500_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__or3_1
X_1145_ _0095_ _0123_ _0152_ _0171_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1076_ _0259_ _0263_ _0336_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__or3_1
X_0929_ net120 net122 net126 net124 VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__and4b_1
Xhold24 net19 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 net35 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0714_ net116 net111 _0687_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1128_ _0066_ _0067_ _0127_ _0420_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1059_ _0084_ _0085_ _0086_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__or3_2
XFILLER_0_7_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput36 net36 VGND VGND VPWR VPWR dout0[4] sky130_fd_sc_hd__buf_2
Xoutput25 net25 VGND VGND VPWR VPWR dout0[23] sky130_fd_sc_hd__buf_2
Xoutput14 net14 VGND VGND VPWR VPWR dout0[13] sky130_fd_sc_hd__buf_2
XFILLER_0_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1393_ net138 net153 net45 _0667_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_19_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0962_ net90 net53 net50 net88 VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__a22o_2
X_0893_ _0185_ _0191_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__or2_1
X_1445_ clknet_2_2__leaf_clk0 _0023_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1376_ _0699_ _0097_ _0201_ _0246_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout82 net84 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout93 _0035_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_2
Xfanout60 net61 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
Xfanout71 _0070_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_47_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1230_ _0103_ _0182_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__or2_1
X_1092_ _0379_ _0380_ _0385_ _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__or4_1
X_1161_ _0703_ _0074_ _0087_ _0451_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0876_ net97 net67 net65 net99 VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__a22o_1
X_0945_ _0237_ _0238_ _0240_ _0241_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_30_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1428_ clknet_2_2__leaf_clk0 _0006_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dfxtp_1
X_1359_ _0086_ _0087_ _0136_ _0139_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__or4_1
Xclkload2 clknet_2_3__leaf_clk0 VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0730_ net111 net105 net103 net116 VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1213_ _0702_ _0705_ _0106_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1144_ _0285_ _0306_ _0308_ _0377_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__or4_1
X_1075_ _0367_ _0368_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__or3_1
X_0928_ _0220_ _0226_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0859_ _0154_ _0156_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__or2_1
Xhold14 net18 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 net10 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0713_ net129 net131 net133 net127 VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__or4b_4
XFILLER_0_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1127_ net48 _0103_ _0111_ net46 VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__or4_1
X_1058_ _0072_ _0138_ _0139_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__or3_2
XFILLER_0_43_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput37 net37 VGND VGND VPWR VPWR dout0[5] sky130_fd_sc_hd__buf_2
Xoutput15 net15 VGND VGND VPWR VPWR dout0[14] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput26 net26 VGND VGND VPWR VPWR dout0[24] sky130_fd_sc_hd__buf_2
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1392_ _0660_ _0663_ _0664_ _0666_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0961_ _0258_ _0259_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0892_ _0186_ _0187_ _0188_ _0189_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__or4_1
X_1444_ clknet_2_1__leaf_clk0 _0022_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfxtp_1
X_1375_ net135 net142 net42 _0650_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__a22o_1
Xfanout50 net51 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_1
Xfanout94 _0034_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_2
XFILLER_0_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout61 _0181_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout72 _0070_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_0_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1091_ _0115_ _0378_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__or2_1
X_1160_ _0147_ _0156_ _0188_ _0195_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__or4_1
X_0944_ _0238_ _0241_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0875_ net107 net66 net65 net109 VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_30_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1427_ clknet_2_1__leaf_clk0 _0005_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dfxtp_1
X_1358_ _0106_ _0107_ _0132_ _0155_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__or4_1
X_1289_ _0132_ _0136_ _0137_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__or3_1
XFILLER_0_33_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1212_ net135 net164 net42 _0499_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__a22o_1
X_1143_ _0205_ _0232_ _0253_ _0434_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1074_ _0193_ _0197_ _0269_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_23_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0927_ _0221_ _0222_ _0224_ _0225_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0858_ _0154_ _0155_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__or2_1
X_0789_ _0084_ _0085_ _0086_ _0087_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__or4_2
Xhold15 net28 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 net12 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_41_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0712_ net118 net116 net114 net111 VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__a22o_2
XFILLER_0_12_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1126_ _0706_ _0101_ _0197_ _0330_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1057_ _0072_ _0139_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput27 net27 VGND VGND VPWR VPWR dout0[25] sky130_fd_sc_hd__buf_2
Xoutput38 net38 VGND VGND VPWR VPWR dout0[6] sky130_fd_sc_hd__buf_2
Xoutput16 net16 VGND VGND VPWR VPWR dout0[15] sky130_fd_sc_hd__buf_2
Xclkbuf_2_3__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_3__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap91 _0037_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_17_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ _0161_ _0313_ _0396_ _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1391_ _0069_ _0178_ _0199_ _0665_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0960_ net93 net53 net49 net95 VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__a22o_2
X_0891_ _0188_ _0189_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__or2_1
X_1443_ clknet_2_2__leaf_clk0 _0021_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfxtp_1
X_1374_ _0641_ _0642_ _0649_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout62 _0167_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
Xfanout73 _0065_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_2
Xfanout95 _0034_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_0_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1090_ _0064_ _0079_ _0384_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__or3_1
X_0874_ net104 net67 net65 net102 VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__a22o_2
X_0943_ _0240_ _0241_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1357_ _0147_ _0176_ _0249_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__or3_1
X_1426_ clknet_2_2__leaf_clk0 _0004_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dfxtp_1
X_1288_ _0565_ _0567_ _0568_ _0569_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1142_ _0077_ net48 _0080_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__or3_1
X_1211_ _0496_ _0497_ _0498_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1073_ _0267_ _0272_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0926_ net93 net58 net54 net95 VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a22o_2
X_0857_ net109 net66 net64 net107 VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__a22o_1
Xhold16 net29 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ _0058_ _0083_ _0227_ _0579_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__or4_1
Xhold27 net25 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dlygate4sd3_1
X_0788_ net104 net73 net70 net102 VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0711_ net126 net124 net122 net120 VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1125_ _0118_ _0187_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__or2_1
X_1056_ _0174_ _0177_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput28 net28 VGND VGND VPWR VPWR dout0[26] sky130_fd_sc_hd__buf_2
X_0909_ _0179_ _0192_ _0207_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__or3_1
Xoutput39 net39 VGND VGND VPWR VPWR dout0[7] sky130_fd_sc_hd__buf_2
Xoutput17 net17 VGND VGND VPWR VPWR dout0[16] sky130_fd_sc_hd__buf_2
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1039_ _0246_ _0248_ _0249_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1108_ _0082_ _0108_ _0351_ _0399_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1390_ net47 _0188_ _0238_ _0252_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0890_ net104 net63 net60 net102 VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_10_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1442_ clknet_2_2__leaf_clk0 _0020_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfxtp_1
X_1373_ _0160_ _0644_ _0646_ _0647_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout52 net53 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_2
Xfanout63 _0167_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_1
Xfanout74 _0065_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
Xfanout96 _0701_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_2
Xfanout85 _0042_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0942_ net88 net59 net55 net90 VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__a22o_2
X_0873_ _0163_ _0164_ _0166_ _0168_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1425_ clknet_2_2__leaf_clk0 _0003_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dfxtp_1
X_1356_ _0124_ _0130_ _0413_ _0631_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__or4_1
X_1287_ _0046_ _0170_ _0278_ _0374_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1141_ _0193_ _0249_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1210_ _0161_ _0492_ _0494_ _0495_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__or4_1
X_1072_ _0084_ _0085_ _0158_ _0220_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__or4_1
X_0925_ net82 net58 net54 net86 VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__a22o_2
X_0856_ net113 net66 net64 net117 VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__a22o_1
X_0787_ net106 net73 net69 net108 VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1408_ net137 net147 net44 _0682_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__a22o_1
Xhold17 net23 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 net13 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dlygate4sd3_1
X_1339_ _0375_ _0610_ _0614_ _0616_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_41_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0710_ net127 net131 net133 net129 VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1055_ _0118_ _0119_ _0122_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__or3_1
X_1124_ _0241_ _0256_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0908_ _0199_ _0200_ _0205_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__or3_1
Xoutput29 net29 VGND VGND VPWR VPWR dout0[27] sky130_fd_sc_hd__buf_2
Xoutput18 net18 VGND VGND VPWR VPWR dout0[17] sky130_fd_sc_hd__buf_2
X_0839_ net80 net71 _0687_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1107_ _0307_ _0311_ _0393_ _0394_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1038_ _0237_ _0241_ _0252_ _0253_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1441_ clknet_2_2__leaf_clk0 _0019_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfxtp_1
X_1372_ _0169_ _0218_ _0463_ _0538_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout97 _0701_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_2
Xfanout86 _0042_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
Xfanout53 _0228_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout75 _0061_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_2
Xfanout42 _0281_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout64 _0146_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_2
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0941_ net86 net59 net55 net82 VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__a22o_2
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0872_ _0164_ _0168_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__or2_1
X_1355_ _0045_ net48 _0080_ _0094_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__or4_1
X_1424_ clknet_2_3__leaf_clk0 _0002_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dfxtp_1
X_1286_ _0204_ _0482_ _0493_ _0552_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1071_ net136 net151 net43 _0366_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__a22o_1
X_1140_ _0104_ _0107_ _0216_ _0431_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__or4_1
X_0924_ _0221_ _0222_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__or2_1
X_0855_ net102 net66 net64 net104 VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__a22o_2
X_0786_ net96 net73 net69 net98 VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__a22o_2
XFILLER_0_11_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold29 net27 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1407_ _0179_ _0679_ _0681_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__or3_1
X_1338_ _0109_ _0317_ _0335_ _0615_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__or4_1
Xhold18 net16 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_41_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1269_ _0048_ _0125_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1054_ _0269_ _0273_ _0349_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__or3b_1
X_1123_ _0182_ _0183_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_11_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0907_ _0200_ _0202_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__or2_1
Xoutput19 net19 VGND VGND VPWR VPWR dout0[18] sky130_fd_sc_hd__buf_2
X_0838_ net73 net69 _0687_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__o21ba_1
X_0769_ _0062_ _0066_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__or2_2
XFILLER_0_34_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap83 net84 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1106_ _0205_ _0395_ _0397_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__or3_1
X_1037_ _0332_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1440_ clknet_2_3__leaf_clk0 _0018_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfxtp_1
X_1371_ _0177_ _0263_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout87 _0038_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_4
Xfanout65 _0146_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_2
Xfanout54 net57 VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_4
Xfanout76 _0061_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout98 net100 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_2
Xfanout43 _0281_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_47_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0940_ _0237_ _0238_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0871_ _0163_ _0166_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__or2_1
X_1354_ _0165_ _0311_ _0550_ _0599_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__or4_1
X_1285_ _0149_ _0183_ _0200_ _0566_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__or4_1
X_1423_ clknet_2_2__leaf_clk0 _0001_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_41_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1070_ _0355_ _0361_ _0362_ _0365_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__or4_1
X_0923_ net90 net59 net54 net88 VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__a22o_2
X_0854_ _0148_ _0149_ _0150_ _0151_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__or4_2
XFILLER_0_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0785_ net117 net74 net70 net113 VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold19 net37 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dlygate4sd3_1
X_1268_ _0232_ _0234_ _0550_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__or3_1
X_1406_ _0698_ _0047_ _0678_ _0680_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__or4_1
X_1337_ _0041_ _0137_ _0148_ _0248_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__or4_1
X_1199_ _0088_ _0147_ _0194_ _0261_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1122_ _0188_ _0247_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__or2_2
X_1053_ _0686_ _0691_ _0694_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__nor3_1
XFILLER_0_28_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0906_ _0201_ _0202_ _0203_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__or3_2
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0837_ net102 net74 net69 net104 VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__a22o_2
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0768_ net89 net77 net75 net87 VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_44_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap51 _0229_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1105_ _0131_ _0132_ _0137_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_16_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1036_ _0090_ _0091_ _0111_ _0114_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1019_ _0084_ _0086_ _0087_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__or3_1
XFILLER_0_40_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1370_ _0049_ _0052_ _0225_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__or3_1
XFILLER_0_10_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout44 _0281_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
Xfanout55 net56 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout99 net101 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_2
Xfanout88 _0038_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout66 _0145_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_2
Xfanout77 _0059_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_2
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0870_ _0163_ _0168_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__or2_2
XFILLER_0_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1422_ clknet_2_3__leaf_clk0 _0000_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfxtp_1
X_1353_ net137 net141 net44 _0629_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__a22o_1
X_1284_ _0091_ net47 _0100_ _0134_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0999_ _0156_ _0164_ _0195_ _0202_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0922_ net99 net59 net55 net97 VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a22o_1
X_0853_ _0150_ _0151_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__or2_2
X_0784_ _0077_ net48 _0080_ _0081_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__or4_1
X_1405_ _0191_ _0266_ _0354_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__or3_1
Xinput1 addr0[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_1198_ _0686_ _0695_ _0485_ _0486_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__or4_1
X_1267_ _0688_ _0694_ _0194_ _0195_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__or4_1
X_1336_ _0152_ _0206_ _0613_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1121_ _0702_ _0137_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__or2_1
X_1052_ _0080_ _0184_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__or2_1
X_0767_ net77 net74 _0050_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__o21ba_1
X_0905_ _0201_ _0203_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__or2_1
X_0836_ _0050_ net70 VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1319_ _0045_ _0080_ _0081_ _0597_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1035_ net46 _0182_ _0187_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__or3_1
X_1104_ _0131_ _0137_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0819_ net94 net77 net75 net92 VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1018_ _0036_ _0044_ net48 _0081_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout45 _0281_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout67 net68 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_1
Xfanout78 _0059_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_24_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout89 net91 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
XFILLER_0_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1421_ clknet_2_0__leaf_clk0 net8 VGND VGND VPWR VPWR addr0_reg\[7\] sky130_fd_sc_hd__dfxtp_1
X_1352_ _0608_ _0623_ _0628_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__or3_1
X_1283_ _0177_ _0190_ _0288_ _0564_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_21_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0998_ _0211_ _0230_ _0233_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0921_ _0211_ _0212_ _0213_ _0215_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__or4_2
X_0852_ net82 net66 net64 net86 VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0783_ _0077_ net48 _0081_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__or3_1
X_1404_ _0109_ _0116_ _0207_ _0669_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__or4_1
X_1335_ _0071_ _0075_ _0136_ _0138_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__or4_1
X_1197_ _0221_ _0222_ _0225_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__or3_1
Xinput2 addr0[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1266_ net136 net156 net43 _0549_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1051_ _0240_ _0253_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__or2_1
X_1120_ _0049_ _0286_ _0412_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__or3_1
X_0904_ net81 net62 net60 net85 VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__a22o_2
XFILLER_0_43_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0766_ net121 net119 net123 net125 VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__and4b_1
X_0835_ net85 net74 net70 net81 VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1318_ _0099_ _0100_ _0202_ _0203_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__or4_1
X_1249_ _0530_ _0531_ _0532_ _0533_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1103_ _0075_ _0294_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__or2_1
X_1034_ _0074_ _0075_ _0132_ _0151_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0749_ net115 net89 net87 net110 VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0818_ _0096_ _0102_ _0109_ _0116_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_39_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1017_ _0247_ _0250_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_18_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout79 _0051_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_2
XFILLER_0_35_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1351_ _0554_ _0600_ _0624_ _0627_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__or4_1
X_1420_ clknet_2_0__leaf_clk0 net7 VGND VGND VPWR VPWR addr0_reg\[6\] sky130_fd_sc_hd__dfxtp_1
X_1282_ _0052_ _0119_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0997_ _0081_ _0138_ _0246_ _0247_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0920_ _0211_ _0215_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__or2_1
X_0851_ net90 net66 net64 net87 VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0782_ net92 net79 net71 net94 VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1403_ _0706_ _0123_ _0184_ _0247_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1334_ _0392_ _0608_ _0611_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__or3_1
X_1265_ _0542_ _0546_ _0548_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__or3_1
X_1196_ _0193_ _0196_ _0258_ _0259_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__or4_1
Xinput3 addr0[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1050_ net136 net146 net43 _0346_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__a22o_1
X_0903_ net98 net62 net60 net96 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__a22o_2
X_0834_ _0131_ _0132_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0765_ _0062_ _0063_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1317_ _0398_ _0415_ _0595_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__or3_1
X_1248_ _0062_ _0085_ _0087_ _0190_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1179_ _0047_ _0127_ _0129_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_30 _0225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1102_ _0130_ _0211_ _0237_ _0261_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__or4_1
X_1033_ _0262_ _0272_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_16_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0817_ _0110_ _0111_ _0113_ _0114_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__or4_1
X_0748_ _0036_ _0039_ _0041_ _0044_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_39_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1016_ _0163_ _0166_ _0168_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout58 _0209_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_4
Xfanout69 _0073_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_2
Xfanout47 _0097_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
XFILLER_0_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1281_ net137 net145 net44 _0563_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__a22o_1
X_1350_ _0355_ _0447_ _0625_ _0626_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0996_ _0125_ _0128_ _0294_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0850_ net92 net66 net64 net94 VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__a22o_2
X_1402_ net138 net154 net45 _0676_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0781_ net98 net80 net72 net96 VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__a22o_2
Xinput4 addr0[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_1264_ _0178_ _0295_ _0547_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__or3_1
X_1333_ _0394_ _0458_ _0482_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__or3_1
X_1195_ _0411_ _0480_ _0481_ _0483_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__or4_1
X_0979_ _0253_ _0256_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_40_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0833_ net108 net73 net69 net106 VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__a22o_2
X_0902_ net89 net62 net60 net87 VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0764_ net81 net78 net76 net85 VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__a22o_1
X_1316_ _0077_ _0224_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__or2_1
X_1178_ _0434_ _0465_ _0466_ _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1247_ _0151_ _0155_ _0156_ _0269_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_31 _0240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_20 _0464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1101_ _0246_ _0247_ _0249_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__or3_1
X_1032_ _0327_ _0328_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0747_ _0036_ _0041_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__or2_2
XFILLER_0_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0816_ _0110_ _0111_ _0114_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__or3_2
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1015_ _0068_ _0099_ _0100_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout59 _0209_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_32_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout48 _0078_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_2
XFILLER_0_35_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1280_ _0558_ _0559_ _0562_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_46_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0995_ _0074_ _0134_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_21_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0780_ _0077_ net48 VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__or2_1
X_1401_ _0673_ _0675_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__or2_1
X_1263_ _0232_ _0253_ _0395_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__or3_1
Xinput5 addr0[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_1194_ net46 _0250_ _0462_ _0482_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__or4_1
X_1332_ _0078_ _0081_ _0169_ _0235_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__or4_1
X_0978_ _0266_ _0276_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_40_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0832_ net113 net73 net69 net117 VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__a22o_2
X_0901_ net92 net63 net61 net94 VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__a22o_2
X_0763_ net92 net77 net75 net94 VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1315_ net135 net160 net42 _0594_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1177_ _0706_ _0055_ _0074_ _0311_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1246_ _0702_ _0039_ _0398_ _0458_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__or4_1
XANTENNA_21 _0534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 _0464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_10 _0149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_cap56 net57 VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1100_ _0222_ _0224_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1031_ _0062_ _0084_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__or2_1
X_0746_ _0041_ _0044_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0815_ net85 net80 net71 net81 VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__a22o_2
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1229_ _0048_ _0049_ _0053_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_2__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_2__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1014_ _0194_ _0267_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0729_ _0699_ _0702_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout49 _0229_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_2
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0994_ _0046_ _0186_ _0188_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1400_ _0179_ _0336_ _0592_ _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__or4_1
X_1331_ _0198_ _0352_ _0377_ _0461_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1193_ _0182_ _0184_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__or2_1
Xinput6 addr0[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_1262_ _0464_ _0543_ _0544_ _0545_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0977_ _0267_ _0268_ _0271_ _0272_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__nand4_2
XFILLER_0_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0193_ _0194_ _0195_ _0196_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0831_ _0125_ _0126_ _0128_ _0129_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__or4_4
X_0762_ net125 net121 net119 net123 VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_47_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1314_ _0591_ _0592_ _0593_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__or3_1
X_1176_ _0174_ _0175_ _0182_ _0200_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1245_ _0056_ net48 _0529_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__or3_1
XANTENNA_22 _0558_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_11 _0169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 _0225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap46 _0180_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
Xmax_cap68 _0145_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1030_ _0067_ _0256_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0814_ net95 net79 net71 net93 VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__a22o_1
X_0745_ net115 net85 net81 net110 VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__a22o_2
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1228_ net135 net166 net42 _0514_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1159_ _0094_ _0270_ _0393_ _0446_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_13_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1013_ _0258_ _0262_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0728_ net115 net98 net96 net110 VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0993_ _0289_ _0290_ _0291_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1330_ _0032_ _0515_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__or2_1
X_1261_ _0083_ _0159_ _0354_ _0412_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__or4_1
X_1192_ _0079_ _0278_ _0479_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__or3_1
Xinput7 addr0[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
X_0976_ _0268_ _0272_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0830_ net78 net76 _0687_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0761_ net126 net124 net120 VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__nand3b_1
X_1313_ _0350_ _0367_ _0584_ _0586_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__or4_1
X_1244_ _0092_ _0103_ _0259_ _0271_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__or4b_1
X_1175_ _0448_ _0460_ _0461_ _0464_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_19_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0959_ net99 net52 net50 net97 VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__a22o_2
XANTENNA_34 _0464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 _0169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_23 _0570_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0813_ _0110_ _0111_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_26_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0744_ net130 net128 net134 net132 VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__nor4b_1
XPHY_EDGE_ROW_10_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1227_ _0504_ _0507_ _0509_ _0513_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__or4_1
X_1158_ _0054_ _0127_ _0129_ _0447_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__or4_1
X_1089_ _0122_ _0131_ _0149_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1012_ _0686_ _0119_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0727_ net132 net133 net130 net128 VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0992_ _0067_ _0110_ _0180_ _0182_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput8 addr0[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
X_1191_ _0103_ _0114_ _0284_ _0373_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__or4_1
X_1260_ _0091_ _0095_ _0112_ _0263_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__or4_1
X_0975_ _0267_ _0271_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1389_ _0217_ _0376_ _0431_ _0624_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0760_ net123 net119 net121 net125 VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__and4b_1
XFILLER_0_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1243_ _0093_ _0460_ _0476_ _0527_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__or4_1
X_1174_ _0118_ _0119_ _0121_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__or3_2
X_1312_ _0047_ _0130_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_19_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_13 _0177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0958_ _0251_ _0254_ _0256_ _0255_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__or4b_1
X_0889_ net106 net62 net61 net108 VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__a22o_2
XANTENNA_24 _0595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0743_ net134 net132 net128 net129 VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__and4b_1
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0812_ net87 net80 net71 net89 VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__a22o_2
X_1157_ _0148_ _0149_ _0151_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__or3_1
X_1226_ _0171_ _0265_ _0510_ _0512_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__or4_1
X_1088_ _0371_ _0372_ _0381_ _0382_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1011_ _0305_ _0306_ _0308_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__or3_1
X_0726_ net128 net132 net134 net130 VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1209_ _0356_ _0390_ _0447_ _0491_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0709_ net125 net123 net119 net121 VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0991_ _0694_ _0039_ _0086_ _0114_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 cs0 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
X_1190_ _0052_ _0053_ _0067_ _0099_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__or4_1
X_0974_ _0271_ _0272_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1388_ _0162_ _0371_ _0661_ _0662_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1311_ _0555_ _0588_ _0589_ _0590_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__or4_1
X_1242_ _0230_ _0254_ _0349_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__or3b_1
X_1173_ _0118_ _0121_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_25 _0603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_14 _0237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0957_ net88 net52 net49 net90 VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__a22o_2
X_0888_ net96 net62 net60 net98 VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0742_ net110 net98 net96 net115 VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0811_ _0050_ _0060_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__nor2_2
X_1087_ _0691_ _0225_ _0374_ _0375_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__or4_1
X_1156_ _0071_ _0138_ _0139_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__or3_1
X_1225_ _0130_ _0511_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_7_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1010_ _0173_ _0175_ _0176_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__or3_1
X_0725_ net116 net113 net110 net117 VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1208_ _0389_ _0432_ _0483_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1139_ _0113_ _0114_ _0222_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1 net33 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_1_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0708_ net129 net127 net131 net133 VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__and4b_1
XFILLER_0_35_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0990_ _0252_ _0256_ _0264_ _0288_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0973_ net118 net58 net54 net114 VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_14_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1387_ _0695_ _0275_ _0619_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1241_ net137 net170 net44 _0526_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1310_ _0112_ _0263_ _0412_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__or3_1
X_1172_ _0119_ _0121_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0956_ net126 net124 net122 _0050_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__or4_1
XANTENNA_15 _0240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _0603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0887_ net117 net62 net60 net113 VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__a22o_2
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1439_ clknet_2_2__leaf_clk0 _0017_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0810_ _0103_ _0104_ _0106_ _0107_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__or4_4
X_0741_ _0036_ _0039_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1224_ _0111_ _0119_ _0173_ _0231_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__or4_1
X_1155_ _0704_ _0164_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__or2_1
X_1086_ _0046_ _0171_ _0294_ _0373_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__or4_1
X_0939_ net95 net58 net54 net93 VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_15_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0724_ _0686_ _0688_ _0691_ _0694_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__or4_2
X_1207_ _0173_ _0188_ _0196_ _0201_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1138_ _0697_ _0040_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__or2_1
X_1069_ _0327_ _0350_ _0363_ _0364_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_26_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 net34 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dlygate4sd3_1
X_0707_ net9 VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0972_ net107 net58 net54 net109 VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_22_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1386_ _0079_ _0120_ _0127_ _0232_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1240_ _0518_ _0523_ _0525_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__or3_1
X_1171_ _0063_ _0067_ _0098_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0955_ _0252_ _0253_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__or2_1
XANTENNA_16 _0288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0886_ net46 _0182_ _0183_ _0184_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__or4_1
XANTENNA_27 _0630_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1438_ clknet_2_3__leaf_clk0 _0016_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1369_ _0696_ _0247_ _0249_ _0643_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0740_ net110 net89 net87 net115 VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__a22o_2
X_1223_ _0071_ _0081_ _0224_ _0225_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__or4_1
X_1154_ _0101_ _0169_ _0232_ _0328_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__or4_1
X_1085_ _0092_ _0094_ _0376_ _0377_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__or4_1
X_0938_ net54 net53 _0050_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0869_ net64 _0167_ _0050_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__o21ba_2
XTAP_TAPCELL_ROW_7_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0723_ _0688_ _0691_ _0694_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1137_ net135 net169 net42 _0429_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__a22o_1
X_1206_ _0127_ _0133_ _0294_ _0493_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1068_ _0216_ _0284_ _0347_ _0348_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_47_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_31_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3 net24 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0971_ _0267_ _0268_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__nand2_1
X_1385_ net46 _0354_ _0416_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ _0221_ _0222_ _0224_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__or3_1
X_0954_ net86 net53 net50 net82 VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__a22o_2
XFILLER_0_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_28 _0644_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 _0300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0885_ net94 net63 net60 net92 VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1437_ clknet_2_2__leaf_clk0 _0015_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1299_ _0165_ _0311_ _0331_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__or3_1
X_1368_ _0036_ _0041_ _0125_ _0128_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1222_ _0315_ _0340_ _0508_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__or3_1
X_1084_ _0173_ _0174_ _0183_ _0184_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__or4_1
X_1153_ net136 net158 net43 _0444_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__a22o_1
X_0937_ _0231_ _0234_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__or2_1
X_0799_ net108 net77 net75 net106 VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__a22o_2
X_0868_ net123 net119 net121 net125 VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_7_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0722_ _0688_ _0691_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1136_ _0424_ _0427_ _0428_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__or3_1
X_1205_ _0066_ net48 VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__or2_1
X_1067_ _0194_ _0195_ _0250_ _0294_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 net26 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1119_ _0221_ _0224_ _0225_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0970_ net97 net58 net55 net99 VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__a22o_2
XFILLER_0_39_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1453_ clknet_2_3__leaf_clk0 _0031_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dfxtp_1
X_1384_ net138 net167 net45 _0659_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_18 _0415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_29 _0056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0953_ net95 net52 net49 net93 VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__a22o_2
X_0884_ net87 net62 net60 net89 VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__a22o_2
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1436_ clknet_2_1__leaf_clk0 _0014_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfxtp_1
X_1367_ _0378_ _0425_ _0543_ _0571_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__or4_1
X_1298_ _0071_ _0274_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_18_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1221_ _0092_ _0094_ _0185_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__or3_1
X_1152_ _0430_ _0432_ _0438_ _0443_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__or4_1
X_1083_ _0231_ _0233_ _0253_ _0256_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__or4_2
X_0936_ _0233_ _0234_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__or2_2
XFILLER_0_15_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0867_ net86 net66 net64 net82 VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0798_ net98 net78 net76 net96 VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__a22o_1
X_1419_ clknet_2_0__leaf_clk0 net6 VGND VGND VPWR VPWR addr0_reg\[5\] sky130_fd_sc_hd__dfxtp_1
Xwire84 _0043_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0721_ _0691_ _0694_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_12_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1204_ _0096_ _0102_ _0285_ _0286_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1135_ _0160_ _0411_ _0413_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__or3_1
X_1066_ _0180_ _0352_ _0354_ _0356_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0919_ _0211_ _0213_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 net22 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1118_ _0202_ _0409_ _0410_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__or3_1
X_1049_ _0338_ _0342_ _0345_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1452_ clknet_2_3__leaf_clk0 _0030_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dfxtp_1
X_1383_ _0478_ _0654_ _0657_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_19 _0452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0952_ _0246_ _0247_ _0248_ _0249_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0883_ net85 net62 net60 net81 VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__a22o_2
X_1435_ clknet_2_3__leaf_clk0 _0013_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1366_ _0334_ _0372_ _0501_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_18_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1297_ _0105_ _0186_ _0189_ _0409_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1220_ _0501_ _0502_ _0505_ _0506_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__or4_1
X_1151_ _0435_ _0436_ _0442_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__or3_1
X_1082_ _0186_ _0187_ _0189_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__or3_1
X_0935_ net107 net52 net49 net109 VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__a22o_1
X_0866_ _0163_ _0164_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0797_ _0090_ _0091_ _0092_ _0093_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__or4_2
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1418_ clknet_2_0__leaf_clk0 net5 VGND VGND VPWR VPWR addr0_reg\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1349_ _0213_ _0215_ _0248_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0720_ net116 net105 net103 net111 VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__a22o_2
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1134_ _0698_ _0300_ _0425_ _0426_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__or4_1
X_1203_ _0243_ _0265_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1065_ _0357_ _0358_ _0359_ _0360_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__or4_1
X_0849_ net99 net67 net65 net97 VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__a22o_2
X_0918_ _0214_ _0215_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_9_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_1__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
Xhold6 net21 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1117_ _0200_ _0203_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1048_ _0329_ _0334_ _0343_ _0344_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_23_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1451_ clknet_2_3__leaf_clk0 _0029_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dfxtp_1
X_1382_ _0264_ _0652_ _0655_ _0656_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0951_ _0248_ _0249_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__or2_1
X_0882_ net125 net119 net121 net123 VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_27_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1296_ _0462_ _0574_ _0575_ _0576_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__or4_1
X_1365_ net135 net165 net42 _0640_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__a22o_1
X_1434_ clknet_2_2__leaf_clk0 _0012_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1150_ _0161_ _0439_ _0440_ _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__or4_1
X_1081_ _0699_ _0702_ _0052_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__or3_1
X_0934_ net105 net52 net49 net103 VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__a22o_1
X_0865_ net95 net66 net64 net93 VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1417_ clknet_2_0__leaf_clk0 net4 VGND VGND VPWR VPWR addr0_reg\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0796_ _0090_ _0092_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__or2_1
X_1279_ _0190_ _0556_ _0560_ _0561_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__or4_1
X_1348_ _0099_ _0106_ _0111_ _0149_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_6_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1202_ net137 net168 net44 _0490_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__a22o_1
X_1133_ _0044_ _0046_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1064_ _0036_ _0077_ net47 _0136_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_25_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0848_ net67 net65 _0687_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__o21ba_2
X_0917_ _0212_ _0215_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__or2_1
X_0779_ net81 net80 net72 net85 VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold7 net17 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1116_ _0211_ _0212_ _0213_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_0_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1047_ _0109_ _0158_ _0260_ _0330_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk0 clk0 VGND VGND VPWR VPWR clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1450_ clknet_2_1__leaf_clk0 _0028_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1381_ _0054_ _0111_ _0458_ _0587_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0950_ net103 net53 net49 net105 VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__a22o_2
X_0881_ net125 net119 _0050_ net123 VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1433_ clknet_2_2__leaf_clk0 _0011_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfxtp_1
X_1295_ _0039_ _0044_ _0085_ _0122_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__or4_1
X_1364_ _0630_ _0632_ _0639_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_18_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1080_ _0121_ _0128_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0864_ net88 net67 net65 net90 VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__a22o_2
X_0933_ _0230_ _0231_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__or2_2
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0795_ _0090_ _0093_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__or2_2
XFILLER_0_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1416_ clknet_2_0__leaf_clk0 net3 VGND VGND VPWR VPWR addr0_reg\[2\] sky130_fd_sc_hd__dfxtp_1
X_1347_ _0039_ _0044_ _0164_ _0166_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1278_ _0214_ _0254_ _0265_ _0446_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__or4_1
Xfanout130 addr0_reg\[2\] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1201_ _0293_ _0478_ _0484_ _0489_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__or4_1
X_1132_ _0080_ _0081_ _0353_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__or3_1
X_1063_ _0107_ _0113_ _0154_ _0203_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__or4_1
X_0916_ net109 net58 net54 net107 VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0847_ net120 net122 net126 net124 VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__and4bb_1
X_0778_ net89 net79 net72 net88 VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__a22o_2
XFILLER_0_38_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_42_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold8 net32 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1115_ net137 net157 net44 _0408_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1046_ _0169_ _0339_ _0340_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_23_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1029_ net136 net144 net43 _0326_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1380_ _0269_ _0273_ _0651_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0880_ _0153_ _0161_ _0172_ _0178_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__or4_1
X_1432_ clknet_2_3__leaf_clk0 _0010_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1363_ _0112_ _0636_ _0637_ _0638_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__or4_1
X_1294_ _0090_ _0128_ _0225_ _0252_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0932_ net118 net52 net49 net114 VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_15_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0863_ _0153_ _0161_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__or2_1
X_0794_ net98 net73 net69 net96 VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1415_ clknet_2_0__leaf_clk0 net2 VGND VGND VPWR VPWR addr0_reg\[1\] sky130_fd_sc_hd__dfxtp_1
X_1346_ _0192_ _0245_ _0620_ _0622_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__or4_1
X_1277_ _0095_ _0140_ _0147_ _0202_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout131 addr0_reg\[1\] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout120 addr0_reg\[7\] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_29_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1200_ _0276_ _0397_ _0487_ _0488_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1131_ _0419_ _0421_ _0422_ _0423_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__or4_1
X_1062_ _0057_ _0230_ _0238_ _0258_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__or4_1
X_0915_ _0212_ _0213_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__or2_1
X_0777_ _0071_ _0072_ _0074_ _0075_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__or4_1
X_0846_ net126 net124 net120 net121 VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__nor4b_1
X_1329_ net135 net143 net42 _0607_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 net30 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1114_ _0400_ _0403_ _0407_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__or3_1
XFILLER_0_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1045_ _0082_ _0331_ _0335_ _0341_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0829_ net106 net77 net75 net108 VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__a22o_2
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1028_ _0309_ _0318_ _0320_ _0325_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1431_ clknet_2_1__leaf_clk0 _0009_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dfxtp_1
X_1293_ net47 _0098_ _0348_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__or3_1
X_1362_ _0068_ _0219_ _0284_ _0368_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0931_ net97 net52 net50 net99 VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_15_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0862_ _0147_ _0154_ _0155_ _0156_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__or4_4
X_0793_ net89 net73 net69 net87 VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__a22o_2
X_1414_ clknet_2_0__leaf_clk0 net1 VGND VGND VPWR VPWR addr0_reg\[0\] sky130_fd_sc_hd__dfxtp_1
X_1345_ _0036_ _0080_ _0152_ _0621_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__or4_1
X_1276_ _0486_ _0503_ _0554_ _0555_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout132 addr0_reg\[1\] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__buf_1
Xfanout110 net112 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__buf_2
Xfanout121 addr0_reg\[6\] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1130_ _0165_ _0414_ _0418_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1061_ _0172_ _0226_ _0339_ _0351_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__or4_1
X_0914_ net114 net58 net54 net118 VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__a22o_1
X_0845_ _0058_ _0089_ _0117_ _0143_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0776_ net94 net74 net70 net92 VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__a22o_2
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1328_ _0603_ _0604_ _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__or3_1
X_1259_ _0197_ _0410_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1113_ _0389_ _0392_ _0401_ _0406_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__or4_1
X_1044_ _0071_ _0072_ _0138_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0828_ _0125_ _0126_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__or2_2
X_0759_ _0698_ _0032_ _0047_ _0057_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1027_ _0299_ _0321_ _0323_ _0324_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1430_ clknet_2_1__leaf_clk0 _0008_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1292_ net135 net152 net42 _0573_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__a22o_1
X_1361_ net47 _0098_ _0204_ _0243_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0930_ net126 net124 net120 net122 VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_15_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0792_ net92 net73 net69 net94 VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__a22o_2
X_0861_ _0153_ _0159_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__or2_1
X_1413_ net140 _0144_ net9 VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1344_ _0202_ _0203_ _0224_ _0225_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__or4_1
X_1275_ _0502_ _0551_ _0553_ _0557_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__or4_1
Xwire57 _0210_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout133 addr0_reg\[0\] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
Xfanout111 net112 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_1
Xfanout122 addr0_reg\[6\] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1060_ _0064_ _0148_ _0149_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0913_ net103 net59 net55 net105 VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__a22o_1
X_0844_ _0124_ _0130_ _0141_ _0142_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__or4_1
X_0775_ net87 net74 net70 net89 VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_3_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1189_ _0168_ _0477_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__or2_1
X_1327_ _0111_ _0391_ _0458_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__or4_1
X_1258_ _0372_ _0430_ _0540_ _0541_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1043_ net47 _0099_ _0100_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__or3_1
X_1112_ _0404_ _0405_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0758_ _0048_ _0049_ _0052_ _0053_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__or4_1
X_0827_ net104 net78 net75 net102 VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_46_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_30_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1026_ _0696_ _0157_ _0206_ _0278_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1009_ _0173_ _0175_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1360_ _0153_ _0633_ _0634_ _0635_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__or4_1
X_1291_ _0033_ _0370_ _0570_ _0572_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0791_ net81 net73 net69 net85 VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_15_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0860_ _0154_ _0155_ _0156_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__or3_1
X_1412_ net9 net139 _0280_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__o21a_1
X_1343_ _0140_ _0312_ _0459_ _0619_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1274_ _0702_ _0039_ _0103_ _0114_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__or4_1
X_0989_ _0150_ _0224_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__or2_1
Xfanout134 addr0_reg\[0\] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_1
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout123 addr0_reg\[5\] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_29_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0912_ net58 net54 _0687_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_11_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0774_ net125 net123 net119 net121 VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__and4bb_1
X_0843_ _0134_ _0135_ _0138_ _0139_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1326_ _0122_ _0126_ _0248_ _0379_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__or4_1
X_1188_ _0094_ _0131_ _0163_ _0476_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__or4_1
X_1257_ _0149_ _0168_ _0214_ _0516_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1042_ _0125_ _0128_ _0129_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__or3_1
X_1111_ _0688_ _0071_ _0085_ _0110_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0757_ _0048_ _0053_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__or2_1
X_0826_ net117 net77 net75 net113 VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1309_ _0091_ _0095_ _0571_ _0587_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1025_ _0096_ _0322_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__or2_1
X_0809_ _0103_ _0104_ _0107_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1 _0039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1008_ _0072_ _0128_ _0129_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1290_ _0111_ _0458_ _0491_ _0571_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0790_ _0069_ _0076_ _0083_ _0088_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1411_ net138 net148 net45 _0684_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__a22o_1
X_1273_ _0069_ _0276_ _0296_ _0332_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__or4_1
X_1342_ _0092_ _0104_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0988_ _0283_ _0285_ _0286_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__or3_1
Xfanout102 _0693_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_4
Xfanout113 _0677_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout135 _0648_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_2
Xfanout124 addr0_reg\[5\] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0911_ net124 net120 net122 net126 VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__nor4b_1
X_0842_ _0131_ _0132_ _0136_ _0137_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0773_ net102 net80 net72 net104 VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__a22o_2
X_1256_ _0414_ _0538_ _0539_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_3_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1325_ _0305_ _0502_ _0596_ _0598_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1187_ _0091_ _0173_ _0174_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1110_ _0049_ _0163_ _0183_ _0193_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1041_ _0232_ _0233_ _0336_ _0337_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__or4_2
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0825_ _0118_ _0119_ _0121_ _0122_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__or4_2
X_0756_ _0048_ _0049_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1239_ _0397_ _0464_ _0515_ _0524_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__or4_1
X_1308_ net47 _0101_ _0285_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1024_ _0074_ _0075_ _0149_ _0196_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0808_ net117 net79 net71 net113 VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__a22o_2
X_0739_ net130 net127 net132 net134 VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_2 _0039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1007_ _0706_ _0056_ _0304_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1410_ _0208_ _0683_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1341_ net135 net155 net42 _0618_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__a22o_1
X_1272_ _0237_ _0242_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__or2_1
X_0987_ _0048_ _0052_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout103 _0693_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__buf_2
Xfanout114 _0677_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
Xfanout125 addr0_reg\[4\] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
Xfanout136 _0648_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__buf_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0910_ net126 net120 net122 net124 VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_7_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0772_ net113 net79 net71 net117 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0841_ _0131_ _0136_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1186_ net137 net161 net44 _0475_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1324_ _0217_ _0599_ _0600_ _0602_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__or4_1
X_1255_ _0049_ _0085_ _0237_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_3_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1040_ _0691_ _0699_ _0055_ _0308_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0824_ _0121_ _0122_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0755_ _0049_ _0052_ _0053_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__or3_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1169_ _0147_ _0154_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__or2_1
X_1307_ _0072_ _0081_ _0182_ _0183_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__or4_1
X_1238_ _0698_ _0130_ _0285_ _0355_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1023_ _0109_ _0220_ _0232_ _0235_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__or4_1
X_0738_ net129 net128 net131 net134 VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_31_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0807_ net104 net79 net71 net102 VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_3 _0044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1006_ _0186_ _0187_ _0237_ _0240_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput40 net40 VGND VGND VPWR VPWR dout0[8] sky130_fd_sc_hd__buf_2
XFILLER_0_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1340_ _0609_ _0612_ _0617_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1271_ _0093_ _0098_ _0129_ _0174_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__or4_2
XFILLER_0_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0986_ _0699_ _0702_ _0705_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__or3_2
Xfanout137 _0648_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_2
Xfanout104 _0692_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_4
Xfanout126 addr0_reg\[4\] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
Xfanout115 _0668_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_2
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0840_ net108 net79 net71 net106 VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__a22o_2
X_0771_ net125 net123 net119 net121 VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__and4b_1
X_1323_ _0341_ _0485_ _0503_ _0601_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__or4_1
X_1185_ _0468_ _0471_ _0474_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__or3_1
X_1254_ _0189_ _0272_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0969_ net97 net58 net55 net99 VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0823_ net85 net78 net76 net81 VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__a22o_2
X_0754_ net110 net85 net81 net115 VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_24_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1306_ _0066_ _0067_ _0152_ _0585_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1237_ _0477_ _0520_ _0521_ _0522_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__or4_1
X_1099_ _0212_ _0225_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__or2_1
X_1168_ _0110_ _0113_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__or2_2
XFILLER_0_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_2_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_45_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1022_ _0115_ _0316_ _0319_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0737_ net115 net94 net92 net110 VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__a22o_2
X_0806_ _0103_ _0104_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 _0044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1005_ net163 net138 net45 _0303_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput41 net41 VGND VGND VPWR VPWR dout0[9] sky130_fd_sc_hd__buf_2
Xoutput30 net30 VGND VGND VPWR VPWR dout0[28] sky130_fd_sc_hd__buf_2
XFILLER_0_37_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
.ends

