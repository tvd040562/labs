assign table_[  0] = 32'H00000000;
assign table_[  1] = 32'H03242abf;
assign table_[  2] = 32'H0647d97c;
assign table_[  3] = 32'H096a9049;
assign table_[  4] = 32'H0c8bd35e;
assign table_[  5] = 32'H0fab272b;
assign table_[  6] = 32'H12c8106e;
assign table_[  7] = 32'H15e21444;
assign table_[  8] = 32'H18f8b83c;
assign table_[  9] = 32'H1c0b826a;
assign table_[ 10] = 32'H1f19f97b;
assign table_[ 11] = 32'H2223a4c5;
assign table_[ 12] = 32'H25280c5d;
assign table_[ 13] = 32'H2826b928;
assign table_[ 14] = 32'H2b1f34eb;
assign table_[ 15] = 32'H2e110a62;
assign table_[ 16] = 32'H30fbc54d;
assign table_[ 17] = 32'H33def287;
assign table_[ 18] = 32'H36ba2013;
assign table_[ 19] = 32'H398cdd32;
assign table_[ 20] = 32'H3c56ba70;
assign table_[ 21] = 32'H3f1749b7;
assign table_[ 22] = 32'H41ce1e64;
assign table_[ 23] = 32'H447acd50;
assign table_[ 24] = 32'H471cece6;
assign table_[ 25] = 32'H49b41533;
assign table_[ 26] = 32'H4c3fdff3;
assign table_[ 27] = 32'H4ebfe8a4;
assign table_[ 28] = 32'H5133cc94;
assign table_[ 29] = 32'H539b2aef;
assign table_[ 30] = 32'H55f5a4d2;
assign table_[ 31] = 32'H5842dd54;
assign table_[ 32] = 32'H5a827999;
assign table_[ 33] = 32'H5cb420df;
assign table_[ 34] = 32'H5ed77c89;
assign table_[ 35] = 32'H60ec382f;
assign table_[ 36] = 32'H62f201ac;
assign table_[ 37] = 32'H64e88925;
assign table_[ 38] = 32'H66cf811f;
assign table_[ 39] = 32'H68a69e80;
assign table_[ 40] = 32'H6a6d98a3;
assign table_[ 41] = 32'H6c24295f;
assign table_[ 42] = 32'H6dca0d14;
assign table_[ 43] = 32'H6f5f02b1;
assign table_[ 44] = 32'H70e2cbc5;
assign table_[ 45] = 32'H72552c84;
assign table_[ 46] = 32'H73b5ebd0;
assign table_[ 47] = 32'H7504d344;
assign table_[ 48] = 32'H7641af3c;
assign table_[ 49] = 32'H776c4eda;
assign table_[ 50] = 32'H78848413;
assign table_[ 51] = 32'H798a23b0;
assign table_[ 52] = 32'H7a7d055a;
assign table_[ 53] = 32'H7b5d039d;
assign table_[ 54] = 32'H7c29fbed;
assign table_[ 55] = 32'H7ce3ceb1;
assign table_[ 56] = 32'H7d8a5f3f;
assign table_[ 57] = 32'H7e1d93e9;
assign table_[ 58] = 32'H7e9d55fb;
assign table_[ 59] = 32'H7f0991c3;
assign table_[ 60] = 32'H7f62368e;
assign table_[ 61] = 32'H7fa736b3;
assign table_[ 62] = 32'H7fd8878d;
assign table_[ 63] = 32'H7ff62181;
assign table_[ 64] = 32'H7fffffff;
assign table_[ 65] = 32'H7ff62181;
assign table_[ 66] = 32'H7fd8878d;
assign table_[ 67] = 32'H7fa736b3;
assign table_[ 68] = 32'H7f62368e;
assign table_[ 69] = 32'H7f0991c3;
assign table_[ 70] = 32'H7e9d55fb;
assign table_[ 71] = 32'H7e1d93e9;
assign table_[ 72] = 32'H7d8a5f3f;
assign table_[ 73] = 32'H7ce3ceb1;
assign table_[ 74] = 32'H7c29fbed;
assign table_[ 75] = 32'H7b5d039d;
assign table_[ 76] = 32'H7a7d055a;
assign table_[ 77] = 32'H798a23b0;
assign table_[ 78] = 32'H78848413;
assign table_[ 79] = 32'H776c4eda;
assign table_[ 80] = 32'H7641af3c;
assign table_[ 81] = 32'H7504d344;
assign table_[ 82] = 32'H73b5ebd0;
assign table_[ 83] = 32'H72552c84;
assign table_[ 84] = 32'H70e2cbc5;
assign table_[ 85] = 32'H6f5f02b1;
assign table_[ 86] = 32'H6dca0d14;
assign table_[ 87] = 32'H6c24295f;
assign table_[ 88] = 32'H6a6d98a3;
assign table_[ 89] = 32'H68a69e80;
assign table_[ 90] = 32'H66cf811f;
assign table_[ 91] = 32'H64e88925;
assign table_[ 92] = 32'H62f201ac;
assign table_[ 93] = 32'H60ec382f;
assign table_[ 94] = 32'H5ed77c89;
assign table_[ 95] = 32'H5cb420df;
assign table_[ 96] = 32'H5a827999;
assign table_[ 97] = 32'H5842dd54;
assign table_[ 98] = 32'H55f5a4d2;
assign table_[ 99] = 32'H539b2aef;
assign table_[100] = 32'H5133cc94;
assign table_[101] = 32'H4ebfe8a4;
assign table_[102] = 32'H4c3fdff3;
assign table_[103] = 32'H49b41533;
assign table_[104] = 32'H471cece6;
assign table_[105] = 32'H447acd50;
assign table_[106] = 32'H41ce1e64;
assign table_[107] = 32'H3f1749b7;
assign table_[108] = 32'H3c56ba70;
assign table_[109] = 32'H398cdd32;
assign table_[110] = 32'H36ba2013;
assign table_[111] = 32'H33def287;
assign table_[112] = 32'H30fbc54d;
assign table_[113] = 32'H2e110a62;
assign table_[114] = 32'H2b1f34eb;
assign table_[115] = 32'H2826b928;
assign table_[116] = 32'H25280c5d;
assign table_[117] = 32'H2223a4c5;
assign table_[118] = 32'H1f19f97b;
assign table_[119] = 32'H1c0b826a;
assign table_[120] = 32'H18f8b83c;
assign table_[121] = 32'H15e21444;
assign table_[122] = 32'H12c8106e;
assign table_[123] = 32'H0fab272b;
assign table_[124] = 32'H0c8bd35e;
assign table_[125] = 32'H096a9049;
assign table_[126] = 32'H0647d97c;
assign table_[127] = 32'H03242abf;
assign table_[128] = 32'H00000000;
assign table_[129] = 32'Hfcdbd541;
assign table_[130] = 32'Hf9b82684;
assign table_[131] = 32'Hf6956fb7;
assign table_[132] = 32'Hf3742ca2;
assign table_[133] = 32'Hf054d8d5;
assign table_[134] = 32'Hed37ef92;
assign table_[135] = 32'Hea1debbc;
assign table_[136] = 32'He70747c4;
assign table_[137] = 32'He3f47d96;
assign table_[138] = 32'He0e60685;
assign table_[139] = 32'Hdddc5b3b;
assign table_[140] = 32'Hdad7f3a3;
assign table_[141] = 32'Hd7d946d8;
assign table_[142] = 32'Hd4e0cb15;
assign table_[143] = 32'Hd1eef59e;
assign table_[144] = 32'Hcf043ab3;
assign table_[145] = 32'Hcc210d79;
assign table_[146] = 32'Hc945dfed;
assign table_[147] = 32'Hc67322ce;
assign table_[148] = 32'Hc3a94590;
assign table_[149] = 32'Hc0e8b649;
assign table_[150] = 32'Hbe31e19c;
assign table_[151] = 32'Hbb8532b0;
assign table_[152] = 32'Hb8e3131a;
assign table_[153] = 32'Hb64beacd;
assign table_[154] = 32'Hb3c0200d;
assign table_[155] = 32'Hb140175c;
assign table_[156] = 32'Haecc336c;
assign table_[157] = 32'Hac64d511;
assign table_[158] = 32'Haa0a5b2e;
assign table_[159] = 32'Ha7bd22ac;
assign table_[160] = 32'Ha57d8667;
assign table_[161] = 32'Ha34bdf21;
assign table_[162] = 32'Ha1288377;
assign table_[163] = 32'H9f13c7d1;
assign table_[164] = 32'H9d0dfe54;
assign table_[165] = 32'H9b1776db;
assign table_[166] = 32'H99307ee1;
assign table_[167] = 32'H97596180;
assign table_[168] = 32'H9592675d;
assign table_[169] = 32'H93dbd6a1;
assign table_[170] = 32'H9235f2ec;
assign table_[171] = 32'H90a0fd4f;
assign table_[172] = 32'H8f1d343b;
assign table_[173] = 32'H8daad37c;
assign table_[174] = 32'H8c4a1430;
assign table_[175] = 32'H8afb2cbc;
assign table_[176] = 32'H89be50c4;
assign table_[177] = 32'H8893b126;
assign table_[178] = 32'H877b7bed;
assign table_[179] = 32'H8675dc50;
assign table_[180] = 32'H8582faa6;
assign table_[181] = 32'H84a2fc63;
assign table_[182] = 32'H83d60413;
assign table_[183] = 32'H831c314f;
assign table_[184] = 32'H8275a0c1;
assign table_[185] = 32'H81e26c17;
assign table_[186] = 32'H8162aa05;
assign table_[187] = 32'H80f66e3d;
assign table_[188] = 32'H809dc972;
assign table_[189] = 32'H8058c94d;
assign table_[190] = 32'H80277873;
assign table_[191] = 32'H8009de7f;
assign table_[192] = 32'H80000001;
assign table_[193] = 32'H8009de7f;
assign table_[194] = 32'H80277873;
assign table_[195] = 32'H8058c94d;
assign table_[196] = 32'H809dc972;
assign table_[197] = 32'H80f66e3d;
assign table_[198] = 32'H8162aa05;
assign table_[199] = 32'H81e26c17;
assign table_[200] = 32'H8275a0c1;
assign table_[201] = 32'H831c314f;
assign table_[202] = 32'H83d60413;
assign table_[203] = 32'H84a2fc63;
assign table_[204] = 32'H8582faa6;
assign table_[205] = 32'H8675dc50;
assign table_[206] = 32'H877b7bed;
assign table_[207] = 32'H8893b126;
assign table_[208] = 32'H89be50c4;
assign table_[209] = 32'H8afb2cbc;
assign table_[210] = 32'H8c4a1430;
assign table_[211] = 32'H8daad37c;
assign table_[212] = 32'H8f1d343b;
assign table_[213] = 32'H90a0fd4f;
assign table_[214] = 32'H9235f2ec;
assign table_[215] = 32'H93dbd6a1;
assign table_[216] = 32'H9592675d;
assign table_[217] = 32'H97596180;
assign table_[218] = 32'H99307ee1;
assign table_[219] = 32'H9b1776db;
assign table_[220] = 32'H9d0dfe54;
assign table_[221] = 32'H9f13c7d1;
assign table_[222] = 32'Ha1288377;
assign table_[223] = 32'Ha34bdf21;
assign table_[224] = 32'Ha57d8667;
assign table_[225] = 32'Ha7bd22ac;
assign table_[226] = 32'Haa0a5b2e;
assign table_[227] = 32'Hac64d511;
assign table_[228] = 32'Haecc336c;
assign table_[229] = 32'Hb140175c;
assign table_[230] = 32'Hb3c0200d;
assign table_[231] = 32'Hb64beacd;
assign table_[232] = 32'Hb8e3131a;
assign table_[233] = 32'Hbb8532b0;
assign table_[234] = 32'Hbe31e19c;
assign table_[235] = 32'Hc0e8b649;
assign table_[236] = 32'Hc3a94590;
assign table_[237] = 32'Hc67322ce;
assign table_[238] = 32'Hc945dfed;
assign table_[239] = 32'Hcc210d79;
assign table_[240] = 32'Hcf043ab3;
assign table_[241] = 32'Hd1eef59e;
assign table_[242] = 32'Hd4e0cb15;
assign table_[243] = 32'Hd7d946d8;
assign table_[244] = 32'Hdad7f3a3;
assign table_[245] = 32'Hdddc5b3b;
assign table_[246] = 32'He0e60685;
assign table_[247] = 32'He3f47d96;
assign table_[248] = 32'He70747c4;
assign table_[249] = 32'Hea1debbc;
assign table_[250] = 32'Hed37ef92;
assign table_[251] = 32'Hf054d8d5;
assign table_[252] = 32'Hf3742ca2;
assign table_[253] = 32'Hf6956fb7;
assign table_[254] = 32'Hf9b82684;
assign table_[255] = 32'Hfcdbd541;
