VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cust_rom
  CLASS BLOCK ;
  FOREIGN cust_rom ;
  ORIGIN 0.000 0.000 ;
  SIZE 152.730 BY 163.450 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 152.560 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 152.560 ;
    END
  END VPWR
  PIN addr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END addr0[7]
  PIN clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END clk0
  PIN cs0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 148.730 20.440 152.730 21.040 ;
    END
  END cs0
  PIN dout0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 159.450 77.650 163.450 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 159.450 84.090 163.450 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 148.730 122.440 152.730 123.040 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 148.730 54.440 152.730 55.040 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 159.450 61.550 163.450 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 148.730 64.640 152.730 65.240 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 159.450 106.630 163.450 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 159.450 71.210 163.450 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 159.450 55.110 163.450 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 159.450 32.570 163.450 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 159.450 45.450 163.450 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 148.730 85.040 152.730 85.640 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 159.450 42.230 163.450 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 159.450 29.350 163.450 ;
    END
  END dout0[31]
  PIN dout0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END dout0[3]
  PIN dout0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 159.450 122.730 163.450 ;
    END
  END dout0[4]
  PIN dout0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 148.730 74.840 152.730 75.440 ;
    END
  END dout0[5]
  PIN dout0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 148.730 105.440 152.730 106.040 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 148.730 95.240 152.730 95.840 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 159.450 93.750 163.450 ;
    END
  END dout0[9]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 147.390 152.405 ;
      LAYER li1 ;
        RECT 5.520 10.795 147.200 152.405 ;
      LAYER met1 ;
        RECT 4.210 10.640 147.500 152.560 ;
      LAYER met2 ;
        RECT 4.230 159.170 28.790 160.210 ;
        RECT 29.630 159.170 32.010 160.210 ;
        RECT 32.850 159.170 41.670 160.210 ;
        RECT 42.510 159.170 44.890 160.210 ;
        RECT 45.730 159.170 54.550 160.210 ;
        RECT 55.390 159.170 60.990 160.210 ;
        RECT 61.830 159.170 70.650 160.210 ;
        RECT 71.490 159.170 77.090 160.210 ;
        RECT 77.930 159.170 83.530 160.210 ;
        RECT 84.370 159.170 93.190 160.210 ;
        RECT 94.030 159.170 106.070 160.210 ;
        RECT 106.910 159.170 122.170 160.210 ;
        RECT 123.010 159.170 146.190 160.210 ;
        RECT 4.230 4.280 146.190 159.170 ;
        RECT 4.230 4.000 22.350 4.280 ;
        RECT 23.190 4.000 57.770 4.280 ;
        RECT 58.610 4.000 73.870 4.280 ;
        RECT 74.710 4.000 83.530 4.280 ;
        RECT 84.370 4.000 93.190 4.280 ;
        RECT 94.030 4.000 106.070 4.280 ;
        RECT 106.910 4.000 146.190 4.280 ;
      LAYER met3 ;
        RECT 3.990 147.240 148.730 152.485 ;
        RECT 4.400 145.840 148.730 147.240 ;
        RECT 3.990 143.840 148.730 145.840 ;
        RECT 4.400 142.440 148.730 143.840 ;
        RECT 3.990 137.040 148.730 142.440 ;
        RECT 4.400 135.640 148.730 137.040 ;
        RECT 3.990 133.640 148.730 135.640 ;
        RECT 4.400 132.240 148.730 133.640 ;
        RECT 3.990 130.240 148.730 132.240 ;
        RECT 4.400 128.840 148.730 130.240 ;
        RECT 3.990 126.840 148.730 128.840 ;
        RECT 4.400 125.440 148.730 126.840 ;
        RECT 3.990 123.440 148.730 125.440 ;
        RECT 3.990 122.040 148.330 123.440 ;
        RECT 3.990 120.040 148.730 122.040 ;
        RECT 4.400 118.640 148.730 120.040 ;
        RECT 3.990 109.840 148.730 118.640 ;
        RECT 4.400 108.440 148.730 109.840 ;
        RECT 3.990 106.440 148.730 108.440 ;
        RECT 3.990 105.040 148.330 106.440 ;
        RECT 3.990 96.240 148.730 105.040 ;
        RECT 3.990 94.840 148.330 96.240 ;
        RECT 3.990 89.440 148.730 94.840 ;
        RECT 4.400 88.040 148.730 89.440 ;
        RECT 3.990 86.040 148.730 88.040 ;
        RECT 3.990 84.640 148.330 86.040 ;
        RECT 3.990 82.640 148.730 84.640 ;
        RECT 4.400 81.240 148.730 82.640 ;
        RECT 3.990 75.840 148.730 81.240 ;
        RECT 3.990 74.440 148.330 75.840 ;
        RECT 3.990 72.440 148.730 74.440 ;
        RECT 4.400 71.040 148.730 72.440 ;
        RECT 3.990 65.640 148.730 71.040 ;
        RECT 4.400 64.240 148.330 65.640 ;
        RECT 3.990 55.440 148.730 64.240 ;
        RECT 4.400 54.040 148.330 55.440 ;
        RECT 3.990 45.240 148.730 54.040 ;
        RECT 4.400 43.840 148.730 45.240 ;
        RECT 3.990 38.440 148.730 43.840 ;
        RECT 4.400 37.040 148.730 38.440 ;
        RECT 3.990 31.640 148.730 37.040 ;
        RECT 4.400 30.240 148.730 31.640 ;
        RECT 3.990 21.440 148.730 30.240 ;
        RECT 3.990 20.040 148.330 21.440 ;
        RECT 3.990 10.715 148.730 20.040 ;
      LAYER met4 ;
        RECT 11.335 23.975 20.640 146.025 ;
        RECT 23.040 23.975 23.940 146.025 ;
        RECT 26.340 23.975 138.625 146.025 ;
      LAYER met5 ;
        RECT 80.620 136.900 131.900 138.500 ;
  END
END cust_rom
END LIBRARY

