assign table3[0] = 32'h80000001;
assign table3[1] = 32'h80009deb;
assign table3[2] = 32'h800277a7;
assign table3[3] = 32'h80058d30;
assign table3[4] = 32'h8009de7f;
assign table3[5] = 32'h800f6b89;
assign table3[6] = 32'h80163441;
assign table3[7] = 32'h801e3896;
assign table3[8] = 32'h80277873;
assign table3[9] = 32'h8031f3c3;
assign table3[10] = 32'h803daa6b;
assign table3[11] = 32'h804a9c4e;
assign table3[12] = 32'h8058c94d;
assign table3[13] = 32'h80683144;
assign table3[14] = 32'h8078d40e;
assign table3[15] = 32'h808ab181;
assign table3[16] = 32'h809dc972;
assign table3[17] = 32'h80b21bb0;
assign table3[18] = 32'h80c7a80b;
assign table3[19] = 32'h80de6e4d;
assign table3[20] = 32'h80f66e3d;
assign table3[21] = 32'h810fa7a1;
assign table3[22] = 32'h812a1a3b;
assign table3[23] = 32'h8145c5c8;
assign table3[24] = 32'h8162aa05;
assign table3[25] = 32'h8180c6aa;
assign table3[26] = 32'h81a01b6e;
assign table3[27] = 32'h81c0a802;
assign table3[28] = 32'h81e26c17;
assign table3[29] = 32'h82056759;
assign table3[30] = 32'h82299972;
assign table3[31] = 32'h824f0209;
assign table3[32] = 32'h8275a0c1;
assign table3[33] = 32'h829d753b;
assign table3[34] = 32'h82c67f15;
assign table3[35] = 32'h82f0bde9;
assign table3[36] = 32'h831c314f;
assign table3[37] = 32'h8348d8dd;
assign table3[38] = 32'h8376b423;
assign table3[39] = 32'h83a5c2b1;
assign table3[40] = 32'h83d60413;
assign table3[41] = 32'h840777d1;
assign table3[42] = 32'h843a1d71;
assign table3[43] = 32'h846df478;
assign table3[44] = 32'h84a2fc63;
assign table3[45] = 32'h84d934b2;
assign table3[46] = 32'h85109cdd;
assign table3[47] = 32'h8549345d;
assign table3[48] = 32'h8582faa6;
assign table3[49] = 32'h85bdef28;
assign table3[50] = 32'h85fa1154;
assign table3[51] = 32'h86376093;
assign table3[52] = 32'h8675dc50;
assign table3[53] = 32'h86b583ef;
assign table3[54] = 32'h86f656d4;
assign table3[55] = 32'h8738545f;
assign table3[56] = 32'h877b7bed;
assign table3[57] = 32'h87bfccd8;
assign table3[58] = 32'h88054678;
assign table3[59] = 32'h884be821;
assign table3[60] = 32'h8893b126;
assign table3[61] = 32'h88dca0d4;
assign table3[62] = 32'h8926b678;
assign table3[63] = 32'h8971f15b;
assign table3[64] = 32'h89be50c4;
assign table3[65] = 32'h8a0bd3f6;
assign table3[66] = 32'h8a5a7a32;
assign table3[67] = 32'h8aaa42b5;
assign table3[68] = 32'h8afb2cbc;
assign table3[69] = 32'h8b4d377d;
assign table3[70] = 32'h8ba06230;
assign table3[71] = 32'h8bf4ac06;
assign table3[72] = 32'h8c4a1430;
assign table3[73] = 32'h8ca099db;
assign table3[74] = 32'h8cf83c31;
assign table3[75] = 32'h8d50fa5a;
assign table3[76] = 32'h8daad37c;
assign table3[77] = 32'h8e05c6b8;
assign table3[78] = 32'h8e61d32f;
assign table3[79] = 32'h8ebef7fc;
assign table3[80] = 32'h8f1d343b;
assign table3[81] = 32'h8f7c8702;
assign table3[82] = 32'h8fdcef67;
assign table3[83] = 32'h903e6c7c;
assign table3[84] = 32'h90a0fd4f;
assign table3[85] = 32'h9104a0ef;
assign table3[86] = 32'h91695664;
assign table3[87] = 32'h91cf1cb7;
assign table3[88] = 32'h9235f2ec;
assign table3[89] = 32'h929dd807;
assign table3[90] = 32'h9306cb05;
assign table3[91] = 32'h9370cae5;
assign table3[92] = 32'h93dbd6a1;
assign table3[93] = 32'h9447ed30;
assign table3[94] = 32'h94b50d88;
assign table3[95] = 32'h9523369c;
assign table3[96] = 32'h9592675d;
assign table3[97] = 32'h96029eb6;
assign table3[98] = 32'h9673db95;
assign table3[99] = 32'h96e61ce1;
assign table3[100] = 32'h97596180;
assign table3[101] = 32'h97cda856;
assign table3[102] = 32'h9842f044;
assign table3[103] = 32'h98b93829;
assign table3[104] = 32'h99307ee1;
assign table3[105] = 32'h99a8c345;
assign table3[106] = 32'h9a22042e;
assign table3[107] = 32'h9a9c406f;
assign table3[108] = 32'h9b1776db;
assign table3[109] = 32'h9b93a641;
assign table3[110] = 32'h9c10cd71;
assign table3[111] = 32'h9c8eeb34;
assign table3[112] = 32'h9d0dfe54;
assign table3[113] = 32'h9d8e0598;
assign table3[114] = 32'h9e0effc2;
assign table3[115] = 32'h9e90eb95;
assign table3[116] = 32'h9f13c7d1;
assign table3[117] = 32'h9f979332;
assign table3[118] = 32'ha01c4c73;
assign table3[119] = 32'ha0a1f24e;
assign table3[120] = 32'ha1288377;
assign table3[121] = 32'ha1affea3;
assign table3[122] = 32'ha2386285;
assign table3[123] = 32'ha2c1adca;
assign table3[124] = 32'ha34bdf21;
assign table3[125] = 32'ha3d6f534;
assign table3[126] = 32'ha462eead;
assign table3[127] = 32'ha4efca32;
assign table3[128] = 32'ha57d8667;
assign table3[129] = 32'ha60c21ee;
assign table3[130] = 32'ha69b9b69;
assign table3[131] = 32'ha72bf174;
assign table3[132] = 32'ha7bd22ac;
assign table3[133] = 32'ha84f2dab;
assign table3[134] = 32'ha8e21107;
assign table3[135] = 32'ha975cb57;
assign table3[136] = 32'haa0a5b2e;
assign table3[137] = 32'haa9fbf1e;
assign table3[138] = 32'hab35f5b6;
assign table3[139] = 32'habccfd83;
assign table3[140] = 32'hac64d511;
assign table3[141] = 32'hacfd7ae9;
assign table3[142] = 32'had96ed92;
assign table3[143] = 32'hae312b92;
assign table3[144] = 32'haecc336c;
assign table3[145] = 32'haf6803a2;
assign table3[146] = 32'hb0049ab4;
assign table3[147] = 32'hb0a1f71e;
assign table3[148] = 32'hb140175c;
assign table3[149] = 32'hb1def9e9;
assign table3[150] = 32'hb27e9d3d;
assign table3[151] = 32'hb31effcc;
assign table3[152] = 32'hb3c0200d;
assign table3[153] = 32'hb461fc71;
assign table3[154] = 32'hb5049369;
assign table3[155] = 32'hb5a7e363;
assign table3[156] = 32'hb64beacd;
assign table3[157] = 32'hb6f0a812;
assign table3[158] = 32'hb796199c;
assign table3[159] = 32'hb83c3dd2;
assign table3[160] = 32'hb8e3131a;
assign table3[161] = 32'hb98a97d9;
assign table3[162] = 32'hba32ca71;
assign table3[163] = 32'hbadba944;
assign table3[164] = 32'hbb8532b0;
assign table3[165] = 32'hbc2f6514;
assign table3[166] = 32'hbcda3ecb;
assign table3[167] = 32'hbd85be30;
assign table3[168] = 32'hbe31e19c;
assign table3[169] = 32'hbedea766;
assign table3[170] = 32'hbf8c0de3;
assign table3[171] = 32'hc03a1369;
assign table3[172] = 32'hc0e8b649;
assign table3[173] = 32'hc197f4d4;
assign table3[174] = 32'hc247cd5b;
assign table3[175] = 32'hc2f83e2b;
assign table3[176] = 32'hc3a94590;
assign table3[177] = 32'hc45ae1d7;
assign table3[178] = 32'hc50d1149;
assign table3[179] = 32'hc5bfd22f;
assign table3[180] = 32'hc67322ce;
assign table3[181] = 32'hc727016d;
assign table3[182] = 32'hc7db6c50;
assign table3[183] = 32'hc89061ba;
assign table3[184] = 32'hc945dfed;
assign table3[185] = 32'hc9fbe527;
assign table3[186] = 32'hcab26faa;
assign table3[187] = 32'hcb697db1;
assign table3[188] = 32'hcc210d79;
assign table3[189] = 32'hccd91d3e;
assign table3[190] = 32'hcd91ab39;
assign table3[191] = 32'hce4ab5a3;
assign table3[192] = 32'hcf043ab3;
assign table3[193] = 32'hcfbe38a0;
assign table3[194] = 32'hd078ad9e;
assign table3[195] = 32'hd13397e2;
assign table3[196] = 32'hd1eef59e;
assign table3[197] = 32'hd2aac505;
assign table3[198] = 32'hd3670446;
assign table3[199] = 32'hd423b191;
assign table3[200] = 32'hd4e0cb15;
assign table3[201] = 32'hd59e4eff;
assign table3[202] = 32'hd65c3b7b;
assign table3[203] = 32'hd71a8eb6;
assign table3[204] = 32'hd7d946d8;
assign table3[205] = 32'hd898620c;
assign table3[206] = 32'hd957de7b;
assign table3[207] = 32'hda17ba4a;
assign table3[208] = 32'hdad7f3a3;
assign table3[209] = 32'hdb9888a9;
assign table3[210] = 32'hdc597782;
assign table3[211] = 32'hdd1abe51;
assign table3[212] = 32'hdddc5b3b;
assign table3[213] = 32'hde9e4c61;
assign table3[214] = 32'hdf608fe4;
assign table3[215] = 32'he02323e5;
assign table3[216] = 32'he0e60685;
assign table3[217] = 32'he1a935e2;
assign table3[218] = 32'he26cb01b;
assign table3[219] = 32'he330734d;
assign table3[220] = 32'he3f47d96;
assign table3[221] = 32'he4b8cd11;
assign table3[222] = 32'he57d5fdb;
assign table3[223] = 32'he642340d;
assign table3[224] = 32'he70747c4;
assign table3[225] = 32'he7cc9918;
assign table3[226] = 32'he8922622;
assign table3[227] = 32'he957ecfb;
assign table3[228] = 32'hea1debbc;
assign table3[229] = 32'heae4207b;
assign table3[230] = 32'hebaa894f;
assign table3[231] = 32'hec71244f;
assign table3[232] = 32'hed37ef92;
assign table3[233] = 32'hedfee92b;
assign table3[234] = 32'heec60f31;
assign table3[235] = 32'hef8d5fb8;
assign table3[236] = 32'hf054d8d5;
assign table3[237] = 32'hf11c789a;
assign table3[238] = 32'hf1e43d1c;
assign table3[239] = 32'hf2ac246e;
assign table3[240] = 32'hf3742ca2;
assign table3[241] = 32'hf43c53cb;
assign table3[242] = 32'hf50497fb;
assign table3[243] = 32'hf5ccf744;
assign table3[244] = 32'hf6956fb7;
assign table3[245] = 32'hf75dff66;
assign table3[246] = 32'hf826a462;
assign table3[247] = 32'hf8ef5cbb;
assign table3[248] = 32'hf9b82684;
assign table3[249] = 32'hfa80ffcb;
assign table3[250] = 32'hfb49e6a3;
assign table3[251] = 32'hfc12d91a;
assign table3[252] = 32'hfcdbd541;
assign table3[253] = 32'hfda4d929;
assign table3[254] = 32'hfe6de2e0;
assign table3[255] = 32'hff36f078;
