assign table0[0] = 32'h00000000;
assign table0[1] = 32'h00c90e90;
assign table0[2] = 32'h0192155f;
assign table0[3] = 32'h025b0caf;
assign table0[4] = 32'h0323ecbe;
assign table0[5] = 32'h03ecadcf;
assign table0[6] = 32'h04b54825;
assign table0[7] = 32'h057db403;
assign table0[8] = 32'h0645e9af;
assign table0[9] = 32'h070de172;
assign table0[10] = 32'h07d59396;
assign table0[11] = 32'h089cf867;
assign table0[12] = 32'h09640837;
assign table0[13] = 32'h0a2abb59;
assign table0[14] = 32'h0af10a22;
assign table0[15] = 32'h0bb6ecef;
assign table0[16] = 32'h0c7c5c1e;
assign table0[17] = 32'h0d415013;
assign table0[18] = 32'h0e05c135;
assign table0[19] = 32'h0ec9a7f3;
assign table0[20] = 32'h0f8cfcbe;
assign table0[21] = 32'h104fb80e;
assign table0[22] = 32'h1111d263;
assign table0[23] = 32'h11d3443f;
assign table0[24] = 32'h1294062f;
assign table0[25] = 32'h135410c3;
assign table0[26] = 32'h14135c94;
assign table0[27] = 32'h14d1e242;
assign table0[28] = 32'h158f9a76;
assign table0[29] = 32'h164c7ddd;
assign table0[30] = 32'h17088531;
assign table0[31] = 32'h17c3a931;
assign table0[32] = 32'h187de2a7;
assign table0[33] = 32'h19372a64;
assign table0[34] = 32'h19ef7944;
assign table0[35] = 32'h1aa6c82b;
assign table0[36] = 32'h1b5d100a;
assign table0[37] = 32'h1c1249d8;
assign table0[38] = 32'h1cc66e99;
assign table0[39] = 32'h1d79775c;
assign table0[40] = 32'h1e2b5d38;
assign table0[41] = 32'h1edc1953;
assign table0[42] = 32'h1f8ba4dc;
assign table0[43] = 32'h2039f90f;
assign table0[44] = 32'h20e70f32;
assign table0[45] = 32'h2192e09b;
assign table0[46] = 32'h223d66a8;
assign table0[47] = 32'h22e69ac8;
assign table0[48] = 32'h238e7673;
assign table0[49] = 32'h2434f332;
assign table0[50] = 32'h24da0a9a;
assign table0[51] = 32'h257db64c;
assign table0[52] = 32'h261feffa;
assign table0[53] = 32'h26c0b162;
assign table0[54] = 32'h275ff452;
assign table0[55] = 32'h27fdb2a7;
assign table0[56] = 32'h2899e64a;
assign table0[57] = 32'h29348937;
assign table0[58] = 32'h29cd9578;
assign table0[59] = 32'h2a650525;
assign table0[60] = 32'h2afad269;
assign table0[61] = 32'h2b8ef77d;
assign table0[62] = 32'h2c216eaa;
assign table0[63] = 32'h2cb2324c;
assign table0[64] = 32'h2d413ccd;
assign table0[65] = 32'h2dce88aa;
assign table0[66] = 32'h2e5a1070;
assign table0[67] = 32'h2ee3cebe;
assign table0[68] = 32'h2f6bbe45;
assign table0[69] = 32'h2ff1d9c7;
assign table0[70] = 32'h30761c18;
assign table0[71] = 32'h30f8801f;
assign table0[72] = 32'h317900d6;
assign table0[73] = 32'h31f79948;
assign table0[74] = 32'h32744493;
assign table0[75] = 32'h32eefdea;
assign table0[76] = 32'h3367c090;
assign table0[77] = 32'h33de87de;
assign table0[78] = 32'h34534f41;
assign table0[79] = 32'h34c61236;
assign table0[80] = 32'h3536cc52;
assign table0[81] = 32'h35a5793c;
assign table0[82] = 32'h361214b0;
assign table0[83] = 32'h367c9a7e;
assign table0[84] = 32'h36e5068a;
assign table0[85] = 32'h374b54ce;
assign table0[86] = 32'h37af8159;
assign table0[87] = 32'h3811884d;
assign table0[88] = 32'h387165e3;
assign table0[89] = 32'h38cf1669;
assign table0[90] = 32'h392a9642;
assign table0[91] = 32'h3983e1e8;
assign table0[92] = 32'h39daf5e8;
assign table0[93] = 32'h3a2fcee8;
assign table0[94] = 32'h3a8269a3;
assign table0[95] = 32'h3ad2c2e8;
assign table0[96] = 32'h3b20d79e;
assign table0[97] = 32'h3b6ca4c4;
assign table0[98] = 32'h3bb6276e;
assign table0[99] = 32'h3bfd5cc4;
assign table0[100] = 32'h3c42420a;
assign table0[101] = 32'h3c84d496;
assign table0[102] = 32'h3cc511d9;
assign table0[103] = 32'h3d02f757;
assign table0[104] = 32'h3d3e82ae;
assign table0[105] = 32'h3d77b192;
assign table0[106] = 32'h3dae81cf;
assign table0[107] = 32'h3de2f148;
assign table0[108] = 32'h3e14fdf7;
assign table0[109] = 32'h3e44a5ef;
assign table0[110] = 32'h3e71e759;
assign table0[111] = 32'h3e9cc076;
assign table0[112] = 32'h3ec52fa0;
assign table0[113] = 32'h3eeb3347;
assign table0[114] = 32'h3f0ec9f5;
assign table0[115] = 32'h3f2ff24a;
assign table0[116] = 32'h3f4eaafe;
assign table0[117] = 32'h3f6af2e3;
assign table0[118] = 32'h3f84c8e2;
assign table0[119] = 32'h3f9c2bfb;
assign table0[120] = 32'h3fb11b48;
assign table0[121] = 32'h3fc395f9;
assign table0[122] = 32'h3fd39b5a;
assign table0[123] = 32'h3fe12acb;
assign table0[124] = 32'h3fec43c7;
assign table0[125] = 32'h3ff4e5e0;
assign table0[126] = 32'h3ffb10c1;
assign table0[127] = 32'h3ffec42d;
assign table0[128] = 32'h40000000;
assign table0[129] = 32'h3ffec42d;
assign table0[130] = 32'h3ffb10c1;
assign table0[131] = 32'h3ff4e5e0;
assign table0[132] = 32'h3fec43c7;
assign table0[133] = 32'h3fe12acb;
assign table0[134] = 32'h3fd39b5a;
assign table0[135] = 32'h3fc395f9;
assign table0[136] = 32'h3fb11b48;
assign table0[137] = 32'h3f9c2bfb;
assign table0[138] = 32'h3f84c8e2;
assign table0[139] = 32'h3f6af2e3;
assign table0[140] = 32'h3f4eaafe;
assign table0[141] = 32'h3f2ff24a;
assign table0[142] = 32'h3f0ec9f5;
assign table0[143] = 32'h3eeb3347;
assign table0[144] = 32'h3ec52fa0;
assign table0[145] = 32'h3e9cc076;
assign table0[146] = 32'h3e71e759;
assign table0[147] = 32'h3e44a5ef;
assign table0[148] = 32'h3e14fdf7;
assign table0[149] = 32'h3de2f148;
assign table0[150] = 32'h3dae81cf;
assign table0[151] = 32'h3d77b192;
assign table0[152] = 32'h3d3e82ae;
assign table0[153] = 32'h3d02f757;
assign table0[154] = 32'h3cc511d9;
assign table0[155] = 32'h3c84d496;
assign table0[156] = 32'h3c42420a;
assign table0[157] = 32'h3bfd5cc4;
assign table0[158] = 32'h3bb6276e;
assign table0[159] = 32'h3b6ca4c4;
assign table0[160] = 32'h3b20d79e;
assign table0[161] = 32'h3ad2c2e8;
assign table0[162] = 32'h3a8269a3;
assign table0[163] = 32'h3a2fcee8;
assign table0[164] = 32'h39daf5e8;
assign table0[165] = 32'h3983e1e8;
assign table0[166] = 32'h392a9642;
assign table0[167] = 32'h38cf1669;
assign table0[168] = 32'h387165e3;
assign table0[169] = 32'h3811884d;
assign table0[170] = 32'h37af8159;
assign table0[171] = 32'h374b54ce;
assign table0[172] = 32'h36e5068a;
assign table0[173] = 32'h367c9a7e;
assign table0[174] = 32'h361214b0;
assign table0[175] = 32'h35a5793c;
assign table0[176] = 32'h3536cc52;
assign table0[177] = 32'h34c61236;
assign table0[178] = 32'h34534f41;
assign table0[179] = 32'h33de87de;
assign table0[180] = 32'h3367c090;
assign table0[181] = 32'h32eefdea;
assign table0[182] = 32'h32744493;
assign table0[183] = 32'h31f79948;
assign table0[184] = 32'h317900d6;
assign table0[185] = 32'h30f8801f;
assign table0[186] = 32'h30761c18;
assign table0[187] = 32'h2ff1d9c7;
assign table0[188] = 32'h2f6bbe45;
assign table0[189] = 32'h2ee3cebe;
assign table0[190] = 32'h2e5a1070;
assign table0[191] = 32'h2dce88aa;
assign table0[192] = 32'h2d413ccd;
assign table0[193] = 32'h2cb2324c;
assign table0[194] = 32'h2c216eaa;
assign table0[195] = 32'h2b8ef77d;
assign table0[196] = 32'h2afad269;
assign table0[197] = 32'h2a650525;
assign table0[198] = 32'h29cd9578;
assign table0[199] = 32'h29348937;
assign table0[200] = 32'h2899e64a;
assign table0[201] = 32'h27fdb2a7;
assign table0[202] = 32'h275ff452;
assign table0[203] = 32'h26c0b162;
assign table0[204] = 32'h261feffa;
assign table0[205] = 32'h257db64c;
assign table0[206] = 32'h24da0a9a;
assign table0[207] = 32'h2434f332;
assign table0[208] = 32'h238e7673;
assign table0[209] = 32'h22e69ac8;
assign table0[210] = 32'h223d66a8;
assign table0[211] = 32'h2192e09b;
assign table0[212] = 32'h20e70f32;
assign table0[213] = 32'h2039f90f;
assign table0[214] = 32'h1f8ba4dc;
assign table0[215] = 32'h1edc1953;
assign table0[216] = 32'h1e2b5d38;
assign table0[217] = 32'h1d79775c;
assign table0[218] = 32'h1cc66e99;
assign table0[219] = 32'h1c1249d8;
assign table0[220] = 32'h1b5d100a;
assign table0[221] = 32'h1aa6c82b;
assign table0[222] = 32'h19ef7944;
assign table0[223] = 32'h19372a64;
assign table0[224] = 32'h187de2a7;
assign table0[225] = 32'h17c3a931;
assign table0[226] = 32'h17088531;
assign table0[227] = 32'h164c7ddd;
assign table0[228] = 32'h158f9a76;
assign table0[229] = 32'h14d1e242;
assign table0[230] = 32'h14135c94;
assign table0[231] = 32'h135410c3;
assign table0[232] = 32'h1294062f;
assign table0[233] = 32'h11d3443f;
assign table0[234] = 32'h1111d263;
assign table0[235] = 32'h104fb80e;
assign table0[236] = 32'h0f8cfcbe;
assign table0[237] = 32'h0ec9a7f3;
assign table0[238] = 32'h0e05c135;
assign table0[239] = 32'h0d415013;
assign table0[240] = 32'h0c7c5c1e;
assign table0[241] = 32'h0bb6ecef;
assign table0[242] = 32'h0af10a22;
assign table0[243] = 32'h0a2abb59;
assign table0[244] = 32'h09640837;
assign table0[245] = 32'h089cf867;
assign table0[246] = 32'h07d59396;
assign table0[247] = 32'h070de172;
assign table0[248] = 32'h0645e9af;
assign table0[249] = 32'h057db403;
assign table0[250] = 32'h04b54825;
assign table0[251] = 32'h03ecadcf;
assign table0[252] = 32'h0323ecbe;
assign table0[253] = 32'h025b0caf;
assign table0[254] = 32'h0192155f;
assign table0[255] = 32'h00c90e90;
