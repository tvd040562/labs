assign table0[0] = 32'h00000000;
assign table0[1] = 32'h00c90f88;
assign table0[2] = 32'h01921d20;
assign table0[3] = 32'h025b26d7;
assign table0[4] = 32'h03242abf;
assign table0[5] = 32'h03ed26e6;
assign table0[6] = 32'h04b6195d;
assign table0[7] = 32'h057f0035;
assign table0[8] = 32'h0647d97c;
assign table0[9] = 32'h0710a345;
assign table0[10] = 32'h07d95b9e;
assign table0[11] = 32'h08a2009a;
assign table0[12] = 32'h096a9049;
assign table0[13] = 32'h0a3308bc;
assign table0[14] = 32'h0afb6805;
assign table0[15] = 32'h0bc3ac35;
assign table0[16] = 32'h0c8bd35e;
assign table0[17] = 32'h0d53db92;
assign table0[18] = 32'h0e1bc2e4;
assign table0[19] = 32'h0ee38766;
assign table0[20] = 32'h0fab272b;
assign table0[21] = 32'h1072a048;
assign table0[22] = 32'h1139f0cf;
assign table0[23] = 32'h120116d5;
assign table0[24] = 32'h12c8106e;
assign table0[25] = 32'h138edbb1;
assign table0[26] = 32'h145576b1;
assign table0[27] = 32'h151bdf85;
assign table0[28] = 32'h15e21444;
assign table0[29] = 32'h16a81305;
assign table0[30] = 32'h176dd9de;
assign table0[31] = 32'h183366e8;
assign table0[32] = 32'h18f8b83c;
assign table0[33] = 32'h19bdcbf3;
assign table0[34] = 32'h1a82a025;
assign table0[35] = 32'h1b4732ef;
assign table0[36] = 32'h1c0b826a;
assign table0[37] = 32'h1ccf8cb3;
assign table0[38] = 32'h1d934fe5;
assign table0[39] = 32'h1e56ca1e;
assign table0[40] = 32'h1f19f97b;
assign table0[41] = 32'h1fdcdc1b;
assign table0[42] = 32'h209f701c;
assign table0[43] = 32'h2161b39f;
assign table0[44] = 32'h2223a4c5;
assign table0[45] = 32'h22e541af;
assign table0[46] = 32'h23a6887e;
assign table0[47] = 32'h24677757;
assign table0[48] = 32'h25280c5d;
assign table0[49] = 32'h25e845b6;
assign table0[50] = 32'h26a82185;
assign table0[51] = 32'h27679df4;
assign table0[52] = 32'h2826b928;
assign table0[53] = 32'h28e5714a;
assign table0[54] = 32'h29a3c485;
assign table0[55] = 32'h2a61b101;
assign table0[56] = 32'h2b1f34eb;
assign table0[57] = 32'h2bdc4e6f;
assign table0[58] = 32'h2c98fbba;
assign table0[59] = 32'h2d553afb;
assign table0[60] = 32'h2e110a62;
assign table0[61] = 32'h2ecc681e;
assign table0[62] = 32'h2f875262;
assign table0[63] = 32'h3041c760;
assign table0[64] = 32'h30fbc54d;
assign table0[65] = 32'h31b54a5d;
assign table0[66] = 32'h326e54c7;
assign table0[67] = 32'h3326e2c2;
assign table0[68] = 32'h33def287;
assign table0[69] = 32'h3496824f;
assign table0[70] = 32'h354d9056;
assign table0[71] = 32'h36041ad9;
assign table0[72] = 32'h36ba2013;
assign table0[73] = 32'h376f9e46;
assign table0[74] = 32'h382493b0;
assign table0[75] = 32'h38d8fe93;
assign table0[76] = 32'h398cdd32;
assign table0[77] = 32'h3a402dd1;
assign table0[78] = 32'h3af2eeb7;
assign table0[79] = 32'h3ba51e29;
assign table0[80] = 32'h3c56ba70;
assign table0[81] = 32'h3d07c1d5;
assign table0[82] = 32'h3db832a5;
assign table0[83] = 32'h3e680b2c;
assign table0[84] = 32'h3f1749b7;
assign table0[85] = 32'h3fc5ec97;
assign table0[86] = 32'h4073f21d;
assign table0[87] = 32'h4121589a;
assign table0[88] = 32'h41ce1e64;
assign table0[89] = 32'h427a41d0;
assign table0[90] = 32'h4325c135;
assign table0[91] = 32'h43d09aec;
assign table0[92] = 32'h447acd50;
assign table0[93] = 32'h452456bc;
assign table0[94] = 32'h45cd358f;
assign table0[95] = 32'h46756827;
assign table0[96] = 32'h471cece6;
assign table0[97] = 32'h47c3c22e;
assign table0[98] = 32'h4869e664;
assign table0[99] = 32'h490f57ee;
assign table0[100] = 32'h49b41533;
assign table0[101] = 32'h4a581c9d;
assign table0[102] = 32'h4afb6c97;
assign table0[103] = 32'h4b9e038f;
assign table0[104] = 32'h4c3fdff3;
assign table0[105] = 32'h4ce10034;
assign table0[106] = 32'h4d8162c3;
assign table0[107] = 32'h4e210617;
assign table0[108] = 32'h4ebfe8a4;
assign table0[109] = 32'h4f5e08e2;
assign table0[110] = 32'h4ffb654c;
assign table0[111] = 32'h5097fc5e;
assign table0[112] = 32'h5133cc94;
assign table0[113] = 32'h51ced46e;
assign table0[114] = 32'h5269126e;
assign table0[115] = 32'h53028517;
assign table0[116] = 32'h539b2aef;
assign table0[117] = 32'h5433027d;
assign table0[118] = 32'h54ca0a4a;
assign table0[119] = 32'h556040e2;
assign table0[120] = 32'h55f5a4d2;
assign table0[121] = 32'h568a34a9;
assign table0[122] = 32'h571deef9;
assign table0[123] = 32'h57b0d255;
assign table0[124] = 32'h5842dd54;
assign table0[125] = 32'h58d40e8c;
assign table0[126] = 32'h59646497;
assign table0[127] = 32'h59f3de12;
assign table0[128] = 32'h5a827999;
assign table0[129] = 32'h5b1035ce;
assign table0[130] = 32'h5b9d1153;
assign table0[131] = 32'h5c290acc;
assign table0[132] = 32'h5cb420df;
assign table0[133] = 32'h5d3e5236;
assign table0[134] = 32'h5dc79d7b;
assign table0[135] = 32'h5e50015d;
assign table0[136] = 32'h5ed77c89;
assign table0[137] = 32'h5f5e0db2;
assign table0[138] = 32'h5fe3b38d;
assign table0[139] = 32'h60686cce;
assign table0[140] = 32'h60ec382f;
assign table0[141] = 32'h616f146b;
assign table0[142] = 32'h61f1003e;
assign table0[143] = 32'h6271fa68;
assign table0[144] = 32'h62f201ac;
assign table0[145] = 32'h637114cc;
assign table0[146] = 32'h63ef328f;
assign table0[147] = 32'h646c59bf;
assign table0[148] = 32'h64e88925;
assign table0[149] = 32'h6563bf91;
assign table0[150] = 32'h65ddfbd2;
assign table0[151] = 32'h66573cbb;
assign table0[152] = 32'h66cf811f;
assign table0[153] = 32'h6746c7d7;
assign table0[154] = 32'h67bd0fbc;
assign table0[155] = 32'h683257aa;
assign table0[156] = 32'h68a69e80;
assign table0[157] = 32'h6919e31f;
assign table0[158] = 32'h698c246b;
assign table0[159] = 32'h69fd614a;
assign table0[160] = 32'h6a6d98a3;
assign table0[161] = 32'h6adcc964;
assign table0[162] = 32'h6b4af278;
assign table0[163] = 32'h6bb812d0;
assign table0[164] = 32'h6c24295f;
assign table0[165] = 32'h6c8f351b;
assign table0[166] = 32'h6cf934fb;
assign table0[167] = 32'h6d6227f9;
assign table0[168] = 32'h6dca0d14;
assign table0[169] = 32'h6e30e349;
assign table0[170] = 32'h6e96a99c;
assign table0[171] = 32'h6efb5f11;
assign table0[172] = 32'h6f5f02b1;
assign table0[173] = 32'h6fc19384;
assign table0[174] = 32'h70231099;
assign table0[175] = 32'h708378fe;
assign table0[176] = 32'h70e2cbc5;
assign table0[177] = 32'h71410804;
assign table0[178] = 32'h719e2cd1;
assign table0[179] = 32'h71fa3948;
assign table0[180] = 32'h72552c84;
assign table0[181] = 32'h72af05a6;
assign table0[182] = 32'h7307c3cf;
assign table0[183] = 32'h735f6625;
assign table0[184] = 32'h73b5ebd0;
assign table0[185] = 32'h740b53fa;
assign table0[186] = 32'h745f9dd0;
assign table0[187] = 32'h74b2c883;
assign table0[188] = 32'h7504d344;
assign table0[189] = 32'h7555bd4b;
assign table0[190] = 32'h75a585ce;
assign table0[191] = 32'h75f42c0a;
assign table0[192] = 32'h7641af3c;
assign table0[193] = 32'h768e0ea5;
assign table0[194] = 32'h76d94988;
assign table0[195] = 32'h77235f2c;
assign table0[196] = 32'h776c4eda;
assign table0[197] = 32'h77b417df;
assign table0[198] = 32'h77fab988;
assign table0[199] = 32'h78403328;
assign table0[200] = 32'h78848413;
assign table0[201] = 32'h78c7aba1;
assign table0[202] = 32'h7909a92c;
assign table0[203] = 32'h794a7c11;
assign table0[204] = 32'h798a23b0;
assign table0[205] = 32'h79c89f6d;
assign table0[206] = 32'h7a05eeac;
assign table0[207] = 32'h7a4210d8;
assign table0[208] = 32'h7a7d055a;
assign table0[209] = 32'h7ab6cba3;
assign table0[210] = 32'h7aef6323;
assign table0[211] = 32'h7b26cb4e;
assign table0[212] = 32'h7b5d039d;
assign table0[213] = 32'h7b920b88;
assign table0[214] = 32'h7bc5e28f;
assign table0[215] = 32'h7bf8882f;
assign table0[216] = 32'h7c29fbed;
assign table0[217] = 32'h7c5a3d4f;
assign table0[218] = 32'h7c894bdd;
assign table0[219] = 32'h7cb72723;
assign table0[220] = 32'h7ce3ceb1;
assign table0[221] = 32'h7d0f4217;
assign table0[222] = 32'h7d3980eb;
assign table0[223] = 32'h7d628ac5;
assign table0[224] = 32'h7d8a5f3f;
assign table0[225] = 32'h7db0fdf7;
assign table0[226] = 32'h7dd6668e;
assign table0[227] = 32'h7dfa98a7;
assign table0[228] = 32'h7e1d93e9;
assign table0[229] = 32'h7e3f57fe;
assign table0[230] = 32'h7e5fe492;
assign table0[231] = 32'h7e7f3956;
assign table0[232] = 32'h7e9d55fb;
assign table0[233] = 32'h7eba3a38;
assign table0[234] = 32'h7ed5e5c5;
assign table0[235] = 32'h7ef0585f;
assign table0[236] = 32'h7f0991c3;
assign table0[237] = 32'h7f2191b3;
assign table0[238] = 32'h7f3857f5;
assign table0[239] = 32'h7f4de450;
assign table0[240] = 32'h7f62368e;
assign table0[241] = 32'h7f754e7f;
assign table0[242] = 32'h7f872bf2;
assign table0[243] = 32'h7f97cebc;
assign table0[244] = 32'h7fa736b3;
assign table0[245] = 32'h7fb563b2;
assign table0[246] = 32'h7fc25595;
assign table0[247] = 32'h7fce0c3d;
assign table0[248] = 32'h7fd8878d;
assign table0[249] = 32'h7fe1c76a;
assign table0[250] = 32'h7fe9cbbf;
assign table0[251] = 32'h7ff09477;
assign table0[252] = 32'h7ff62181;
assign table0[253] = 32'h7ffa72d0;
assign table0[254] = 32'h7ffd8859;
assign table0[255] = 32'h7fff6215;
